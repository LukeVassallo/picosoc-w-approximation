magic
tech gf180mcuD
magscale 1 10
timestamp 1702204434
<< metal1 >>
rect 69010 77198 69022 77250
rect 69074 77247 69086 77250
rect 70242 77247 70254 77250
rect 69074 77201 70254 77247
rect 69074 77198 69086 77201
rect 70242 77198 70254 77201
rect 70306 77198 70318 77250
rect 75058 77198 75070 77250
rect 75122 77247 75134 77250
rect 75842 77247 75854 77250
rect 75122 77201 75854 77247
rect 75122 77198 75134 77201
rect 75842 77198 75854 77201
rect 75906 77247 75918 77250
rect 76402 77247 76414 77250
rect 75906 77201 76414 77247
rect 75906 77198 75918 77201
rect 76402 77198 76414 77201
rect 76466 77198 76478 77250
rect 50866 77086 50878 77138
rect 50930 77135 50942 77138
rect 51762 77135 51774 77138
rect 50930 77089 51774 77135
rect 50930 77086 50942 77089
rect 51762 77086 51774 77089
rect 51826 77135 51838 77138
rect 52098 77135 52110 77138
rect 51826 77089 52110 77135
rect 51826 77086 51838 77089
rect 52098 77086 52110 77089
rect 52162 77086 52174 77138
rect 66322 77086 66334 77138
rect 66386 77135 66398 77138
rect 67106 77135 67118 77138
rect 66386 77089 67118 77135
rect 66386 77086 66398 77089
rect 67106 77086 67118 77089
rect 67170 77086 67182 77138
rect 67442 77086 67454 77138
rect 67506 77135 67518 77138
rect 68674 77135 68686 77138
rect 67506 77089 68686 77135
rect 67506 77086 67518 77089
rect 68674 77086 68686 77089
rect 68738 77086 68750 77138
rect 42802 76974 42814 77026
rect 42866 77023 42878 77026
rect 43586 77023 43598 77026
rect 42866 76977 43598 77023
rect 42866 76974 42878 76977
rect 43586 76974 43598 76977
rect 43650 76974 43662 77026
rect 45490 76974 45502 77026
rect 45554 77023 45566 77026
rect 46274 77023 46286 77026
rect 45554 76977 46286 77023
rect 45554 76974 45566 76977
rect 46274 76974 46286 76977
rect 46338 76974 46350 77026
rect 47506 76974 47518 77026
rect 47570 77023 47582 77026
rect 48290 77023 48302 77026
rect 47570 76977 48302 77023
rect 47570 76974 47582 76977
rect 48290 76974 48302 76977
rect 48354 76974 48366 77026
rect 48850 76974 48862 77026
rect 48914 77023 48926 77026
rect 50082 77023 50094 77026
rect 48914 76977 50094 77023
rect 48914 76974 48926 76977
rect 50082 76974 50094 76977
rect 50146 76974 50158 77026
rect 51538 76974 51550 77026
rect 51602 77023 51614 77026
rect 52994 77023 53006 77026
rect 51602 76977 53006 77023
rect 51602 76974 51614 76977
rect 52994 76974 53006 76977
rect 53058 76974 53070 77026
rect 60946 76974 60958 77026
rect 61010 77023 61022 77026
rect 61842 77023 61854 77026
rect 61010 76977 61854 77023
rect 61010 76974 61022 76977
rect 61842 76974 61854 76977
rect 61906 76974 61918 77026
rect 62290 76974 62302 77026
rect 62354 77023 62366 77026
rect 63298 77023 63310 77026
rect 62354 76977 63310 77023
rect 62354 76974 62366 76977
rect 63298 76974 63310 76977
rect 63362 76974 63374 77026
rect 64306 76974 64318 77026
rect 64370 77023 64382 77026
rect 65314 77023 65326 77026
rect 64370 76977 65326 77023
rect 64370 76974 64382 76977
rect 65314 76974 65326 76977
rect 65378 76974 65390 77026
rect 65650 76974 65662 77026
rect 65714 77023 65726 77026
rect 66434 77023 66446 77026
rect 65714 76977 66446 77023
rect 65714 76974 65726 76977
rect 66434 76974 66446 76977
rect 66498 76974 66510 77026
rect 67666 76974 67678 77026
rect 67730 77023 67742 77026
rect 68450 77023 68462 77026
rect 67730 76977 68462 77023
rect 67730 76974 67742 76977
rect 68450 76974 68462 76977
rect 68514 76974 68526 77026
rect 71026 76974 71038 77026
rect 71090 77023 71102 77026
rect 71922 77023 71934 77026
rect 71090 76977 71934 77023
rect 71090 76974 71102 76977
rect 71922 76974 71934 76977
rect 71986 77023 71998 77026
rect 72594 77023 72606 77026
rect 71986 76977 72606 77023
rect 71986 76974 71998 76977
rect 72594 76974 72606 76977
rect 72658 76974 72670 77026
rect 74386 76974 74398 77026
rect 74450 77023 74462 77026
rect 75058 77023 75070 77026
rect 74450 76977 75070 77023
rect 74450 76974 74462 76977
rect 75058 76974 75070 76977
rect 75122 77023 75134 77026
rect 75730 77023 75742 77026
rect 75122 76977 75742 77023
rect 75122 76974 75134 76977
rect 75730 76974 75742 76977
rect 75794 76974 75806 77026
rect 76626 76974 76638 77026
rect 76690 77023 76702 77026
rect 77186 77023 77198 77026
rect 76690 76977 77198 77023
rect 76690 76974 76702 76977
rect 77186 76974 77198 76977
rect 77250 76974 77262 77026
rect 1344 76858 78624 76892
rect 1344 76806 19838 76858
rect 19890 76806 19942 76858
rect 19994 76806 20046 76858
rect 20098 76806 50558 76858
rect 50610 76806 50662 76858
rect 50714 76806 50766 76858
rect 50818 76806 78624 76858
rect 1344 76772 78624 76806
rect 4622 76690 4674 76702
rect 4622 76626 4674 76638
rect 15374 76690 15426 76702
rect 15374 76626 15426 76638
rect 19182 76690 19234 76702
rect 19182 76626 19234 76638
rect 21086 76690 21138 76702
rect 21086 76626 21138 76638
rect 24894 76690 24946 76702
rect 24894 76626 24946 76638
rect 25566 76690 25618 76702
rect 25566 76626 25618 76638
rect 26238 76690 26290 76702
rect 26238 76626 26290 76638
rect 26910 76690 26962 76702
rect 26910 76626 26962 76638
rect 27582 76690 27634 76702
rect 27582 76626 27634 76638
rect 28366 76690 28418 76702
rect 28366 76626 28418 76638
rect 28926 76690 28978 76702
rect 28926 76626 28978 76638
rect 29598 76690 29650 76702
rect 29598 76626 29650 76638
rect 30270 76690 30322 76702
rect 30270 76626 30322 76638
rect 30942 76690 30994 76702
rect 30942 76626 30994 76638
rect 31502 76690 31554 76702
rect 31502 76626 31554 76638
rect 32286 76690 32338 76702
rect 32286 76626 32338 76638
rect 36766 76690 36818 76702
rect 36766 76626 36818 76638
rect 37662 76690 37714 76702
rect 37662 76626 37714 76638
rect 39230 76690 39282 76702
rect 39230 76626 39282 76638
rect 40126 76690 40178 76702
rect 40126 76626 40178 76638
rect 41022 76690 41074 76702
rect 41022 76626 41074 76638
rect 42030 76690 42082 76702
rect 42030 76626 42082 76638
rect 42366 76690 42418 76702
rect 42366 76626 42418 76638
rect 43598 76690 43650 76702
rect 43598 76626 43650 76638
rect 44494 76690 44546 76702
rect 44494 76626 44546 76638
rect 45390 76690 45442 76702
rect 45390 76626 45442 76638
rect 46286 76690 46338 76702
rect 46286 76626 46338 76638
rect 47406 76690 47458 76702
rect 47406 76626 47458 76638
rect 48302 76690 48354 76702
rect 48302 76626 48354 76638
rect 49198 76690 49250 76702
rect 49198 76626 49250 76638
rect 50094 76690 50146 76702
rect 50094 76626 50146 76638
rect 51214 76690 51266 76702
rect 51214 76626 51266 76638
rect 52110 76690 52162 76702
rect 52110 76626 52162 76638
rect 53006 76690 53058 76702
rect 53006 76626 53058 76638
rect 53902 76690 53954 76702
rect 53902 76626 53954 76638
rect 55134 76690 55186 76702
rect 55134 76626 55186 76638
rect 59838 76690 59890 76702
rect 59838 76626 59890 76638
rect 63310 76690 63362 76702
rect 63310 76626 63362 76638
rect 63982 76690 64034 76702
rect 63982 76626 64034 76638
rect 64654 76690 64706 76702
rect 64654 76626 64706 76638
rect 65326 76690 65378 76702
rect 65326 76626 65378 76638
rect 66446 76690 66498 76702
rect 66446 76626 66498 76638
rect 67118 76690 67170 76702
rect 67118 76626 67170 76638
rect 67790 76690 67842 76702
rect 67790 76626 67842 76638
rect 68462 76690 68514 76702
rect 68462 76626 68514 76638
rect 69134 76690 69186 76702
rect 69134 76626 69186 76638
rect 72606 76690 72658 76702
rect 72606 76626 72658 76638
rect 74062 76690 74114 76702
rect 74062 76626 74114 76638
rect 75406 76690 75458 76702
rect 75406 76626 75458 76638
rect 76414 76690 76466 76702
rect 76414 76626 76466 76638
rect 4958 76578 5010 76590
rect 4958 76514 5010 76526
rect 5518 76578 5570 76590
rect 62638 76578 62690 76590
rect 36082 76526 36094 76578
rect 36146 76526 36158 76578
rect 61730 76526 61742 76578
rect 61794 76526 61806 76578
rect 5518 76514 5570 76526
rect 62638 76514 62690 76526
rect 62974 76578 63026 76590
rect 70254 76578 70306 76590
rect 63634 76526 63646 76578
rect 63698 76526 63710 76578
rect 64306 76526 64318 76578
rect 64370 76526 64382 76578
rect 64978 76526 64990 76578
rect 65042 76526 65054 76578
rect 65650 76526 65662 76578
rect 65714 76526 65726 76578
rect 66770 76526 66782 76578
rect 66834 76526 66846 76578
rect 67442 76526 67454 76578
rect 67506 76526 67518 76578
rect 68114 76526 68126 76578
rect 68178 76526 68190 76578
rect 68786 76526 68798 76578
rect 68850 76526 68862 76578
rect 69458 76526 69470 76578
rect 69522 76526 69534 76578
rect 62974 76514 63026 76526
rect 70254 76514 70306 76526
rect 70590 76578 70642 76590
rect 70590 76514 70642 76526
rect 70926 76578 70978 76590
rect 70926 76514 70978 76526
rect 71262 76578 71314 76590
rect 71262 76514 71314 76526
rect 71598 76578 71650 76590
rect 72942 76578 72994 76590
rect 74734 76578 74786 76590
rect 72258 76526 72270 76578
rect 72322 76526 72334 76578
rect 74386 76526 74398 76578
rect 74450 76526 74462 76578
rect 71598 76514 71650 76526
rect 72942 76514 72994 76526
rect 74734 76514 74786 76526
rect 75742 76578 75794 76590
rect 78206 76578 78258 76590
rect 76066 76526 76078 76578
rect 76130 76526 76142 76578
rect 75742 76514 75794 76526
rect 78206 76514 78258 76526
rect 62078 76466 62130 76478
rect 77870 76466 77922 76478
rect 4274 76414 4286 76466
rect 4338 76414 4350 76466
rect 5730 76414 5742 76466
rect 5794 76414 5806 76466
rect 12114 76414 12126 76466
rect 12178 76414 12190 76466
rect 16370 76414 16382 76466
rect 16434 76414 16446 76466
rect 19730 76414 19742 76466
rect 19794 76414 19806 76466
rect 23874 76414 23886 76466
rect 23938 76414 23950 76466
rect 35074 76414 35086 76466
rect 35138 76414 35150 76466
rect 36306 76414 36318 76466
rect 36370 76414 36382 76466
rect 58258 76414 58270 76466
rect 58322 76414 58334 76466
rect 58818 76414 58830 76466
rect 58882 76414 58894 76466
rect 71810 76414 71822 76466
rect 71874 76414 71886 76466
rect 73154 76414 73166 76466
rect 73218 76414 73230 76466
rect 74946 76414 74958 76466
rect 75010 76414 75022 76466
rect 77186 76414 77198 76466
rect 77250 76414 77262 76466
rect 62078 76402 62130 76414
rect 77870 76402 77922 76414
rect 13358 76354 13410 76366
rect 13358 76290 13410 76302
rect 17166 76354 17218 76366
rect 17166 76290 17218 76302
rect 21646 76354 21698 76366
rect 37326 76354 37378 76366
rect 38670 76354 38722 76366
rect 33394 76302 33406 76354
rect 33458 76302 33470 76354
rect 38098 76302 38110 76354
rect 38162 76302 38174 76354
rect 21646 76290 21698 76302
rect 37326 76290 37378 76302
rect 38670 76290 38722 76302
rect 40686 76354 40738 76366
rect 40686 76290 40738 76302
rect 41582 76354 41634 76366
rect 44158 76354 44210 76366
rect 42802 76302 42814 76354
rect 42866 76302 42878 76354
rect 41582 76290 41634 76302
rect 44158 76290 44210 76302
rect 45054 76354 45106 76366
rect 45054 76290 45106 76302
rect 45950 76354 46002 76366
rect 45950 76290 46002 76302
rect 46846 76354 46898 76366
rect 48862 76354 48914 76366
rect 47842 76302 47854 76354
rect 47906 76302 47918 76354
rect 46846 76290 46898 76302
rect 48862 76290 48914 76302
rect 49758 76354 49810 76366
rect 52670 76354 52722 76366
rect 55918 76354 55970 76366
rect 50530 76302 50542 76354
rect 50594 76302 50606 76354
rect 51650 76302 51662 76354
rect 51714 76302 51726 76354
rect 53442 76302 53454 76354
rect 53506 76302 53518 76354
rect 54338 76302 54350 76354
rect 54402 76302 54414 76354
rect 49758 76290 49810 76302
rect 52670 76290 52722 76302
rect 55918 76290 55970 76302
rect 76750 76354 76802 76366
rect 76750 76290 76802 76302
rect 1934 76242 1986 76254
rect 1934 76178 1986 76190
rect 11566 76242 11618 76254
rect 11566 76178 11618 76190
rect 1344 76074 78624 76108
rect 1344 76022 4478 76074
rect 4530 76022 4582 76074
rect 4634 76022 4686 76074
rect 4738 76022 35198 76074
rect 35250 76022 35302 76074
rect 35354 76022 35406 76074
rect 35458 76022 65918 76074
rect 65970 76022 66022 76074
rect 66074 76022 66126 76074
rect 66178 76022 78624 76074
rect 1344 75988 78624 76022
rect 11902 75906 11954 75918
rect 11902 75842 11954 75854
rect 16830 75906 16882 75918
rect 16830 75842 16882 75854
rect 21534 75906 21586 75918
rect 21534 75842 21586 75854
rect 56702 75906 56754 75918
rect 62626 75854 62638 75906
rect 62690 75903 62702 75906
rect 63074 75903 63086 75906
rect 62690 75857 63086 75903
rect 62690 75854 62702 75857
rect 63074 75854 63086 75857
rect 63138 75854 63150 75906
rect 71362 75854 71374 75906
rect 71426 75903 71438 75906
rect 71810 75903 71822 75906
rect 71426 75857 71822 75903
rect 71426 75854 71438 75857
rect 71810 75854 71822 75857
rect 71874 75854 71886 75906
rect 56702 75842 56754 75854
rect 1934 75794 1986 75806
rect 24782 75794 24834 75806
rect 18610 75742 18622 75794
rect 18674 75742 18686 75794
rect 1934 75730 1986 75742
rect 24782 75730 24834 75742
rect 32734 75794 32786 75806
rect 32734 75730 32786 75742
rect 34078 75794 34130 75806
rect 34078 75730 34130 75742
rect 35422 75794 35474 75806
rect 35422 75730 35474 75742
rect 36430 75794 36482 75806
rect 36430 75730 36482 75742
rect 37326 75794 37378 75806
rect 37326 75730 37378 75742
rect 37886 75794 37938 75806
rect 40014 75794 40066 75806
rect 38546 75742 38558 75794
rect 38610 75742 38622 75794
rect 37886 75730 37938 75742
rect 40014 75730 40066 75742
rect 41470 75794 41522 75806
rect 41470 75730 41522 75742
rect 42478 75794 42530 75806
rect 42478 75730 42530 75742
rect 43374 75794 43426 75806
rect 43374 75730 43426 75742
rect 43934 75794 43986 75806
rect 43934 75730 43986 75742
rect 44382 75794 44434 75806
rect 44382 75730 44434 75742
rect 46062 75794 46114 75806
rect 46062 75730 46114 75742
rect 46510 75794 46562 75806
rect 46510 75730 46562 75742
rect 48078 75794 48130 75806
rect 48078 75730 48130 75742
rect 48526 75794 48578 75806
rect 48526 75730 48578 75742
rect 49086 75794 49138 75806
rect 49086 75730 49138 75742
rect 49534 75794 49586 75806
rect 50766 75794 50818 75806
rect 50194 75742 50206 75794
rect 50258 75742 50270 75794
rect 49534 75730 49586 75742
rect 50766 75730 50818 75742
rect 51214 75794 51266 75806
rect 51214 75730 51266 75742
rect 51774 75794 51826 75806
rect 51774 75730 51826 75742
rect 52222 75794 52274 75806
rect 63086 75794 63138 75806
rect 54226 75742 54238 75794
rect 54290 75742 54302 75794
rect 55122 75742 55134 75794
rect 55186 75742 55198 75794
rect 56018 75742 56030 75794
rect 56082 75742 56094 75794
rect 52222 75730 52274 75742
rect 63086 75730 63138 75742
rect 63534 75794 63586 75806
rect 63534 75730 63586 75742
rect 63982 75794 64034 75806
rect 63982 75730 64034 75742
rect 64542 75794 64594 75806
rect 64542 75730 64594 75742
rect 64990 75794 65042 75806
rect 64990 75730 65042 75742
rect 65998 75794 66050 75806
rect 65998 75730 66050 75742
rect 66446 75794 66498 75806
rect 66446 75730 66498 75742
rect 67006 75794 67058 75806
rect 67006 75730 67058 75742
rect 67566 75794 67618 75806
rect 67566 75730 67618 75742
rect 68462 75794 68514 75806
rect 68462 75730 68514 75742
rect 69022 75794 69074 75806
rect 69022 75730 69074 75742
rect 70030 75794 70082 75806
rect 70030 75730 70082 75742
rect 70702 75794 70754 75806
rect 70702 75730 70754 75742
rect 71374 75794 71426 75806
rect 71374 75730 71426 75742
rect 71934 75794 71986 75806
rect 71934 75730 71986 75742
rect 72382 75794 72434 75806
rect 72382 75730 72434 75742
rect 73390 75794 73442 75806
rect 73390 75730 73442 75742
rect 73950 75794 74002 75806
rect 73950 75730 74002 75742
rect 74510 75794 74562 75806
rect 74510 75730 74562 75742
rect 75070 75794 75122 75806
rect 75070 75730 75122 75742
rect 4958 75682 5010 75694
rect 13582 75682 13634 75694
rect 25230 75682 25282 75694
rect 4274 75630 4286 75682
rect 4338 75630 4350 75682
rect 12674 75630 12686 75682
rect 12738 75630 12750 75682
rect 17826 75630 17838 75682
rect 17890 75630 17902 75682
rect 20290 75630 20302 75682
rect 20354 75630 20366 75682
rect 23650 75630 23662 75682
rect 23714 75630 23726 75682
rect 4958 75618 5010 75630
rect 13582 75618 13634 75630
rect 25230 75618 25282 75630
rect 32958 75682 33010 75694
rect 32958 75618 33010 75630
rect 33518 75682 33570 75694
rect 33518 75618 33570 75630
rect 34302 75682 34354 75694
rect 34302 75618 34354 75630
rect 34862 75682 34914 75694
rect 34862 75618 34914 75630
rect 35646 75682 35698 75694
rect 39006 75682 39058 75694
rect 38210 75630 38222 75682
rect 38274 75630 38286 75682
rect 35646 75618 35698 75630
rect 39006 75618 39058 75630
rect 39566 75682 39618 75694
rect 39566 75618 39618 75630
rect 40910 75682 40962 75694
rect 40910 75618 40962 75630
rect 41694 75682 41746 75694
rect 45614 75682 45666 75694
rect 45154 75630 45166 75682
rect 45218 75630 45230 75682
rect 41694 75618 41746 75630
rect 45614 75618 45666 75630
rect 47070 75682 47122 75694
rect 47070 75618 47122 75630
rect 47630 75682 47682 75694
rect 47630 75618 47682 75630
rect 49758 75682 49810 75694
rect 49758 75618 49810 75630
rect 52670 75682 52722 75694
rect 52670 75618 52722 75630
rect 53230 75682 53282 75694
rect 53230 75618 53282 75630
rect 53790 75682 53842 75694
rect 53790 75618 53842 75630
rect 54686 75682 54738 75694
rect 54686 75618 54738 75630
rect 55582 75682 55634 75694
rect 61854 75682 61906 75694
rect 59042 75630 59054 75682
rect 59106 75630 59118 75682
rect 55582 75618 55634 75630
rect 61854 75618 61906 75630
rect 62638 75682 62690 75694
rect 62638 75618 62690 75630
rect 65214 75682 65266 75694
rect 65214 75618 65266 75630
rect 72606 75682 72658 75694
rect 76190 75682 76242 75694
rect 75394 75630 75406 75682
rect 75458 75630 75470 75682
rect 72606 75618 72658 75630
rect 76190 75618 76242 75630
rect 76862 75682 76914 75694
rect 78082 75630 78094 75682
rect 78146 75630 78158 75682
rect 76862 75618 76914 75630
rect 4622 75570 4674 75582
rect 4622 75506 4674 75518
rect 24222 75570 24274 75582
rect 24222 75506 24274 75518
rect 59390 75570 59442 75582
rect 59390 75506 59442 75518
rect 61182 75570 61234 75582
rect 61182 75506 61234 75518
rect 75630 75570 75682 75582
rect 76514 75518 76526 75570
rect 76578 75518 76590 75570
rect 77858 75518 77870 75570
rect 77922 75518 77934 75570
rect 75630 75506 75682 75518
rect 14254 75458 14306 75470
rect 14254 75394 14306 75406
rect 14702 75458 14754 75470
rect 60510 75458 60562 75470
rect 62190 75458 62242 75470
rect 77198 75458 77250 75470
rect 35970 75406 35982 75458
rect 36034 75406 36046 75458
rect 42018 75406 42030 75458
rect 42082 75406 42094 75458
rect 59714 75406 59726 75458
rect 59778 75406 59790 75458
rect 60834 75406 60846 75458
rect 60898 75406 60910 75458
rect 61506 75406 61518 75458
rect 61570 75406 61582 75458
rect 65538 75406 65550 75458
rect 65602 75406 65614 75458
rect 72930 75406 72942 75458
rect 72994 75406 73006 75458
rect 14702 75394 14754 75406
rect 60510 75394 60562 75406
rect 62190 75394 62242 75406
rect 77198 75394 77250 75406
rect 1344 75290 78624 75324
rect 1344 75238 19838 75290
rect 19890 75238 19942 75290
rect 19994 75238 20046 75290
rect 20098 75238 50558 75290
rect 50610 75238 50662 75290
rect 50714 75238 50766 75290
rect 50818 75238 78624 75290
rect 1344 75204 78624 75238
rect 4622 75122 4674 75134
rect 4622 75058 4674 75070
rect 12910 75122 12962 75134
rect 12910 75058 12962 75070
rect 15262 75122 15314 75134
rect 15262 75058 15314 75070
rect 23102 75122 23154 75134
rect 23102 75058 23154 75070
rect 23550 75122 23602 75134
rect 23550 75058 23602 75070
rect 34750 75122 34802 75134
rect 34750 75058 34802 75070
rect 37438 75122 37490 75134
rect 37438 75058 37490 75070
rect 38894 75122 38946 75134
rect 38894 75058 38946 75070
rect 46846 75122 46898 75134
rect 46846 75058 46898 75070
rect 52782 75122 52834 75134
rect 52782 75058 52834 75070
rect 53566 75122 53618 75134
rect 53566 75058 53618 75070
rect 54462 75122 54514 75134
rect 54462 75058 54514 75070
rect 55358 75122 55410 75134
rect 55358 75058 55410 75070
rect 57486 75122 57538 75134
rect 57486 75058 57538 75070
rect 61294 75122 61346 75134
rect 61294 75058 61346 75070
rect 61742 75122 61794 75134
rect 61742 75058 61794 75070
rect 62190 75122 62242 75134
rect 62190 75058 62242 75070
rect 74062 75122 74114 75134
rect 74062 75058 74114 75070
rect 74510 75122 74562 75134
rect 74510 75058 74562 75070
rect 74958 75122 75010 75134
rect 74958 75058 75010 75070
rect 75406 75122 75458 75134
rect 75406 75058 75458 75070
rect 76862 75122 76914 75134
rect 76862 75058 76914 75070
rect 75630 75010 75682 75022
rect 34962 74958 34974 75010
rect 35026 74958 35038 75010
rect 75630 74946 75682 74958
rect 75966 75010 76018 75022
rect 75966 74946 76018 74958
rect 77534 75010 77586 75022
rect 77534 74946 77586 74958
rect 77870 75010 77922 75022
rect 77870 74946 77922 74958
rect 60846 74898 60898 74910
rect 4162 74846 4174 74898
rect 4226 74846 4238 74898
rect 4834 74846 4846 74898
rect 4898 74846 4910 74898
rect 13458 74846 13470 74898
rect 13522 74846 13534 74898
rect 14690 74846 14702 74898
rect 14754 74846 14766 74898
rect 22754 74846 22766 74898
rect 22818 74846 22830 74898
rect 35186 74846 35198 74898
rect 35250 74846 35262 74898
rect 60386 74846 60398 74898
rect 60450 74846 60462 74898
rect 77298 74846 77310 74898
rect 77362 74846 77374 74898
rect 78082 74846 78094 74898
rect 78146 74846 78158 74898
rect 60846 74834 60898 74846
rect 17950 74786 18002 74798
rect 2146 74734 2158 74786
rect 2210 74734 2222 74786
rect 17950 74722 18002 74734
rect 18286 74786 18338 74798
rect 18286 74722 18338 74734
rect 19406 74786 19458 74798
rect 19406 74722 19458 74734
rect 19854 74786 19906 74798
rect 19854 74722 19906 74734
rect 20414 74786 20466 74798
rect 20414 74722 20466 74734
rect 35758 74786 35810 74798
rect 35758 74722 35810 74734
rect 58046 74786 58098 74798
rect 58046 74722 58098 74734
rect 76302 74786 76354 74798
rect 76302 74722 76354 74734
rect 1344 74506 78624 74540
rect 1344 74454 4478 74506
rect 4530 74454 4582 74506
rect 4634 74454 4686 74506
rect 4738 74454 35198 74506
rect 35250 74454 35302 74506
rect 35354 74454 35406 74506
rect 35458 74454 65918 74506
rect 65970 74454 66022 74506
rect 66074 74454 66126 74506
rect 66178 74454 78624 74506
rect 1344 74420 78624 74454
rect 19182 74338 19234 74350
rect 77746 74286 77758 74338
rect 77810 74335 77822 74338
rect 77970 74335 77982 74338
rect 77810 74289 77982 74335
rect 77810 74286 77822 74289
rect 77970 74286 77982 74289
rect 78034 74286 78046 74338
rect 19182 74274 19234 74286
rect 1934 74226 1986 74238
rect 58494 74226 58546 74238
rect 11218 74174 11230 74226
rect 11282 74174 11294 74226
rect 16034 74174 16046 74226
rect 16098 74174 16110 74226
rect 1934 74162 1986 74174
rect 58494 74162 58546 74174
rect 59166 74226 59218 74238
rect 59166 74162 59218 74174
rect 75294 74226 75346 74238
rect 75294 74162 75346 74174
rect 75742 74226 75794 74238
rect 75742 74162 75794 74174
rect 76414 74226 76466 74238
rect 76414 74162 76466 74174
rect 77982 74226 78034 74238
rect 77982 74162 78034 74174
rect 14030 74114 14082 74126
rect 76974 74114 77026 74126
rect 4274 74062 4286 74114
rect 4338 74062 4350 74114
rect 4834 74062 4846 74114
rect 4898 74062 4910 74114
rect 12898 74062 12910 74114
rect 12962 74062 12974 74114
rect 17826 74062 17838 74114
rect 17890 74062 17902 74114
rect 18162 74062 18174 74114
rect 18226 74062 18238 74114
rect 14030 74050 14082 74062
rect 76974 74050 77026 74062
rect 77534 74114 77586 74126
rect 77534 74050 77586 74062
rect 4622 74002 4674 74014
rect 4622 73938 4674 73950
rect 14366 74002 14418 74014
rect 14366 73938 14418 73950
rect 22990 74002 23042 74014
rect 22990 73938 23042 73950
rect 59502 73890 59554 73902
rect 59502 73826 59554 73838
rect 1344 73722 78624 73756
rect 1344 73670 19838 73722
rect 19890 73670 19942 73722
rect 19994 73670 20046 73722
rect 20098 73670 50558 73722
rect 50610 73670 50662 73722
rect 50714 73670 50766 73722
rect 50818 73670 78624 73722
rect 1344 73636 78624 73670
rect 76078 73554 76130 73566
rect 76078 73490 76130 73502
rect 76526 73554 76578 73566
rect 76526 73490 76578 73502
rect 76974 73554 77026 73566
rect 76974 73490 77026 73502
rect 77422 73554 77474 73566
rect 77422 73490 77474 73502
rect 78206 73554 78258 73566
rect 78206 73490 78258 73502
rect 4622 73442 4674 73454
rect 12114 73390 12126 73442
rect 12178 73390 12190 73442
rect 4622 73378 4674 73390
rect 4274 73278 4286 73330
rect 4338 73278 4350 73330
rect 4834 73278 4846 73330
rect 4898 73278 4910 73330
rect 13906 73278 13918 73330
rect 13970 73278 13982 73330
rect 16370 73278 16382 73330
rect 16434 73278 16446 73330
rect 18062 73218 18114 73230
rect 14578 73166 14590 73218
rect 14642 73166 14654 73218
rect 18062 73154 18114 73166
rect 77646 73218 77698 73230
rect 77646 73154 77698 73166
rect 1934 73106 1986 73118
rect 76626 73054 76638 73106
rect 76690 73103 76702 73106
rect 77186 73103 77198 73106
rect 76690 73057 77198 73103
rect 76690 73054 76702 73057
rect 77186 73054 77198 73057
rect 77250 73054 77262 73106
rect 1934 73042 1986 73054
rect 1344 72938 78624 72972
rect 1344 72886 4478 72938
rect 4530 72886 4582 72938
rect 4634 72886 4686 72938
rect 4738 72886 35198 72938
rect 35250 72886 35302 72938
rect 35354 72886 35406 72938
rect 35458 72886 65918 72938
rect 65970 72886 66022 72938
rect 66074 72886 66126 72938
rect 66178 72886 78624 72938
rect 1344 72852 78624 72886
rect 1934 72658 1986 72670
rect 1934 72594 1986 72606
rect 77198 72658 77250 72670
rect 77198 72594 77250 72606
rect 4958 72546 5010 72558
rect 3826 72494 3838 72546
rect 3890 72494 3902 72546
rect 4958 72482 5010 72494
rect 77646 72434 77698 72446
rect 77646 72370 77698 72382
rect 78206 72434 78258 72446
rect 78206 72370 78258 72382
rect 4622 72322 4674 72334
rect 4622 72258 4674 72270
rect 14142 72322 14194 72334
rect 14142 72258 14194 72270
rect 77870 72322 77922 72334
rect 77870 72258 77922 72270
rect 1344 72154 78624 72188
rect 1344 72102 19838 72154
rect 19890 72102 19942 72154
rect 19994 72102 20046 72154
rect 20098 72102 50558 72154
rect 50610 72102 50662 72154
rect 50714 72102 50766 72154
rect 50818 72102 78624 72154
rect 1344 72068 78624 72102
rect 2494 71986 2546 71998
rect 2494 71922 2546 71934
rect 3166 71986 3218 71998
rect 3166 71922 3218 71934
rect 3502 71986 3554 71998
rect 3502 71922 3554 71934
rect 3838 71874 3890 71886
rect 77858 71822 77870 71874
rect 77922 71822 77934 71874
rect 3838 71810 3890 71822
rect 2158 71762 2210 71774
rect 77646 71762 77698 71774
rect 2930 71710 2942 71762
rect 2994 71710 3006 71762
rect 2158 71698 2210 71710
rect 77646 71698 77698 71710
rect 78206 71762 78258 71774
rect 78206 71698 78258 71710
rect 1934 71650 1986 71662
rect 1934 71586 1986 71598
rect 1344 71370 78624 71404
rect 1344 71318 4478 71370
rect 4530 71318 4582 71370
rect 4634 71318 4686 71370
rect 4738 71318 35198 71370
rect 35250 71318 35302 71370
rect 35354 71318 35406 71370
rect 35458 71318 65918 71370
rect 65970 71318 66022 71370
rect 66074 71318 66126 71370
rect 66178 71318 78624 71370
rect 1344 71284 78624 71318
rect 1934 71090 1986 71102
rect 77746 71038 77758 71090
rect 77810 71038 77822 71090
rect 1934 71026 1986 71038
rect 3938 70926 3950 70978
rect 4002 70926 4014 70978
rect 77422 70754 77474 70766
rect 77422 70690 77474 70702
rect 78206 70754 78258 70766
rect 78206 70690 78258 70702
rect 1344 70586 78624 70620
rect 1344 70534 19838 70586
rect 19890 70534 19942 70586
rect 19994 70534 20046 70586
rect 20098 70534 50558 70586
rect 50610 70534 50662 70586
rect 50714 70534 50766 70586
rect 50818 70534 78624 70586
rect 1344 70500 78624 70534
rect 3826 70142 3838 70194
rect 3890 70142 3902 70194
rect 1934 69970 1986 69982
rect 1934 69906 1986 69918
rect 1344 69802 78624 69836
rect 1344 69750 4478 69802
rect 4530 69750 4582 69802
rect 4634 69750 4686 69802
rect 4738 69750 35198 69802
rect 35250 69750 35302 69802
rect 35354 69750 35406 69802
rect 35458 69750 65918 69802
rect 65970 69750 66022 69802
rect 66074 69750 66126 69802
rect 66178 69750 78624 69802
rect 1344 69716 78624 69750
rect 2930 69358 2942 69410
rect 2994 69358 3006 69410
rect 2382 69298 2434 69310
rect 2382 69234 2434 69246
rect 2718 69298 2770 69310
rect 2718 69234 2770 69246
rect 2046 69186 2098 69198
rect 2046 69122 2098 69134
rect 77646 69186 77698 69198
rect 78206 69186 78258 69198
rect 77858 69134 77870 69186
rect 77922 69134 77934 69186
rect 77646 69122 77698 69134
rect 78206 69122 78258 69134
rect 1344 69018 78624 69052
rect 1344 68966 19838 69018
rect 19890 68966 19942 69018
rect 19994 68966 20046 69018
rect 20098 68966 50558 69018
rect 50610 68966 50662 69018
rect 50714 68966 50766 69018
rect 50818 68966 78624 69018
rect 1344 68932 78624 68966
rect 78206 68626 78258 68638
rect 2034 68574 2046 68626
rect 2098 68574 2110 68626
rect 78206 68562 78258 68574
rect 77422 68514 77474 68526
rect 77422 68450 77474 68462
rect 77646 68514 77698 68526
rect 77646 68450 77698 68462
rect 2718 68402 2770 68414
rect 2718 68338 2770 68350
rect 1344 68234 78624 68268
rect 1344 68182 4478 68234
rect 4530 68182 4582 68234
rect 4634 68182 4686 68234
rect 4738 68182 35198 68234
rect 35250 68182 35302 68234
rect 35354 68182 35406 68234
rect 35458 68182 65918 68234
rect 65970 68182 66022 68234
rect 66074 68182 66126 68234
rect 66178 68182 78624 68234
rect 1344 68148 78624 68182
rect 1934 67954 1986 67966
rect 1934 67890 1986 67902
rect 4050 67790 4062 67842
rect 4114 67790 4126 67842
rect 1344 67450 78624 67484
rect 1344 67398 19838 67450
rect 19890 67398 19942 67450
rect 19994 67398 20046 67450
rect 20098 67398 50558 67450
rect 50610 67398 50662 67450
rect 50714 67398 50766 67450
rect 50818 67398 78624 67450
rect 1344 67364 78624 67398
rect 4062 67282 4114 67294
rect 4062 67218 4114 67230
rect 2046 67170 2098 67182
rect 2046 67106 2098 67118
rect 2718 67170 2770 67182
rect 2718 67106 2770 67118
rect 3054 67170 3106 67182
rect 3054 67106 3106 67118
rect 3726 67170 3778 67182
rect 77858 67118 77870 67170
rect 77922 67118 77934 67170
rect 3726 67106 3778 67118
rect 2382 67058 2434 67070
rect 2382 66994 2434 67006
rect 3390 67058 3442 67070
rect 78206 67058 78258 67070
rect 4274 67006 4286 67058
rect 4338 67006 4350 67058
rect 3390 66994 3442 67006
rect 78206 66994 78258 67006
rect 77646 66946 77698 66958
rect 77646 66882 77698 66894
rect 1344 66666 78624 66700
rect 1344 66614 4478 66666
rect 4530 66614 4582 66666
rect 4634 66614 4686 66666
rect 4738 66614 35198 66666
rect 35250 66614 35302 66666
rect 35354 66614 35406 66666
rect 35458 66614 65918 66666
rect 65970 66614 66022 66666
rect 66074 66614 66126 66666
rect 66178 66614 78624 66666
rect 1344 66580 78624 66614
rect 1934 66386 1986 66398
rect 1934 66322 1986 66334
rect 77646 66274 77698 66286
rect 3826 66222 3838 66274
rect 3890 66222 3902 66274
rect 77646 66210 77698 66222
rect 77422 66050 77474 66062
rect 77422 65986 77474 65998
rect 78206 66050 78258 66062
rect 78206 65986 78258 65998
rect 1344 65882 78624 65916
rect 1344 65830 19838 65882
rect 19890 65830 19942 65882
rect 19994 65830 20046 65882
rect 20098 65830 50558 65882
rect 50610 65830 50662 65882
rect 50714 65830 50766 65882
rect 50818 65830 78624 65882
rect 1344 65796 78624 65830
rect 2034 65438 2046 65490
rect 2098 65438 2110 65490
rect 2718 65266 2770 65278
rect 2718 65202 2770 65214
rect 1344 65098 78624 65132
rect 1344 65046 4478 65098
rect 4530 65046 4582 65098
rect 4634 65046 4686 65098
rect 4738 65046 35198 65098
rect 35250 65046 35302 65098
rect 35354 65046 35406 65098
rect 35458 65046 65918 65098
rect 65970 65046 66022 65098
rect 66074 65046 66126 65098
rect 66178 65046 78624 65098
rect 1344 65012 78624 65046
rect 1934 64818 1986 64830
rect 1934 64754 1986 64766
rect 77646 64706 77698 64718
rect 3826 64654 3838 64706
rect 3890 64654 3902 64706
rect 77646 64642 77698 64654
rect 77422 64594 77474 64606
rect 77422 64530 77474 64542
rect 78206 64594 78258 64606
rect 78206 64530 78258 64542
rect 1344 64314 78624 64348
rect 1344 64262 19838 64314
rect 19890 64262 19942 64314
rect 19994 64262 20046 64314
rect 20098 64262 50558 64314
rect 50610 64262 50662 64314
rect 50714 64262 50766 64314
rect 50818 64262 78624 64314
rect 1344 64228 78624 64262
rect 2494 64146 2546 64158
rect 2494 64082 2546 64094
rect 3502 64146 3554 64158
rect 3502 64082 3554 64094
rect 2830 64034 2882 64046
rect 2830 63970 2882 63982
rect 3166 64034 3218 64046
rect 77858 63982 77870 64034
rect 77922 63982 77934 64034
rect 3166 63970 3218 63982
rect 77646 63922 77698 63934
rect 2258 63870 2270 63922
rect 2322 63870 2334 63922
rect 3714 63870 3726 63922
rect 3778 63870 3790 63922
rect 77646 63858 77698 63870
rect 78206 63922 78258 63934
rect 78206 63858 78258 63870
rect 1344 63530 78624 63564
rect 1344 63478 4478 63530
rect 4530 63478 4582 63530
rect 4634 63478 4686 63530
rect 4738 63478 35198 63530
rect 35250 63478 35302 63530
rect 35354 63478 35406 63530
rect 35458 63478 65918 63530
rect 65970 63478 66022 63530
rect 66074 63478 66126 63530
rect 66178 63478 78624 63530
rect 1344 63444 78624 63478
rect 1934 63250 1986 63262
rect 1934 63186 1986 63198
rect 77646 63138 77698 63150
rect 3826 63086 3838 63138
rect 3890 63086 3902 63138
rect 77646 63074 77698 63086
rect 77422 62914 77474 62926
rect 77422 62850 77474 62862
rect 78206 62914 78258 62926
rect 78206 62850 78258 62862
rect 1344 62746 78624 62780
rect 1344 62694 19838 62746
rect 19890 62694 19942 62746
rect 19994 62694 20046 62746
rect 20098 62694 50558 62746
rect 50610 62694 50662 62746
rect 50714 62694 50766 62746
rect 50818 62694 78624 62746
rect 1344 62660 78624 62694
rect 3826 62302 3838 62354
rect 3890 62302 3902 62354
rect 1934 62130 1986 62142
rect 1934 62066 1986 62078
rect 1344 61962 78624 61996
rect 1344 61910 4478 61962
rect 4530 61910 4582 61962
rect 4634 61910 4686 61962
rect 4738 61910 35198 61962
rect 35250 61910 35302 61962
rect 35354 61910 35406 61962
rect 35458 61910 65918 61962
rect 65970 61910 66022 61962
rect 66074 61910 66126 61962
rect 66178 61910 78624 61962
rect 1344 61876 78624 61910
rect 2258 61518 2270 61570
rect 2322 61518 2334 61570
rect 3602 61518 3614 61570
rect 3666 61518 3678 61570
rect 2718 61458 2770 61470
rect 2718 61394 2770 61406
rect 3054 61458 3106 61470
rect 3054 61394 3106 61406
rect 3390 61458 3442 61470
rect 3390 61394 3442 61406
rect 2046 61346 2098 61358
rect 2046 61282 2098 61294
rect 4286 61346 4338 61358
rect 4286 61282 4338 61294
rect 77646 61346 77698 61358
rect 78206 61346 78258 61358
rect 77858 61294 77870 61346
rect 77922 61294 77934 61346
rect 77646 61282 77698 61294
rect 78206 61282 78258 61294
rect 1344 61178 78624 61212
rect 1344 61126 19838 61178
rect 19890 61126 19942 61178
rect 19994 61126 20046 61178
rect 20098 61126 50558 61178
rect 50610 61126 50662 61178
rect 50714 61126 50766 61178
rect 50818 61126 78624 61178
rect 1344 61092 78624 61126
rect 77870 60898 77922 60910
rect 77870 60834 77922 60846
rect 77646 60786 77698 60798
rect 2034 60734 2046 60786
rect 2098 60734 2110 60786
rect 77646 60722 77698 60734
rect 78206 60786 78258 60798
rect 78206 60722 78258 60734
rect 2718 60562 2770 60574
rect 2718 60498 2770 60510
rect 1344 60394 78624 60428
rect 1344 60342 4478 60394
rect 4530 60342 4582 60394
rect 4634 60342 4686 60394
rect 4738 60342 35198 60394
rect 35250 60342 35302 60394
rect 35354 60342 35406 60394
rect 35458 60342 65918 60394
rect 65970 60342 66022 60394
rect 66074 60342 66126 60394
rect 66178 60342 78624 60394
rect 1344 60308 78624 60342
rect 1934 60114 1986 60126
rect 1934 60050 1986 60062
rect 3826 59950 3838 60002
rect 3890 59950 3902 60002
rect 1344 59610 78624 59644
rect 1344 59558 19838 59610
rect 19890 59558 19942 59610
rect 19994 59558 20046 59610
rect 20098 59558 50558 59610
rect 50610 59558 50662 59610
rect 50714 59558 50766 59610
rect 50818 59558 78624 59610
rect 1344 59524 78624 59558
rect 2718 59442 2770 59454
rect 2718 59378 2770 59390
rect 2046 59330 2098 59342
rect 2046 59266 2098 59278
rect 2382 59218 2434 59230
rect 3502 59218 3554 59230
rect 2930 59166 2942 59218
rect 2994 59166 3006 59218
rect 2382 59154 2434 59166
rect 3502 59154 3554 59166
rect 78206 59218 78258 59230
rect 78206 59154 78258 59166
rect 77422 59106 77474 59118
rect 77422 59042 77474 59054
rect 77646 59106 77698 59118
rect 77646 59042 77698 59054
rect 1344 58826 78624 58860
rect 1344 58774 4478 58826
rect 4530 58774 4582 58826
rect 4634 58774 4686 58826
rect 4738 58774 35198 58826
rect 35250 58774 35302 58826
rect 35354 58774 35406 58826
rect 35458 58774 65918 58826
rect 65970 58774 66022 58826
rect 66074 58774 66126 58826
rect 66178 58774 78624 58826
rect 1344 58740 78624 58774
rect 2034 58382 2046 58434
rect 2098 58382 2110 58434
rect 2718 58210 2770 58222
rect 2718 58146 2770 58158
rect 77646 58210 77698 58222
rect 78206 58210 78258 58222
rect 77858 58158 77870 58210
rect 77922 58158 77934 58210
rect 77646 58146 77698 58158
rect 78206 58146 78258 58158
rect 1344 58042 78624 58076
rect 1344 57990 19838 58042
rect 19890 57990 19942 58042
rect 19994 57990 20046 58042
rect 20098 57990 50558 58042
rect 50610 57990 50662 58042
rect 50714 57990 50766 58042
rect 50818 57990 78624 58042
rect 1344 57956 78624 57990
rect 4274 57598 4286 57650
rect 4338 57598 4350 57650
rect 1934 57426 1986 57438
rect 1934 57362 1986 57374
rect 1344 57258 78624 57292
rect 1344 57206 4478 57258
rect 4530 57206 4582 57258
rect 4634 57206 4686 57258
rect 4738 57206 35198 57258
rect 35250 57206 35302 57258
rect 35354 57206 35406 57258
rect 35458 57206 65918 57258
rect 65970 57206 66022 57258
rect 66074 57206 66126 57258
rect 66178 57206 78624 57258
rect 1344 57172 78624 57206
rect 1934 56978 1986 56990
rect 1934 56914 1986 56926
rect 3826 56814 3838 56866
rect 3890 56814 3902 56866
rect 4834 56814 4846 56866
rect 4898 56814 4910 56866
rect 4622 56754 4674 56766
rect 4622 56690 4674 56702
rect 77646 56754 77698 56766
rect 77646 56690 77698 56702
rect 78206 56754 78258 56766
rect 78206 56690 78258 56702
rect 77858 56590 77870 56642
rect 77922 56590 77934 56642
rect 1344 56474 78624 56508
rect 1344 56422 19838 56474
rect 19890 56422 19942 56474
rect 19994 56422 20046 56474
rect 20098 56422 50558 56474
rect 50610 56422 50662 56474
rect 50714 56422 50766 56474
rect 50818 56422 78624 56474
rect 1344 56388 78624 56422
rect 2718 56306 2770 56318
rect 2718 56242 2770 56254
rect 3726 56306 3778 56318
rect 3726 56242 3778 56254
rect 2046 56194 2098 56206
rect 2046 56130 2098 56142
rect 2382 56194 2434 56206
rect 2382 56130 2434 56142
rect 3390 56194 3442 56206
rect 3390 56130 3442 56142
rect 78206 56082 78258 56094
rect 2930 56030 2942 56082
rect 2994 56030 3006 56082
rect 78206 56018 78258 56030
rect 77422 55970 77474 55982
rect 77422 55906 77474 55918
rect 77646 55970 77698 55982
rect 77646 55906 77698 55918
rect 1344 55690 78624 55724
rect 1344 55638 4478 55690
rect 4530 55638 4582 55690
rect 4634 55638 4686 55690
rect 4738 55638 35198 55690
rect 35250 55638 35302 55690
rect 35354 55638 35406 55690
rect 35458 55638 65918 55690
rect 65970 55638 66022 55690
rect 66074 55638 66126 55690
rect 66178 55638 78624 55690
rect 1344 55604 78624 55638
rect 2034 55246 2046 55298
rect 2098 55246 2110 55298
rect 77646 55186 77698 55198
rect 77646 55122 77698 55134
rect 78206 55186 78258 55198
rect 78206 55122 78258 55134
rect 2718 55074 2770 55086
rect 2718 55010 2770 55022
rect 77870 55074 77922 55086
rect 77870 55010 77922 55022
rect 1344 54906 78624 54940
rect 1344 54854 19838 54906
rect 19890 54854 19942 54906
rect 19994 54854 20046 54906
rect 20098 54854 50558 54906
rect 50610 54854 50662 54906
rect 50714 54854 50766 54906
rect 50818 54854 78624 54906
rect 1344 54820 78624 54854
rect 3826 54462 3838 54514
rect 3890 54462 3902 54514
rect 1934 54290 1986 54302
rect 1934 54226 1986 54238
rect 1344 54122 78624 54156
rect 1344 54070 4478 54122
rect 4530 54070 4582 54122
rect 4634 54070 4686 54122
rect 4738 54070 35198 54122
rect 35250 54070 35302 54122
rect 35354 54070 35406 54122
rect 35458 54070 65918 54122
rect 65970 54070 66022 54122
rect 66074 54070 66126 54122
rect 66178 54070 78624 54122
rect 1344 54036 78624 54070
rect 2258 53678 2270 53730
rect 2322 53678 2334 53730
rect 2930 53678 2942 53730
rect 2994 53678 3006 53730
rect 1934 53618 1986 53630
rect 1934 53554 1986 53566
rect 3166 53618 3218 53630
rect 3166 53554 3218 53566
rect 3502 53618 3554 53630
rect 3502 53554 3554 53566
rect 3838 53618 3890 53630
rect 3838 53554 3890 53566
rect 78206 53618 78258 53630
rect 78206 53554 78258 53566
rect 2494 53506 2546 53518
rect 2494 53442 2546 53454
rect 77646 53506 77698 53518
rect 77646 53442 77698 53454
rect 77870 53506 77922 53518
rect 77870 53442 77922 53454
rect 1344 53338 78624 53372
rect 1344 53286 19838 53338
rect 19890 53286 19942 53338
rect 19994 53286 20046 53338
rect 20098 53286 50558 53338
rect 50610 53286 50662 53338
rect 50714 53286 50766 53338
rect 50818 53286 78624 53338
rect 1344 53252 78624 53286
rect 77870 53058 77922 53070
rect 77870 52994 77922 53006
rect 78206 52946 78258 52958
rect 3938 52894 3950 52946
rect 4002 52894 4014 52946
rect 78206 52882 78258 52894
rect 77646 52834 77698 52846
rect 77646 52770 77698 52782
rect 1934 52722 1986 52734
rect 1934 52658 1986 52670
rect 1344 52554 78624 52588
rect 1344 52502 4478 52554
rect 4530 52502 4582 52554
rect 4634 52502 4686 52554
rect 4738 52502 35198 52554
rect 35250 52502 35302 52554
rect 35354 52502 35406 52554
rect 35458 52502 65918 52554
rect 65970 52502 66022 52554
rect 66074 52502 66126 52554
rect 66178 52502 78624 52554
rect 1344 52468 78624 52502
rect 1934 52274 1986 52286
rect 1934 52210 1986 52222
rect 3826 52110 3838 52162
rect 3890 52110 3902 52162
rect 1344 51770 78624 51804
rect 1344 51718 19838 51770
rect 19890 51718 19942 51770
rect 19994 51718 20046 51770
rect 20098 51718 50558 51770
rect 50610 51718 50662 51770
rect 50714 51718 50766 51770
rect 50818 51718 78624 51770
rect 1344 51684 78624 51718
rect 2494 51602 2546 51614
rect 2494 51538 2546 51550
rect 3502 51602 3554 51614
rect 3502 51538 3554 51550
rect 2830 51490 2882 51502
rect 2830 51426 2882 51438
rect 3838 51490 3890 51502
rect 3838 51426 3890 51438
rect 77870 51490 77922 51502
rect 77870 51426 77922 51438
rect 3166 51378 3218 51390
rect 2258 51326 2270 51378
rect 2322 51326 2334 51378
rect 3166 51314 3218 51326
rect 78206 51378 78258 51390
rect 78206 51314 78258 51326
rect 77646 51266 77698 51278
rect 77646 51202 77698 51214
rect 1344 50986 78624 51020
rect 1344 50934 4478 50986
rect 4530 50934 4582 50986
rect 4634 50934 4686 50986
rect 4738 50934 35198 50986
rect 35250 50934 35302 50986
rect 35354 50934 35406 50986
rect 35458 50934 65918 50986
rect 65970 50934 66022 50986
rect 66074 50934 66126 50986
rect 66178 50934 78624 50986
rect 1344 50900 78624 50934
rect 1934 50706 1986 50718
rect 1934 50642 1986 50654
rect 3826 50542 3838 50594
rect 3890 50542 3902 50594
rect 77646 50482 77698 50494
rect 77646 50418 77698 50430
rect 78206 50482 78258 50494
rect 78206 50418 78258 50430
rect 77870 50370 77922 50382
rect 77870 50306 77922 50318
rect 1344 50202 78624 50236
rect 1344 50150 19838 50202
rect 19890 50150 19942 50202
rect 19994 50150 20046 50202
rect 20098 50150 50558 50202
rect 50610 50150 50662 50202
rect 50714 50150 50766 50202
rect 50818 50150 78624 50202
rect 1344 50116 78624 50150
rect 3826 49758 3838 49810
rect 3890 49758 3902 49810
rect 1934 49586 1986 49598
rect 1934 49522 1986 49534
rect 1344 49418 78624 49452
rect 1344 49366 4478 49418
rect 4530 49366 4582 49418
rect 4634 49366 4686 49418
rect 4738 49366 35198 49418
rect 35250 49366 35302 49418
rect 35354 49366 35406 49418
rect 35458 49366 65918 49418
rect 65970 49366 66022 49418
rect 66074 49366 66126 49418
rect 66178 49366 78624 49418
rect 1344 49332 78624 49366
rect 1934 49138 1986 49150
rect 1934 49074 1986 49086
rect 3826 48974 3838 49026
rect 3890 48974 3902 49026
rect 77646 48914 77698 48926
rect 77646 48850 77698 48862
rect 78206 48914 78258 48926
rect 78206 48850 78258 48862
rect 77870 48802 77922 48814
rect 77870 48738 77922 48750
rect 1344 48634 78624 48668
rect 1344 48582 19838 48634
rect 19890 48582 19942 48634
rect 19994 48582 20046 48634
rect 20098 48582 50558 48634
rect 50610 48582 50662 48634
rect 50714 48582 50766 48634
rect 50818 48582 78624 48634
rect 1344 48548 78624 48582
rect 2718 48466 2770 48478
rect 2718 48402 2770 48414
rect 3390 48466 3442 48478
rect 3390 48402 3442 48414
rect 2046 48354 2098 48366
rect 2046 48290 2098 48302
rect 77870 48354 77922 48366
rect 77870 48290 77922 48302
rect 2382 48242 2434 48254
rect 77646 48242 77698 48254
rect 2930 48190 2942 48242
rect 2994 48190 3006 48242
rect 3602 48190 3614 48242
rect 3666 48190 3678 48242
rect 2382 48178 2434 48190
rect 77646 48178 77698 48190
rect 78206 48242 78258 48254
rect 78206 48178 78258 48190
rect 1344 47850 78624 47884
rect 1344 47798 4478 47850
rect 4530 47798 4582 47850
rect 4634 47798 4686 47850
rect 4738 47798 35198 47850
rect 35250 47798 35302 47850
rect 35354 47798 35406 47850
rect 35458 47798 65918 47850
rect 65970 47798 66022 47850
rect 66074 47798 66126 47850
rect 66178 47798 78624 47850
rect 1344 47764 78624 47798
rect 2034 47406 2046 47458
rect 2098 47406 2110 47458
rect 78206 47346 78258 47358
rect 78206 47282 78258 47294
rect 2718 47234 2770 47246
rect 2718 47170 2770 47182
rect 77646 47234 77698 47246
rect 77646 47170 77698 47182
rect 77870 47234 77922 47246
rect 77870 47170 77922 47182
rect 1344 47066 78624 47100
rect 1344 47014 19838 47066
rect 19890 47014 19942 47066
rect 19994 47014 20046 47066
rect 20098 47014 50558 47066
rect 50610 47014 50662 47066
rect 50714 47014 50766 47066
rect 50818 47014 78624 47066
rect 1344 46980 78624 47014
rect 3826 46622 3838 46674
rect 3890 46622 3902 46674
rect 1934 46450 1986 46462
rect 1934 46386 1986 46398
rect 1344 46282 78624 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 65918 46282
rect 65970 46230 66022 46282
rect 66074 46230 66126 46282
rect 66178 46230 78624 46282
rect 1344 46196 78624 46230
rect 2382 45890 2434 45902
rect 2382 45826 2434 45838
rect 2718 45890 2770 45902
rect 4286 45890 4338 45902
rect 3602 45838 3614 45890
rect 3666 45838 3678 45890
rect 2718 45826 2770 45838
rect 4286 45826 4338 45838
rect 3054 45778 3106 45790
rect 3054 45714 3106 45726
rect 3390 45778 3442 45790
rect 3390 45714 3442 45726
rect 78206 45778 78258 45790
rect 78206 45714 78258 45726
rect 2046 45666 2098 45678
rect 2046 45602 2098 45614
rect 77646 45666 77698 45678
rect 77646 45602 77698 45614
rect 77870 45666 77922 45678
rect 77870 45602 77922 45614
rect 1344 45498 78624 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 50558 45498
rect 50610 45446 50662 45498
rect 50714 45446 50766 45498
rect 50818 45446 78624 45498
rect 1344 45412 78624 45446
rect 77870 45218 77922 45230
rect 77870 45154 77922 45166
rect 78206 45106 78258 45118
rect 2034 45054 2046 45106
rect 2098 45054 2110 45106
rect 78206 45042 78258 45054
rect 77646 44994 77698 45006
rect 77646 44930 77698 44942
rect 2718 44882 2770 44894
rect 2718 44818 2770 44830
rect 1344 44714 78624 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 65918 44714
rect 65970 44662 66022 44714
rect 66074 44662 66126 44714
rect 66178 44662 78624 44714
rect 1344 44628 78624 44662
rect 2034 44270 2046 44322
rect 2098 44270 2110 44322
rect 2718 44098 2770 44110
rect 2718 44034 2770 44046
rect 78318 44098 78370 44110
rect 78318 44034 78370 44046
rect 1344 43930 78624 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 50558 43930
rect 50610 43878 50662 43930
rect 50714 43878 50766 43930
rect 50818 43878 78624 43930
rect 1344 43844 78624 43878
rect 2046 43762 2098 43774
rect 2046 43698 2098 43710
rect 2718 43650 2770 43662
rect 2718 43586 2770 43598
rect 3054 43538 3106 43550
rect 2258 43486 2270 43538
rect 2322 43486 2334 43538
rect 3054 43474 3106 43486
rect 56590 43538 56642 43550
rect 56590 43474 56642 43486
rect 77086 43538 77138 43550
rect 77086 43474 77138 43486
rect 77422 43538 77474 43550
rect 77422 43474 77474 43486
rect 77646 43538 77698 43550
rect 77646 43474 77698 43486
rect 76974 43426 77026 43438
rect 57026 43374 57038 43426
rect 57090 43374 57102 43426
rect 76974 43362 77026 43374
rect 77310 43426 77362 43438
rect 77310 43362 77362 43374
rect 78206 43426 78258 43438
rect 78206 43362 78258 43374
rect 76626 43262 76638 43314
rect 76690 43311 76702 43314
rect 76962 43311 76974 43314
rect 76690 43265 76974 43311
rect 76690 43262 76702 43265
rect 76962 43262 76974 43265
rect 77026 43262 77038 43314
rect 1344 43146 78624 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 65918 43146
rect 65970 43094 66022 43146
rect 66074 43094 66126 43146
rect 66178 43094 78624 43146
rect 1344 43060 78624 43094
rect 1934 42866 1986 42878
rect 1934 42802 1986 42814
rect 56030 42866 56082 42878
rect 56030 42802 56082 42814
rect 57262 42866 57314 42878
rect 57262 42802 57314 42814
rect 58158 42866 58210 42878
rect 58158 42802 58210 42814
rect 62302 42866 62354 42878
rect 62302 42802 62354 42814
rect 75742 42866 75794 42878
rect 75742 42802 75794 42814
rect 77534 42754 77586 42766
rect 3826 42702 3838 42754
rect 3890 42702 3902 42754
rect 55570 42702 55582 42754
rect 55634 42702 55646 42754
rect 76514 42702 76526 42754
rect 76578 42702 76590 42754
rect 78082 42702 78094 42754
rect 78146 42702 78158 42754
rect 77534 42690 77586 42702
rect 76974 42642 77026 42654
rect 76974 42578 77026 42590
rect 77310 42642 77362 42654
rect 77310 42578 77362 42590
rect 56702 42530 56754 42542
rect 56702 42466 56754 42478
rect 57598 42530 57650 42542
rect 57598 42466 57650 42478
rect 76302 42530 76354 42542
rect 76302 42466 76354 42478
rect 77198 42530 77250 42542
rect 77198 42466 77250 42478
rect 77870 42530 77922 42542
rect 77870 42466 77922 42478
rect 1344 42362 78624 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 50558 42362
rect 50610 42310 50662 42362
rect 50714 42310 50766 42362
rect 50818 42310 78624 42362
rect 1344 42276 78624 42310
rect 55682 42142 55694 42194
rect 55746 42142 55758 42194
rect 56578 42142 56590 42194
rect 56642 42142 56654 42194
rect 57474 42142 57486 42194
rect 57538 42142 57550 42194
rect 75294 42082 75346 42094
rect 75294 42018 75346 42030
rect 4734 41970 4786 41982
rect 3826 41918 3838 41970
rect 3890 41918 3902 41970
rect 4734 41906 4786 41918
rect 60622 41970 60674 41982
rect 60622 41906 60674 41918
rect 61070 41970 61122 41982
rect 62526 41970 62578 41982
rect 61618 41918 61630 41970
rect 61682 41918 61694 41970
rect 61070 41906 61122 41918
rect 62526 41906 62578 41918
rect 62862 41970 62914 41982
rect 62862 41906 62914 41918
rect 63198 41970 63250 41982
rect 63198 41906 63250 41918
rect 64430 41970 64482 41982
rect 64430 41906 64482 41918
rect 65438 41970 65490 41982
rect 65438 41906 65490 41918
rect 65886 41970 65938 41982
rect 65886 41906 65938 41918
rect 74062 41970 74114 41982
rect 74062 41906 74114 41918
rect 74958 41970 75010 41982
rect 75618 41918 75630 41970
rect 75682 41918 75694 41970
rect 74958 41906 75010 41918
rect 54910 41858 54962 41870
rect 54910 41794 54962 41806
rect 55134 41858 55186 41870
rect 55134 41794 55186 41806
rect 57150 41858 57202 41870
rect 57150 41794 57202 41806
rect 58046 41858 58098 41870
rect 62078 41858 62130 41870
rect 60162 41806 60174 41858
rect 60226 41806 60238 41858
rect 58046 41794 58098 41806
rect 62078 41794 62130 41806
rect 62750 41858 62802 41870
rect 62750 41794 62802 41806
rect 64990 41858 65042 41870
rect 64990 41794 65042 41806
rect 69806 41858 69858 41870
rect 69806 41794 69858 41806
rect 70254 41858 70306 41870
rect 70254 41794 70306 41806
rect 70702 41858 70754 41870
rect 70702 41794 70754 41806
rect 71150 41858 71202 41870
rect 71150 41794 71202 41806
rect 74734 41858 74786 41870
rect 74734 41794 74786 41806
rect 77982 41858 78034 41870
rect 77982 41794 78034 41806
rect 1934 41746 1986 41758
rect 1934 41682 1986 41694
rect 55358 41746 55410 41758
rect 55358 41682 55410 41694
rect 56926 41746 56978 41758
rect 56926 41682 56978 41694
rect 57822 41746 57874 41758
rect 69794 41694 69806 41746
rect 69858 41743 69870 41746
rect 70130 41743 70142 41746
rect 69858 41697 70142 41743
rect 69858 41694 69870 41697
rect 70130 41694 70142 41697
rect 70194 41743 70206 41746
rect 71026 41743 71038 41746
rect 70194 41697 71038 41743
rect 70194 41694 70206 41697
rect 71026 41694 71038 41697
rect 71090 41694 71102 41746
rect 57822 41682 57874 41694
rect 1344 41578 78624 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 65918 41578
rect 65970 41526 66022 41578
rect 66074 41526 66126 41578
rect 66178 41526 78624 41578
rect 1344 41492 78624 41526
rect 55582 41410 55634 41422
rect 71150 41410 71202 41422
rect 55906 41358 55918 41410
rect 55970 41358 55982 41410
rect 55582 41346 55634 41358
rect 71150 41346 71202 41358
rect 71598 41410 71650 41422
rect 71598 41346 71650 41358
rect 71710 41410 71762 41422
rect 71710 41346 71762 41358
rect 74398 41410 74450 41422
rect 74722 41358 74734 41410
rect 74786 41358 74798 41410
rect 74398 41346 74450 41358
rect 1934 41298 1986 41310
rect 1934 41234 1986 41246
rect 4734 41298 4786 41310
rect 4734 41234 4786 41246
rect 56366 41298 56418 41310
rect 64990 41298 65042 41310
rect 71374 41298 71426 41310
rect 58930 41246 58942 41298
rect 58994 41246 59006 41298
rect 60610 41246 60622 41298
rect 60674 41246 60686 41298
rect 62402 41246 62414 41298
rect 62466 41246 62478 41298
rect 70466 41246 70478 41298
rect 70530 41246 70542 41298
rect 56366 41234 56418 41246
rect 64990 41234 65042 41246
rect 71374 41234 71426 41246
rect 74174 41298 74226 41310
rect 74174 41234 74226 41246
rect 75070 41298 75122 41310
rect 75070 41234 75122 41246
rect 75294 41298 75346 41310
rect 75294 41234 75346 41246
rect 78094 41298 78146 41310
rect 78094 41234 78146 41246
rect 55358 41186 55410 41198
rect 4162 41134 4174 41186
rect 4226 41134 4238 41186
rect 55358 41122 55410 41134
rect 58494 41186 58546 41198
rect 73614 41186 73666 41198
rect 59378 41134 59390 41186
rect 59442 41134 59454 41186
rect 59938 41134 59950 41186
rect 60002 41134 60014 41186
rect 60498 41134 60510 41186
rect 60562 41134 60574 41186
rect 61618 41134 61630 41186
rect 61682 41134 61694 41186
rect 62514 41134 62526 41186
rect 62578 41134 62590 41186
rect 62850 41134 62862 41186
rect 62914 41134 62926 41186
rect 63410 41134 63422 41186
rect 63474 41134 63486 41186
rect 64306 41134 64318 41186
rect 64370 41134 64382 41186
rect 65650 41134 65662 41186
rect 65714 41134 65726 41186
rect 66770 41134 66782 41186
rect 66834 41134 66846 41186
rect 70130 41134 70142 41186
rect 70194 41134 70206 41186
rect 70914 41134 70926 41186
rect 70978 41134 70990 41186
rect 58494 41122 58546 41134
rect 73614 41122 73666 41134
rect 76078 41186 76130 41198
rect 76078 41122 76130 41134
rect 76526 41186 76578 41198
rect 76526 41122 76578 41134
rect 76974 41186 77026 41198
rect 76974 41122 77026 41134
rect 77534 41186 77586 41198
rect 77534 41122 77586 41134
rect 58158 41074 58210 41086
rect 73278 41074 73330 41086
rect 59154 41022 59166 41074
rect 59218 41022 59230 41074
rect 60946 41022 60958 41074
rect 61010 41022 61022 41074
rect 61954 41022 61966 41074
rect 62018 41022 62030 41074
rect 63522 41022 63534 41074
rect 63586 41022 63598 41074
rect 65762 41022 65774 41074
rect 65826 41022 65838 41074
rect 69570 41022 69582 41074
rect 69634 41022 69646 41074
rect 58158 41010 58210 41022
rect 73278 41010 73330 41022
rect 73838 41074 73890 41086
rect 73838 41010 73890 41022
rect 76750 41074 76802 41086
rect 76750 41010 76802 41022
rect 77422 41074 77474 41086
rect 77422 41010 77474 41022
rect 55022 40962 55074 40974
rect 55022 40898 55074 40910
rect 57150 40962 57202 40974
rect 69022 40962 69074 40974
rect 64306 40910 64318 40962
rect 64370 40910 64382 40962
rect 66546 40910 66558 40962
rect 66610 40910 66622 40962
rect 57150 40898 57202 40910
rect 69022 40898 69074 40910
rect 69246 40962 69298 40974
rect 69246 40898 69298 40910
rect 73390 40962 73442 40974
rect 76302 40962 76354 40974
rect 75618 40910 75630 40962
rect 75682 40910 75694 40962
rect 73390 40898 73442 40910
rect 76302 40898 76354 40910
rect 77198 40962 77250 40974
rect 77198 40898 77250 40910
rect 1344 40794 78624 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 50558 40794
rect 50610 40742 50662 40794
rect 50714 40742 50766 40794
rect 50818 40742 78624 40794
rect 1344 40708 78624 40742
rect 2270 40626 2322 40638
rect 2270 40562 2322 40574
rect 5406 40626 5458 40638
rect 61518 40626 61570 40638
rect 67454 40626 67506 40638
rect 71374 40626 71426 40638
rect 59938 40574 59950 40626
rect 60002 40574 60014 40626
rect 64642 40574 64654 40626
rect 64706 40574 64718 40626
rect 66882 40574 66894 40626
rect 66946 40574 66958 40626
rect 67890 40574 67902 40626
rect 67954 40574 67966 40626
rect 5406 40562 5458 40574
rect 61518 40562 61570 40574
rect 67454 40562 67506 40574
rect 71374 40562 71426 40574
rect 72942 40626 72994 40638
rect 72942 40562 72994 40574
rect 73950 40626 74002 40638
rect 73950 40562 74002 40574
rect 74622 40626 74674 40638
rect 74622 40562 74674 40574
rect 75182 40626 75234 40638
rect 75182 40562 75234 40574
rect 4062 40514 4114 40526
rect 4062 40450 4114 40462
rect 4510 40514 4562 40526
rect 62974 40514 63026 40526
rect 70926 40514 70978 40526
rect 60722 40462 60734 40514
rect 60786 40462 60798 40514
rect 63522 40462 63534 40514
rect 63586 40462 63598 40514
rect 65090 40462 65102 40514
rect 65154 40462 65166 40514
rect 66322 40462 66334 40514
rect 66386 40462 66398 40514
rect 69346 40462 69358 40514
rect 69410 40462 69422 40514
rect 4510 40450 4562 40462
rect 62974 40450 63026 40462
rect 70926 40450 70978 40462
rect 73614 40514 73666 40526
rect 73614 40450 73666 40462
rect 74286 40514 74338 40526
rect 76626 40462 76638 40514
rect 76690 40462 76702 40514
rect 74286 40450 74338 40462
rect 1710 40402 1762 40414
rect 1710 40338 1762 40350
rect 2606 40402 2658 40414
rect 2606 40338 2658 40350
rect 3166 40402 3218 40414
rect 3166 40338 3218 40350
rect 3502 40402 3554 40414
rect 3502 40338 3554 40350
rect 4958 40402 5010 40414
rect 61742 40402 61794 40414
rect 60050 40350 60062 40402
rect 60114 40350 60126 40402
rect 60498 40350 60510 40402
rect 60562 40350 60574 40402
rect 4958 40338 5010 40350
rect 61742 40338 61794 40350
rect 62302 40402 62354 40414
rect 62302 40338 62354 40350
rect 62638 40402 62690 40414
rect 62638 40338 62690 40350
rect 63198 40402 63250 40414
rect 68238 40402 68290 40414
rect 70142 40402 70194 40414
rect 73390 40402 73442 40414
rect 63746 40350 63758 40402
rect 63810 40350 63822 40402
rect 64418 40350 64430 40402
rect 64482 40350 64494 40402
rect 65538 40350 65550 40402
rect 65602 40350 65614 40402
rect 65874 40350 65886 40402
rect 65938 40350 65950 40402
rect 66770 40350 66782 40402
rect 66834 40350 66846 40402
rect 68562 40350 68574 40402
rect 68626 40350 68638 40402
rect 69682 40350 69694 40402
rect 69746 40350 69758 40402
rect 70690 40350 70702 40402
rect 70754 40350 70766 40402
rect 77858 40350 77870 40402
rect 77922 40350 77934 40402
rect 63198 40338 63250 40350
rect 68238 40338 68290 40350
rect 70142 40338 70194 40350
rect 73390 40338 73442 40350
rect 62750 40290 62802 40302
rect 72494 40290 72546 40302
rect 69458 40238 69470 40290
rect 69522 40238 69534 40290
rect 62750 40226 62802 40238
rect 72494 40226 72546 40238
rect 74958 40178 75010 40190
rect 74958 40114 75010 40126
rect 75294 40178 75346 40190
rect 75294 40114 75346 40126
rect 1344 40010 78624 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 65918 40010
rect 65970 39958 66022 40010
rect 66074 39958 66126 40010
rect 66178 39958 78624 40010
rect 1344 39924 78624 39958
rect 1934 39730 1986 39742
rect 1934 39666 1986 39678
rect 61294 39730 61346 39742
rect 61294 39666 61346 39678
rect 61854 39730 61906 39742
rect 61854 39666 61906 39678
rect 63422 39730 63474 39742
rect 63422 39666 63474 39678
rect 67118 39730 67170 39742
rect 67118 39666 67170 39678
rect 71934 39730 71986 39742
rect 74622 39730 74674 39742
rect 72930 39678 72942 39730
rect 72994 39678 73006 39730
rect 76738 39678 76750 39730
rect 76802 39678 76814 39730
rect 71934 39666 71986 39678
rect 74622 39666 74674 39678
rect 4734 39618 4786 39630
rect 3826 39566 3838 39618
rect 3890 39566 3902 39618
rect 4734 39554 4786 39566
rect 65214 39618 65266 39630
rect 70366 39618 70418 39630
rect 65538 39566 65550 39618
rect 65602 39566 65614 39618
rect 66658 39566 66670 39618
rect 66722 39566 66734 39618
rect 68338 39566 68350 39618
rect 68402 39566 68414 39618
rect 69234 39566 69246 39618
rect 69298 39566 69310 39618
rect 65214 39554 65266 39566
rect 70366 39554 70418 39566
rect 70590 39618 70642 39630
rect 70590 39554 70642 39566
rect 71374 39618 71426 39630
rect 71374 39554 71426 39566
rect 72382 39618 72434 39630
rect 75070 39618 75122 39630
rect 73154 39566 73166 39618
rect 73218 39566 73230 39618
rect 73602 39566 73614 39618
rect 73666 39566 73678 39618
rect 74050 39566 74062 39618
rect 74114 39566 74126 39618
rect 72382 39554 72434 39566
rect 75070 39554 75122 39566
rect 75406 39618 75458 39630
rect 75406 39554 75458 39566
rect 75518 39618 75570 39630
rect 76514 39566 76526 39618
rect 76578 39566 76590 39618
rect 77298 39566 77310 39618
rect 77362 39566 77374 39618
rect 78082 39566 78094 39618
rect 78146 39566 78158 39618
rect 75518 39554 75570 39566
rect 70030 39506 70082 39518
rect 65762 39454 65774 39506
rect 65826 39454 65838 39506
rect 68450 39454 68462 39506
rect 68514 39454 68526 39506
rect 70030 39442 70082 39454
rect 70926 39506 70978 39518
rect 70926 39442 70978 39454
rect 71262 39506 71314 39518
rect 77870 39506 77922 39518
rect 76402 39454 76414 39506
rect 76466 39454 76478 39506
rect 71262 39442 71314 39454
rect 77870 39442 77922 39454
rect 64654 39394 64706 39406
rect 67566 39394 67618 39406
rect 70254 39394 70306 39406
rect 66434 39342 66446 39394
rect 66498 39342 66510 39394
rect 69346 39342 69358 39394
rect 69410 39342 69422 39394
rect 64654 39330 64706 39342
rect 67566 39330 67618 39342
rect 70254 39330 70306 39342
rect 71150 39394 71202 39406
rect 71150 39330 71202 39342
rect 75294 39394 75346 39406
rect 75294 39330 75346 39342
rect 1344 39226 78624 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 50558 39226
rect 50610 39174 50662 39226
rect 50714 39174 50766 39226
rect 50818 39174 78624 39226
rect 1344 39140 78624 39174
rect 43598 39058 43650 39070
rect 42018 39006 42030 39058
rect 42082 39006 42094 39058
rect 43598 38994 43650 39006
rect 62190 39058 62242 39070
rect 62190 38994 62242 39006
rect 65326 39058 65378 39070
rect 65326 38994 65378 39006
rect 69246 39058 69298 39070
rect 69246 38994 69298 39006
rect 71374 39058 71426 39070
rect 71374 38994 71426 39006
rect 73502 39058 73554 39070
rect 73502 38994 73554 39006
rect 74398 39058 74450 39070
rect 74398 38994 74450 39006
rect 41246 38946 41298 38958
rect 41246 38882 41298 38894
rect 41470 38946 41522 38958
rect 43038 38946 43090 38958
rect 42578 38894 42590 38946
rect 42642 38894 42654 38946
rect 41470 38882 41522 38894
rect 43038 38882 43090 38894
rect 43262 38946 43314 38958
rect 43262 38882 43314 38894
rect 61854 38946 61906 38958
rect 69694 38946 69746 38958
rect 67106 38894 67118 38946
rect 67170 38894 67182 38946
rect 68002 38894 68014 38946
rect 68066 38894 68078 38946
rect 61854 38882 61906 38894
rect 69694 38882 69746 38894
rect 70926 38946 70978 38958
rect 70926 38882 70978 38894
rect 72718 38946 72770 38958
rect 72718 38882 72770 38894
rect 73054 38946 73106 38958
rect 73054 38882 73106 38894
rect 73278 38946 73330 38958
rect 73278 38882 73330 38894
rect 75182 38946 75234 38958
rect 75182 38882 75234 38894
rect 76190 38946 76242 38958
rect 77634 38894 77646 38946
rect 77698 38894 77710 38946
rect 76190 38882 76242 38894
rect 41582 38834 41634 38846
rect 42926 38834 42978 38846
rect 2034 38782 2046 38834
rect 2098 38782 2110 38834
rect 42018 38782 42030 38834
rect 42082 38782 42094 38834
rect 41582 38770 41634 38782
rect 42926 38770 42978 38782
rect 44046 38834 44098 38846
rect 44046 38770 44098 38782
rect 62526 38834 62578 38846
rect 62526 38770 62578 38782
rect 65886 38834 65938 38846
rect 70366 38834 70418 38846
rect 66322 38782 66334 38834
rect 66386 38782 66398 38834
rect 67330 38782 67342 38834
rect 67394 38782 67406 38834
rect 68226 38782 68238 38834
rect 68290 38782 68302 38834
rect 68562 38782 68574 38834
rect 68626 38782 68638 38834
rect 65886 38770 65938 38782
rect 70366 38770 70418 38782
rect 70702 38834 70754 38846
rect 73726 38834 73778 38846
rect 74846 38834 74898 38846
rect 72482 38782 72494 38834
rect 72546 38782 72558 38834
rect 74162 38782 74174 38834
rect 74226 38782 74238 38834
rect 70702 38770 70754 38782
rect 73726 38770 73778 38782
rect 74846 38770 74898 38782
rect 75630 38834 75682 38846
rect 75630 38770 75682 38782
rect 75966 38834 76018 38846
rect 75966 38770 76018 38782
rect 76638 38834 76690 38846
rect 77074 38782 77086 38834
rect 77138 38782 77150 38834
rect 77522 38782 77534 38834
rect 77586 38782 77598 38834
rect 78082 38782 78094 38834
rect 78146 38782 78158 38834
rect 76638 38770 76690 38782
rect 41134 38722 41186 38734
rect 70478 38722 70530 38734
rect 3378 38670 3390 38722
rect 3442 38670 3454 38722
rect 66658 38670 66670 38722
rect 66722 38670 66734 38722
rect 67890 38670 67902 38722
rect 67954 38670 67966 38722
rect 41134 38658 41186 38670
rect 70478 38658 70530 38670
rect 76414 38722 76466 38734
rect 76414 38658 76466 38670
rect 1344 38442 78624 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 65918 38442
rect 65970 38390 66022 38442
rect 66074 38390 66126 38442
rect 66178 38390 78624 38442
rect 1344 38356 78624 38390
rect 2942 38162 2994 38174
rect 2034 38110 2046 38162
rect 2098 38110 2110 38162
rect 2942 38098 2994 38110
rect 67230 38162 67282 38174
rect 67230 38098 67282 38110
rect 70590 38162 70642 38174
rect 70590 38098 70642 38110
rect 72942 38162 72994 38174
rect 72942 38098 72994 38110
rect 75630 38162 75682 38174
rect 75630 38098 75682 38110
rect 77534 38162 77586 38174
rect 77534 38098 77586 38110
rect 78206 38162 78258 38174
rect 78206 38098 78258 38110
rect 2494 38050 2546 38062
rect 69806 38050 69858 38062
rect 68338 37998 68350 38050
rect 68402 37998 68414 38050
rect 69234 37998 69246 38050
rect 69298 37998 69310 38050
rect 2494 37986 2546 37998
rect 69806 37986 69858 37998
rect 71038 38050 71090 38062
rect 71038 37986 71090 37998
rect 71262 38050 71314 38062
rect 71262 37986 71314 37998
rect 72158 38050 72210 38062
rect 72158 37986 72210 37998
rect 73166 38050 73218 38062
rect 73166 37986 73218 37998
rect 73278 38050 73330 38062
rect 73278 37986 73330 37998
rect 74286 38050 74338 38062
rect 74286 37986 74338 37998
rect 74622 38050 74674 38062
rect 74622 37986 74674 37998
rect 75070 38050 75122 38062
rect 75070 37986 75122 37998
rect 76190 38050 76242 38062
rect 76190 37986 76242 37998
rect 76638 38050 76690 38062
rect 76638 37986 76690 37998
rect 77086 38050 77138 38062
rect 77086 37986 77138 37998
rect 70142 37938 70194 37950
rect 68450 37886 68462 37938
rect 68514 37886 68526 37938
rect 70142 37874 70194 37886
rect 71598 37938 71650 37950
rect 71598 37874 71650 37886
rect 72830 37938 72882 37950
rect 72830 37874 72882 37886
rect 73726 37938 73778 37950
rect 73726 37874 73778 37886
rect 73950 37938 74002 37950
rect 73950 37874 74002 37886
rect 74958 37938 75010 37950
rect 74958 37874 75010 37886
rect 76526 37938 76578 37950
rect 76526 37874 76578 37886
rect 77310 37938 77362 37950
rect 77310 37874 77362 37886
rect 77646 37938 77698 37950
rect 77646 37874 77698 37886
rect 67790 37826 67842 37838
rect 71486 37826 71538 37838
rect 69234 37774 69246 37826
rect 69298 37774 69310 37826
rect 67790 37762 67842 37774
rect 71486 37762 71538 37774
rect 72494 37826 72546 37838
rect 72494 37762 72546 37774
rect 74062 37826 74114 37838
rect 74062 37762 74114 37774
rect 74734 37826 74786 37838
rect 74734 37762 74786 37774
rect 76302 37826 76354 37838
rect 76302 37762 76354 37774
rect 1344 37658 78624 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 50558 37658
rect 50610 37606 50662 37658
rect 50714 37606 50766 37658
rect 50818 37606 78624 37658
rect 1344 37572 78624 37606
rect 68126 37490 68178 37502
rect 68126 37426 68178 37438
rect 68686 37490 68738 37502
rect 69694 37490 69746 37502
rect 69010 37438 69022 37490
rect 69074 37438 69086 37490
rect 68686 37426 68738 37438
rect 69694 37426 69746 37438
rect 70926 37490 70978 37502
rect 75070 37490 75122 37502
rect 71586 37438 71598 37490
rect 71650 37438 71662 37490
rect 70926 37426 70978 37438
rect 75070 37426 75122 37438
rect 76414 37490 76466 37502
rect 76414 37426 76466 37438
rect 70590 37378 70642 37390
rect 2034 37326 2046 37378
rect 2098 37326 2110 37378
rect 70590 37314 70642 37326
rect 71262 37378 71314 37390
rect 71262 37314 71314 37326
rect 72270 37378 72322 37390
rect 72270 37314 72322 37326
rect 74510 37378 74562 37390
rect 74510 37314 74562 37326
rect 74846 37378 74898 37390
rect 74846 37314 74898 37326
rect 75406 37378 75458 37390
rect 75406 37314 75458 37326
rect 75966 37378 76018 37390
rect 75966 37314 76018 37326
rect 1710 37266 1762 37278
rect 1710 37202 1762 37214
rect 69358 37266 69410 37278
rect 69358 37202 69410 37214
rect 72494 37266 72546 37278
rect 72494 37202 72546 37214
rect 72718 37266 72770 37278
rect 72718 37202 72770 37214
rect 73054 37266 73106 37278
rect 73054 37202 73106 37214
rect 73390 37266 73442 37278
rect 73390 37202 73442 37214
rect 73614 37266 73666 37278
rect 75182 37266 75234 37278
rect 74274 37214 74286 37266
rect 74338 37214 74350 37266
rect 73614 37202 73666 37214
rect 75182 37202 75234 37214
rect 76190 37266 76242 37278
rect 76190 37202 76242 37214
rect 76638 37266 76690 37278
rect 77186 37214 77198 37266
rect 77250 37214 77262 37266
rect 77858 37214 77870 37266
rect 77922 37214 77934 37266
rect 76638 37202 76690 37214
rect 2494 37154 2546 37166
rect 2494 37090 2546 37102
rect 72382 37154 72434 37166
rect 72382 37090 72434 37102
rect 73278 37154 73330 37166
rect 77298 37102 77310 37154
rect 77362 37102 77374 37154
rect 73278 37090 73330 37102
rect 77410 36990 77422 37042
rect 77474 36990 77486 37042
rect 1344 36874 78624 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 65918 36874
rect 65970 36822 66022 36874
rect 66074 36822 66126 36874
rect 66178 36822 78624 36874
rect 1344 36788 78624 36822
rect 74958 36706 75010 36718
rect 72482 36654 72494 36706
rect 72546 36703 72558 36706
rect 73266 36703 73278 36706
rect 72546 36657 73278 36703
rect 72546 36654 72558 36657
rect 73266 36654 73278 36657
rect 73330 36654 73342 36706
rect 74958 36642 75010 36654
rect 77870 36706 77922 36718
rect 77870 36642 77922 36654
rect 71262 36594 71314 36606
rect 71262 36530 71314 36542
rect 71934 36594 71986 36606
rect 71934 36530 71986 36542
rect 72942 36594 72994 36606
rect 72942 36530 72994 36542
rect 73278 36594 73330 36606
rect 73278 36530 73330 36542
rect 74846 36594 74898 36606
rect 77982 36594 78034 36606
rect 76402 36542 76414 36594
rect 76466 36542 76478 36594
rect 76738 36542 76750 36594
rect 76802 36542 76814 36594
rect 74846 36530 74898 36542
rect 77982 36530 78034 36542
rect 72494 36482 72546 36494
rect 74610 36430 74622 36482
rect 74674 36430 74686 36482
rect 75394 36430 75406 36482
rect 75458 36430 75470 36482
rect 76178 36430 76190 36482
rect 76242 36430 76254 36482
rect 76850 36430 76862 36482
rect 76914 36430 76926 36482
rect 78194 36430 78206 36482
rect 78258 36430 78270 36482
rect 72494 36418 72546 36430
rect 1710 36370 1762 36382
rect 1710 36306 1762 36318
rect 44830 36370 44882 36382
rect 44830 36306 44882 36318
rect 45390 36370 45442 36382
rect 45390 36306 45442 36318
rect 73950 36370 74002 36382
rect 73950 36306 74002 36318
rect 74398 36370 74450 36382
rect 74398 36306 74450 36318
rect 2046 36258 2098 36270
rect 2046 36194 2098 36206
rect 2494 36258 2546 36270
rect 2494 36194 2546 36206
rect 44942 36258 44994 36270
rect 44942 36194 44994 36206
rect 69022 36258 69074 36270
rect 69022 36194 69074 36206
rect 75630 36258 75682 36270
rect 75630 36194 75682 36206
rect 1344 36090 78624 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 50558 36090
rect 50610 36038 50662 36090
rect 50714 36038 50766 36090
rect 50818 36038 78624 36090
rect 1344 36004 78624 36038
rect 44270 35922 44322 35934
rect 44270 35858 44322 35870
rect 54350 35922 54402 35934
rect 54350 35858 54402 35870
rect 72942 35922 72994 35934
rect 72942 35858 72994 35870
rect 77646 35922 77698 35934
rect 77646 35858 77698 35870
rect 78206 35922 78258 35934
rect 78206 35858 78258 35870
rect 44606 35810 44658 35822
rect 44606 35746 44658 35758
rect 45838 35810 45890 35822
rect 45838 35746 45890 35758
rect 46622 35810 46674 35822
rect 46622 35746 46674 35758
rect 46958 35810 47010 35822
rect 46958 35746 47010 35758
rect 73278 35810 73330 35822
rect 73278 35746 73330 35758
rect 73614 35810 73666 35822
rect 73614 35746 73666 35758
rect 74174 35810 74226 35822
rect 74174 35746 74226 35758
rect 74510 35810 74562 35822
rect 74510 35746 74562 35758
rect 75182 35810 75234 35822
rect 76526 35810 76578 35822
rect 76066 35758 76078 35810
rect 76130 35758 76142 35810
rect 75182 35746 75234 35758
rect 76526 35746 76578 35758
rect 76862 35810 76914 35822
rect 76862 35746 76914 35758
rect 44718 35698 44770 35710
rect 44718 35634 44770 35646
rect 45390 35698 45442 35710
rect 45390 35634 45442 35646
rect 45950 35698 46002 35710
rect 45950 35634 46002 35646
rect 46398 35698 46450 35710
rect 46398 35634 46450 35646
rect 72606 35698 72658 35710
rect 72606 35634 72658 35646
rect 73950 35698 74002 35710
rect 73950 35634 74002 35646
rect 74734 35698 74786 35710
rect 74734 35634 74786 35646
rect 75294 35698 75346 35710
rect 75294 35634 75346 35646
rect 75742 35698 75794 35710
rect 75742 35634 75794 35646
rect 76974 35698 77026 35710
rect 76974 35634 77026 35646
rect 77870 35698 77922 35710
rect 77870 35634 77922 35646
rect 45614 35586 45666 35598
rect 45614 35522 45666 35534
rect 46846 35586 46898 35598
rect 46846 35522 46898 35534
rect 71710 35586 71762 35598
rect 71710 35522 71762 35534
rect 74398 35586 74450 35598
rect 74398 35522 74450 35534
rect 74958 35586 75010 35598
rect 74958 35522 75010 35534
rect 76638 35586 76690 35598
rect 76638 35522 76690 35534
rect 54002 35422 54014 35474
rect 54066 35471 54078 35474
rect 54338 35471 54350 35474
rect 54066 35425 54350 35471
rect 54066 35422 54078 35425
rect 54338 35422 54350 35425
rect 54402 35422 54414 35474
rect 1344 35306 78624 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 65918 35306
rect 65970 35254 66022 35306
rect 66074 35254 66126 35306
rect 66178 35254 78624 35306
rect 1344 35220 78624 35254
rect 77870 35138 77922 35150
rect 77870 35074 77922 35086
rect 55582 35026 55634 35038
rect 55582 34962 55634 34974
rect 75406 35026 75458 35038
rect 76514 34974 76526 35026
rect 76578 34974 76590 35026
rect 76738 34974 76750 35026
rect 76802 34974 76814 35026
rect 78082 34974 78094 35026
rect 78146 34974 78158 35026
rect 75406 34962 75458 34974
rect 44942 34914 44994 34926
rect 44942 34850 44994 34862
rect 45390 34914 45442 34926
rect 45390 34850 45442 34862
rect 45614 34914 45666 34926
rect 45614 34850 45666 34862
rect 45838 34914 45890 34926
rect 45838 34850 45890 34862
rect 45950 34914 46002 34926
rect 71262 34914 71314 34926
rect 53554 34862 53566 34914
rect 53618 34862 53630 34914
rect 54450 34862 54462 34914
rect 54514 34862 54526 34914
rect 45950 34850 46002 34862
rect 71262 34850 71314 34862
rect 71598 34914 71650 34926
rect 71598 34850 71650 34862
rect 71822 34914 71874 34926
rect 71822 34850 71874 34862
rect 72158 34914 72210 34926
rect 72158 34850 72210 34862
rect 72830 34914 72882 34926
rect 72830 34850 72882 34862
rect 73054 34914 73106 34926
rect 73054 34850 73106 34862
rect 73278 34914 73330 34926
rect 73278 34850 73330 34862
rect 73502 34914 73554 34926
rect 73502 34850 73554 34862
rect 73838 34914 73890 34926
rect 73838 34850 73890 34862
rect 74062 34914 74114 34926
rect 74722 34862 74734 34914
rect 74786 34862 74798 34914
rect 76066 34862 76078 34914
rect 76130 34862 76142 34914
rect 76850 34862 76862 34914
rect 76914 34862 76926 34914
rect 78194 34862 78206 34914
rect 78258 34862 78270 34914
rect 74062 34850 74114 34862
rect 1710 34802 1762 34814
rect 1710 34738 1762 34750
rect 2494 34802 2546 34814
rect 2494 34738 2546 34750
rect 44830 34802 44882 34814
rect 70926 34802 70978 34814
rect 54002 34750 54014 34802
rect 54066 34750 54078 34802
rect 54786 34750 54798 34802
rect 54850 34750 54862 34802
rect 44830 34738 44882 34750
rect 70926 34738 70978 34750
rect 72382 34802 72434 34814
rect 72382 34738 72434 34750
rect 75294 34802 75346 34814
rect 75294 34738 75346 34750
rect 2046 34690 2098 34702
rect 2046 34626 2098 34638
rect 44382 34690 44434 34702
rect 71374 34690 71426 34702
rect 53554 34638 53566 34690
rect 53618 34638 53630 34690
rect 55010 34638 55022 34690
rect 55074 34638 55086 34690
rect 44382 34626 44434 34638
rect 71374 34626 71426 34638
rect 71934 34690 71986 34702
rect 71934 34626 71986 34638
rect 73054 34690 73106 34702
rect 73054 34626 73106 34638
rect 73726 34690 73778 34702
rect 73726 34626 73778 34638
rect 74958 34690 75010 34702
rect 74958 34626 75010 34638
rect 75518 34690 75570 34702
rect 75518 34626 75570 34638
rect 1344 34522 78624 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 50558 34522
rect 50610 34470 50662 34522
rect 50714 34470 50766 34522
rect 50818 34470 78624 34522
rect 1344 34436 78624 34470
rect 55470 34354 55522 34366
rect 55470 34290 55522 34302
rect 71822 34354 71874 34366
rect 71822 34290 71874 34302
rect 72494 34354 72546 34366
rect 72494 34290 72546 34302
rect 73390 34354 73442 34366
rect 73390 34290 73442 34302
rect 73838 34354 73890 34366
rect 73838 34290 73890 34302
rect 75966 34354 76018 34366
rect 75966 34290 76018 34302
rect 78206 34354 78258 34366
rect 78206 34290 78258 34302
rect 2046 34242 2098 34254
rect 2046 34178 2098 34190
rect 44158 34242 44210 34254
rect 44158 34178 44210 34190
rect 44382 34242 44434 34254
rect 71374 34242 71426 34254
rect 53330 34190 53342 34242
rect 53394 34190 53406 34242
rect 54562 34190 54574 34242
rect 54626 34190 54638 34242
rect 44382 34178 44434 34190
rect 71374 34178 71426 34190
rect 76302 34242 76354 34254
rect 76302 34178 76354 34190
rect 76638 34242 76690 34254
rect 76638 34178 76690 34190
rect 77534 34242 77586 34254
rect 77534 34178 77586 34190
rect 1710 34130 1762 34142
rect 76414 34130 76466 34142
rect 52994 34078 53006 34130
rect 53058 34078 53070 34130
rect 54226 34078 54238 34130
rect 54290 34078 54302 34130
rect 72706 34078 72718 34130
rect 72770 34078 72782 34130
rect 73042 34078 73054 34130
rect 73106 34078 73118 34130
rect 74722 34078 74734 34130
rect 74786 34078 74798 34130
rect 75058 34078 75070 34130
rect 75122 34078 75134 34130
rect 1710 34066 1762 34078
rect 2494 34018 2546 34030
rect 54562 33966 54574 34018
rect 54626 33966 54638 34018
rect 2494 33954 2546 33966
rect 44494 33906 44546 33918
rect 44494 33842 44546 33854
rect 53118 33906 53170 33918
rect 73057 33903 73103 34078
rect 76414 34066 76466 34078
rect 76862 34130 76914 34142
rect 76862 34066 76914 34078
rect 77086 34130 77138 34142
rect 77086 34066 77138 34078
rect 77646 34130 77698 34142
rect 77646 34066 77698 34078
rect 77310 34018 77362 34030
rect 74834 33966 74846 34018
rect 74898 33966 74910 34018
rect 77310 33954 77362 33966
rect 73602 33903 73614 33906
rect 73057 33857 73614 33903
rect 73602 33854 73614 33857
rect 73666 33854 73678 33906
rect 74722 33854 74734 33906
rect 74786 33854 74798 33906
rect 53118 33842 53170 33854
rect 1344 33738 78624 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 65918 33738
rect 65970 33686 66022 33738
rect 66074 33686 66126 33738
rect 66178 33686 78624 33738
rect 1344 33652 78624 33686
rect 76750 33570 76802 33582
rect 76750 33506 76802 33518
rect 54014 33458 54066 33470
rect 54014 33394 54066 33406
rect 72718 33458 72770 33470
rect 72718 33394 72770 33406
rect 73390 33458 73442 33470
rect 76526 33458 76578 33470
rect 74386 33406 74398 33458
rect 74450 33406 74462 33458
rect 74834 33406 74846 33458
rect 74898 33406 74910 33458
rect 73390 33394 73442 33406
rect 76526 33394 76578 33406
rect 78206 33458 78258 33470
rect 78206 33394 78258 33406
rect 45390 33346 45442 33358
rect 45390 33282 45442 33294
rect 45838 33346 45890 33358
rect 45838 33282 45890 33294
rect 72046 33346 72098 33358
rect 72046 33282 72098 33294
rect 72158 33346 72210 33358
rect 72158 33282 72210 33294
rect 73614 33346 73666 33358
rect 74610 33294 74622 33346
rect 74674 33294 74686 33346
rect 75282 33294 75294 33346
rect 75346 33294 75358 33346
rect 77522 33294 77534 33346
rect 77586 33294 77598 33346
rect 73614 33282 73666 33294
rect 46062 33234 46114 33246
rect 71710 33234 71762 33246
rect 46386 33182 46398 33234
rect 46450 33182 46462 33234
rect 46062 33170 46114 33182
rect 71710 33170 71762 33182
rect 76862 33234 76914 33246
rect 76862 33170 76914 33182
rect 77086 33234 77138 33246
rect 77746 33182 77758 33234
rect 77810 33182 77822 33234
rect 77086 33170 77138 33182
rect 1710 33122 1762 33134
rect 2494 33122 2546 33134
rect 2034 33070 2046 33122
rect 2098 33070 2110 33122
rect 1710 33058 1762 33070
rect 2494 33058 2546 33070
rect 45726 33122 45778 33134
rect 45726 33058 45778 33070
rect 46734 33122 46786 33134
rect 46734 33058 46786 33070
rect 71822 33122 71874 33134
rect 71822 33058 71874 33070
rect 73950 33122 74002 33134
rect 73950 33058 74002 33070
rect 1344 32954 78624 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 50558 32954
rect 50610 32902 50662 32954
rect 50714 32902 50766 32954
rect 50818 32902 78624 32954
rect 1344 32868 78624 32902
rect 46062 32786 46114 32798
rect 46062 32722 46114 32734
rect 74846 32786 74898 32798
rect 76750 32786 76802 32798
rect 75618 32734 75630 32786
rect 75682 32734 75694 32786
rect 74846 32722 74898 32734
rect 76750 32722 76802 32734
rect 77870 32786 77922 32798
rect 77870 32722 77922 32734
rect 45390 32674 45442 32686
rect 45390 32610 45442 32622
rect 46734 32674 46786 32686
rect 46734 32610 46786 32622
rect 71374 32674 71426 32686
rect 71374 32610 71426 32622
rect 72606 32674 72658 32686
rect 72606 32610 72658 32622
rect 73166 32674 73218 32686
rect 73166 32610 73218 32622
rect 74286 32674 74338 32686
rect 74286 32610 74338 32622
rect 74958 32674 75010 32686
rect 74958 32610 75010 32622
rect 76862 32674 76914 32686
rect 76862 32610 76914 32622
rect 71262 32562 71314 32574
rect 45826 32510 45838 32562
rect 45890 32510 45902 32562
rect 46498 32510 46510 32562
rect 46562 32510 46574 32562
rect 71262 32498 71314 32510
rect 71710 32562 71762 32574
rect 71710 32498 71762 32510
rect 72158 32562 72210 32574
rect 72158 32498 72210 32510
rect 72830 32562 72882 32574
rect 75294 32562 75346 32574
rect 73378 32510 73390 32562
rect 73442 32510 73454 32562
rect 74050 32510 74062 32562
rect 74114 32510 74126 32562
rect 74610 32510 74622 32562
rect 74674 32510 74686 32562
rect 72830 32498 72882 32510
rect 75294 32498 75346 32510
rect 76414 32562 76466 32574
rect 76414 32498 76466 32510
rect 76974 32562 77026 32574
rect 76974 32498 77026 32510
rect 77646 32562 77698 32574
rect 77646 32498 77698 32510
rect 78206 32562 78258 32574
rect 78206 32498 78258 32510
rect 45054 32450 45106 32462
rect 45054 32386 45106 32398
rect 71598 32450 71650 32462
rect 71598 32386 71650 32398
rect 72382 32450 72434 32462
rect 72382 32386 72434 32398
rect 76078 32450 76130 32462
rect 76078 32386 76130 32398
rect 1344 32170 78624 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 65918 32170
rect 65970 32118 66022 32170
rect 66074 32118 66126 32170
rect 66178 32118 78624 32170
rect 1344 32084 78624 32118
rect 77534 32002 77586 32014
rect 72594 31950 72606 32002
rect 72658 31999 72670 32002
rect 73154 31999 73166 32002
rect 72658 31953 73166 31999
rect 72658 31950 72670 31953
rect 73154 31950 73166 31953
rect 73218 31950 73230 32002
rect 76962 31950 76974 32002
rect 77026 31999 77038 32002
rect 77186 31999 77198 32002
rect 77026 31953 77198 31999
rect 77026 31950 77038 31953
rect 77186 31950 77198 31953
rect 77250 31950 77262 32002
rect 77534 31938 77586 31950
rect 77870 32002 77922 32014
rect 77870 31938 77922 31950
rect 45278 31890 45330 31902
rect 45278 31826 45330 31838
rect 73166 31890 73218 31902
rect 73166 31826 73218 31838
rect 74734 31890 74786 31902
rect 74734 31826 74786 31838
rect 77310 31890 77362 31902
rect 77310 31826 77362 31838
rect 44942 31778 44994 31790
rect 44942 31714 44994 31726
rect 45726 31778 45778 31790
rect 45726 31714 45778 31726
rect 45950 31778 46002 31790
rect 45950 31714 46002 31726
rect 46286 31778 46338 31790
rect 52782 31778 52834 31790
rect 51426 31726 51438 31778
rect 51490 31726 51502 31778
rect 46286 31714 46338 31726
rect 52782 31714 52834 31726
rect 72046 31778 72098 31790
rect 72046 31714 72098 31726
rect 73278 31778 73330 31790
rect 73278 31714 73330 31726
rect 75070 31778 75122 31790
rect 75070 31714 75122 31726
rect 76190 31778 76242 31790
rect 76190 31714 76242 31726
rect 76414 31778 76466 31790
rect 76414 31714 76466 31726
rect 76638 31778 76690 31790
rect 76638 31714 76690 31726
rect 1710 31666 1762 31678
rect 1710 31602 1762 31614
rect 2046 31666 2098 31678
rect 2046 31602 2098 31614
rect 44382 31666 44434 31678
rect 44382 31602 44434 31614
rect 44830 31666 44882 31678
rect 44830 31602 44882 31614
rect 45390 31666 45442 31678
rect 45390 31602 45442 31614
rect 46174 31666 46226 31678
rect 72718 31666 72770 31678
rect 51538 31614 51550 31666
rect 51602 31614 51614 31666
rect 46174 31602 46226 31614
rect 72718 31602 72770 31614
rect 2494 31554 2546 31566
rect 73726 31554 73778 31566
rect 51762 31502 51774 31554
rect 51826 31502 51838 31554
rect 2494 31490 2546 31502
rect 73726 31490 73778 31502
rect 73838 31554 73890 31566
rect 73838 31490 73890 31502
rect 73950 31554 74002 31566
rect 73950 31490 74002 31502
rect 75406 31554 75458 31566
rect 75406 31490 75458 31502
rect 76302 31554 76354 31566
rect 76302 31490 76354 31502
rect 77758 31554 77810 31566
rect 77758 31490 77810 31502
rect 1344 31386 78624 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 50558 31386
rect 50610 31334 50662 31386
rect 50714 31334 50766 31386
rect 50818 31334 78624 31386
rect 1344 31300 78624 31334
rect 53678 31218 53730 31230
rect 53678 31154 53730 31166
rect 73390 31218 73442 31230
rect 73390 31154 73442 31166
rect 74062 31218 74114 31230
rect 74062 31154 74114 31166
rect 74846 31218 74898 31230
rect 74846 31154 74898 31166
rect 75182 31218 75234 31230
rect 75182 31154 75234 31166
rect 77310 31218 77362 31230
rect 77310 31154 77362 31166
rect 77534 31218 77586 31230
rect 77534 31154 77586 31166
rect 2046 31106 2098 31118
rect 2046 31042 2098 31054
rect 44158 31106 44210 31118
rect 44158 31042 44210 31054
rect 44382 31106 44434 31118
rect 44382 31042 44434 31054
rect 45502 31106 45554 31118
rect 45502 31042 45554 31054
rect 46174 31106 46226 31118
rect 72606 31106 72658 31118
rect 47058 31054 47070 31106
rect 47122 31054 47134 31106
rect 51762 31054 51774 31106
rect 51826 31054 51838 31106
rect 52546 31054 52558 31106
rect 52610 31054 52622 31106
rect 46174 31042 46226 31054
rect 72606 31042 72658 31054
rect 74174 31106 74226 31118
rect 74174 31042 74226 31054
rect 75854 31106 75906 31118
rect 75854 31042 75906 31054
rect 76414 31106 76466 31118
rect 76414 31042 76466 31054
rect 77870 31106 77922 31118
rect 77870 31042 77922 31054
rect 1710 30994 1762 31006
rect 45726 30994 45778 31006
rect 45266 30942 45278 30994
rect 45330 30942 45342 30994
rect 1710 30930 1762 30942
rect 45726 30930 45778 30942
rect 46286 30994 46338 31006
rect 72270 30994 72322 31006
rect 46834 30942 46846 30994
rect 46898 30942 46910 30994
rect 51426 30942 51438 30994
rect 51490 30942 51502 30994
rect 52434 30942 52446 30994
rect 52498 30942 52510 30994
rect 46286 30930 46338 30942
rect 72270 30930 72322 30942
rect 72718 30994 72770 31006
rect 72718 30930 72770 30942
rect 73614 30994 73666 31006
rect 73614 30930 73666 30942
rect 74286 30994 74338 31006
rect 74286 30930 74338 30942
rect 75518 30994 75570 31006
rect 75518 30930 75570 30942
rect 76078 30994 76130 31006
rect 76078 30930 76130 30942
rect 76750 30994 76802 31006
rect 76750 30930 76802 30942
rect 2494 30882 2546 30894
rect 2494 30818 2546 30830
rect 45950 30882 46002 30894
rect 72382 30882 72434 30894
rect 51986 30830 51998 30882
rect 52050 30830 52062 30882
rect 52882 30830 52894 30882
rect 52946 30830 52958 30882
rect 45950 30818 46002 30830
rect 72382 30818 72434 30830
rect 75630 30882 75682 30894
rect 75630 30818 75682 30830
rect 44494 30770 44546 30782
rect 44494 30706 44546 30718
rect 1344 30602 78624 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 65918 30602
rect 65970 30550 66022 30602
rect 66074 30550 66126 30602
rect 66178 30550 78624 30602
rect 1344 30516 78624 30550
rect 72830 30434 72882 30446
rect 72830 30370 72882 30382
rect 52894 30322 52946 30334
rect 52894 30258 52946 30270
rect 71934 30322 71986 30334
rect 74622 30322 74674 30334
rect 73602 30270 73614 30322
rect 73666 30270 73678 30322
rect 71934 30258 71986 30270
rect 74622 30258 74674 30270
rect 45726 30210 45778 30222
rect 45726 30146 45778 30158
rect 46174 30210 46226 30222
rect 46174 30146 46226 30158
rect 46286 30210 46338 30222
rect 46286 30146 46338 30158
rect 46734 30210 46786 30222
rect 46734 30146 46786 30158
rect 46958 30210 47010 30222
rect 46958 30146 47010 30158
rect 47182 30210 47234 30222
rect 72046 30210 72098 30222
rect 50866 30158 50878 30210
rect 50930 30158 50942 30210
rect 47182 30146 47234 30158
rect 72046 30146 72098 30158
rect 72494 30210 72546 30222
rect 75070 30210 75122 30222
rect 76078 30210 76130 30222
rect 72930 30158 72942 30210
rect 72994 30158 73006 30210
rect 73714 30158 73726 30210
rect 73778 30158 73790 30210
rect 75394 30158 75406 30210
rect 75458 30158 75470 30210
rect 72494 30146 72546 30158
rect 75070 30146 75122 30158
rect 76078 30146 76130 30158
rect 76638 30210 76690 30222
rect 76638 30146 76690 30158
rect 77086 30210 77138 30222
rect 77086 30146 77138 30158
rect 78206 30210 78258 30222
rect 78206 30146 78258 30158
rect 47294 30098 47346 30110
rect 51998 30098 52050 30110
rect 76526 30098 76578 30110
rect 51202 30046 51214 30098
rect 51266 30046 51278 30098
rect 71474 30046 71486 30098
rect 71538 30046 71550 30098
rect 47294 30034 47346 30046
rect 51998 30034 52050 30046
rect 76526 30034 76578 30046
rect 77422 30098 77474 30110
rect 77422 30034 77474 30046
rect 77870 30098 77922 30110
rect 77870 30034 77922 30046
rect 46062 29986 46114 29998
rect 71150 29986 71202 29998
rect 51426 29934 51438 29986
rect 51490 29934 51502 29986
rect 46062 29922 46114 29934
rect 71150 29922 71202 29934
rect 71822 29986 71874 29998
rect 71822 29922 71874 29934
rect 75630 29986 75682 29998
rect 75630 29922 75682 29934
rect 76302 29986 76354 29998
rect 76302 29922 76354 29934
rect 1344 29818 78624 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 50558 29818
rect 50610 29766 50662 29818
rect 50714 29766 50766 29818
rect 50818 29766 78624 29818
rect 1344 29732 78624 29766
rect 44942 29650 44994 29662
rect 44942 29586 44994 29598
rect 71374 29650 71426 29662
rect 71374 29586 71426 29598
rect 71822 29650 71874 29662
rect 77646 29650 77698 29662
rect 76290 29598 76302 29650
rect 76354 29598 76366 29650
rect 71822 29586 71874 29598
rect 2046 29538 2098 29550
rect 2046 29474 2098 29486
rect 44606 29538 44658 29550
rect 44606 29474 44658 29486
rect 44830 29538 44882 29550
rect 44830 29474 44882 29486
rect 73166 29538 73218 29550
rect 73166 29474 73218 29486
rect 75854 29538 75906 29550
rect 75854 29474 75906 29486
rect 76078 29538 76130 29550
rect 76078 29474 76130 29486
rect 1710 29426 1762 29438
rect 1710 29362 1762 29374
rect 72718 29426 72770 29438
rect 72718 29362 72770 29374
rect 72830 29426 72882 29438
rect 75518 29426 75570 29438
rect 73490 29374 73502 29426
rect 73554 29374 73566 29426
rect 74386 29374 74398 29426
rect 74450 29374 74462 29426
rect 74834 29374 74846 29426
rect 74898 29374 74910 29426
rect 72830 29362 72882 29374
rect 75518 29362 75570 29374
rect 75630 29426 75682 29438
rect 75630 29362 75682 29374
rect 2494 29314 2546 29326
rect 2494 29250 2546 29262
rect 70926 29314 70978 29326
rect 70926 29250 70978 29262
rect 73054 29314 73106 29326
rect 73054 29250 73106 29262
rect 74062 29202 74114 29214
rect 76305 29202 76351 29598
rect 77646 29586 77698 29598
rect 77758 29650 77810 29662
rect 77758 29586 77810 29598
rect 76638 29538 76690 29550
rect 76638 29474 76690 29486
rect 76974 29538 77026 29550
rect 76974 29474 77026 29486
rect 77086 29426 77138 29438
rect 77086 29362 77138 29374
rect 76750 29314 76802 29326
rect 76750 29250 76802 29262
rect 77534 29202 77586 29214
rect 72146 29150 72158 29202
rect 72210 29199 72222 29202
rect 72482 29199 72494 29202
rect 72210 29153 72494 29199
rect 72210 29150 72222 29153
rect 72482 29150 72494 29153
rect 72546 29150 72558 29202
rect 76290 29150 76302 29202
rect 76354 29150 76366 29202
rect 74062 29138 74114 29150
rect 77534 29138 77586 29150
rect 1344 29034 78624 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 65918 29034
rect 65970 28982 66022 29034
rect 66074 28982 66126 29034
rect 66178 28982 78624 29034
rect 1344 28948 78624 28982
rect 70802 28814 70814 28866
rect 70866 28814 70878 28866
rect 37102 28754 37154 28766
rect 73502 28754 73554 28766
rect 70578 28702 70590 28754
rect 70642 28702 70654 28754
rect 37102 28690 37154 28702
rect 73502 28690 73554 28702
rect 76302 28754 76354 28766
rect 76302 28690 76354 28702
rect 78206 28754 78258 28766
rect 78206 28690 78258 28702
rect 1710 28642 1762 28654
rect 1710 28578 1762 28590
rect 2494 28642 2546 28654
rect 72494 28642 72546 28654
rect 70354 28590 70366 28642
rect 70418 28590 70430 28642
rect 70690 28590 70702 28642
rect 70754 28590 70766 28642
rect 2494 28578 2546 28590
rect 72494 28578 72546 28590
rect 73726 28642 73778 28654
rect 73726 28578 73778 28590
rect 74398 28642 74450 28654
rect 74398 28578 74450 28590
rect 75070 28642 75122 28654
rect 75070 28578 75122 28590
rect 76078 28642 76130 28654
rect 76078 28578 76130 28590
rect 76526 28642 76578 28654
rect 76526 28578 76578 28590
rect 76974 28642 77026 28654
rect 76974 28578 77026 28590
rect 77422 28642 77474 28654
rect 77422 28578 77474 28590
rect 77646 28642 77698 28654
rect 77646 28578 77698 28590
rect 71822 28530 71874 28542
rect 2034 28478 2046 28530
rect 2098 28478 2110 28530
rect 71822 28466 71874 28478
rect 72158 28530 72210 28542
rect 72158 28466 72210 28478
rect 72830 28530 72882 28542
rect 76750 28530 76802 28542
rect 74722 28478 74734 28530
rect 74786 28478 74798 28530
rect 72830 28466 72882 28478
rect 76750 28466 76802 28478
rect 74062 28418 74114 28430
rect 77198 28418 77250 28430
rect 75394 28366 75406 28418
rect 75458 28366 75470 28418
rect 74062 28354 74114 28366
rect 77198 28354 77250 28366
rect 1344 28250 78624 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 50558 28250
rect 50610 28198 50662 28250
rect 50714 28198 50766 28250
rect 50818 28198 78624 28250
rect 1344 28164 78624 28198
rect 36990 28082 37042 28094
rect 36990 28018 37042 28030
rect 37438 28082 37490 28094
rect 39342 28082 39394 28094
rect 42478 28082 42530 28094
rect 38658 28030 38670 28082
rect 38722 28030 38734 28082
rect 41010 28030 41022 28082
rect 41074 28030 41086 28082
rect 37438 28018 37490 28030
rect 39342 28018 39394 28030
rect 42478 28018 42530 28030
rect 44718 28082 44770 28094
rect 44718 28018 44770 28030
rect 72606 28082 72658 28094
rect 72606 28018 72658 28030
rect 77646 28082 77698 28094
rect 77646 28018 77698 28030
rect 35086 27970 35138 27982
rect 45054 27970 45106 27982
rect 36418 27918 36430 27970
rect 36482 27918 36494 27970
rect 38210 27918 38222 27970
rect 38274 27918 38286 27970
rect 41570 27918 41582 27970
rect 41634 27918 41646 27970
rect 35086 27906 35138 27918
rect 45054 27906 45106 27918
rect 72830 27970 72882 27982
rect 72830 27906 72882 27918
rect 73726 27970 73778 27982
rect 73726 27906 73778 27918
rect 75182 27970 75234 27982
rect 75182 27906 75234 27918
rect 75854 27970 75906 27982
rect 75854 27906 75906 27918
rect 76414 27970 76466 27982
rect 76414 27906 76466 27918
rect 76638 27970 76690 27982
rect 76638 27906 76690 27918
rect 76750 27970 76802 27982
rect 76750 27906 76802 27918
rect 77534 27970 77586 27982
rect 77534 27906 77586 27918
rect 77758 27970 77810 27982
rect 77758 27906 77810 27918
rect 40350 27858 40402 27870
rect 70254 27858 70306 27870
rect 35522 27806 35534 27858
rect 35586 27806 35598 27858
rect 35970 27806 35982 27858
rect 36034 27806 36046 27858
rect 37762 27806 37774 27858
rect 37826 27806 37838 27858
rect 38770 27806 38782 27858
rect 38834 27806 38846 27858
rect 41010 27806 41022 27858
rect 41074 27806 41086 27858
rect 41458 27806 41470 27858
rect 41522 27806 41534 27858
rect 40350 27794 40402 27806
rect 70254 27794 70306 27806
rect 70702 27858 70754 27870
rect 70702 27794 70754 27806
rect 70926 27858 70978 27870
rect 70926 27794 70978 27806
rect 73166 27858 73218 27870
rect 73166 27794 73218 27806
rect 73390 27858 73442 27870
rect 73390 27794 73442 27806
rect 73950 27858 74002 27870
rect 73950 27794 74002 27806
rect 74286 27858 74338 27870
rect 74286 27794 74338 27806
rect 74734 27858 74786 27870
rect 74734 27794 74786 27806
rect 74958 27858 75010 27870
rect 76862 27858 76914 27870
rect 75618 27806 75630 27858
rect 75682 27806 75694 27858
rect 74958 27794 75010 27806
rect 76862 27794 76914 27806
rect 77086 27858 77138 27870
rect 77086 27794 77138 27806
rect 70142 27746 70194 27758
rect 36082 27694 36094 27746
rect 36146 27694 36158 27746
rect 70142 27682 70194 27694
rect 70814 27746 70866 27758
rect 70814 27682 70866 27694
rect 71486 27746 71538 27758
rect 71486 27682 71538 27694
rect 72942 27746 72994 27758
rect 72942 27682 72994 27694
rect 73838 27746 73890 27758
rect 73838 27682 73890 27694
rect 75070 27746 75122 27758
rect 75070 27682 75122 27694
rect 45166 27634 45218 27646
rect 45166 27570 45218 27582
rect 1344 27466 78624 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 65918 27466
rect 65970 27414 66022 27466
rect 66074 27414 66126 27466
rect 66178 27414 78624 27466
rect 1344 27380 78624 27414
rect 49646 27298 49698 27310
rect 45154 27246 45166 27298
rect 45218 27295 45230 27298
rect 46274 27295 46286 27298
rect 45218 27249 46286 27295
rect 45218 27246 45230 27249
rect 46274 27246 46286 27249
rect 46338 27246 46350 27298
rect 49646 27234 49698 27246
rect 76862 27298 76914 27310
rect 76862 27234 76914 27246
rect 77198 27298 77250 27310
rect 77198 27234 77250 27246
rect 42590 27186 42642 27198
rect 35858 27134 35870 27186
rect 35922 27134 35934 27186
rect 38546 27134 38558 27186
rect 38610 27134 38622 27186
rect 39666 27134 39678 27186
rect 39730 27134 39742 27186
rect 42590 27122 42642 27134
rect 43038 27186 43090 27198
rect 43038 27122 43090 27134
rect 44830 27186 44882 27198
rect 44830 27122 44882 27134
rect 45390 27186 45442 27198
rect 45390 27122 45442 27134
rect 45838 27186 45890 27198
rect 45838 27122 45890 27134
rect 46622 27186 46674 27198
rect 46622 27122 46674 27134
rect 50206 27186 50258 27198
rect 50206 27122 50258 27134
rect 71822 27186 71874 27198
rect 71822 27122 71874 27134
rect 72270 27186 72322 27198
rect 72270 27122 72322 27134
rect 72718 27186 72770 27198
rect 75394 27134 75406 27186
rect 75458 27134 75470 27186
rect 72718 27122 72770 27134
rect 37550 27074 37602 27086
rect 46398 27074 46450 27086
rect 33842 27022 33854 27074
rect 33906 27022 33918 27074
rect 34850 27022 34862 27074
rect 34914 27022 34926 27074
rect 35522 27022 35534 27074
rect 35586 27022 35598 27074
rect 36194 27022 36206 27074
rect 36258 27022 36270 27074
rect 38098 27022 38110 27074
rect 38162 27022 38174 27074
rect 38770 27022 38782 27074
rect 38834 27022 38846 27074
rect 39778 27022 39790 27074
rect 39842 27022 39854 27074
rect 40674 27022 40686 27074
rect 40738 27022 40750 27074
rect 41010 27022 41022 27074
rect 41074 27022 41086 27074
rect 42130 27022 42142 27074
rect 42194 27022 42206 27074
rect 37550 27010 37602 27022
rect 46398 27010 46450 27022
rect 47294 27074 47346 27086
rect 47294 27010 47346 27022
rect 47518 27074 47570 27086
rect 47518 27010 47570 27022
rect 47854 27074 47906 27086
rect 47854 27010 47906 27022
rect 48974 27074 49026 27086
rect 48974 27010 49026 27022
rect 49534 27074 49586 27086
rect 49534 27010 49586 27022
rect 70702 27074 70754 27086
rect 73166 27074 73218 27086
rect 71026 27022 71038 27074
rect 71090 27022 71102 27074
rect 70702 27010 70754 27022
rect 73166 27010 73218 27022
rect 73502 27074 73554 27086
rect 73502 27010 73554 27022
rect 74062 27074 74114 27086
rect 77870 27074 77922 27086
rect 75282 27022 75294 27074
rect 75346 27022 75358 27074
rect 76402 27022 76414 27074
rect 76466 27022 76478 27074
rect 74062 27010 74114 27022
rect 77870 27010 77922 27022
rect 1710 26962 1762 26974
rect 1710 26898 1762 26910
rect 2046 26962 2098 26974
rect 2046 26898 2098 26910
rect 2494 26962 2546 26974
rect 36990 26962 37042 26974
rect 44942 26962 44994 26974
rect 34290 26910 34302 26962
rect 34354 26910 34366 26962
rect 36418 26910 36430 26962
rect 36482 26910 36494 26962
rect 38210 26910 38222 26962
rect 38274 26910 38286 26962
rect 40002 26910 40014 26962
rect 40066 26910 40078 26962
rect 42018 26910 42030 26962
rect 42082 26910 42094 26962
rect 2494 26898 2546 26910
rect 36990 26898 37042 26910
rect 44942 26898 44994 26910
rect 46846 26962 46898 26974
rect 46846 26898 46898 26910
rect 47070 26962 47122 26974
rect 47070 26898 47122 26910
rect 47742 26962 47794 26974
rect 47742 26898 47794 26910
rect 49086 26962 49138 26974
rect 49086 26898 49138 26910
rect 49646 26962 49698 26974
rect 49646 26898 49698 26910
rect 50654 26962 50706 26974
rect 50654 26898 50706 26910
rect 70590 26962 70642 26974
rect 70590 26898 70642 26910
rect 72942 26962 72994 26974
rect 72942 26898 72994 26910
rect 74622 26962 74674 26974
rect 74622 26898 74674 26910
rect 74958 26962 75010 26974
rect 74958 26898 75010 26910
rect 75630 26962 75682 26974
rect 75630 26898 75682 26910
rect 76190 26962 76242 26974
rect 76190 26898 76242 26910
rect 77534 26962 77586 26974
rect 77534 26898 77586 26910
rect 49310 26850 49362 26862
rect 34850 26798 34862 26850
rect 34914 26798 34926 26850
rect 41122 26798 41134 26850
rect 41186 26798 41198 26850
rect 49310 26786 49362 26798
rect 70478 26850 70530 26862
rect 70478 26786 70530 26798
rect 73166 26850 73218 26862
rect 73166 26786 73218 26798
rect 76974 26850 77026 26862
rect 76974 26786 77026 26798
rect 1344 26682 78624 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 50558 26682
rect 50610 26630 50662 26682
rect 50714 26630 50766 26682
rect 50818 26630 78624 26682
rect 1344 26596 78624 26630
rect 42366 26514 42418 26526
rect 48862 26514 48914 26526
rect 36642 26462 36654 26514
rect 36706 26462 36718 26514
rect 44482 26462 44494 26514
rect 44546 26462 44558 26514
rect 42366 26450 42418 26462
rect 48862 26450 48914 26462
rect 50094 26514 50146 26526
rect 50094 26450 50146 26462
rect 50542 26514 50594 26526
rect 50542 26450 50594 26462
rect 72494 26514 72546 26526
rect 72494 26450 72546 26462
rect 76190 26514 76242 26526
rect 76190 26450 76242 26462
rect 76750 26514 76802 26526
rect 76750 26450 76802 26462
rect 77310 26514 77362 26526
rect 77310 26450 77362 26462
rect 77758 26514 77810 26526
rect 77758 26450 77810 26462
rect 2046 26402 2098 26414
rect 46846 26402 46898 26414
rect 35522 26350 35534 26402
rect 35586 26350 35598 26402
rect 37986 26350 37998 26402
rect 38050 26350 38062 26402
rect 39106 26350 39118 26402
rect 39170 26350 39182 26402
rect 42018 26350 42030 26402
rect 42082 26350 42094 26402
rect 43474 26350 43486 26402
rect 43538 26350 43550 26402
rect 46162 26350 46174 26402
rect 46226 26350 46238 26402
rect 2046 26338 2098 26350
rect 46846 26338 46898 26350
rect 47742 26402 47794 26414
rect 47742 26338 47794 26350
rect 49422 26402 49474 26414
rect 74610 26350 74622 26402
rect 74674 26350 74686 26402
rect 75506 26350 75518 26402
rect 75570 26350 75582 26402
rect 49422 26338 49474 26350
rect 1710 26290 1762 26302
rect 1710 26226 1762 26238
rect 33742 26290 33794 26302
rect 33742 26226 33794 26238
rect 34302 26290 34354 26302
rect 34302 26226 34354 26238
rect 35198 26290 35250 26302
rect 42926 26290 42978 26302
rect 45054 26290 45106 26302
rect 46398 26290 46450 26302
rect 36082 26238 36094 26290
rect 36146 26238 36158 26290
rect 37650 26238 37662 26290
rect 37714 26238 37726 26290
rect 39666 26238 39678 26290
rect 39730 26238 39742 26290
rect 40002 26238 40014 26290
rect 40066 26238 40078 26290
rect 40898 26238 40910 26290
rect 40962 26238 40974 26290
rect 41906 26238 41918 26290
rect 41970 26238 41982 26290
rect 44034 26238 44046 26290
rect 44098 26238 44110 26290
rect 44370 26238 44382 26290
rect 44434 26238 44446 26290
rect 45938 26238 45950 26290
rect 46002 26238 46014 26290
rect 35198 26226 35250 26238
rect 42926 26226 42978 26238
rect 45054 26226 45106 26238
rect 46398 26226 46450 26238
rect 46622 26290 46674 26302
rect 46622 26226 46674 26238
rect 46958 26290 47010 26302
rect 46958 26226 47010 26238
rect 47294 26290 47346 26302
rect 47294 26226 47346 26238
rect 47854 26290 47906 26302
rect 47854 26226 47906 26238
rect 48750 26290 48802 26302
rect 48750 26226 48802 26238
rect 49310 26290 49362 26302
rect 49310 26226 49362 26238
rect 49646 26290 49698 26302
rect 77534 26290 77586 26302
rect 73378 26238 73390 26290
rect 73442 26238 73454 26290
rect 74162 26238 74174 26290
rect 74226 26238 74238 26290
rect 74722 26238 74734 26290
rect 74786 26238 74798 26290
rect 75282 26238 75294 26290
rect 75346 26238 75358 26290
rect 76514 26238 76526 26290
rect 76578 26238 76590 26290
rect 49646 26226 49698 26238
rect 77534 26226 77586 26238
rect 77646 26290 77698 26302
rect 77646 26226 77698 26238
rect 2494 26178 2546 26190
rect 44942 26178 44994 26190
rect 34738 26126 34750 26178
rect 34802 26126 34814 26178
rect 39778 26126 39790 26178
rect 39842 26126 39854 26178
rect 41458 26126 41470 26178
rect 41522 26126 41534 26178
rect 2494 26114 2546 26126
rect 44942 26114 44994 26126
rect 45502 26178 45554 26190
rect 45502 26114 45554 26126
rect 47518 26178 47570 26190
rect 47518 26114 47570 26126
rect 71374 26178 71426 26190
rect 71374 26114 71426 26126
rect 71822 26178 71874 26190
rect 71822 26114 71874 26126
rect 73166 26178 73218 26190
rect 73166 26114 73218 26126
rect 48862 26066 48914 26078
rect 48862 26002 48914 26014
rect 1344 25898 78624 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 65918 25898
rect 65970 25846 66022 25898
rect 66074 25846 66126 25898
rect 66178 25846 78624 25898
rect 1344 25812 78624 25846
rect 47070 25730 47122 25742
rect 39666 25678 39678 25730
rect 39730 25727 39742 25730
rect 40114 25727 40126 25730
rect 39730 25681 40126 25727
rect 39730 25678 39742 25681
rect 40114 25678 40126 25681
rect 40178 25678 40190 25730
rect 47070 25666 47122 25678
rect 71262 25730 71314 25742
rect 74386 25678 74398 25730
rect 74450 25727 74462 25730
rect 74722 25727 74734 25730
rect 74450 25681 74734 25727
rect 74450 25678 74462 25681
rect 74722 25678 74734 25681
rect 74786 25678 74798 25730
rect 71262 25666 71314 25678
rect 40126 25618 40178 25630
rect 41918 25618 41970 25630
rect 35970 25566 35982 25618
rect 36034 25566 36046 25618
rect 40898 25566 40910 25618
rect 40962 25566 40974 25618
rect 40126 25554 40178 25566
rect 41918 25554 41970 25566
rect 44270 25618 44322 25630
rect 74734 25618 74786 25630
rect 45266 25566 45278 25618
rect 45330 25566 45342 25618
rect 72034 25566 72046 25618
rect 72098 25566 72110 25618
rect 72930 25566 72942 25618
rect 72994 25566 73006 25618
rect 73714 25566 73726 25618
rect 73778 25566 73790 25618
rect 44270 25554 44322 25566
rect 74734 25554 74786 25566
rect 37214 25506 37266 25518
rect 34962 25454 34974 25506
rect 35026 25454 35038 25506
rect 35522 25454 35534 25506
rect 35586 25454 35598 25506
rect 37214 25442 37266 25454
rect 37774 25506 37826 25518
rect 40462 25506 40514 25518
rect 38322 25454 38334 25506
rect 38386 25454 38398 25506
rect 38658 25454 38670 25506
rect 38722 25454 38734 25506
rect 37774 25442 37826 25454
rect 40462 25442 40514 25454
rect 41358 25506 41410 25518
rect 43710 25506 43762 25518
rect 46286 25506 46338 25518
rect 42802 25454 42814 25506
rect 42866 25454 42878 25506
rect 43362 25454 43374 25506
rect 43426 25454 43438 25506
rect 44930 25454 44942 25506
rect 44994 25454 45006 25506
rect 45826 25454 45838 25506
rect 45890 25454 45902 25506
rect 41358 25442 41410 25454
rect 43710 25442 43762 25454
rect 46286 25442 46338 25454
rect 70926 25506 70978 25518
rect 77422 25506 77474 25518
rect 71026 25454 71038 25506
rect 71090 25454 71102 25506
rect 71810 25454 71822 25506
rect 71874 25454 71886 25506
rect 72706 25454 72718 25506
rect 72770 25454 72782 25506
rect 73490 25454 73502 25506
rect 73554 25454 73566 25506
rect 75394 25454 75406 25506
rect 75458 25454 75470 25506
rect 70926 25442 70978 25454
rect 77422 25442 77474 25454
rect 78206 25506 78258 25518
rect 78206 25442 78258 25454
rect 46622 25394 46674 25406
rect 2034 25342 2046 25394
rect 2098 25342 2110 25394
rect 35746 25342 35758 25394
rect 35810 25342 35822 25394
rect 39106 25342 39118 25394
rect 39170 25342 39182 25394
rect 42690 25342 42702 25394
rect 42754 25342 42766 25394
rect 45490 25342 45502 25394
rect 45554 25342 45566 25394
rect 46622 25330 46674 25342
rect 46958 25394 47010 25406
rect 46958 25330 47010 25342
rect 47518 25394 47570 25406
rect 47518 25330 47570 25342
rect 70478 25394 70530 25406
rect 70478 25330 70530 25342
rect 76190 25394 76242 25406
rect 76190 25330 76242 25342
rect 76526 25394 76578 25406
rect 76526 25330 76578 25342
rect 77870 25394 77922 25406
rect 77870 25330 77922 25342
rect 1710 25282 1762 25294
rect 1710 25218 1762 25230
rect 2494 25282 2546 25294
rect 2494 25218 2546 25230
rect 34750 25282 34802 25294
rect 39678 25282 39730 25294
rect 75630 25282 75682 25294
rect 38210 25230 38222 25282
rect 38274 25230 38286 25282
rect 43250 25230 43262 25282
rect 43314 25230 43326 25282
rect 34750 25218 34802 25230
rect 39678 25218 39730 25230
rect 75630 25218 75682 25230
rect 77086 25282 77138 25294
rect 77086 25218 77138 25230
rect 1344 25114 78624 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 50558 25114
rect 50610 25062 50662 25114
rect 50714 25062 50766 25114
rect 50818 25062 78624 25114
rect 1344 25028 78624 25062
rect 25566 24946 25618 24958
rect 25566 24882 25618 24894
rect 26574 24946 26626 24958
rect 40910 24946 40962 24958
rect 44606 24946 44658 24958
rect 36866 24894 36878 24946
rect 36930 24894 36942 24946
rect 42018 24894 42030 24946
rect 42082 24894 42094 24946
rect 44034 24894 44046 24946
rect 44098 24894 44110 24946
rect 26574 24882 26626 24894
rect 40910 24882 40962 24894
rect 44606 24882 44658 24894
rect 45502 24946 45554 24958
rect 45502 24882 45554 24894
rect 46622 24946 46674 24958
rect 46622 24882 46674 24894
rect 63086 24946 63138 24958
rect 63086 24882 63138 24894
rect 63310 24946 63362 24958
rect 63310 24882 63362 24894
rect 64654 24946 64706 24958
rect 64654 24882 64706 24894
rect 71710 24946 71762 24958
rect 71710 24882 71762 24894
rect 75854 24946 75906 24958
rect 75854 24882 75906 24894
rect 76526 24946 76578 24958
rect 76526 24882 76578 24894
rect 77646 24946 77698 24958
rect 77646 24882 77698 24894
rect 17502 24834 17554 24846
rect 17502 24770 17554 24782
rect 19742 24834 19794 24846
rect 35310 24834 35362 24846
rect 20962 24782 20974 24834
rect 21026 24782 21038 24834
rect 19742 24770 19794 24782
rect 35310 24770 35362 24782
rect 35534 24834 35586 24846
rect 39342 24834 39394 24846
rect 36194 24782 36206 24834
rect 36258 24782 36270 24834
rect 37986 24782 37998 24834
rect 38050 24782 38062 24834
rect 35534 24770 35586 24782
rect 39342 24770 39394 24782
rect 40350 24834 40402 24846
rect 40350 24770 40402 24782
rect 41246 24834 41298 24846
rect 45166 24834 45218 24846
rect 75742 24834 75794 24846
rect 43026 24782 43038 24834
rect 43090 24782 43102 24834
rect 46162 24782 46174 24834
rect 46226 24782 46238 24834
rect 41246 24770 41298 24782
rect 45166 24770 45218 24782
rect 75742 24770 75794 24782
rect 77198 24834 77250 24846
rect 77198 24770 77250 24782
rect 77534 24834 77586 24846
rect 77534 24770 77586 24782
rect 17390 24722 17442 24734
rect 17390 24658 17442 24670
rect 17726 24722 17778 24734
rect 17726 24658 17778 24670
rect 19630 24722 19682 24734
rect 25118 24722 25170 24734
rect 20290 24670 20302 24722
rect 20354 24670 20366 24722
rect 19630 24658 19682 24670
rect 25118 24658 25170 24670
rect 25790 24722 25842 24734
rect 25790 24658 25842 24670
rect 26686 24722 26738 24734
rect 30270 24722 30322 24734
rect 27122 24670 27134 24722
rect 27186 24670 27198 24722
rect 26686 24658 26738 24670
rect 30270 24658 30322 24670
rect 34974 24722 35026 24734
rect 34974 24658 35026 24670
rect 35198 24722 35250 24734
rect 39678 24722 39730 24734
rect 42366 24722 42418 24734
rect 63534 24722 63586 24734
rect 35970 24670 35982 24722
rect 36034 24670 36046 24722
rect 37874 24670 37886 24722
rect 37938 24670 37950 24722
rect 40114 24670 40126 24722
rect 40178 24670 40190 24722
rect 43586 24670 43598 24722
rect 43650 24670 43662 24722
rect 44146 24670 44158 24722
rect 44210 24670 44222 24722
rect 45938 24670 45950 24722
rect 46002 24670 46014 24722
rect 72146 24670 72158 24722
rect 72210 24670 72222 24722
rect 72930 24670 72942 24722
rect 72994 24670 73006 24722
rect 73490 24670 73502 24722
rect 73554 24670 73566 24722
rect 73826 24670 73838 24722
rect 73890 24670 73902 24722
rect 74610 24670 74622 24722
rect 74674 24670 74686 24722
rect 75170 24670 75182 24722
rect 75234 24670 75246 24722
rect 76850 24670 76862 24722
rect 76914 24670 76926 24722
rect 77858 24670 77870 24722
rect 77922 24670 77934 24722
rect 35198 24658 35250 24670
rect 39678 24658 39730 24670
rect 42366 24658 42418 24670
rect 63534 24658 63586 24670
rect 18062 24610 18114 24622
rect 18062 24546 18114 24558
rect 19294 24610 19346 24622
rect 23438 24610 23490 24622
rect 25678 24610 25730 24622
rect 30382 24610 30434 24622
rect 23090 24558 23102 24610
rect 23154 24558 23166 24610
rect 23762 24558 23774 24610
rect 23826 24558 23838 24610
rect 27794 24558 27806 24610
rect 27858 24558 27870 24610
rect 29922 24558 29934 24610
rect 29986 24558 29998 24610
rect 19294 24546 19346 24558
rect 23438 24546 23490 24558
rect 25678 24546 25730 24558
rect 30382 24546 30434 24558
rect 41694 24610 41746 24622
rect 41694 24546 41746 24558
rect 47070 24610 47122 24622
rect 47070 24546 47122 24558
rect 63422 24610 63474 24622
rect 63422 24546 63474 24558
rect 71374 24610 71426 24622
rect 74050 24558 74062 24610
rect 74114 24558 74126 24610
rect 71374 24546 71426 24558
rect 19742 24498 19794 24510
rect 19742 24434 19794 24446
rect 72382 24498 72434 24510
rect 72382 24434 72434 24446
rect 75966 24498 76018 24510
rect 75966 24434 76018 24446
rect 76862 24498 76914 24510
rect 76862 24434 76914 24446
rect 1344 24330 78624 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 65918 24330
rect 65970 24278 66022 24330
rect 66074 24278 66126 24330
rect 66178 24278 78624 24330
rect 1344 24244 78624 24278
rect 77534 24162 77586 24174
rect 42578 24110 42590 24162
rect 42642 24159 42654 24162
rect 43362 24159 43374 24162
rect 42642 24113 43374 24159
rect 42642 24110 42654 24113
rect 43362 24110 43374 24113
rect 43426 24110 43438 24162
rect 74050 24110 74062 24162
rect 74114 24110 74126 24162
rect 77534 24098 77586 24110
rect 19966 24050 20018 24062
rect 19618 23998 19630 24050
rect 19682 23998 19694 24050
rect 19966 23986 20018 23998
rect 21422 24050 21474 24062
rect 21422 23986 21474 23998
rect 23102 24050 23154 24062
rect 27918 24050 27970 24062
rect 24770 23998 24782 24050
rect 24834 23998 24846 24050
rect 26898 23998 26910 24050
rect 26962 23998 26974 24050
rect 23102 23986 23154 23998
rect 27918 23986 27970 23998
rect 34078 24050 34130 24062
rect 34078 23986 34130 23998
rect 41806 24050 41858 24062
rect 41806 23986 41858 23998
rect 44942 24050 44994 24062
rect 44942 23986 44994 23998
rect 48078 24050 48130 24062
rect 48078 23986 48130 23998
rect 62862 24050 62914 24062
rect 62862 23986 62914 23998
rect 63534 24050 63586 24062
rect 63534 23986 63586 23998
rect 64094 24050 64146 24062
rect 64094 23986 64146 23998
rect 73166 24050 73218 24062
rect 73166 23986 73218 23998
rect 74510 24050 74562 24062
rect 75282 23998 75294 24050
rect 75346 23998 75358 24050
rect 76402 23998 76414 24050
rect 76466 23998 76478 24050
rect 74510 23986 74562 23998
rect 34526 23938 34578 23950
rect 16818 23886 16830 23938
rect 16882 23886 16894 23938
rect 21858 23886 21870 23938
rect 21922 23886 21934 23938
rect 23986 23886 23998 23938
rect 24050 23886 24062 23938
rect 34526 23874 34578 23886
rect 35646 23938 35698 23950
rect 35646 23874 35698 23886
rect 35982 23938 36034 23950
rect 35982 23874 36034 23886
rect 37662 23938 37714 23950
rect 45726 23938 45778 23950
rect 38434 23886 38446 23938
rect 38498 23886 38510 23938
rect 40338 23886 40350 23938
rect 40402 23886 40414 23938
rect 37662 23874 37714 23886
rect 45726 23874 45778 23886
rect 46062 23938 46114 23950
rect 46062 23874 46114 23886
rect 46734 23938 46786 23950
rect 46734 23874 46786 23886
rect 48526 23938 48578 23950
rect 48526 23874 48578 23886
rect 62974 23938 63026 23950
rect 62974 23874 63026 23886
rect 63422 23938 63474 23950
rect 63422 23874 63474 23886
rect 72158 23938 72210 23950
rect 72158 23874 72210 23886
rect 72718 23938 72770 23950
rect 73266 23886 73278 23938
rect 73330 23886 73342 23938
rect 74386 23886 74398 23938
rect 74450 23886 74462 23938
rect 77074 23886 77086 23938
rect 77138 23886 77150 23938
rect 72718 23874 72770 23886
rect 23550 23826 23602 23838
rect 2034 23774 2046 23826
rect 2098 23774 2110 23826
rect 17490 23774 17502 23826
rect 17554 23774 17566 23826
rect 20290 23774 20302 23826
rect 20354 23774 20366 23826
rect 23550 23762 23602 23774
rect 23662 23826 23714 23838
rect 23662 23762 23714 23774
rect 27806 23826 27858 23838
rect 27806 23762 27858 23774
rect 35758 23826 35810 23838
rect 35758 23762 35810 23774
rect 36206 23826 36258 23838
rect 36206 23762 36258 23774
rect 36318 23826 36370 23838
rect 36318 23762 36370 23774
rect 37102 23826 37154 23838
rect 37102 23762 37154 23774
rect 37214 23826 37266 23838
rect 37214 23762 37266 23774
rect 37774 23826 37826 23838
rect 37774 23762 37826 23774
rect 37998 23826 38050 23838
rect 46398 23826 46450 23838
rect 38546 23774 38558 23826
rect 38610 23774 38622 23826
rect 40450 23774 40462 23826
rect 40514 23774 40526 23826
rect 37998 23762 38050 23774
rect 46398 23762 46450 23774
rect 47406 23826 47458 23838
rect 47406 23762 47458 23774
rect 47518 23826 47570 23838
rect 47518 23762 47570 23774
rect 75630 23826 75682 23838
rect 75630 23762 75682 23774
rect 76190 23826 76242 23838
rect 76190 23762 76242 23774
rect 77758 23826 77810 23838
rect 77758 23762 77810 23774
rect 1710 23714 1762 23726
rect 1710 23650 1762 23662
rect 2494 23714 2546 23726
rect 2494 23650 2546 23662
rect 21310 23714 21362 23726
rect 21310 23650 21362 23662
rect 21534 23714 21586 23726
rect 21534 23650 21586 23662
rect 22318 23714 22370 23726
rect 22318 23650 22370 23662
rect 23326 23714 23378 23726
rect 23326 23650 23378 23662
rect 27582 23714 27634 23726
rect 27582 23650 27634 23662
rect 28030 23714 28082 23726
rect 28030 23650 28082 23662
rect 34862 23714 34914 23726
rect 34862 23650 34914 23662
rect 35422 23714 35474 23726
rect 35422 23650 35474 23662
rect 36542 23714 36594 23726
rect 36542 23650 36594 23662
rect 37438 23714 37490 23726
rect 42366 23714 42418 23726
rect 40226 23662 40238 23714
rect 40290 23662 40302 23714
rect 37438 23650 37490 23662
rect 42366 23650 42418 23662
rect 42814 23714 42866 23726
rect 42814 23650 42866 23662
rect 43262 23714 43314 23726
rect 43262 23650 43314 23662
rect 44270 23714 44322 23726
rect 44270 23650 44322 23662
rect 45390 23714 45442 23726
rect 45390 23650 45442 23662
rect 46062 23714 46114 23726
rect 46062 23650 46114 23662
rect 47070 23714 47122 23726
rect 47070 23650 47122 23662
rect 47742 23714 47794 23726
rect 47742 23650 47794 23662
rect 48974 23714 49026 23726
rect 48974 23650 49026 23662
rect 49534 23714 49586 23726
rect 49534 23650 49586 23662
rect 63646 23714 63698 23726
rect 63646 23650 63698 23662
rect 75406 23714 75458 23726
rect 75406 23650 75458 23662
rect 76414 23714 76466 23726
rect 76414 23650 76466 23662
rect 76862 23714 76914 23726
rect 76862 23650 76914 23662
rect 77646 23714 77698 23726
rect 77646 23650 77698 23662
rect 1344 23546 78624 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 50558 23546
rect 50610 23494 50662 23546
rect 50714 23494 50766 23546
rect 50818 23494 78624 23546
rect 1344 23460 78624 23494
rect 17502 23378 17554 23390
rect 17502 23314 17554 23326
rect 17614 23378 17666 23390
rect 17614 23314 17666 23326
rect 17838 23378 17890 23390
rect 17838 23314 17890 23326
rect 18398 23378 18450 23390
rect 21870 23378 21922 23390
rect 19282 23326 19294 23378
rect 19346 23326 19358 23378
rect 18398 23314 18450 23326
rect 21870 23314 21922 23326
rect 24670 23378 24722 23390
rect 28030 23378 28082 23390
rect 45166 23378 45218 23390
rect 26114 23326 26126 23378
rect 26178 23326 26190 23378
rect 38210 23326 38222 23378
rect 38274 23326 38286 23378
rect 24670 23314 24722 23326
rect 28030 23314 28082 23326
rect 45166 23314 45218 23326
rect 46286 23378 46338 23390
rect 46286 23314 46338 23326
rect 46846 23378 46898 23390
rect 46846 23314 46898 23326
rect 47406 23378 47458 23390
rect 47406 23314 47458 23326
rect 48974 23378 49026 23390
rect 48974 23314 49026 23326
rect 50318 23378 50370 23390
rect 50318 23314 50370 23326
rect 50766 23378 50818 23390
rect 50766 23314 50818 23326
rect 71710 23378 71762 23390
rect 71710 23314 71762 23326
rect 75742 23378 75794 23390
rect 75742 23314 75794 23326
rect 76526 23378 76578 23390
rect 76526 23314 76578 23326
rect 77646 23378 77698 23390
rect 77646 23314 77698 23326
rect 19966 23266 20018 23278
rect 2034 23214 2046 23266
rect 2098 23214 2110 23266
rect 19966 23202 20018 23214
rect 20078 23266 20130 23278
rect 20078 23202 20130 23214
rect 24334 23266 24386 23278
rect 24334 23202 24386 23214
rect 24446 23266 24498 23278
rect 24446 23202 24498 23214
rect 25230 23266 25282 23278
rect 25230 23202 25282 23214
rect 25342 23266 25394 23278
rect 45054 23266 45106 23278
rect 36418 23214 36430 23266
rect 36482 23214 36494 23266
rect 37538 23214 37550 23266
rect 37602 23214 37614 23266
rect 39666 23214 39678 23266
rect 39730 23214 39742 23266
rect 41682 23214 41694 23266
rect 41746 23214 41758 23266
rect 25342 23202 25394 23214
rect 45054 23202 45106 23214
rect 46734 23266 46786 23278
rect 46734 23202 46786 23214
rect 47966 23266 48018 23278
rect 47966 23202 48018 23214
rect 49422 23266 49474 23278
rect 49422 23202 49474 23214
rect 75630 23266 75682 23278
rect 75630 23202 75682 23214
rect 76750 23266 76802 23278
rect 76750 23202 76802 23214
rect 77086 23266 77138 23278
rect 77086 23202 77138 23214
rect 77534 23266 77586 23278
rect 77534 23202 77586 23214
rect 1710 23154 1762 23166
rect 1710 23090 1762 23102
rect 17390 23154 17442 23166
rect 20302 23154 20354 23166
rect 19506 23102 19518 23154
rect 19570 23102 19582 23154
rect 17390 23090 17442 23102
rect 20302 23090 20354 23102
rect 21198 23154 21250 23166
rect 21198 23090 21250 23102
rect 21646 23154 21698 23166
rect 21646 23090 21698 23102
rect 23550 23154 23602 23166
rect 23550 23090 23602 23102
rect 25566 23154 25618 23166
rect 27358 23154 27410 23166
rect 25890 23102 25902 23154
rect 25954 23102 25966 23154
rect 25566 23090 25618 23102
rect 27358 23090 27410 23102
rect 27806 23154 27858 23166
rect 31614 23154 31666 23166
rect 28354 23102 28366 23154
rect 28418 23102 28430 23154
rect 27806 23090 27858 23102
rect 31614 23090 31666 23102
rect 31726 23154 31778 23166
rect 45950 23154 46002 23166
rect 34066 23102 34078 23154
rect 34130 23102 34142 23154
rect 34962 23102 34974 23154
rect 35026 23102 35038 23154
rect 36530 23102 36542 23154
rect 36594 23102 36606 23154
rect 37314 23102 37326 23154
rect 37378 23102 37390 23154
rect 39218 23102 39230 23154
rect 39282 23102 39294 23154
rect 41010 23102 41022 23154
rect 41074 23102 41086 23154
rect 44258 23102 44270 23154
rect 44322 23102 44334 23154
rect 31726 23090 31778 23102
rect 45950 23090 46002 23102
rect 46174 23154 46226 23166
rect 46174 23090 46226 23102
rect 46510 23154 46562 23166
rect 46510 23090 46562 23102
rect 47294 23154 47346 23166
rect 47294 23090 47346 23102
rect 47854 23154 47906 23166
rect 72146 23102 72158 23154
rect 72210 23102 72222 23154
rect 72930 23102 72942 23154
rect 72994 23102 73006 23154
rect 73938 23102 73950 23154
rect 74002 23102 74014 23154
rect 74946 23102 74958 23154
rect 75010 23102 75022 23154
rect 75954 23102 75966 23154
rect 76018 23102 76030 23154
rect 77858 23102 77870 23154
rect 77922 23102 77934 23154
rect 47854 23090 47906 23102
rect 2494 23042 2546 23054
rect 2494 22978 2546 22990
rect 20638 23042 20690 23054
rect 21758 23042 21810 23054
rect 21186 22990 21198 23042
rect 21250 22990 21262 23042
rect 20638 22978 20690 22990
rect 20402 22878 20414 22930
rect 20466 22927 20478 22930
rect 21201 22927 21247 22990
rect 21758 22978 21810 22990
rect 23998 23042 24050 23054
rect 23998 22978 24050 22990
rect 27918 23042 27970 23054
rect 33854 23042 33906 23054
rect 44718 23042 44770 23054
rect 29138 22990 29150 23042
rect 29202 22990 29214 23042
rect 31266 22990 31278 23042
rect 31330 22990 31342 23042
rect 43810 22990 43822 23042
rect 43874 22990 43886 23042
rect 27918 22978 27970 22990
rect 33854 22978 33906 22990
rect 44718 22978 44770 22990
rect 49758 23042 49810 23054
rect 72370 22990 72382 23042
rect 72434 22990 72446 23042
rect 73266 22990 73278 23042
rect 73330 22990 73342 23042
rect 74722 22990 74734 23042
rect 74786 22990 74798 23042
rect 49758 22978 49810 22990
rect 20466 22881 21247 22927
rect 46846 22930 46898 22942
rect 20466 22878 20478 22881
rect 46846 22866 46898 22878
rect 47406 22930 47458 22942
rect 47406 22866 47458 22878
rect 47966 22930 48018 22942
rect 74062 22930 74114 22942
rect 49858 22878 49870 22930
rect 49922 22927 49934 22930
rect 50194 22927 50206 22930
rect 49922 22881 50206 22927
rect 49922 22878 49934 22881
rect 50194 22878 50206 22881
rect 50258 22878 50270 22930
rect 47966 22866 48018 22878
rect 74062 22866 74114 22878
rect 1344 22762 78624 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 65918 22762
rect 65970 22710 66022 22762
rect 66074 22710 66126 22762
rect 66178 22710 78624 22762
rect 1344 22676 78624 22710
rect 35758 22594 35810 22606
rect 35758 22530 35810 22542
rect 46734 22594 46786 22606
rect 46734 22530 46786 22542
rect 74286 22594 74338 22606
rect 74286 22530 74338 22542
rect 76862 22594 76914 22606
rect 76862 22530 76914 22542
rect 77198 22594 77250 22606
rect 77198 22530 77250 22542
rect 77534 22594 77586 22606
rect 77534 22530 77586 22542
rect 15598 22482 15650 22494
rect 19742 22482 19794 22494
rect 24558 22482 24610 22494
rect 29150 22482 29202 22494
rect 19394 22430 19406 22482
rect 19458 22430 19470 22482
rect 20066 22430 20078 22482
rect 20130 22430 20142 22482
rect 22082 22430 22094 22482
rect 22146 22430 22158 22482
rect 24210 22430 24222 22482
rect 24274 22430 24286 22482
rect 28354 22430 28366 22482
rect 28418 22430 28430 22482
rect 15598 22418 15650 22430
rect 19742 22418 19794 22430
rect 24558 22418 24610 22430
rect 29150 22418 29202 22430
rect 34414 22482 34466 22494
rect 46286 22482 46338 22494
rect 37314 22430 37326 22482
rect 37378 22430 37390 22482
rect 42130 22430 42142 22482
rect 42194 22430 42206 22482
rect 34414 22418 34466 22430
rect 46286 22418 46338 22430
rect 51774 22482 51826 22494
rect 51774 22418 51826 22430
rect 52782 22482 52834 22494
rect 52782 22418 52834 22430
rect 71934 22482 71986 22494
rect 77646 22482 77698 22494
rect 72258 22430 72270 22482
rect 72322 22430 72334 22482
rect 71934 22418 71986 22430
rect 77646 22418 77698 22430
rect 16158 22370 16210 22382
rect 43374 22370 43426 22382
rect 16594 22318 16606 22370
rect 16658 22318 16670 22370
rect 21298 22318 21310 22370
rect 21362 22318 21374 22370
rect 25554 22318 25566 22370
rect 25618 22318 25630 22370
rect 38322 22318 38334 22370
rect 38386 22318 38398 22370
rect 40338 22318 40350 22370
rect 40402 22318 40414 22370
rect 42466 22318 42478 22370
rect 42530 22318 42542 22370
rect 16158 22306 16210 22318
rect 43374 22306 43426 22318
rect 45166 22370 45218 22382
rect 45166 22306 45218 22318
rect 45950 22370 46002 22382
rect 45950 22306 46002 22318
rect 46174 22370 46226 22382
rect 46174 22306 46226 22318
rect 47182 22370 47234 22382
rect 47182 22306 47234 22318
rect 48078 22370 48130 22382
rect 48078 22306 48130 22318
rect 48638 22370 48690 22382
rect 51326 22370 51378 22382
rect 76190 22370 76242 22382
rect 48962 22318 48974 22370
rect 49026 22318 49038 22370
rect 50082 22318 50094 22370
rect 50146 22318 50158 22370
rect 50866 22318 50878 22370
rect 50930 22318 50942 22370
rect 72034 22318 72046 22370
rect 72098 22318 72110 22370
rect 72818 22318 72830 22370
rect 72882 22318 72894 22370
rect 73378 22318 73390 22370
rect 73442 22318 73454 22370
rect 74050 22318 74062 22370
rect 74114 22318 74126 22370
rect 74834 22318 74846 22370
rect 74898 22318 74910 22370
rect 75394 22318 75406 22370
rect 75458 22318 75470 22370
rect 48638 22306 48690 22318
rect 51326 22306 51378 22318
rect 76190 22306 76242 22318
rect 16046 22258 16098 22270
rect 35198 22258 35250 22270
rect 17266 22206 17278 22258
rect 17330 22206 17342 22258
rect 20402 22206 20414 22258
rect 20466 22206 20478 22258
rect 26226 22206 26238 22258
rect 26290 22206 26302 22258
rect 16046 22194 16098 22206
rect 35198 22194 35250 22206
rect 35310 22258 35362 22270
rect 35310 22194 35362 22206
rect 35870 22258 35922 22270
rect 35870 22194 35922 22206
rect 36206 22258 36258 22270
rect 36206 22194 36258 22206
rect 36318 22258 36370 22270
rect 43710 22258 43762 22270
rect 38434 22206 38446 22258
rect 38498 22206 38510 22258
rect 40450 22206 40462 22258
rect 40514 22206 40526 22258
rect 42354 22206 42366 22258
rect 42418 22206 42430 22258
rect 36318 22194 36370 22206
rect 43710 22194 43762 22206
rect 43822 22258 43874 22270
rect 43822 22194 43874 22206
rect 46398 22258 46450 22270
rect 46398 22194 46450 22206
rect 46846 22258 46898 22270
rect 76526 22258 76578 22270
rect 49858 22206 49870 22258
rect 49922 22206 49934 22258
rect 46846 22194 46898 22206
rect 76526 22194 76578 22206
rect 15822 22146 15874 22158
rect 15822 22082 15874 22094
rect 20750 22146 20802 22158
rect 20750 22082 20802 22094
rect 24670 22146 24722 22158
rect 24670 22082 24722 22094
rect 29262 22146 29314 22158
rect 29262 22082 29314 22094
rect 33966 22146 34018 22158
rect 33966 22082 34018 22094
rect 34750 22146 34802 22158
rect 34750 22082 34802 22094
rect 34974 22146 35026 22158
rect 34974 22082 35026 22094
rect 35758 22146 35810 22158
rect 35758 22082 35810 22094
rect 36542 22146 36594 22158
rect 36542 22082 36594 22094
rect 37774 22146 37826 22158
rect 44046 22146 44098 22158
rect 40002 22094 40014 22146
rect 40066 22094 40078 22146
rect 43026 22094 43038 22146
rect 43090 22094 43102 22146
rect 37774 22082 37826 22094
rect 44046 22082 44098 22094
rect 45502 22146 45554 22158
rect 45502 22082 45554 22094
rect 47742 22146 47794 22158
rect 76974 22146 77026 22158
rect 49074 22094 49086 22146
rect 49138 22094 49150 22146
rect 47742 22082 47794 22094
rect 76974 22082 77026 22094
rect 77758 22146 77810 22158
rect 77758 22082 77810 22094
rect 1344 21978 78624 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 50558 21978
rect 50610 21926 50662 21978
rect 50714 21926 50766 21978
rect 50818 21926 78624 21978
rect 1344 21892 78624 21926
rect 17502 21810 17554 21822
rect 17502 21746 17554 21758
rect 17726 21810 17778 21822
rect 17726 21746 17778 21758
rect 17838 21810 17890 21822
rect 17838 21746 17890 21758
rect 17950 21810 18002 21822
rect 17950 21746 18002 21758
rect 18510 21810 18562 21822
rect 26462 21810 26514 21822
rect 23874 21758 23886 21810
rect 23938 21758 23950 21810
rect 18510 21746 18562 21758
rect 26462 21746 26514 21758
rect 26574 21810 26626 21822
rect 48078 21810 48130 21822
rect 39218 21758 39230 21810
rect 39282 21758 39294 21810
rect 45714 21758 45726 21810
rect 45778 21758 45790 21810
rect 26574 21746 26626 21758
rect 48078 21746 48130 21758
rect 53790 21810 53842 21822
rect 55918 21810 55970 21822
rect 55346 21758 55358 21810
rect 55410 21758 55422 21810
rect 53790 21746 53842 21758
rect 55918 21746 55970 21758
rect 25230 21698 25282 21710
rect 2034 21646 2046 21698
rect 2098 21646 2110 21698
rect 25230 21634 25282 21646
rect 25342 21698 25394 21710
rect 25342 21634 25394 21646
rect 35198 21698 35250 21710
rect 36878 21698 36930 21710
rect 43262 21698 43314 21710
rect 47182 21698 47234 21710
rect 35970 21646 35982 21698
rect 36034 21646 36046 21698
rect 39890 21646 39902 21698
rect 39954 21646 39966 21698
rect 44258 21646 44270 21698
rect 44322 21646 44334 21698
rect 46386 21646 46398 21698
rect 46450 21646 46462 21698
rect 35198 21634 35250 21646
rect 36878 21634 36930 21646
rect 43262 21634 43314 21646
rect 47182 21634 47234 21646
rect 47406 21698 47458 21710
rect 47406 21634 47458 21646
rect 47630 21698 47682 21710
rect 47630 21634 47682 21646
rect 48190 21698 48242 21710
rect 71710 21698 71762 21710
rect 76078 21698 76130 21710
rect 49858 21646 49870 21698
rect 49922 21646 49934 21698
rect 51314 21646 51326 21698
rect 51378 21646 51390 21698
rect 54338 21646 54350 21698
rect 54402 21646 54414 21698
rect 73938 21646 73950 21698
rect 74002 21646 74014 21698
rect 48190 21634 48242 21646
rect 71710 21634 71762 21646
rect 76078 21634 76130 21646
rect 76638 21698 76690 21710
rect 76638 21634 76690 21646
rect 76974 21698 77026 21710
rect 76974 21634 77026 21646
rect 77534 21698 77586 21710
rect 77534 21634 77586 21646
rect 77758 21698 77810 21710
rect 77758 21634 77810 21646
rect 1710 21586 1762 21598
rect 24222 21586 24274 21598
rect 18834 21534 18846 21586
rect 18898 21534 18910 21586
rect 1710 21522 1762 21534
rect 24222 21522 24274 21534
rect 25566 21586 25618 21598
rect 25566 21522 25618 21534
rect 25902 21586 25954 21598
rect 25902 21522 25954 21534
rect 26350 21586 26402 21598
rect 32398 21586 32450 21598
rect 29138 21534 29150 21586
rect 29202 21534 29214 21586
rect 26350 21522 26402 21534
rect 32398 21522 32450 21534
rect 34974 21586 35026 21598
rect 34974 21522 35026 21534
rect 35422 21586 35474 21598
rect 35422 21522 35474 21534
rect 35646 21586 35698 21598
rect 35646 21522 35698 21534
rect 36318 21586 36370 21598
rect 41358 21586 41410 21598
rect 37650 21534 37662 21586
rect 37714 21534 37726 21586
rect 38546 21534 38558 21586
rect 38610 21534 38622 21586
rect 39106 21534 39118 21586
rect 39170 21534 39182 21586
rect 36318 21522 36370 21534
rect 41358 21522 41410 21534
rect 42478 21586 42530 21598
rect 47854 21586 47906 21598
rect 50206 21586 50258 21598
rect 52782 21586 52834 21598
rect 44146 21534 44158 21586
rect 44210 21534 44222 21586
rect 45602 21534 45614 21586
rect 45666 21534 45678 21586
rect 48962 21534 48974 21586
rect 49026 21534 49038 21586
rect 49522 21534 49534 21586
rect 49586 21534 49598 21586
rect 51874 21534 51886 21586
rect 51938 21534 51950 21586
rect 52434 21534 52446 21586
rect 52498 21534 52510 21586
rect 42478 21522 42530 21534
rect 47854 21522 47906 21534
rect 50206 21522 50258 21534
rect 52782 21522 52834 21534
rect 53342 21586 53394 21598
rect 75742 21586 75794 21598
rect 54898 21534 54910 21586
rect 54962 21534 54974 21586
rect 55458 21534 55470 21586
rect 55522 21534 55534 21586
rect 72146 21534 72158 21586
rect 72210 21534 72222 21586
rect 72930 21534 72942 21586
rect 72994 21534 73006 21586
rect 73490 21534 73502 21586
rect 73554 21534 73566 21586
rect 74274 21534 74286 21586
rect 74338 21534 74350 21586
rect 74946 21534 74958 21586
rect 75010 21534 75022 21586
rect 53342 21522 53394 21534
rect 75742 21522 75794 21534
rect 2494 21474 2546 21486
rect 24670 21474 24722 21486
rect 34862 21474 34914 21486
rect 19618 21422 19630 21474
rect 19682 21422 19694 21474
rect 21746 21422 21758 21474
rect 21810 21422 21822 21474
rect 29922 21422 29934 21474
rect 29986 21422 29998 21474
rect 32050 21422 32062 21474
rect 32114 21422 32126 21474
rect 2494 21410 2546 21422
rect 24670 21410 24722 21422
rect 34862 21410 34914 21422
rect 41022 21474 41074 21486
rect 49186 21422 49198 21474
rect 49250 21422 49262 21474
rect 50642 21422 50654 21474
rect 50706 21422 50718 21474
rect 51986 21422 51998 21474
rect 52050 21422 52062 21474
rect 74610 21422 74622 21474
rect 74674 21422 74686 21474
rect 77858 21422 77870 21474
rect 77922 21422 77934 21474
rect 41022 21410 41074 21422
rect 32510 21362 32562 21374
rect 32510 21298 32562 21310
rect 42142 21362 42194 21374
rect 42142 21298 42194 21310
rect 72382 21362 72434 21374
rect 72382 21298 72434 21310
rect 1344 21194 78624 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 65918 21194
rect 65970 21142 66022 21194
rect 66074 21142 66126 21194
rect 66178 21142 78624 21194
rect 1344 21108 78624 21142
rect 38782 21026 38834 21038
rect 32498 20974 32510 21026
rect 32562 21023 32574 21026
rect 32946 21023 32958 21026
rect 32562 20977 32958 21023
rect 32562 20974 32574 20977
rect 32946 20974 32958 20977
rect 33010 20974 33022 21026
rect 38782 20962 38834 20974
rect 75294 21026 75346 21038
rect 75294 20962 75346 20974
rect 76526 21026 76578 21038
rect 76526 20962 76578 20974
rect 76862 21026 76914 21038
rect 76862 20962 76914 20974
rect 77198 21026 77250 21038
rect 77198 20962 77250 20974
rect 19518 20914 19570 20926
rect 19518 20850 19570 20862
rect 29822 20914 29874 20926
rect 29822 20850 29874 20862
rect 33182 20914 33234 20926
rect 33182 20850 33234 20862
rect 35310 20914 35362 20926
rect 35310 20850 35362 20862
rect 37214 20914 37266 20926
rect 37214 20850 37266 20862
rect 51886 20914 51938 20926
rect 56926 20914 56978 20926
rect 54114 20862 54126 20914
rect 54178 20862 54190 20914
rect 55010 20862 55022 20914
rect 55074 20862 55086 20914
rect 51886 20850 51938 20862
rect 56926 20850 56978 20862
rect 71262 20914 71314 20926
rect 71262 20850 71314 20862
rect 74286 20914 74338 20926
rect 74286 20850 74338 20862
rect 75070 20914 75122 20926
rect 75070 20850 75122 20862
rect 77310 20914 77362 20926
rect 77310 20850 77362 20862
rect 20078 20802 20130 20814
rect 20078 20738 20130 20750
rect 26574 20802 26626 20814
rect 26574 20738 26626 20750
rect 35086 20802 35138 20814
rect 35086 20738 35138 20750
rect 35534 20802 35586 20814
rect 35534 20738 35586 20750
rect 35646 20802 35698 20814
rect 35646 20738 35698 20750
rect 36430 20802 36482 20814
rect 36430 20738 36482 20750
rect 38110 20802 38162 20814
rect 45054 20802 45106 20814
rect 56478 20802 56530 20814
rect 78206 20802 78258 20814
rect 39442 20750 39454 20802
rect 39506 20750 39518 20802
rect 40114 20750 40126 20802
rect 40178 20750 40190 20802
rect 41234 20750 41246 20802
rect 41298 20750 41310 20802
rect 43138 20750 43150 20802
rect 43202 20750 43214 20802
rect 45490 20750 45502 20802
rect 45554 20750 45566 20802
rect 45938 20750 45950 20802
rect 46002 20750 46014 20802
rect 47058 20750 47070 20802
rect 47122 20750 47134 20802
rect 47618 20750 47630 20802
rect 47682 20750 47694 20802
rect 48402 20750 48414 20802
rect 48466 20750 48478 20802
rect 48962 20750 48974 20802
rect 49026 20750 49038 20802
rect 49522 20750 49534 20802
rect 49586 20750 49598 20802
rect 50306 20750 50318 20802
rect 50370 20750 50382 20802
rect 51426 20750 51438 20802
rect 51490 20750 51502 20802
rect 53554 20750 53566 20802
rect 53618 20750 53630 20802
rect 54002 20750 54014 20802
rect 54066 20750 54078 20802
rect 55122 20750 55134 20802
rect 55186 20750 55198 20802
rect 55794 20750 55806 20802
rect 55858 20750 55870 20802
rect 71362 20750 71374 20802
rect 71426 20750 71438 20802
rect 72482 20750 72494 20802
rect 72546 20750 72558 20802
rect 72706 20750 72718 20802
rect 72770 20750 72782 20802
rect 73042 20750 73054 20802
rect 73106 20750 73118 20802
rect 73938 20750 73950 20802
rect 74002 20750 74014 20802
rect 75282 20750 75294 20802
rect 75346 20750 75358 20802
rect 77522 20750 77534 20802
rect 77586 20750 77598 20802
rect 38110 20738 38162 20750
rect 45054 20738 45106 20750
rect 56478 20738 56530 20750
rect 78206 20738 78258 20750
rect 24446 20690 24498 20702
rect 25230 20690 25282 20702
rect 2034 20638 2046 20690
rect 2098 20638 2110 20690
rect 24770 20638 24782 20690
rect 24834 20638 24846 20690
rect 24446 20626 24498 20638
rect 25230 20626 25282 20638
rect 25790 20690 25842 20702
rect 34302 20690 34354 20702
rect 33506 20638 33518 20690
rect 33570 20638 33582 20690
rect 25790 20626 25842 20638
rect 34302 20626 34354 20638
rect 34638 20690 34690 20702
rect 34638 20626 34690 20638
rect 34862 20690 34914 20702
rect 34862 20626 34914 20638
rect 36094 20690 36146 20702
rect 75630 20690 75682 20702
rect 41122 20638 41134 20690
rect 41186 20638 41198 20690
rect 42914 20638 42926 20690
rect 42978 20638 42990 20690
rect 46386 20638 46398 20690
rect 46450 20638 46462 20690
rect 48514 20638 48526 20690
rect 48578 20638 48590 20690
rect 49970 20638 49982 20690
rect 50034 20638 50046 20690
rect 50978 20638 50990 20690
rect 51042 20638 51054 20690
rect 54338 20638 54350 20690
rect 54402 20638 54414 20690
rect 55010 20638 55022 20690
rect 55074 20638 55086 20690
rect 72258 20638 72270 20690
rect 72322 20638 72334 20690
rect 74050 20638 74062 20690
rect 74114 20638 74126 20690
rect 36094 20626 36146 20638
rect 75630 20626 75682 20638
rect 77870 20690 77922 20702
rect 77870 20626 77922 20638
rect 1710 20578 1762 20590
rect 1710 20514 1762 20526
rect 2494 20578 2546 20590
rect 2494 20514 2546 20526
rect 19406 20578 19458 20590
rect 19406 20514 19458 20526
rect 19630 20578 19682 20590
rect 19630 20514 19682 20526
rect 20526 20578 20578 20590
rect 20526 20514 20578 20526
rect 22990 20578 23042 20590
rect 22990 20514 23042 20526
rect 23662 20578 23714 20590
rect 23662 20514 23714 20526
rect 24110 20578 24162 20590
rect 24110 20514 24162 20526
rect 25342 20578 25394 20590
rect 25342 20514 25394 20526
rect 25566 20578 25618 20590
rect 25566 20514 25618 20526
rect 25902 20578 25954 20590
rect 25902 20514 25954 20526
rect 26126 20578 26178 20590
rect 29486 20578 29538 20590
rect 26898 20526 26910 20578
rect 26962 20526 26974 20578
rect 26126 20514 26178 20526
rect 29486 20514 29538 20526
rect 29710 20578 29762 20590
rect 29710 20514 29762 20526
rect 29934 20578 29986 20590
rect 29934 20514 29986 20526
rect 30494 20578 30546 20590
rect 30494 20514 30546 20526
rect 32398 20578 32450 20590
rect 32398 20514 32450 20526
rect 32958 20578 33010 20590
rect 32958 20514 33010 20526
rect 34078 20578 34130 20590
rect 34078 20514 34130 20526
rect 34526 20578 34578 20590
rect 34526 20514 34578 20526
rect 37438 20578 37490 20590
rect 38446 20578 38498 20590
rect 37762 20526 37774 20578
rect 37826 20526 37838 20578
rect 37438 20514 37490 20526
rect 38446 20514 38498 20526
rect 39902 20578 39954 20590
rect 39902 20514 39954 20526
rect 40686 20578 40738 20590
rect 52782 20578 52834 20590
rect 42130 20526 42142 20578
rect 42194 20526 42206 20578
rect 46834 20526 46846 20578
rect 46898 20526 46910 20578
rect 47618 20526 47630 20578
rect 47682 20526 47694 20578
rect 48962 20526 48974 20578
rect 49026 20526 49038 20578
rect 50418 20526 50430 20578
rect 50482 20526 50494 20578
rect 40686 20514 40738 20526
rect 52782 20514 52834 20526
rect 76638 20578 76690 20590
rect 76638 20514 76690 20526
rect 1344 20410 78624 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 50558 20410
rect 50610 20358 50662 20410
rect 50714 20358 50766 20410
rect 50818 20358 78624 20410
rect 1344 20324 78624 20358
rect 19070 20242 19122 20254
rect 19070 20178 19122 20190
rect 19854 20242 19906 20254
rect 19854 20178 19906 20190
rect 33406 20242 33458 20254
rect 33406 20178 33458 20190
rect 33854 20242 33906 20254
rect 33854 20178 33906 20190
rect 34302 20242 34354 20254
rect 39902 20242 39954 20254
rect 48078 20242 48130 20254
rect 72942 20242 72994 20254
rect 37538 20190 37550 20242
rect 37602 20190 37614 20242
rect 42802 20190 42814 20242
rect 42866 20190 42878 20242
rect 51538 20190 51550 20242
rect 51602 20190 51614 20242
rect 52322 20190 52334 20242
rect 52386 20190 52398 20242
rect 34302 20178 34354 20190
rect 39902 20178 39954 20190
rect 48078 20178 48130 20190
rect 72942 20178 72994 20190
rect 73950 20242 74002 20254
rect 73950 20178 74002 20190
rect 18622 20130 18674 20142
rect 18622 20066 18674 20078
rect 19630 20130 19682 20142
rect 19630 20066 19682 20078
rect 21310 20130 21362 20142
rect 21310 20066 21362 20078
rect 25566 20130 25618 20142
rect 25566 20066 25618 20078
rect 35086 20130 35138 20142
rect 35086 20066 35138 20078
rect 35534 20130 35586 20142
rect 47406 20130 47458 20142
rect 35858 20078 35870 20130
rect 35922 20078 35934 20130
rect 40898 20078 40910 20130
rect 40962 20078 40974 20130
rect 42914 20078 42926 20130
rect 42978 20078 42990 20130
rect 44482 20078 44494 20130
rect 44546 20078 44558 20130
rect 35534 20066 35586 20078
rect 47406 20066 47458 20078
rect 48190 20130 48242 20142
rect 57598 20130 57650 20142
rect 49410 20078 49422 20130
rect 49474 20078 49486 20130
rect 51090 20078 51102 20130
rect 51154 20078 51166 20130
rect 53218 20078 53230 20130
rect 53282 20078 53294 20130
rect 54338 20078 54350 20130
rect 54402 20078 54414 20130
rect 48190 20066 48242 20078
rect 57598 20066 57650 20078
rect 75070 20130 75122 20142
rect 75070 20066 75122 20078
rect 75630 20130 75682 20142
rect 76750 20130 76802 20142
rect 76066 20078 76078 20130
rect 76130 20078 76142 20130
rect 75630 20066 75682 20078
rect 76750 20066 76802 20078
rect 77646 20130 77698 20142
rect 77646 20066 77698 20078
rect 78318 20130 78370 20142
rect 78318 20066 78370 20078
rect 18958 20018 19010 20030
rect 18958 19954 19010 19966
rect 19518 20018 19570 20030
rect 19518 19954 19570 19966
rect 20190 20018 20242 20030
rect 25230 20018 25282 20030
rect 33742 20018 33794 20030
rect 21634 19966 21646 20018
rect 21698 19966 21710 20018
rect 26450 19966 26462 20018
rect 26514 19966 26526 20018
rect 29586 19966 29598 20018
rect 29650 19966 29662 20018
rect 20190 19954 20242 19966
rect 25230 19954 25282 19966
rect 33742 19954 33794 19966
rect 34862 20018 34914 20030
rect 34862 19954 34914 19966
rect 35198 20018 35250 20030
rect 39454 20018 39506 20030
rect 36306 19966 36318 20018
rect 36370 19966 36382 20018
rect 37650 19966 37662 20018
rect 37714 19966 37726 20018
rect 37986 19966 37998 20018
rect 38050 19966 38062 20018
rect 35198 19954 35250 19966
rect 39454 19954 39506 19966
rect 39678 20018 39730 20030
rect 39678 19954 39730 19966
rect 40014 20018 40066 20030
rect 55022 20018 55074 20030
rect 41122 19966 41134 20018
rect 41186 19966 41198 20018
rect 43026 19966 43038 20018
rect 43090 19966 43102 20018
rect 44706 19966 44718 20018
rect 44770 19966 44782 20018
rect 46274 19966 46286 20018
rect 46338 19966 46350 20018
rect 46722 19966 46734 20018
rect 46786 19966 46798 20018
rect 48738 19966 48750 20018
rect 48802 19966 48814 20018
rect 49298 19966 49310 20018
rect 49362 19966 49374 20018
rect 50866 19966 50878 20018
rect 50930 19966 50942 20018
rect 51762 19966 51774 20018
rect 51826 19966 51838 20018
rect 52098 19966 52110 20018
rect 52162 19966 52174 20018
rect 52882 19966 52894 20018
rect 52946 19966 52958 20018
rect 53554 19966 53566 20018
rect 53618 19966 53630 20018
rect 54226 19966 54238 20018
rect 54290 19966 54302 20018
rect 40014 19954 40066 19966
rect 55022 19954 55074 19966
rect 56702 20018 56754 20030
rect 77422 20018 77474 20030
rect 74834 19966 74846 20018
rect 74898 19966 74910 20018
rect 76290 19966 76302 20018
rect 76354 19966 76366 20018
rect 77074 19966 77086 20018
rect 77138 19966 77150 20018
rect 56702 19954 56754 19966
rect 77422 19954 77474 19966
rect 26014 19906 26066 19918
rect 33294 19906 33346 19918
rect 20962 19854 20974 19906
rect 21026 19854 21038 19906
rect 22418 19854 22430 19906
rect 22482 19854 22494 19906
rect 24546 19854 24558 19906
rect 24610 19854 24622 19906
rect 27122 19854 27134 19906
rect 27186 19854 27198 19906
rect 29250 19854 29262 19906
rect 29314 19854 29326 19906
rect 30370 19854 30382 19906
rect 30434 19854 30446 19906
rect 32498 19854 32510 19906
rect 32562 19854 32574 19906
rect 26014 19842 26066 19854
rect 33294 19842 33346 19854
rect 34190 19906 34242 19918
rect 50318 19906 50370 19918
rect 56030 19906 56082 19918
rect 49522 19854 49534 19906
rect 49586 19854 49598 19906
rect 54002 19854 54014 19906
rect 54066 19854 54078 19906
rect 55458 19854 55470 19906
rect 55522 19854 55534 19906
rect 34190 19842 34242 19854
rect 50318 19842 50370 19854
rect 56030 19842 56082 19854
rect 57150 19906 57202 19918
rect 57150 19842 57202 19854
rect 75406 19906 75458 19918
rect 75730 19854 75742 19906
rect 75794 19854 75806 19906
rect 76962 19854 76974 19906
rect 77026 19854 77038 19906
rect 77634 19854 77646 19906
rect 77698 19854 77710 19906
rect 75406 19842 75458 19854
rect 19070 19794 19122 19806
rect 19070 19730 19122 19742
rect 1344 19626 78624 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 65918 19626
rect 65970 19574 66022 19626
rect 66074 19574 66126 19626
rect 66178 19574 78624 19626
rect 1344 19540 78624 19574
rect 33966 19458 34018 19470
rect 32162 19406 32174 19458
rect 32226 19455 32238 19458
rect 32834 19455 32846 19458
rect 32226 19409 32846 19455
rect 32226 19406 32238 19409
rect 32834 19406 32846 19409
rect 32898 19406 32910 19458
rect 33966 19394 34018 19406
rect 22654 19346 22706 19358
rect 22654 19282 22706 19294
rect 27470 19346 27522 19358
rect 27470 19282 27522 19294
rect 28590 19346 28642 19358
rect 30382 19346 30434 19358
rect 29026 19294 29038 19346
rect 29090 19343 29102 19346
rect 29250 19343 29262 19346
rect 29090 19297 29262 19343
rect 29090 19294 29102 19297
rect 29250 19294 29262 19297
rect 29314 19294 29326 19346
rect 28590 19282 28642 19294
rect 30382 19282 30434 19294
rect 31278 19346 31330 19358
rect 31278 19282 31330 19294
rect 33070 19346 33122 19358
rect 33070 19282 33122 19294
rect 35422 19346 35474 19358
rect 35422 19282 35474 19294
rect 38110 19346 38162 19358
rect 38110 19282 38162 19294
rect 48526 19346 48578 19358
rect 75070 19346 75122 19358
rect 53666 19294 53678 19346
rect 53730 19294 53742 19346
rect 48526 19282 48578 19294
rect 75070 19282 75122 19294
rect 22094 19234 22146 19246
rect 19282 19182 19294 19234
rect 19346 19182 19358 19234
rect 21746 19182 21758 19234
rect 21810 19182 21822 19234
rect 22094 19170 22146 19182
rect 22542 19234 22594 19246
rect 22542 19170 22594 19182
rect 26910 19234 26962 19246
rect 26910 19170 26962 19182
rect 27582 19234 27634 19246
rect 27582 19170 27634 19182
rect 29934 19234 29986 19246
rect 29934 19170 29986 19182
rect 30270 19234 30322 19246
rect 30270 19170 30322 19182
rect 30494 19234 30546 19246
rect 30494 19170 30546 19182
rect 34638 19234 34690 19246
rect 34638 19170 34690 19182
rect 35646 19234 35698 19246
rect 35646 19170 35698 19182
rect 36430 19234 36482 19246
rect 37998 19234 38050 19246
rect 37314 19182 37326 19234
rect 37378 19182 37390 19234
rect 36430 19170 36482 19182
rect 37998 19170 38050 19182
rect 38334 19234 38386 19246
rect 38334 19170 38386 19182
rect 38446 19234 38498 19246
rect 38446 19170 38498 19182
rect 39118 19234 39170 19246
rect 39118 19170 39170 19182
rect 39342 19234 39394 19246
rect 39342 19170 39394 19182
rect 40238 19234 40290 19246
rect 40238 19170 40290 19182
rect 40798 19234 40850 19246
rect 40798 19170 40850 19182
rect 41022 19234 41074 19246
rect 44830 19234 44882 19246
rect 78206 19234 78258 19246
rect 41682 19182 41694 19234
rect 41746 19182 41758 19234
rect 43362 19182 43374 19234
rect 43426 19182 43438 19234
rect 45378 19182 45390 19234
rect 45442 19182 45454 19234
rect 46610 19182 46622 19234
rect 46674 19182 46686 19234
rect 47170 19182 47182 19234
rect 47234 19182 47246 19234
rect 49746 19182 49758 19234
rect 49810 19182 49822 19234
rect 50978 19182 50990 19234
rect 51042 19182 51054 19234
rect 52658 19182 52670 19234
rect 52722 19182 52734 19234
rect 53330 19182 53342 19234
rect 53394 19182 53406 19234
rect 54562 19182 54574 19234
rect 54626 19182 54638 19234
rect 56130 19182 56142 19234
rect 56194 19182 56206 19234
rect 57026 19182 57038 19234
rect 57090 19182 57102 19234
rect 76850 19182 76862 19234
rect 76914 19182 76926 19234
rect 41022 19170 41074 19182
rect 44830 19170 44882 19182
rect 78206 19170 78258 19182
rect 1710 19122 1762 19134
rect 1710 19058 1762 19070
rect 2046 19122 2098 19134
rect 2046 19058 2098 19070
rect 2494 19122 2546 19134
rect 2494 19058 2546 19070
rect 19070 19122 19122 19134
rect 22766 19122 22818 19134
rect 21522 19070 21534 19122
rect 21586 19070 21598 19122
rect 19070 19058 19122 19070
rect 22766 19058 22818 19070
rect 23102 19122 23154 19134
rect 23102 19058 23154 19070
rect 23326 19122 23378 19134
rect 23326 19058 23378 19070
rect 24446 19122 24498 19134
rect 24446 19058 24498 19070
rect 24782 19122 24834 19134
rect 25566 19122 25618 19134
rect 25106 19070 25118 19122
rect 25170 19070 25182 19122
rect 24782 19058 24834 19070
rect 25566 19058 25618 19070
rect 25902 19122 25954 19134
rect 25902 19058 25954 19070
rect 26238 19122 26290 19134
rect 26238 19058 26290 19070
rect 29710 19122 29762 19134
rect 33854 19122 33906 19134
rect 35310 19122 35362 19134
rect 33394 19070 33406 19122
rect 33458 19070 33470 19122
rect 34962 19070 34974 19122
rect 35026 19070 35038 19122
rect 29710 19058 29762 19070
rect 33854 19058 33906 19070
rect 35310 19058 35362 19070
rect 35870 19122 35922 19134
rect 35870 19058 35922 19070
rect 36318 19122 36370 19134
rect 36318 19058 36370 19070
rect 37102 19122 37154 19134
rect 37102 19058 37154 19070
rect 38894 19122 38946 19134
rect 38894 19058 38946 19070
rect 39902 19122 39954 19134
rect 39902 19058 39954 19070
rect 40462 19122 40514 19134
rect 40462 19058 40514 19070
rect 40574 19122 40626 19134
rect 76526 19122 76578 19134
rect 42914 19070 42926 19122
rect 42978 19070 42990 19122
rect 49298 19070 49310 19122
rect 49362 19070 49374 19122
rect 51090 19070 51102 19122
rect 51154 19070 51166 19122
rect 53442 19070 53454 19122
rect 53506 19070 53518 19122
rect 54786 19070 54798 19122
rect 54850 19070 54862 19122
rect 40574 19058 40626 19070
rect 76526 19058 76578 19070
rect 77198 19122 77250 19134
rect 77198 19058 77250 19070
rect 77534 19122 77586 19134
rect 77534 19058 77586 19070
rect 23214 19010 23266 19022
rect 23214 18946 23266 18958
rect 23550 19010 23602 19022
rect 23550 18946 23602 18958
rect 24110 19010 24162 19022
rect 24110 18946 24162 18958
rect 24334 19010 24386 19022
rect 24334 18946 24386 18958
rect 26350 19010 26402 19022
rect 26350 18946 26402 18958
rect 26574 19010 26626 19022
rect 26574 18946 26626 18958
rect 27358 19010 27410 19022
rect 27358 18946 27410 18958
rect 28478 19010 28530 19022
rect 28478 18946 28530 18958
rect 29486 19010 29538 19022
rect 29486 18946 29538 18958
rect 29822 19010 29874 19022
rect 29822 18946 29874 18958
rect 30718 19010 30770 19022
rect 30718 18946 30770 18958
rect 31950 19010 32002 19022
rect 31950 18946 32002 18958
rect 32286 19010 32338 19022
rect 32286 18946 32338 18958
rect 32734 19010 32786 19022
rect 32734 18946 32786 18958
rect 39118 19010 39170 19022
rect 39118 18946 39170 18958
rect 40014 19010 40066 19022
rect 75406 19010 75458 19022
rect 43026 18958 43038 19010
rect 43090 18958 43102 19010
rect 46610 18958 46622 19010
rect 46674 18958 46686 19010
rect 49970 18958 49982 19010
rect 50034 18958 50046 19010
rect 56354 18958 56366 19010
rect 56418 18958 56430 19010
rect 40014 18946 40066 18958
rect 75406 18946 75458 18958
rect 76638 19010 76690 19022
rect 76638 18946 76690 18958
rect 77870 19010 77922 19022
rect 77870 18946 77922 18958
rect 1344 18842 78624 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 50558 18842
rect 50610 18790 50662 18842
rect 50714 18790 50766 18842
rect 50818 18790 78624 18842
rect 1344 18756 78624 18790
rect 17838 18674 17890 18686
rect 17838 18610 17890 18622
rect 41358 18674 41410 18686
rect 41358 18610 41410 18622
rect 41918 18674 41970 18686
rect 41918 18610 41970 18622
rect 42366 18674 42418 18686
rect 76750 18674 76802 18686
rect 49858 18622 49870 18674
rect 49922 18622 49934 18674
rect 54786 18622 54798 18674
rect 54850 18622 54862 18674
rect 71250 18622 71262 18674
rect 71314 18622 71326 18674
rect 42366 18610 42418 18622
rect 76750 18610 76802 18622
rect 2046 18562 2098 18574
rect 2046 18498 2098 18510
rect 17950 18562 18002 18574
rect 17950 18498 18002 18510
rect 24334 18562 24386 18574
rect 41806 18562 41858 18574
rect 77422 18562 77474 18574
rect 30034 18510 30046 18562
rect 30098 18510 30110 18562
rect 44034 18510 44046 18562
rect 44098 18510 44110 18562
rect 48850 18510 48862 18562
rect 48914 18510 48926 18562
rect 51090 18510 51102 18562
rect 51154 18510 51166 18562
rect 53218 18510 53230 18562
rect 53282 18510 53294 18562
rect 55122 18510 55134 18562
rect 55186 18510 55198 18562
rect 24334 18498 24386 18510
rect 41806 18498 41858 18510
rect 77422 18498 77474 18510
rect 1710 18450 1762 18462
rect 24670 18450 24722 18462
rect 23426 18398 23438 18450
rect 23490 18398 23502 18450
rect 1710 18386 1762 18398
rect 24670 18386 24722 18398
rect 25342 18450 25394 18462
rect 39230 18450 39282 18462
rect 25778 18398 25790 18450
rect 25842 18398 25854 18450
rect 29362 18398 29374 18450
rect 29426 18398 29438 18450
rect 33618 18398 33630 18450
rect 33682 18398 33694 18450
rect 25342 18386 25394 18398
rect 39230 18386 39282 18398
rect 39342 18450 39394 18462
rect 39342 18386 39394 18398
rect 39790 18450 39842 18462
rect 39790 18386 39842 18398
rect 40014 18450 40066 18462
rect 40014 18386 40066 18398
rect 41246 18450 41298 18462
rect 41246 18386 41298 18398
rect 42702 18450 42754 18462
rect 56702 18450 56754 18462
rect 44258 18398 44270 18450
rect 44322 18398 44334 18450
rect 45602 18398 45614 18450
rect 45666 18398 45678 18450
rect 47842 18398 47854 18450
rect 47906 18398 47918 18450
rect 49970 18398 49982 18450
rect 50034 18398 50046 18450
rect 50866 18398 50878 18450
rect 50930 18398 50942 18450
rect 52994 18398 53006 18450
rect 53058 18398 53070 18450
rect 54898 18398 54910 18450
rect 54962 18398 54974 18450
rect 42702 18386 42754 18398
rect 56702 18386 56754 18398
rect 70926 18450 70978 18462
rect 70926 18386 70978 18398
rect 77198 18450 77250 18462
rect 78318 18450 78370 18462
rect 77746 18398 77758 18450
rect 77810 18398 77822 18450
rect 77198 18386 77250 18398
rect 78318 18386 78370 18398
rect 2494 18338 2546 18350
rect 23998 18338 24050 18350
rect 39566 18338 39618 18350
rect 18834 18286 18846 18338
rect 18898 18286 18910 18338
rect 26450 18286 26462 18338
rect 26514 18286 26526 18338
rect 28578 18286 28590 18338
rect 28642 18286 28654 18338
rect 32162 18286 32174 18338
rect 32226 18286 32238 18338
rect 38210 18286 38222 18338
rect 38274 18286 38286 18338
rect 2494 18274 2546 18286
rect 23998 18274 24050 18286
rect 39566 18274 39618 18286
rect 43038 18338 43090 18350
rect 43038 18274 43090 18286
rect 43150 18338 43202 18350
rect 52558 18338 52610 18350
rect 45490 18286 45502 18338
rect 45554 18286 45566 18338
rect 43150 18274 43202 18286
rect 52558 18274 52610 18286
rect 57150 18338 57202 18350
rect 57150 18274 57202 18286
rect 70590 18338 70642 18350
rect 70590 18274 70642 18286
rect 17838 18226 17890 18238
rect 17838 18162 17890 18174
rect 41358 18226 41410 18238
rect 41358 18162 41410 18174
rect 41918 18226 41970 18238
rect 47182 18226 47234 18238
rect 44034 18174 44046 18226
rect 44098 18174 44110 18226
rect 41918 18162 41970 18174
rect 47182 18162 47234 18174
rect 77758 18226 77810 18238
rect 77758 18162 77810 18174
rect 1344 18058 78624 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 65918 18058
rect 65970 18006 66022 18058
rect 66074 18006 66126 18058
rect 66178 18006 78624 18058
rect 1344 17972 78624 18006
rect 17726 17778 17778 17790
rect 17726 17714 17778 17726
rect 18174 17778 18226 17790
rect 27918 17778 27970 17790
rect 22306 17726 22318 17778
rect 22370 17726 22382 17778
rect 18174 17714 18226 17726
rect 27918 17714 27970 17726
rect 28590 17778 28642 17790
rect 28590 17714 28642 17726
rect 36318 17778 36370 17790
rect 36318 17714 36370 17726
rect 37102 17778 37154 17790
rect 37102 17714 37154 17726
rect 39118 17778 39170 17790
rect 39118 17714 39170 17726
rect 47742 17778 47794 17790
rect 47742 17714 47794 17726
rect 48526 17778 48578 17790
rect 48526 17714 48578 17726
rect 18846 17666 18898 17678
rect 18846 17602 18898 17614
rect 19182 17666 19234 17678
rect 19182 17602 19234 17614
rect 19854 17666 19906 17678
rect 19854 17602 19906 17614
rect 19966 17666 20018 17678
rect 35646 17666 35698 17678
rect 27234 17614 27246 17666
rect 27298 17614 27310 17666
rect 33618 17614 33630 17666
rect 33682 17614 33694 17666
rect 19966 17602 20018 17614
rect 35646 17602 35698 17614
rect 35870 17666 35922 17678
rect 35870 17602 35922 17614
rect 37214 17666 37266 17678
rect 37214 17602 37266 17614
rect 37998 17666 38050 17678
rect 37998 17602 38050 17614
rect 38446 17666 38498 17678
rect 38446 17602 38498 17614
rect 38670 17666 38722 17678
rect 38670 17602 38722 17614
rect 39342 17666 39394 17678
rect 39342 17602 39394 17614
rect 39790 17666 39842 17678
rect 39790 17602 39842 17614
rect 40014 17666 40066 17678
rect 40014 17602 40066 17614
rect 40686 17666 40738 17678
rect 42926 17666 42978 17678
rect 44830 17666 44882 17678
rect 56590 17666 56642 17678
rect 78206 17666 78258 17678
rect 41346 17614 41358 17666
rect 41410 17614 41422 17666
rect 43138 17614 43150 17666
rect 43202 17614 43214 17666
rect 45378 17614 45390 17666
rect 45442 17614 45454 17666
rect 46946 17614 46958 17666
rect 47010 17614 47022 17666
rect 49634 17614 49646 17666
rect 49698 17614 49710 17666
rect 51314 17614 51326 17666
rect 51378 17614 51390 17666
rect 53218 17614 53230 17666
rect 53282 17614 53294 17666
rect 55458 17614 55470 17666
rect 55522 17614 55534 17666
rect 56802 17614 56814 17666
rect 56866 17614 56878 17666
rect 58706 17614 58718 17666
rect 58770 17614 58782 17666
rect 40686 17602 40738 17614
rect 42926 17602 42978 17614
rect 44830 17602 44882 17614
rect 56590 17602 56642 17614
rect 78206 17602 78258 17614
rect 1710 17554 1762 17566
rect 1710 17490 1762 17502
rect 2046 17554 2098 17566
rect 2046 17490 2098 17502
rect 19518 17554 19570 17566
rect 19518 17490 19570 17502
rect 21310 17554 21362 17566
rect 35310 17554 35362 17566
rect 21634 17502 21646 17554
rect 21698 17502 21710 17554
rect 29586 17502 29598 17554
rect 29650 17502 29662 17554
rect 21310 17490 21362 17502
rect 35310 17490 35362 17502
rect 36990 17554 37042 17566
rect 36990 17490 37042 17502
rect 37550 17554 37602 17566
rect 37550 17490 37602 17502
rect 40350 17554 40402 17566
rect 51774 17554 51826 17566
rect 76974 17554 77026 17566
rect 41458 17502 41470 17554
rect 41522 17502 41534 17554
rect 47058 17502 47070 17554
rect 47122 17502 47134 17554
rect 49186 17502 49198 17554
rect 49250 17502 49262 17554
rect 51090 17502 51102 17554
rect 51154 17502 51166 17554
rect 53442 17502 53454 17554
rect 53506 17502 53518 17554
rect 55122 17502 55134 17554
rect 55186 17502 55198 17554
rect 58818 17502 58830 17554
rect 58882 17502 58894 17554
rect 40350 17490 40402 17502
rect 51774 17490 51826 17502
rect 76974 17490 77026 17502
rect 77198 17554 77250 17566
rect 77198 17490 77250 17502
rect 77534 17554 77586 17566
rect 77534 17490 77586 17502
rect 77870 17554 77922 17566
rect 77870 17490 77922 17502
rect 2494 17442 2546 17454
rect 2494 17378 2546 17390
rect 18958 17442 19010 17454
rect 18958 17378 19010 17390
rect 19742 17442 19794 17454
rect 19742 17378 19794 17390
rect 20414 17442 20466 17454
rect 20414 17378 20466 17390
rect 28478 17442 28530 17454
rect 28478 17378 28530 17390
rect 35534 17442 35586 17454
rect 35534 17378 35586 17390
rect 38222 17442 38274 17454
rect 38222 17378 38274 17390
rect 39678 17442 39730 17454
rect 43026 17390 43038 17442
rect 43090 17390 43102 17442
rect 54114 17390 54126 17442
rect 54178 17390 54190 17442
rect 57698 17390 57710 17442
rect 57762 17390 57774 17442
rect 39678 17378 39730 17390
rect 1344 17274 78624 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 50558 17274
rect 50610 17222 50662 17274
rect 50714 17222 50766 17274
rect 50818 17222 78624 17274
rect 1344 17188 78624 17222
rect 26350 17106 26402 17118
rect 26350 17042 26402 17054
rect 26686 17106 26738 17118
rect 26686 17042 26738 17054
rect 26798 17106 26850 17118
rect 26798 17042 26850 17054
rect 27582 17106 27634 17118
rect 27582 17042 27634 17054
rect 28142 17106 28194 17118
rect 28142 17042 28194 17054
rect 32510 17106 32562 17118
rect 32510 17042 32562 17054
rect 33854 17106 33906 17118
rect 33854 17042 33906 17054
rect 34302 17106 34354 17118
rect 34302 17042 34354 17054
rect 35198 17106 35250 17118
rect 35198 17042 35250 17054
rect 35982 17106 36034 17118
rect 35982 17042 36034 17054
rect 37102 17106 37154 17118
rect 37102 17042 37154 17054
rect 37550 17106 37602 17118
rect 37550 17042 37602 17054
rect 37998 17106 38050 17118
rect 37998 17042 38050 17054
rect 39006 17106 39058 17118
rect 39006 17042 39058 17054
rect 39790 17106 39842 17118
rect 39790 17042 39842 17054
rect 41134 17106 41186 17118
rect 41134 17042 41186 17054
rect 41694 17106 41746 17118
rect 41694 17042 41746 17054
rect 42142 17106 42194 17118
rect 42142 17042 42194 17054
rect 42590 17106 42642 17118
rect 42590 17042 42642 17054
rect 44270 17106 44322 17118
rect 57150 17106 57202 17118
rect 48066 17054 48078 17106
rect 48130 17054 48142 17106
rect 49970 17054 49982 17106
rect 50034 17054 50046 17106
rect 44270 17042 44322 17054
rect 57150 17042 57202 17054
rect 77646 17106 77698 17118
rect 77646 17042 77698 17054
rect 77870 17106 77922 17118
rect 77870 17042 77922 17054
rect 27022 16994 27074 17006
rect 36094 16994 36146 17006
rect 19282 16942 19294 16994
rect 19346 16942 19358 16994
rect 22530 16942 22542 16994
rect 22594 16942 22606 16994
rect 32050 16942 32062 16994
rect 32114 16942 32126 16994
rect 27022 16930 27074 16942
rect 36094 16930 36146 16942
rect 39902 16994 39954 17006
rect 39902 16930 39954 16942
rect 41358 16994 41410 17006
rect 41358 16930 41410 16942
rect 41470 16994 41522 17006
rect 45614 16994 45666 17006
rect 42914 16942 42926 16994
rect 42978 16942 42990 16994
rect 47394 16942 47406 16994
rect 47458 16942 47470 16994
rect 49298 16942 49310 16994
rect 49362 16942 49374 16994
rect 51090 16942 51102 16994
rect 51154 16942 51166 16994
rect 52434 16942 52446 16994
rect 52498 16942 52510 16994
rect 41470 16930 41522 16942
rect 45614 16930 45666 16942
rect 26574 16882 26626 16894
rect 33518 16882 33570 16894
rect 18610 16830 18622 16882
rect 18674 16830 18686 16882
rect 21858 16830 21870 16882
rect 21922 16830 21934 16882
rect 28578 16830 28590 16882
rect 28642 16830 28654 16882
rect 26574 16818 26626 16830
rect 33518 16818 33570 16830
rect 34638 16882 34690 16894
rect 34638 16818 34690 16830
rect 34750 16882 34802 16894
rect 34750 16818 34802 16830
rect 35646 16882 35698 16894
rect 35646 16818 35698 16830
rect 36206 16882 36258 16894
rect 36206 16818 36258 16830
rect 37438 16882 37490 16894
rect 37438 16818 37490 16830
rect 38670 16882 38722 16894
rect 38670 16818 38722 16830
rect 38894 16882 38946 16894
rect 38894 16818 38946 16830
rect 39230 16882 39282 16894
rect 39230 16818 39282 16830
rect 39454 16882 39506 16894
rect 39454 16818 39506 16830
rect 40126 16882 40178 16894
rect 40126 16818 40178 16830
rect 44606 16882 44658 16894
rect 54350 16882 54402 16894
rect 56702 16882 56754 16894
rect 46722 16830 46734 16882
rect 46786 16830 46798 16882
rect 47058 16830 47070 16882
rect 47122 16830 47134 16882
rect 48178 16830 48190 16882
rect 48242 16830 48254 16882
rect 49074 16830 49086 16882
rect 49138 16830 49150 16882
rect 50978 16830 50990 16882
rect 51042 16830 51054 16882
rect 52658 16830 52670 16882
rect 52722 16830 52734 16882
rect 54562 16830 54574 16882
rect 54626 16830 54638 16882
rect 44606 16818 44658 16830
rect 54350 16818 54402 16830
rect 56702 16818 56754 16830
rect 77198 16882 77250 16894
rect 78082 16830 78094 16882
rect 78146 16830 78158 16882
rect 77198 16818 77250 16830
rect 31726 16770 31778 16782
rect 21410 16718 21422 16770
rect 21474 16718 21486 16770
rect 24658 16718 24670 16770
rect 24722 16718 24734 16770
rect 29250 16718 29262 16770
rect 29314 16718 29326 16770
rect 31378 16718 31390 16770
rect 31442 16718 31454 16770
rect 31726 16706 31778 16718
rect 33742 16770 33794 16782
rect 33742 16706 33794 16718
rect 34190 16770 34242 16782
rect 34190 16706 34242 16718
rect 37886 16770 37938 16782
rect 37886 16706 37938 16718
rect 55358 16770 55410 16782
rect 55358 16706 55410 16718
rect 1344 16490 78624 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 65918 16490
rect 65970 16438 66022 16490
rect 66074 16438 66126 16490
rect 66178 16438 78624 16490
rect 1344 16404 78624 16438
rect 37102 16322 37154 16334
rect 37102 16258 37154 16270
rect 37998 16322 38050 16334
rect 37998 16258 38050 16270
rect 38446 16322 38498 16334
rect 38446 16258 38498 16270
rect 44046 16322 44098 16334
rect 44046 16258 44098 16270
rect 51102 16322 51154 16334
rect 51102 16258 51154 16270
rect 23774 16210 23826 16222
rect 28254 16210 28306 16222
rect 27906 16158 27918 16210
rect 27970 16158 27982 16210
rect 23774 16146 23826 16158
rect 28254 16146 28306 16158
rect 29262 16210 29314 16222
rect 29262 16146 29314 16158
rect 30158 16210 30210 16222
rect 36094 16210 36146 16222
rect 34962 16158 34974 16210
rect 35026 16158 35038 16210
rect 30158 16146 30210 16158
rect 36094 16146 36146 16158
rect 36542 16210 36594 16222
rect 36542 16146 36594 16158
rect 36990 16210 37042 16222
rect 36990 16146 37042 16158
rect 39678 16210 39730 16222
rect 39678 16146 39730 16158
rect 40462 16210 40514 16222
rect 40462 16146 40514 16158
rect 40910 16210 40962 16222
rect 40910 16146 40962 16158
rect 41470 16210 41522 16222
rect 41470 16146 41522 16158
rect 41918 16210 41970 16222
rect 41918 16146 41970 16158
rect 44942 16210 44994 16222
rect 44942 16146 44994 16158
rect 51998 16210 52050 16222
rect 51998 16146 52050 16158
rect 56478 16210 56530 16222
rect 56478 16146 56530 16158
rect 29374 16098 29426 16110
rect 35310 16098 35362 16110
rect 24994 16046 25006 16098
rect 25058 16046 25070 16098
rect 32162 16046 32174 16098
rect 32226 16046 32238 16098
rect 29374 16034 29426 16046
rect 35310 16034 35362 16046
rect 38894 16098 38946 16110
rect 38894 16034 38946 16046
rect 43038 16098 43090 16110
rect 43038 16034 43090 16046
rect 43374 16098 43426 16110
rect 43374 16034 43426 16046
rect 43710 16098 43762 16110
rect 43710 16034 43762 16046
rect 43934 16098 43986 16110
rect 46062 16098 46114 16110
rect 52670 16098 52722 16110
rect 45490 16046 45502 16098
rect 45554 16046 45566 16098
rect 47282 16046 47294 16098
rect 47346 16046 47358 16098
rect 48962 16046 48974 16098
rect 49026 16046 49038 16098
rect 50418 16046 50430 16098
rect 50482 16046 50494 16098
rect 52882 16046 52894 16098
rect 52946 16046 52958 16098
rect 54450 16046 54462 16098
rect 54514 16046 54526 16098
rect 54786 16046 54798 16098
rect 54850 16046 54862 16098
rect 43934 16034 43986 16046
rect 46062 16034 46114 16046
rect 52670 16034 52722 16046
rect 1710 15986 1762 15998
rect 1710 15922 1762 15934
rect 2046 15986 2098 15998
rect 37550 15986 37602 15998
rect 25778 15934 25790 15986
rect 25842 15934 25854 15986
rect 32834 15934 32846 15986
rect 32898 15934 32910 15986
rect 2046 15922 2098 15934
rect 37550 15922 37602 15934
rect 37886 15986 37938 15998
rect 37886 15922 37938 15934
rect 38334 15986 38386 15998
rect 42142 15986 42194 15998
rect 39218 15934 39230 15986
rect 39282 15934 39294 15986
rect 38334 15922 38386 15934
rect 42142 15922 42194 15934
rect 43486 15986 43538 15998
rect 77870 15986 77922 15998
rect 47730 15934 47742 15986
rect 47794 15934 47806 15986
rect 49522 15934 49534 15986
rect 49586 15934 49598 15986
rect 43486 15922 43538 15934
rect 77870 15922 77922 15934
rect 78206 15986 78258 15998
rect 78206 15922 78258 15934
rect 2494 15874 2546 15886
rect 2494 15810 2546 15822
rect 28366 15874 28418 15886
rect 28366 15810 28418 15822
rect 29150 15874 29202 15886
rect 29150 15810 29202 15822
rect 29598 15874 29650 15886
rect 29598 15810 29650 15822
rect 35422 15874 35474 15886
rect 35422 15810 35474 15822
rect 37438 15874 37490 15886
rect 37438 15810 37490 15822
rect 42254 15874 42306 15886
rect 42254 15810 42306 15822
rect 44046 15874 44098 15886
rect 51438 15874 51490 15886
rect 77646 15874 77698 15886
rect 45714 15822 45726 15874
rect 45778 15822 45790 15874
rect 46386 15822 46398 15874
rect 46450 15822 46462 15874
rect 47954 15822 47966 15874
rect 48018 15822 48030 15874
rect 53778 15822 53790 15874
rect 53842 15822 53854 15874
rect 44046 15810 44098 15822
rect 51438 15810 51490 15822
rect 77646 15810 77698 15822
rect 1344 15706 78624 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 50558 15706
rect 50610 15654 50662 15706
rect 50714 15654 50766 15706
rect 50818 15654 78624 15706
rect 1344 15620 78624 15654
rect 33518 15538 33570 15550
rect 33518 15474 33570 15486
rect 34078 15538 34130 15550
rect 34078 15474 34130 15486
rect 34526 15538 34578 15550
rect 34526 15474 34578 15486
rect 38558 15538 38610 15550
rect 38558 15474 38610 15486
rect 39006 15538 39058 15550
rect 39006 15474 39058 15486
rect 39454 15538 39506 15550
rect 39454 15474 39506 15486
rect 40126 15538 40178 15550
rect 46498 15486 46510 15538
rect 46562 15486 46574 15538
rect 40126 15474 40178 15486
rect 2046 15426 2098 15438
rect 33406 15426 33458 15438
rect 27234 15374 27246 15426
rect 27298 15374 27310 15426
rect 2046 15362 2098 15374
rect 33406 15362 33458 15374
rect 38894 15426 38946 15438
rect 47730 15374 47742 15426
rect 47794 15374 47806 15426
rect 48850 15374 48862 15426
rect 48914 15374 48926 15426
rect 50642 15374 50654 15426
rect 50706 15374 50718 15426
rect 52322 15374 52334 15426
rect 52386 15374 52398 15426
rect 38894 15362 38946 15374
rect 1710 15314 1762 15326
rect 32958 15314 33010 15326
rect 30818 15262 30830 15314
rect 30882 15262 30894 15314
rect 1710 15250 1762 15262
rect 32958 15250 33010 15262
rect 33630 15314 33682 15326
rect 39678 15314 39730 15326
rect 35186 15262 35198 15314
rect 35250 15262 35262 15314
rect 33630 15250 33682 15262
rect 39678 15250 39730 15262
rect 40350 15314 40402 15326
rect 54238 15314 54290 15326
rect 41682 15262 41694 15314
rect 41746 15262 41758 15314
rect 45490 15262 45502 15314
rect 45554 15262 45566 15314
rect 46386 15262 46398 15314
rect 46450 15262 46462 15314
rect 47170 15262 47182 15314
rect 47234 15262 47246 15314
rect 48962 15262 48974 15314
rect 49026 15262 49038 15314
rect 50866 15262 50878 15314
rect 50930 15262 50942 15314
rect 52546 15262 52558 15314
rect 52610 15262 52622 15314
rect 54450 15262 54462 15314
rect 54514 15262 54526 15314
rect 40350 15250 40402 15262
rect 54238 15250 54290 15262
rect 2494 15202 2546 15214
rect 2494 15138 2546 15150
rect 31390 15202 31442 15214
rect 31390 15138 31442 15150
rect 32510 15202 32562 15214
rect 40238 15202 40290 15214
rect 51662 15202 51714 15214
rect 35970 15150 35982 15202
rect 36034 15150 36046 15202
rect 38098 15150 38110 15202
rect 38162 15150 38174 15202
rect 42466 15150 42478 15202
rect 42530 15150 42542 15202
rect 44594 15150 44606 15202
rect 44658 15150 44670 15202
rect 32510 15138 32562 15150
rect 40238 15138 40290 15150
rect 51662 15138 51714 15150
rect 55246 15202 55298 15214
rect 55246 15138 55298 15150
rect 1344 14922 78624 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 65918 14922
rect 65970 14870 66022 14922
rect 66074 14870 66126 14922
rect 66178 14870 78624 14922
rect 1344 14836 78624 14870
rect 45166 14754 45218 14766
rect 43922 14702 43934 14754
rect 43986 14751 43998 14754
rect 44258 14751 44270 14754
rect 43986 14705 44270 14751
rect 43986 14702 43998 14705
rect 44258 14702 44270 14705
rect 44322 14702 44334 14754
rect 45166 14690 45218 14702
rect 53454 14754 53506 14766
rect 53454 14690 53506 14702
rect 26686 14642 26738 14654
rect 34526 14642 34578 14654
rect 35982 14642 36034 14654
rect 42590 14642 42642 14654
rect 34178 14590 34190 14642
rect 34242 14590 34254 14642
rect 34850 14590 34862 14642
rect 34914 14590 34926 14642
rect 40002 14590 40014 14642
rect 40066 14590 40078 14642
rect 42130 14590 42142 14642
rect 42194 14590 42206 14642
rect 26686 14578 26738 14590
rect 34526 14578 34578 14590
rect 35982 14578 36034 14590
rect 42590 14578 42642 14590
rect 43934 14642 43986 14654
rect 43934 14578 43986 14590
rect 44382 14642 44434 14654
rect 44382 14578 44434 14590
rect 45726 14642 45778 14654
rect 45726 14578 45778 14590
rect 50094 14642 50146 14654
rect 50094 14578 50146 14590
rect 50654 14642 50706 14654
rect 50654 14578 50706 14590
rect 26126 14530 26178 14542
rect 35422 14530 35474 14542
rect 31378 14478 31390 14530
rect 31442 14478 31454 14530
rect 26126 14466 26178 14478
rect 35422 14466 35474 14478
rect 35870 14530 35922 14542
rect 42702 14530 42754 14542
rect 39218 14478 39230 14530
rect 39282 14478 39294 14530
rect 35870 14466 35922 14478
rect 42702 14466 42754 14478
rect 45054 14530 45106 14542
rect 52670 14530 52722 14542
rect 47506 14478 47518 14530
rect 47570 14478 47582 14530
rect 48178 14478 48190 14530
rect 48242 14478 48254 14530
rect 48738 14478 48750 14530
rect 48802 14478 48814 14530
rect 51314 14478 51326 14530
rect 51378 14478 51390 14530
rect 45054 14466 45106 14478
rect 52670 14466 52722 14478
rect 26798 14418 26850 14430
rect 29150 14418 29202 14430
rect 28242 14366 28254 14418
rect 28306 14366 28318 14418
rect 26798 14354 26850 14366
rect 29150 14354 29202 14366
rect 30942 14418 30994 14430
rect 42926 14418 42978 14430
rect 77870 14418 77922 14430
rect 32050 14366 32062 14418
rect 32114 14366 32126 14418
rect 46834 14366 46846 14418
rect 46898 14366 46910 14418
rect 30942 14354 30994 14366
rect 42926 14354 42978 14366
rect 77870 14354 77922 14366
rect 78206 14418 78258 14430
rect 78206 14354 78258 14366
rect 26574 14306 26626 14318
rect 26574 14242 26626 14254
rect 27246 14306 27298 14318
rect 27246 14242 27298 14254
rect 28590 14306 28642 14318
rect 28590 14242 28642 14254
rect 29262 14306 29314 14318
rect 29262 14242 29314 14254
rect 29374 14306 29426 14318
rect 29374 14242 29426 14254
rect 29598 14306 29650 14318
rect 29598 14242 29650 14254
rect 30158 14306 30210 14318
rect 30158 14242 30210 14254
rect 30830 14306 30882 14318
rect 30830 14242 30882 14254
rect 36094 14306 36146 14318
rect 36094 14242 36146 14254
rect 42478 14306 42530 14318
rect 51998 14306 52050 14318
rect 48402 14254 48414 14306
rect 48466 14254 48478 14306
rect 42478 14242 42530 14254
rect 51998 14242 52050 14254
rect 77646 14306 77698 14318
rect 77646 14242 77698 14254
rect 1344 14138 78624 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 50558 14138
rect 50610 14086 50662 14138
rect 50714 14086 50766 14138
rect 50818 14086 78624 14138
rect 1344 14052 78624 14086
rect 2046 13970 2098 13982
rect 2046 13906 2098 13918
rect 25902 13970 25954 13982
rect 25902 13906 25954 13918
rect 27022 13970 27074 13982
rect 27022 13906 27074 13918
rect 28142 13970 28194 13982
rect 28142 13906 28194 13918
rect 33406 13970 33458 13982
rect 33406 13906 33458 13918
rect 33518 13970 33570 13982
rect 33518 13906 33570 13918
rect 33630 13970 33682 13982
rect 33630 13906 33682 13918
rect 34190 13970 34242 13982
rect 34190 13906 34242 13918
rect 34414 13970 34466 13982
rect 40238 13970 40290 13982
rect 39330 13918 39342 13970
rect 39394 13918 39406 13970
rect 34414 13906 34466 13918
rect 40238 13906 40290 13918
rect 41582 13970 41634 13982
rect 41582 13906 41634 13918
rect 48302 13970 48354 13982
rect 48302 13906 48354 13918
rect 48974 13970 49026 13982
rect 48974 13906 49026 13918
rect 49422 13970 49474 13982
rect 77870 13970 77922 13982
rect 52210 13918 52222 13970
rect 52274 13918 52286 13970
rect 49422 13906 49474 13918
rect 77870 13906 77922 13918
rect 26126 13858 26178 13870
rect 26126 13794 26178 13806
rect 26686 13858 26738 13870
rect 26686 13794 26738 13806
rect 27246 13858 27298 13870
rect 27246 13794 27298 13806
rect 27918 13858 27970 13870
rect 40014 13858 40066 13870
rect 29138 13806 29150 13858
rect 29202 13806 29214 13858
rect 34738 13806 34750 13858
rect 34802 13806 34814 13858
rect 51986 13806 51998 13858
rect 52050 13806 52062 13858
rect 53890 13806 53902 13858
rect 53954 13806 53966 13858
rect 27918 13794 27970 13806
rect 40014 13794 40066 13806
rect 1710 13746 1762 13758
rect 26238 13746 26290 13758
rect 19618 13694 19630 13746
rect 19682 13694 19694 13746
rect 23426 13694 23438 13746
rect 23490 13694 23502 13746
rect 1710 13682 1762 13694
rect 26238 13682 26290 13694
rect 26574 13746 26626 13758
rect 26574 13682 26626 13694
rect 27358 13746 27410 13758
rect 27358 13682 27410 13694
rect 27806 13746 27858 13758
rect 38334 13746 38386 13758
rect 28466 13694 28478 13746
rect 28530 13694 28542 13746
rect 33058 13694 33070 13746
rect 33122 13694 33134 13746
rect 35074 13694 35086 13746
rect 35138 13694 35150 13746
rect 27806 13682 27858 13694
rect 38334 13682 38386 13694
rect 39006 13746 39058 13758
rect 39006 13682 39058 13694
rect 39566 13746 39618 13758
rect 45278 13746 45330 13758
rect 42018 13694 42030 13746
rect 42082 13694 42094 13746
rect 39566 13682 39618 13694
rect 45278 13682 45330 13694
rect 45390 13746 45442 13758
rect 51314 13694 51326 13746
rect 51378 13694 51390 13746
rect 53554 13694 53566 13746
rect 53618 13694 53630 13746
rect 78082 13694 78094 13746
rect 78146 13694 78158 13746
rect 45390 13682 45442 13694
rect 2494 13634 2546 13646
rect 22542 13634 22594 13646
rect 20402 13582 20414 13634
rect 20466 13582 20478 13634
rect 2494 13570 2546 13582
rect 22542 13570 22594 13582
rect 23662 13634 23714 13646
rect 40126 13634 40178 13646
rect 31266 13582 31278 13634
rect 31330 13582 31342 13634
rect 35858 13582 35870 13634
rect 35922 13582 35934 13634
rect 37986 13582 37998 13634
rect 38050 13582 38062 13634
rect 23662 13570 23714 13582
rect 40126 13570 40178 13582
rect 41694 13634 41746 13646
rect 46958 13634 47010 13646
rect 42802 13582 42814 13634
rect 42866 13582 42878 13634
rect 44930 13582 44942 13634
rect 44994 13582 45006 13634
rect 41694 13570 41746 13582
rect 46958 13570 47010 13582
rect 77646 13634 77698 13646
rect 77646 13570 77698 13582
rect 23774 13522 23826 13534
rect 23774 13458 23826 13470
rect 26686 13522 26738 13534
rect 26686 13458 26738 13470
rect 38446 13522 38498 13534
rect 38446 13458 38498 13470
rect 1344 13354 78624 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 65918 13354
rect 65970 13302 66022 13354
rect 66074 13302 66126 13354
rect 66178 13302 78624 13354
rect 1344 13268 78624 13302
rect 32510 13186 32562 13198
rect 32510 13122 32562 13134
rect 33070 13186 33122 13198
rect 33070 13122 33122 13134
rect 33966 13186 34018 13198
rect 33966 13122 34018 13134
rect 21422 13074 21474 13086
rect 26574 13074 26626 13086
rect 19506 13022 19518 13074
rect 19570 13022 19582 13074
rect 23650 13022 23662 13074
rect 23714 13022 23726 13074
rect 25778 13022 25790 13074
rect 25842 13022 25854 13074
rect 21422 13010 21474 13022
rect 26574 13010 26626 13022
rect 35870 13074 35922 13086
rect 42926 13074 42978 13086
rect 39890 13022 39902 13074
rect 39954 13022 39966 13074
rect 42018 13022 42030 13074
rect 42082 13022 42094 13074
rect 35870 13010 35922 13022
rect 42926 13010 42978 13022
rect 19966 12962 20018 12974
rect 16594 12910 16606 12962
rect 16658 12910 16670 12962
rect 19966 12898 20018 12910
rect 20078 12962 20130 12974
rect 26462 12962 26514 12974
rect 22978 12910 22990 12962
rect 23042 12910 23054 12962
rect 20078 12898 20130 12910
rect 26462 12898 26514 12910
rect 32622 12962 32674 12974
rect 32622 12898 32674 12910
rect 33182 12962 33234 12974
rect 33182 12898 33234 12910
rect 33854 12962 33906 12974
rect 33854 12898 33906 12910
rect 34414 12962 34466 12974
rect 34414 12898 34466 12910
rect 34750 12962 34802 12974
rect 35758 12962 35810 12974
rect 35410 12910 35422 12962
rect 35474 12910 35486 12962
rect 34750 12898 34802 12910
rect 35758 12898 35810 12910
rect 35982 12962 36034 12974
rect 35982 12898 36034 12910
rect 37662 12962 37714 12974
rect 37662 12898 37714 12910
rect 38446 12962 38498 12974
rect 42366 12962 42418 12974
rect 39218 12910 39230 12962
rect 39282 12910 39294 12962
rect 38446 12898 38498 12910
rect 42366 12898 42418 12910
rect 43038 12962 43090 12974
rect 43038 12898 43090 12910
rect 1710 12850 1762 12862
rect 1710 12786 1762 12798
rect 2046 12850 2098 12862
rect 27806 12850 27858 12862
rect 17266 12798 17278 12850
rect 17330 12798 17342 12850
rect 2046 12786 2098 12798
rect 27806 12786 27858 12798
rect 28142 12850 28194 12862
rect 28142 12786 28194 12798
rect 29150 12850 29202 12862
rect 29150 12786 29202 12798
rect 29486 12850 29538 12862
rect 29486 12786 29538 12798
rect 37326 12850 37378 12862
rect 37326 12786 37378 12798
rect 42814 12850 42866 12862
rect 42814 12786 42866 12798
rect 2494 12738 2546 12750
rect 2494 12674 2546 12686
rect 20190 12738 20242 12750
rect 20190 12674 20242 12686
rect 20414 12738 20466 12750
rect 20414 12674 20466 12686
rect 26238 12738 26290 12750
rect 26238 12674 26290 12686
rect 26686 12738 26738 12750
rect 26686 12674 26738 12686
rect 32510 12738 32562 12750
rect 32510 12674 32562 12686
rect 33070 12738 33122 12750
rect 33070 12674 33122 12686
rect 33966 12738 34018 12750
rect 33966 12674 34018 12686
rect 34526 12738 34578 12750
rect 34526 12674 34578 12686
rect 37438 12738 37490 12750
rect 38770 12686 38782 12738
rect 38834 12686 38846 12738
rect 37438 12674 37490 12686
rect 1344 12570 78624 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 50558 12570
rect 50610 12518 50662 12570
rect 50714 12518 50766 12570
rect 50818 12518 78624 12570
rect 1344 12484 78624 12518
rect 19182 12402 19234 12414
rect 12562 12350 12574 12402
rect 12626 12350 12638 12402
rect 19182 12338 19234 12350
rect 19406 12402 19458 12414
rect 19406 12338 19458 12350
rect 20974 12402 21026 12414
rect 20974 12338 21026 12350
rect 25454 12402 25506 12414
rect 25454 12338 25506 12350
rect 28254 12402 28306 12414
rect 28254 12338 28306 12350
rect 33742 12402 33794 12414
rect 33742 12338 33794 12350
rect 36206 12402 36258 12414
rect 36206 12338 36258 12350
rect 37214 12402 37266 12414
rect 37214 12338 37266 12350
rect 41694 12402 41746 12414
rect 41694 12338 41746 12350
rect 42366 12402 42418 12414
rect 42366 12338 42418 12350
rect 74622 12402 74674 12414
rect 74622 12338 74674 12350
rect 75966 12402 76018 12414
rect 75966 12338 76018 12350
rect 77870 12402 77922 12414
rect 77870 12338 77922 12350
rect 17726 12290 17778 12302
rect 17726 12226 17778 12238
rect 20078 12290 20130 12302
rect 20078 12226 20130 12238
rect 20302 12290 20354 12302
rect 20302 12226 20354 12238
rect 36430 12290 36482 12302
rect 36430 12226 36482 12238
rect 36990 12290 37042 12302
rect 36990 12226 37042 12238
rect 19854 12178 19906 12190
rect 25230 12178 25282 12190
rect 9650 12126 9662 12178
rect 9714 12126 9726 12178
rect 21746 12126 21758 12178
rect 21810 12126 21822 12178
rect 19854 12114 19906 12126
rect 25230 12114 25282 12126
rect 25902 12178 25954 12190
rect 25902 12114 25954 12126
rect 27918 12178 27970 12190
rect 36542 12178 36594 12190
rect 29250 12126 29262 12178
rect 29314 12126 29326 12178
rect 33954 12126 33966 12178
rect 34018 12126 34030 12178
rect 27918 12114 27970 12126
rect 36542 12114 36594 12126
rect 36878 12178 36930 12190
rect 41582 12178 41634 12190
rect 37538 12126 37550 12178
rect 37602 12126 37614 12178
rect 36878 12114 36930 12126
rect 41582 12114 41634 12126
rect 74958 12178 75010 12190
rect 74958 12114 75010 12126
rect 75182 12178 75234 12190
rect 75182 12114 75234 12126
rect 78206 12178 78258 12190
rect 78206 12114 78258 12126
rect 17950 12066 18002 12078
rect 10322 12014 10334 12066
rect 10386 12014 10398 12066
rect 17602 12014 17614 12066
rect 17666 12014 17678 12066
rect 17950 12002 18002 12014
rect 19294 12066 19346 12078
rect 25342 12066 25394 12078
rect 41022 12066 41074 12078
rect 20402 12014 20414 12066
rect 20466 12014 20478 12066
rect 22418 12014 22430 12066
rect 22482 12014 22494 12066
rect 24546 12014 24558 12066
rect 24610 12014 24622 12066
rect 29922 12014 29934 12066
rect 29986 12014 29998 12066
rect 32050 12014 32062 12066
rect 32114 12014 32126 12066
rect 38210 12014 38222 12066
rect 38274 12014 38286 12066
rect 40338 12014 40350 12066
rect 40402 12014 40414 12066
rect 19294 12002 19346 12014
rect 25342 12002 25394 12014
rect 41022 12002 41074 12014
rect 77646 12066 77698 12078
rect 77646 12002 77698 12014
rect 40910 11954 40962 11966
rect 75506 11902 75518 11954
rect 75570 11902 75582 11954
rect 40910 11890 40962 11902
rect 1344 11786 78624 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 65918 11786
rect 65970 11734 66022 11786
rect 66074 11734 66126 11786
rect 66178 11734 78624 11786
rect 1344 11700 78624 11734
rect 22430 11618 22482 11630
rect 22430 11554 22482 11566
rect 37998 11618 38050 11630
rect 37998 11554 38050 11566
rect 9438 11506 9490 11518
rect 9438 11442 9490 11454
rect 12462 11506 12514 11518
rect 20638 11506 20690 11518
rect 13458 11454 13470 11506
rect 13522 11454 13534 11506
rect 18386 11454 18398 11506
rect 18450 11454 18462 11506
rect 12462 11442 12514 11454
rect 20638 11442 20690 11454
rect 22318 11506 22370 11518
rect 29934 11506 29986 11518
rect 28242 11454 28254 11506
rect 28306 11454 28318 11506
rect 35970 11454 35982 11506
rect 36034 11454 36046 11506
rect 22318 11442 22370 11454
rect 29934 11442 29986 11454
rect 11678 11394 11730 11406
rect 19630 11394 19682 11406
rect 9202 11342 9214 11394
rect 9266 11342 9278 11394
rect 15362 11342 15374 11394
rect 15426 11342 15438 11394
rect 11678 11330 11730 11342
rect 19630 11330 19682 11342
rect 19854 11394 19906 11406
rect 31502 11394 31554 11406
rect 20178 11342 20190 11394
rect 20242 11342 20254 11394
rect 22082 11342 22094 11394
rect 22146 11342 22158 11394
rect 25330 11342 25342 11394
rect 25394 11342 25406 11394
rect 19854 11330 19906 11342
rect 31502 11330 31554 11342
rect 31950 11394 32002 11406
rect 31950 11330 32002 11342
rect 32398 11394 32450 11406
rect 36990 11394 37042 11406
rect 33170 11342 33182 11394
rect 33234 11342 33246 11394
rect 38770 11342 38782 11394
rect 38834 11342 38846 11394
rect 76402 11342 76414 11394
rect 76466 11342 76478 11394
rect 32398 11330 32450 11342
rect 36990 11330 37042 11342
rect 1710 11282 1762 11294
rect 1710 11218 1762 11230
rect 2046 11282 2098 11294
rect 2046 11218 2098 11230
rect 9550 11282 9602 11294
rect 9550 11218 9602 11230
rect 11566 11282 11618 11294
rect 11566 11218 11618 11230
rect 13806 11282 13858 11294
rect 24894 11282 24946 11294
rect 16146 11230 16158 11282
rect 16210 11230 16222 11282
rect 13806 11218 13858 11230
rect 24894 11218 24946 11230
rect 25006 11282 25058 11294
rect 30046 11282 30098 11294
rect 26114 11230 26126 11282
rect 26178 11230 26190 11282
rect 25006 11218 25058 11230
rect 30046 11218 30098 11230
rect 31390 11282 31442 11294
rect 31390 11218 31442 11230
rect 32622 11282 32674 11294
rect 37326 11282 37378 11294
rect 33842 11230 33854 11282
rect 33906 11230 33918 11282
rect 32622 11218 32674 11230
rect 37326 11218 37378 11230
rect 37886 11282 37938 11294
rect 44830 11282 44882 11294
rect 77870 11282 77922 11294
rect 41458 11230 41470 11282
rect 41522 11230 41534 11282
rect 45154 11230 45166 11282
rect 45218 11230 45230 11282
rect 37886 11218 37938 11230
rect 44830 11218 44882 11230
rect 77870 11218 77922 11230
rect 78206 11282 78258 11294
rect 78206 11218 78258 11230
rect 2494 11170 2546 11182
rect 2494 11106 2546 11118
rect 11454 11170 11506 11182
rect 11454 11106 11506 11118
rect 11902 11170 11954 11182
rect 11902 11106 11954 11118
rect 13582 11170 13634 11182
rect 13582 11106 13634 11118
rect 19742 11170 19794 11182
rect 19742 11106 19794 11118
rect 24782 11170 24834 11182
rect 24782 11106 24834 11118
rect 29822 11170 29874 11182
rect 29822 11106 29874 11118
rect 31278 11170 31330 11182
rect 31278 11106 31330 11118
rect 32174 11170 32226 11182
rect 32174 11106 32226 11118
rect 32286 11170 32338 11182
rect 32286 11106 32338 11118
rect 36430 11170 36482 11182
rect 36430 11106 36482 11118
rect 37998 11170 38050 11182
rect 37998 11106 38050 11118
rect 76190 11170 76242 11182
rect 76190 11106 76242 11118
rect 77198 11170 77250 11182
rect 77198 11106 77250 11118
rect 77646 11170 77698 11182
rect 77646 11106 77698 11118
rect 1344 11002 78624 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 50558 11002
rect 50610 10950 50662 11002
rect 50714 10950 50766 11002
rect 50818 10950 78624 11002
rect 1344 10916 78624 10950
rect 11118 10834 11170 10846
rect 11118 10770 11170 10782
rect 11566 10834 11618 10846
rect 24110 10834 24162 10846
rect 21746 10782 21758 10834
rect 21810 10782 21822 10834
rect 11566 10770 11618 10782
rect 24110 10770 24162 10782
rect 24334 10834 24386 10846
rect 24334 10770 24386 10782
rect 25678 10834 25730 10846
rect 25678 10770 25730 10782
rect 25790 10834 25842 10846
rect 25790 10770 25842 10782
rect 25902 10834 25954 10846
rect 25902 10770 25954 10782
rect 26798 10834 26850 10846
rect 26798 10770 26850 10782
rect 31502 10834 31554 10846
rect 31502 10770 31554 10782
rect 32510 10834 32562 10846
rect 32510 10770 32562 10782
rect 39566 10834 39618 10846
rect 39566 10770 39618 10782
rect 39678 10834 39730 10846
rect 39678 10770 39730 10782
rect 39790 10834 39842 10846
rect 39790 10770 39842 10782
rect 40350 10834 40402 10846
rect 40350 10770 40402 10782
rect 2046 10722 2098 10734
rect 18174 10722 18226 10734
rect 13346 10670 13358 10722
rect 13410 10670 13422 10722
rect 2046 10658 2098 10670
rect 18174 10658 18226 10670
rect 18398 10722 18450 10734
rect 38782 10722 38834 10734
rect 33282 10670 33294 10722
rect 33346 10670 33358 10722
rect 18398 10658 18450 10670
rect 38782 10658 38834 10670
rect 39006 10722 39058 10734
rect 39006 10658 39058 10670
rect 1710 10610 1762 10622
rect 1710 10546 1762 10558
rect 11342 10610 11394 10622
rect 24782 10610 24834 10622
rect 31278 10610 31330 10622
rect 11890 10558 11902 10610
rect 11954 10558 11966 10610
rect 12674 10558 12686 10610
rect 12738 10558 12750 10610
rect 18834 10558 18846 10610
rect 18898 10558 18910 10610
rect 22194 10558 22206 10610
rect 22258 10558 22270 10610
rect 26226 10558 26238 10610
rect 26290 10558 26302 10610
rect 28130 10558 28142 10610
rect 28194 10558 28206 10610
rect 11342 10546 11394 10558
rect 24782 10546 24834 10558
rect 31278 10546 31330 10558
rect 31950 10610 32002 10622
rect 38670 10610 38722 10622
rect 38322 10558 38334 10610
rect 38386 10558 38398 10610
rect 31950 10546 32002 10558
rect 38670 10546 38722 10558
rect 39118 10610 39170 10622
rect 41458 10558 41470 10610
rect 41522 10558 41534 10610
rect 78194 10558 78206 10610
rect 78258 10558 78270 10610
rect 39118 10546 39170 10558
rect 2494 10498 2546 10510
rect 2494 10434 2546 10446
rect 11454 10498 11506 10510
rect 11454 10434 11506 10446
rect 15486 10498 15538 10510
rect 15486 10434 15538 10446
rect 18286 10498 18338 10510
rect 22542 10498 22594 10510
rect 19506 10446 19518 10498
rect 19570 10446 19582 10498
rect 22306 10446 22318 10498
rect 22370 10446 22382 10498
rect 18286 10434 18338 10446
rect 22542 10434 22594 10446
rect 24222 10498 24274 10510
rect 24222 10434 24274 10446
rect 27806 10498 27858 10510
rect 31390 10498 31442 10510
rect 28802 10446 28814 10498
rect 28866 10446 28878 10498
rect 30930 10446 30942 10498
rect 30994 10446 31006 10498
rect 42130 10446 42142 10498
rect 42194 10446 42206 10498
rect 44258 10446 44270 10498
rect 44322 10446 44334 10498
rect 27806 10434 27858 10446
rect 31390 10434 31442 10446
rect 75854 10386 75906 10398
rect 75854 10322 75906 10334
rect 1344 10218 78624 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 65918 10218
rect 65970 10166 66022 10218
rect 66074 10166 66126 10218
rect 66178 10166 78624 10218
rect 1344 10132 78624 10166
rect 8206 10050 8258 10062
rect 8206 9986 8258 9998
rect 29150 10050 29202 10062
rect 29150 9986 29202 9998
rect 29486 10050 29538 10062
rect 33070 10050 33122 10062
rect 30258 9998 30270 10050
rect 30322 10047 30334 10050
rect 31378 10047 31390 10050
rect 30322 10001 31390 10047
rect 30322 9998 30334 10001
rect 31378 9998 31390 10001
rect 31442 9998 31454 10050
rect 32386 9998 32398 10050
rect 32450 10047 32462 10050
rect 32834 10047 32846 10050
rect 32450 10001 32846 10047
rect 32450 9998 32462 10001
rect 32834 9998 32846 10001
rect 32898 9998 32910 10050
rect 29486 9986 29538 9998
rect 33070 9986 33122 9998
rect 35198 10050 35250 10062
rect 35198 9986 35250 9998
rect 13582 9938 13634 9950
rect 11554 9886 11566 9938
rect 11618 9886 11630 9938
rect 13582 9874 13634 9886
rect 14478 9938 14530 9950
rect 20750 9938 20802 9950
rect 15362 9886 15374 9938
rect 15426 9886 15438 9938
rect 14478 9874 14530 9886
rect 20750 9874 20802 9886
rect 31726 9938 31778 9950
rect 31726 9874 31778 9886
rect 33182 9938 33234 9950
rect 33182 9874 33234 9886
rect 34862 9938 34914 9950
rect 34862 9874 34914 9886
rect 41806 9938 41858 9950
rect 41806 9874 41858 9886
rect 42478 9938 42530 9950
rect 42478 9874 42530 9886
rect 76302 9938 76354 9950
rect 76302 9874 76354 9886
rect 12238 9826 12290 9838
rect 31838 9826 31890 9838
rect 8642 9774 8654 9826
rect 8706 9774 8718 9826
rect 12562 9774 12574 9826
rect 12626 9774 12638 9826
rect 14018 9774 14030 9826
rect 14082 9774 14094 9826
rect 20178 9774 20190 9826
rect 20242 9774 20254 9826
rect 22754 9774 22766 9826
rect 22818 9774 22830 9826
rect 12238 9762 12290 9774
rect 31838 9762 31890 9774
rect 32286 9826 32338 9838
rect 32286 9762 32338 9774
rect 35086 9826 35138 9838
rect 35086 9762 35138 9774
rect 36990 9826 37042 9838
rect 36990 9762 37042 9774
rect 37662 9826 37714 9838
rect 37662 9762 37714 9774
rect 38222 9826 38274 9838
rect 38222 9762 38274 9774
rect 38782 9826 38834 9838
rect 38782 9762 38834 9774
rect 42366 9826 42418 9838
rect 42366 9762 42418 9774
rect 42590 9826 42642 9838
rect 42590 9762 42642 9774
rect 42926 9826 42978 9838
rect 42926 9762 42978 9774
rect 1710 9714 1762 9726
rect 1710 9650 1762 9662
rect 2046 9714 2098 9726
rect 2046 9650 2098 9662
rect 8094 9714 8146 9726
rect 13694 9714 13746 9726
rect 37326 9714 37378 9726
rect 9314 9662 9326 9714
rect 9378 9662 9390 9714
rect 23538 9662 23550 9714
rect 23602 9662 23614 9714
rect 26898 9662 26910 9714
rect 26962 9662 26974 9714
rect 33730 9662 33742 9714
rect 33794 9662 33806 9714
rect 8094 9650 8146 9662
rect 13694 9650 13746 9662
rect 37326 9650 37378 9662
rect 39454 9714 39506 9726
rect 39454 9650 39506 9662
rect 40798 9714 40850 9726
rect 40798 9650 40850 9662
rect 77646 9714 77698 9726
rect 77646 9650 77698 9662
rect 77870 9714 77922 9726
rect 77870 9650 77922 9662
rect 78206 9714 78258 9726
rect 78206 9650 78258 9662
rect 2494 9602 2546 9614
rect 2494 9538 2546 9550
rect 7982 9602 8034 9614
rect 7982 9538 8034 9550
rect 12014 9602 12066 9614
rect 12014 9538 12066 9550
rect 12126 9602 12178 9614
rect 12126 9538 12178 9550
rect 13470 9602 13522 9614
rect 13470 9538 13522 9550
rect 27246 9602 27298 9614
rect 27246 9538 27298 9550
rect 27806 9602 27858 9614
rect 27806 9538 27858 9550
rect 28254 9602 28306 9614
rect 28254 9538 28306 9550
rect 28702 9602 28754 9614
rect 28702 9538 28754 9550
rect 29262 9602 29314 9614
rect 29262 9538 29314 9550
rect 30046 9602 30098 9614
rect 30046 9538 30098 9550
rect 30494 9602 30546 9614
rect 30494 9538 30546 9550
rect 30942 9602 30994 9614
rect 30942 9538 30994 9550
rect 31278 9602 31330 9614
rect 31278 9538 31330 9550
rect 31614 9602 31666 9614
rect 31614 9538 31666 9550
rect 32846 9602 32898 9614
rect 32846 9538 32898 9550
rect 33294 9602 33346 9614
rect 33294 9538 33346 9550
rect 34078 9602 34130 9614
rect 34078 9538 34130 9550
rect 37774 9602 37826 9614
rect 37774 9538 37826 9550
rect 37998 9602 38050 9614
rect 37998 9538 38050 9550
rect 38334 9602 38386 9614
rect 38334 9538 38386 9550
rect 38558 9602 38610 9614
rect 38558 9538 38610 9550
rect 38894 9602 38946 9614
rect 38894 9538 38946 9550
rect 39118 9602 39170 9614
rect 39118 9538 39170 9550
rect 40014 9602 40066 9614
rect 40014 9538 40066 9550
rect 40910 9602 40962 9614
rect 40910 9538 40962 9550
rect 42142 9602 42194 9614
rect 42142 9538 42194 9550
rect 43038 9602 43090 9614
rect 43038 9538 43090 9550
rect 43150 9602 43202 9614
rect 43150 9538 43202 9550
rect 43374 9602 43426 9614
rect 43374 9538 43426 9550
rect 43934 9602 43986 9614
rect 43934 9538 43986 9550
rect 74846 9602 74898 9614
rect 74846 9538 74898 9550
rect 75294 9602 75346 9614
rect 75294 9538 75346 9550
rect 75630 9602 75682 9614
rect 75630 9538 75682 9550
rect 77198 9602 77250 9614
rect 77198 9538 77250 9550
rect 1344 9434 78624 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 50558 9434
rect 50610 9382 50662 9434
rect 50714 9382 50766 9434
rect 50818 9382 78624 9434
rect 1344 9348 78624 9382
rect 13806 9266 13858 9278
rect 14478 9266 14530 9278
rect 13458 9214 13470 9266
rect 13522 9214 13534 9266
rect 14130 9214 14142 9266
rect 14194 9214 14206 9266
rect 13806 9202 13858 9214
rect 14478 9202 14530 9214
rect 14926 9266 14978 9278
rect 14926 9202 14978 9214
rect 16158 9266 16210 9278
rect 16158 9202 16210 9214
rect 18286 9266 18338 9278
rect 18286 9202 18338 9214
rect 19182 9266 19234 9278
rect 24670 9266 24722 9278
rect 22530 9214 22542 9266
rect 22594 9214 22606 9266
rect 25218 9214 25230 9266
rect 25282 9214 25294 9266
rect 19182 9202 19234 9214
rect 24670 9202 24722 9214
rect 8766 9154 8818 9166
rect 8766 9090 8818 9102
rect 15374 9154 15426 9166
rect 42578 9102 42590 9154
rect 42642 9102 42654 9154
rect 15374 9090 15426 9102
rect 18062 9042 18114 9054
rect 9650 8990 9662 9042
rect 9714 8990 9726 9042
rect 15922 8990 15934 9042
rect 15986 8990 15998 9042
rect 18062 8978 18114 8990
rect 18734 9042 18786 9054
rect 41470 9042 41522 9054
rect 19506 8990 19518 9042
rect 19570 8990 19582 9042
rect 25442 8990 25454 9042
rect 25506 8990 25518 9042
rect 26114 8990 26126 9042
rect 26178 8990 26190 9042
rect 29362 8990 29374 9042
rect 29426 8990 29438 9042
rect 33282 8990 33294 9042
rect 33346 8990 33358 9042
rect 33954 8990 33966 9042
rect 34018 8990 34030 9042
rect 37538 8990 37550 9042
rect 37602 8990 37614 9042
rect 41794 8990 41806 9042
rect 41858 8990 41870 9042
rect 75170 8990 75182 9042
rect 75234 8990 75246 9042
rect 76066 8990 76078 9042
rect 76130 8990 76142 9042
rect 18734 8978 18786 8990
rect 41470 8978 41522 8990
rect 8878 8930 8930 8942
rect 12462 8930 12514 8942
rect 10322 8878 10334 8930
rect 10386 8878 10398 8930
rect 8878 8866 8930 8878
rect 12462 8866 12514 8878
rect 13246 8930 13298 8942
rect 16270 8930 16322 8942
rect 15362 8878 15374 8930
rect 15426 8878 15438 8930
rect 13246 8866 13298 8878
rect 16270 8866 16322 8878
rect 17726 8930 17778 8942
rect 17726 8866 17778 8878
rect 18174 8930 18226 8942
rect 23438 8930 23490 8942
rect 20290 8878 20302 8930
rect 20354 8878 20366 8930
rect 18174 8866 18226 8878
rect 23438 8866 23490 8878
rect 23886 8930 23938 8942
rect 23886 8866 23938 8878
rect 24334 8930 24386 8942
rect 33518 8930 33570 8942
rect 45054 8930 45106 8942
rect 26898 8878 26910 8930
rect 26962 8878 26974 8930
rect 29026 8878 29038 8930
rect 29090 8878 29102 8930
rect 30146 8878 30158 8930
rect 30210 8878 30222 8930
rect 32274 8878 32286 8930
rect 32338 8878 32350 8930
rect 34738 8878 34750 8930
rect 34802 8878 34814 8930
rect 36866 8878 36878 8930
rect 36930 8878 36942 8930
rect 38210 8878 38222 8930
rect 38274 8878 38286 8930
rect 40338 8878 40350 8930
rect 40402 8878 40414 8930
rect 41010 8878 41022 8930
rect 41074 8878 41086 8930
rect 44706 8878 44718 8930
rect 44770 8878 44782 8930
rect 45266 8878 45278 8930
rect 45330 8878 45342 8930
rect 77858 8878 77870 8930
rect 77922 8878 77934 8930
rect 24334 8866 24386 8878
rect 33518 8866 33570 8878
rect 45054 8866 45106 8878
rect 8990 8818 9042 8830
rect 8990 8754 9042 8766
rect 15598 8818 15650 8830
rect 15598 8754 15650 8766
rect 33630 8818 33682 8830
rect 73826 8766 73838 8818
rect 73890 8766 73902 8818
rect 33630 8754 33682 8766
rect 1344 8650 78624 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 65918 8650
rect 65970 8598 66022 8650
rect 66074 8598 66126 8650
rect 66178 8598 78624 8650
rect 1344 8564 78624 8598
rect 19294 8482 19346 8494
rect 19294 8418 19346 8430
rect 28142 8482 28194 8494
rect 28142 8418 28194 8430
rect 30270 8482 30322 8494
rect 30270 8418 30322 8430
rect 41694 8482 41746 8494
rect 41694 8418 41746 8430
rect 18174 8370 18226 8382
rect 19854 8370 19906 8382
rect 15362 8318 15374 8370
rect 15426 8318 15438 8370
rect 17602 8318 17614 8370
rect 17666 8318 17678 8370
rect 19058 8318 19070 8370
rect 19122 8318 19134 8370
rect 18174 8306 18226 8318
rect 19854 8306 19906 8318
rect 20750 8370 20802 8382
rect 26910 8370 26962 8382
rect 22418 8318 22430 8370
rect 22482 8318 22494 8370
rect 24546 8318 24558 8370
rect 24610 8318 24622 8370
rect 20750 8306 20802 8318
rect 26910 8306 26962 8318
rect 27358 8370 27410 8382
rect 30158 8370 30210 8382
rect 27570 8318 27582 8370
rect 27634 8318 27646 8370
rect 27358 8306 27410 8318
rect 30158 8306 30210 8318
rect 32286 8370 32338 8382
rect 32286 8306 32338 8318
rect 34190 8370 34242 8382
rect 34190 8306 34242 8318
rect 18286 8258 18338 8270
rect 9762 8206 9774 8258
rect 9826 8206 9838 8258
rect 14018 8206 14030 8258
rect 14082 8206 14094 8258
rect 14690 8206 14702 8258
rect 14754 8206 14766 8258
rect 18286 8194 18338 8206
rect 18734 8258 18786 8270
rect 18734 8194 18786 8206
rect 19966 8258 20018 8270
rect 19966 8194 20018 8206
rect 20414 8258 20466 8270
rect 26350 8258 26402 8270
rect 21634 8206 21646 8258
rect 21698 8206 21710 8258
rect 20414 8194 20466 8206
rect 26350 8194 26402 8206
rect 26798 8258 26850 8270
rect 26798 8194 26850 8206
rect 29038 8258 29090 8270
rect 29038 8194 29090 8206
rect 32622 8258 32674 8270
rect 32622 8194 32674 8206
rect 34302 8258 34354 8270
rect 38670 8258 38722 8270
rect 34626 8206 34638 8258
rect 34690 8206 34702 8258
rect 35298 8206 35310 8258
rect 35362 8206 35374 8258
rect 38098 8206 38110 8258
rect 38162 8206 38174 8258
rect 34302 8194 34354 8206
rect 38670 8194 38722 8206
rect 39566 8258 39618 8270
rect 40798 8258 40850 8270
rect 44718 8258 44770 8270
rect 78206 8258 78258 8270
rect 39890 8206 39902 8258
rect 39954 8206 39966 8258
rect 41346 8206 41358 8258
rect 41410 8206 41422 8258
rect 42466 8206 42478 8258
rect 42530 8206 42542 8258
rect 43026 8206 43038 8258
rect 43090 8206 43102 8258
rect 75282 8206 75294 8258
rect 75346 8206 75358 8258
rect 39566 8194 39618 8206
rect 40798 8194 40850 8206
rect 44718 8194 44770 8206
rect 78206 8194 78258 8206
rect 1710 8146 1762 8158
rect 1710 8082 1762 8094
rect 2046 8146 2098 8158
rect 19742 8146 19794 8158
rect 10546 8094 10558 8146
rect 10610 8094 10622 8146
rect 14242 8094 14254 8146
rect 14306 8094 14318 8146
rect 2046 8082 2098 8094
rect 19742 8082 19794 8094
rect 28254 8146 28306 8158
rect 28254 8082 28306 8094
rect 29262 8146 29314 8158
rect 29262 8082 29314 8094
rect 29374 8146 29426 8158
rect 34974 8146 35026 8158
rect 31490 8094 31502 8146
rect 31554 8094 31566 8146
rect 29374 8082 29426 8094
rect 34974 8082 35026 8094
rect 39118 8146 39170 8158
rect 39118 8082 39170 8094
rect 40910 8146 40962 8158
rect 40910 8082 40962 8094
rect 41022 8146 41074 8158
rect 44046 8146 44098 8158
rect 42354 8094 42366 8146
rect 42418 8094 42430 8146
rect 43698 8094 43710 8146
rect 43762 8094 43774 8146
rect 41022 8082 41074 8094
rect 44046 8082 44098 8094
rect 45054 8146 45106 8158
rect 45054 8082 45106 8094
rect 76862 8146 76914 8158
rect 76862 8082 76914 8094
rect 77198 8146 77250 8158
rect 77198 8082 77250 8094
rect 77534 8146 77586 8158
rect 77534 8082 77586 8094
rect 77870 8146 77922 8158
rect 77870 8082 77922 8094
rect 2494 8034 2546 8046
rect 13694 8034 13746 8046
rect 12786 7982 12798 8034
rect 12850 7982 12862 8034
rect 2494 7970 2546 7982
rect 13694 7970 13746 7982
rect 18062 8034 18114 8046
rect 18062 7970 18114 7982
rect 19070 8034 19122 8046
rect 19070 7970 19122 7982
rect 25342 8034 25394 8046
rect 25342 7970 25394 7982
rect 25790 8034 25842 8046
rect 25790 7970 25842 7982
rect 26238 8034 26290 8046
rect 26238 7970 26290 7982
rect 27022 8034 27074 8046
rect 27022 7970 27074 7982
rect 27582 8034 27634 8046
rect 27582 7970 27634 7982
rect 28142 8034 28194 8046
rect 28142 7970 28194 7982
rect 30046 8034 30098 8046
rect 30046 7970 30098 7982
rect 30830 8034 30882 8046
rect 30830 7970 30882 7982
rect 31278 8034 31330 8046
rect 31278 7970 31330 7982
rect 31838 8034 31890 8046
rect 33518 8034 33570 8046
rect 32946 7982 32958 8034
rect 33010 7982 33022 8034
rect 31838 7970 31890 7982
rect 33518 7970 33570 7982
rect 34078 8034 34130 8046
rect 34078 7970 34130 7982
rect 35086 8034 35138 8046
rect 35086 7970 35138 7982
rect 35870 8034 35922 8046
rect 35870 7970 35922 7982
rect 37102 8034 37154 8046
rect 37102 7970 37154 7982
rect 37662 8034 37714 8046
rect 37662 7970 37714 7982
rect 37886 8034 37938 8046
rect 37886 7970 37938 7982
rect 38782 8034 38834 8046
rect 38782 7970 38834 7982
rect 38894 8034 38946 8046
rect 38894 7970 38946 7982
rect 39678 8034 39730 8046
rect 44942 8034 44994 8046
rect 42914 7982 42926 8034
rect 42978 7982 42990 8034
rect 39678 7970 39730 7982
rect 44942 7970 44994 7982
rect 45502 8034 45554 8046
rect 45502 7970 45554 7982
rect 45950 8034 46002 8046
rect 45950 7970 46002 7982
rect 74622 8034 74674 8046
rect 74622 7970 74674 7982
rect 76526 8034 76578 8046
rect 76526 7970 76578 7982
rect 1344 7866 78624 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 50558 7866
rect 50610 7814 50662 7866
rect 50714 7814 50766 7866
rect 50818 7814 78624 7866
rect 1344 7780 78624 7814
rect 2046 7698 2098 7710
rect 2046 7634 2098 7646
rect 8542 7698 8594 7710
rect 8542 7634 8594 7646
rect 13134 7698 13186 7710
rect 13134 7634 13186 7646
rect 13582 7698 13634 7710
rect 13582 7634 13634 7646
rect 16942 7698 16994 7710
rect 16942 7634 16994 7646
rect 18622 7698 18674 7710
rect 18622 7634 18674 7646
rect 18846 7698 18898 7710
rect 20414 7698 20466 7710
rect 19282 7646 19294 7698
rect 19346 7646 19358 7698
rect 20066 7646 20078 7698
rect 20130 7646 20142 7698
rect 18846 7634 18898 7646
rect 20414 7634 20466 7646
rect 20862 7698 20914 7710
rect 20862 7634 20914 7646
rect 23102 7698 23154 7710
rect 23102 7634 23154 7646
rect 24782 7698 24834 7710
rect 24782 7634 24834 7646
rect 25678 7698 25730 7710
rect 25678 7634 25730 7646
rect 25902 7698 25954 7710
rect 25902 7634 25954 7646
rect 27806 7698 27858 7710
rect 30046 7698 30098 7710
rect 28354 7646 28366 7698
rect 28418 7646 28430 7698
rect 29250 7646 29262 7698
rect 29314 7646 29326 7698
rect 27806 7634 27858 7646
rect 30046 7634 30098 7646
rect 30270 7698 30322 7710
rect 30270 7634 30322 7646
rect 31726 7698 31778 7710
rect 31726 7634 31778 7646
rect 33966 7698 34018 7710
rect 33966 7634 34018 7646
rect 38110 7698 38162 7710
rect 71710 7698 71762 7710
rect 39666 7646 39678 7698
rect 39730 7646 39742 7698
rect 42018 7646 42030 7698
rect 42082 7646 42094 7698
rect 38110 7634 38162 7646
rect 71710 7634 71762 7646
rect 11006 7586 11058 7598
rect 15598 7586 15650 7598
rect 18398 7586 18450 7598
rect 30382 7586 30434 7598
rect 14242 7534 14254 7586
rect 14306 7534 14318 7586
rect 18050 7534 18062 7586
rect 18114 7534 18126 7586
rect 26562 7534 26574 7586
rect 26626 7534 26638 7586
rect 11006 7522 11058 7534
rect 15598 7522 15650 7534
rect 18398 7522 18450 7534
rect 30382 7522 30434 7534
rect 31054 7586 31106 7598
rect 33854 7586 33906 7598
rect 43038 7586 43090 7598
rect 32498 7534 32510 7586
rect 32562 7534 32574 7586
rect 35186 7534 35198 7586
rect 35250 7534 35262 7586
rect 38658 7534 38670 7586
rect 38722 7534 38734 7586
rect 39218 7534 39230 7586
rect 39282 7534 39294 7586
rect 40898 7534 40910 7586
rect 40962 7534 40974 7586
rect 31054 7522 31106 7534
rect 33854 7522 33906 7534
rect 43038 7522 43090 7534
rect 44494 7586 44546 7598
rect 44494 7522 44546 7534
rect 66670 7586 66722 7598
rect 66670 7522 66722 7534
rect 1710 7474 1762 7486
rect 13358 7474 13410 7486
rect 17726 7474 17778 7486
rect 8306 7422 8318 7474
rect 8370 7422 8382 7474
rect 13906 7422 13918 7474
rect 13970 7422 13982 7474
rect 14466 7422 14478 7474
rect 14530 7422 14542 7474
rect 1710 7410 1762 7422
rect 13358 7410 13410 7422
rect 17726 7410 17778 7422
rect 19630 7474 19682 7486
rect 25342 7474 25394 7486
rect 23426 7422 23438 7474
rect 23490 7422 23502 7474
rect 19630 7410 19682 7422
rect 25342 7410 25394 7422
rect 26350 7474 26402 7486
rect 26350 7410 26402 7422
rect 26910 7474 26962 7486
rect 26910 7410 26962 7422
rect 28926 7474 28978 7486
rect 28926 7410 28978 7422
rect 29822 7474 29874 7486
rect 29822 7410 29874 7422
rect 30718 7474 30770 7486
rect 30718 7410 30770 7422
rect 32174 7474 32226 7486
rect 32174 7410 32226 7422
rect 33406 7474 33458 7486
rect 33406 7410 33458 7422
rect 34078 7474 34130 7486
rect 40014 7474 40066 7486
rect 34402 7422 34414 7474
rect 34466 7422 34478 7474
rect 41234 7422 41246 7474
rect 41298 7422 41310 7474
rect 41906 7422 41918 7474
rect 41970 7422 41982 7474
rect 43922 7422 43934 7474
rect 43986 7422 43998 7474
rect 46498 7422 46510 7474
rect 46562 7422 46574 7474
rect 66994 7422 67006 7474
rect 67058 7422 67070 7474
rect 72370 7422 72382 7474
rect 72434 7422 72446 7474
rect 75282 7422 75294 7474
rect 75346 7422 75358 7474
rect 34078 7410 34130 7422
rect 40014 7410 40066 7422
rect 2494 7362 2546 7374
rect 2494 7298 2546 7310
rect 10222 7362 10274 7374
rect 11230 7362 11282 7374
rect 10882 7310 10894 7362
rect 10946 7310 10958 7362
rect 10222 7298 10274 7310
rect 11230 7298 11282 7310
rect 11790 7362 11842 7374
rect 11790 7298 11842 7310
rect 12686 7362 12738 7374
rect 12686 7298 12738 7310
rect 13470 7362 13522 7374
rect 13470 7298 13522 7310
rect 15262 7362 15314 7374
rect 15262 7298 15314 7310
rect 15710 7362 15762 7374
rect 15710 7298 15762 7310
rect 15822 7362 15874 7374
rect 15822 7298 15874 7310
rect 16494 7362 16546 7374
rect 16494 7298 16546 7310
rect 18510 7362 18562 7374
rect 18510 7298 18562 7310
rect 21422 7362 21474 7374
rect 21422 7298 21474 7310
rect 21870 7362 21922 7374
rect 21870 7298 21922 7310
rect 22318 7362 22370 7374
rect 22318 7298 22370 7310
rect 22766 7362 22818 7374
rect 22766 7298 22818 7310
rect 23774 7362 23826 7374
rect 23774 7298 23826 7310
rect 24334 7362 24386 7374
rect 24334 7298 24386 7310
rect 25790 7362 25842 7374
rect 25790 7298 25842 7310
rect 27470 7362 27522 7374
rect 33294 7362 33346 7374
rect 47070 7362 47122 7374
rect 31826 7310 31838 7362
rect 31890 7310 31902 7362
rect 37314 7310 37326 7362
rect 37378 7310 37390 7362
rect 41570 7310 41582 7362
rect 41634 7310 41646 7362
rect 46162 7310 46174 7362
rect 46226 7310 46238 7362
rect 27470 7298 27522 7310
rect 33294 7298 33346 7310
rect 47070 7298 47122 7310
rect 47630 7362 47682 7374
rect 47630 7298 47682 7310
rect 60174 7362 60226 7374
rect 73938 7310 73950 7362
rect 74002 7310 74014 7362
rect 60174 7298 60226 7310
rect 8654 7250 8706 7262
rect 23438 7250 23490 7262
rect 21858 7198 21870 7250
rect 21922 7247 21934 7250
rect 22082 7247 22094 7250
rect 21922 7201 22094 7247
rect 21922 7198 21934 7201
rect 22082 7198 22094 7201
rect 22146 7198 22158 7250
rect 22418 7198 22430 7250
rect 22482 7247 22494 7250
rect 23202 7247 23214 7250
rect 22482 7201 23214 7247
rect 22482 7198 22494 7201
rect 23202 7198 23214 7201
rect 23266 7198 23278 7250
rect 8654 7186 8706 7198
rect 23438 7186 23490 7198
rect 28702 7250 28754 7262
rect 28702 7186 28754 7198
rect 29598 7250 29650 7262
rect 29598 7186 29650 7198
rect 31502 7250 31554 7262
rect 31502 7186 31554 7198
rect 38446 7250 38498 7262
rect 38446 7186 38498 7198
rect 68014 7250 68066 7262
rect 68014 7186 68066 7198
rect 76302 7250 76354 7262
rect 76302 7186 76354 7198
rect 1344 7082 78624 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 65918 7082
rect 65970 7030 66022 7082
rect 66074 7030 66126 7082
rect 66178 7030 78624 7082
rect 1344 6996 78624 7030
rect 8206 6914 8258 6926
rect 8206 6850 8258 6862
rect 8878 6914 8930 6926
rect 8878 6850 8930 6862
rect 9214 6914 9266 6926
rect 9214 6850 9266 6862
rect 8766 6802 8818 6814
rect 7970 6750 7982 6802
rect 8034 6750 8046 6802
rect 8766 6738 8818 6750
rect 9326 6802 9378 6814
rect 9326 6738 9378 6750
rect 13582 6802 13634 6814
rect 17838 6802 17890 6814
rect 26238 6802 26290 6814
rect 15698 6750 15710 6802
rect 15762 6750 15774 6802
rect 25554 6750 25566 6802
rect 25618 6750 25630 6802
rect 13582 6738 13634 6750
rect 17838 6738 17890 6750
rect 26238 6738 26290 6750
rect 28478 6802 28530 6814
rect 31838 6802 31890 6814
rect 31490 6750 31502 6802
rect 31554 6750 31566 6802
rect 28478 6738 28530 6750
rect 31838 6738 31890 6750
rect 32734 6802 32786 6814
rect 74734 6802 74786 6814
rect 36418 6750 36430 6802
rect 36482 6750 36494 6802
rect 37986 6750 37998 6802
rect 38050 6750 38062 6802
rect 40114 6750 40126 6802
rect 40178 6750 40190 6802
rect 32734 6738 32786 6750
rect 74734 6738 74786 6750
rect 76414 6802 76466 6814
rect 76414 6738 76466 6750
rect 78094 6802 78146 6814
rect 78094 6738 78146 6750
rect 12126 6690 12178 6702
rect 12126 6626 12178 6638
rect 13694 6690 13746 6702
rect 19966 6690 20018 6702
rect 14914 6638 14926 6690
rect 14978 6638 14990 6690
rect 13694 6626 13746 6638
rect 19966 6626 20018 6638
rect 21870 6690 21922 6702
rect 26126 6690 26178 6702
rect 22642 6638 22654 6690
rect 22706 6638 22718 6690
rect 23426 6638 23438 6690
rect 23490 6638 23502 6690
rect 21870 6626 21922 6638
rect 26126 6626 26178 6638
rect 26350 6690 26402 6702
rect 26350 6626 26402 6638
rect 26798 6690 26850 6702
rect 28254 6690 28306 6702
rect 30606 6690 30658 6702
rect 27234 6638 27246 6690
rect 27298 6638 27310 6690
rect 27906 6638 27918 6690
rect 27970 6638 27982 6690
rect 29362 6638 29374 6690
rect 29426 6638 29438 6690
rect 30034 6638 30046 6690
rect 30098 6638 30110 6690
rect 26798 6626 26850 6638
rect 28254 6626 28306 6638
rect 30606 6626 30658 6638
rect 30830 6690 30882 6702
rect 30830 6626 30882 6638
rect 32622 6690 32674 6702
rect 32622 6626 32674 6638
rect 32846 6690 32898 6702
rect 32846 6626 32898 6638
rect 33294 6690 33346 6702
rect 49982 6690 50034 6702
rect 51438 6690 51490 6702
rect 33618 6638 33630 6690
rect 33682 6638 33694 6690
rect 37314 6638 37326 6690
rect 37378 6638 37390 6690
rect 40450 6638 40462 6690
rect 40514 6638 40526 6690
rect 44258 6638 44270 6690
rect 44322 6638 44334 6690
rect 46610 6638 46622 6690
rect 46674 6638 46686 6690
rect 47058 6638 47070 6690
rect 47122 6638 47134 6690
rect 50978 6638 50990 6690
rect 51042 6638 51054 6690
rect 33294 6626 33346 6638
rect 49982 6626 50034 6638
rect 51438 6626 51490 6638
rect 59502 6690 59554 6702
rect 59502 6626 59554 6638
rect 60062 6690 60114 6702
rect 67902 6690 67954 6702
rect 74958 6690 75010 6702
rect 60498 6638 60510 6690
rect 60562 6638 60574 6690
rect 63410 6638 63422 6690
rect 63474 6638 63486 6690
rect 68338 6638 68350 6690
rect 68402 6638 68414 6690
rect 71250 6638 71262 6690
rect 71314 6638 71326 6690
rect 60062 6626 60114 6638
rect 67902 6626 67954 6638
rect 74958 6626 75010 6638
rect 75182 6690 75234 6702
rect 75182 6626 75234 6638
rect 76190 6690 76242 6702
rect 76190 6626 76242 6638
rect 77086 6690 77138 6702
rect 77086 6626 77138 6638
rect 77310 6690 77362 6702
rect 77310 6626 77362 6638
rect 9438 6578 9490 6590
rect 21534 6578 21586 6590
rect 30270 6578 30322 6590
rect 41582 6578 41634 6590
rect 19618 6526 19630 6578
rect 19682 6526 19694 6578
rect 22194 6526 22206 6578
rect 22258 6526 22270 6578
rect 27010 6526 27022 6578
rect 27074 6526 27086 6578
rect 31154 6526 31166 6578
rect 31218 6526 31230 6578
rect 34290 6526 34302 6578
rect 34354 6526 34366 6578
rect 9438 6514 9490 6526
rect 21534 6514 21586 6526
rect 30270 6514 30322 6526
rect 41582 6514 41634 6526
rect 43598 6578 43650 6590
rect 43598 6514 43650 6526
rect 46062 6578 46114 6590
rect 50542 6578 50594 6590
rect 48626 6526 48638 6578
rect 48690 6526 48702 6578
rect 46062 6514 46114 6526
rect 50542 6514 50594 6526
rect 6638 6466 6690 6478
rect 6638 6402 6690 6414
rect 7086 6466 7138 6478
rect 7086 6402 7138 6414
rect 7646 6466 7698 6478
rect 7646 6402 7698 6414
rect 7982 6466 8034 6478
rect 7982 6402 8034 6414
rect 8654 6466 8706 6478
rect 8654 6402 8706 6414
rect 10222 6466 10274 6478
rect 10222 6402 10274 6414
rect 10894 6466 10946 6478
rect 10894 6402 10946 6414
rect 11678 6466 11730 6478
rect 11678 6402 11730 6414
rect 12574 6466 12626 6478
rect 12574 6402 12626 6414
rect 13022 6466 13074 6478
rect 13022 6402 13074 6414
rect 13470 6466 13522 6478
rect 13470 6402 13522 6414
rect 13918 6466 13970 6478
rect 13918 6402 13970 6414
rect 14702 6466 14754 6478
rect 14702 6402 14754 6414
rect 18958 6466 19010 6478
rect 18958 6402 19010 6414
rect 19406 6466 19458 6478
rect 19406 6402 19458 6414
rect 20862 6466 20914 6478
rect 31614 6466 31666 6478
rect 29586 6414 29598 6466
rect 29650 6414 29662 6466
rect 20862 6402 20914 6414
rect 31614 6402 31666 6414
rect 32398 6466 32450 6478
rect 49086 6466 49138 6478
rect 40674 6414 40686 6466
rect 40738 6414 40750 6466
rect 47058 6414 47070 6466
rect 47122 6414 47134 6466
rect 32398 6402 32450 6414
rect 49086 6402 49138 6414
rect 49646 6466 49698 6478
rect 49646 6402 49698 6414
rect 51886 6466 51938 6478
rect 51886 6402 51938 6414
rect 56814 6466 56866 6478
rect 56814 6402 56866 6414
rect 61518 6466 61570 6478
rect 61518 6402 61570 6414
rect 64430 6466 64482 6478
rect 64430 6402 64482 6414
rect 67342 6466 67394 6478
rect 67342 6402 67394 6414
rect 69358 6466 69410 6478
rect 69358 6402 69410 6414
rect 72270 6466 72322 6478
rect 75506 6414 75518 6466
rect 75570 6414 75582 6466
rect 76738 6414 76750 6466
rect 76802 6414 76814 6466
rect 77634 6414 77646 6466
rect 77698 6414 77710 6466
rect 72270 6402 72322 6414
rect 1344 6298 78624 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 50558 6298
rect 50610 6246 50662 6298
rect 50714 6246 50766 6298
rect 50818 6246 78624 6298
rect 1344 6212 78624 6246
rect 8318 6130 8370 6142
rect 2034 6078 2046 6130
rect 2098 6078 2110 6130
rect 8318 6066 8370 6078
rect 8654 6130 8706 6142
rect 8654 6066 8706 6078
rect 13918 6130 13970 6142
rect 13918 6066 13970 6078
rect 14366 6130 14418 6142
rect 15150 6130 15202 6142
rect 14802 6078 14814 6130
rect 14866 6078 14878 6130
rect 14366 6066 14418 6078
rect 15150 6066 15202 6078
rect 15598 6130 15650 6142
rect 15598 6066 15650 6078
rect 18062 6130 18114 6142
rect 18062 6066 18114 6078
rect 18286 6130 18338 6142
rect 18286 6066 18338 6078
rect 21534 6130 21586 6142
rect 21534 6066 21586 6078
rect 26350 6130 26402 6142
rect 28926 6130 28978 6142
rect 27906 6078 27918 6130
rect 27970 6078 27982 6130
rect 26350 6066 26402 6078
rect 28926 6066 28978 6078
rect 34190 6130 34242 6142
rect 34190 6066 34242 6078
rect 34414 6130 34466 6142
rect 34414 6066 34466 6078
rect 34638 6130 34690 6142
rect 41134 6130 41186 6142
rect 47966 6130 48018 6142
rect 36082 6078 36094 6130
rect 36146 6078 36158 6130
rect 40226 6078 40238 6130
rect 40290 6078 40302 6130
rect 44034 6078 44046 6130
rect 44098 6078 44110 6130
rect 46722 6078 46734 6130
rect 46786 6078 46798 6130
rect 34638 6066 34690 6078
rect 41134 6066 41186 6078
rect 47966 6066 48018 6078
rect 49646 6130 49698 6142
rect 49646 6066 49698 6078
rect 50766 6130 50818 6142
rect 50766 6066 50818 6078
rect 53902 6130 53954 6142
rect 53902 6066 53954 6078
rect 56030 6130 56082 6142
rect 56030 6066 56082 6078
rect 63870 6130 63922 6142
rect 63870 6066 63922 6078
rect 71038 6130 71090 6142
rect 71038 6066 71090 6078
rect 78206 6130 78258 6142
rect 78206 6066 78258 6078
rect 6638 6018 6690 6030
rect 6638 5954 6690 5966
rect 8990 6018 9042 6030
rect 8990 5954 9042 5966
rect 13694 6018 13746 6030
rect 13694 5954 13746 5966
rect 14142 6018 14194 6030
rect 14142 5954 14194 5966
rect 15710 6018 15762 6030
rect 15710 5954 15762 5966
rect 16494 6018 16546 6030
rect 16494 5954 16546 5966
rect 16830 6018 16882 6030
rect 16830 5954 16882 5966
rect 22654 6018 22706 6030
rect 22654 5954 22706 5966
rect 23326 6018 23378 6030
rect 23326 5954 23378 5966
rect 23662 6018 23714 6030
rect 23662 5954 23714 5966
rect 23998 6018 24050 6030
rect 23998 5954 24050 5966
rect 24334 6018 24386 6030
rect 24334 5954 24386 5966
rect 24670 6018 24722 6030
rect 24670 5954 24722 5966
rect 25566 6018 25618 6030
rect 25566 5954 25618 5966
rect 26126 6018 26178 6030
rect 26126 5954 26178 5966
rect 27470 6018 27522 6030
rect 35646 6018 35698 6030
rect 30370 5966 30382 6018
rect 30434 5966 30446 6018
rect 27470 5954 27522 5966
rect 35646 5954 35698 5966
rect 37662 6018 37714 6030
rect 42254 6018 42306 6030
rect 39554 5966 39566 6018
rect 39618 5966 39630 6018
rect 40002 5966 40014 6018
rect 40066 5966 40078 6018
rect 37662 5954 37714 5966
rect 42254 5954 42306 5966
rect 43150 6018 43202 6030
rect 43150 5954 43202 5966
rect 45166 6018 45218 6030
rect 45166 5954 45218 5966
rect 48750 6018 48802 6030
rect 48750 5954 48802 5966
rect 63198 6018 63250 6030
rect 63198 5954 63250 5966
rect 1710 5906 1762 5918
rect 1710 5842 1762 5854
rect 7982 5906 8034 5918
rect 14030 5906 14082 5918
rect 17726 5906 17778 5918
rect 9874 5854 9886 5906
rect 9938 5854 9950 5906
rect 17378 5854 17390 5906
rect 17442 5854 17454 5906
rect 7982 5842 8034 5854
rect 14030 5842 14082 5854
rect 17726 5842 17778 5854
rect 18174 5906 18226 5918
rect 18174 5842 18226 5854
rect 18734 5906 18786 5918
rect 22318 5906 22370 5918
rect 26798 5906 26850 5918
rect 21746 5854 21758 5906
rect 21810 5854 21822 5906
rect 22978 5854 22990 5906
rect 23042 5854 23054 5906
rect 18734 5842 18786 5854
rect 22318 5842 22370 5854
rect 26798 5842 26850 5854
rect 28254 5906 28306 5918
rect 28254 5842 28306 5854
rect 28478 5906 28530 5918
rect 28478 5842 28530 5854
rect 29262 5906 29314 5918
rect 41806 5906 41858 5918
rect 29698 5854 29710 5906
rect 29762 5854 29774 5906
rect 33842 5854 33854 5906
rect 33906 5854 33918 5906
rect 35074 5854 35086 5906
rect 35138 5854 35150 5906
rect 37090 5854 37102 5906
rect 37154 5854 37166 5906
rect 39330 5854 39342 5906
rect 39394 5854 39406 5906
rect 29262 5842 29314 5854
rect 41806 5842 41858 5854
rect 44270 5906 44322 5918
rect 47070 5906 47122 5918
rect 46386 5854 46398 5906
rect 46450 5854 46462 5906
rect 44270 5842 44322 5854
rect 47070 5842 47122 5854
rect 47630 5906 47682 5918
rect 47630 5842 47682 5854
rect 49086 5906 49138 5918
rect 71710 5906 71762 5918
rect 49858 5854 49870 5906
rect 49922 5854 49934 5906
rect 56914 5854 56926 5906
rect 56978 5854 56990 5906
rect 59826 5854 59838 5906
rect 59890 5854 59902 5906
rect 64418 5854 64430 5906
rect 64482 5854 64494 5906
rect 67330 5854 67342 5906
rect 67394 5854 67406 5906
rect 72258 5854 72270 5906
rect 72322 5854 72334 5906
rect 77298 5854 77310 5906
rect 77362 5854 77374 5906
rect 49086 5842 49138 5854
rect 71710 5842 71762 5854
rect 2494 5794 2546 5806
rect 2494 5730 2546 5742
rect 5294 5794 5346 5806
rect 5294 5730 5346 5742
rect 5742 5794 5794 5806
rect 5742 5730 5794 5742
rect 6190 5794 6242 5806
rect 6190 5730 6242 5742
rect 7086 5794 7138 5806
rect 7086 5730 7138 5742
rect 7534 5794 7586 5806
rect 12798 5794 12850 5806
rect 10658 5742 10670 5794
rect 10722 5742 10734 5794
rect 7534 5730 7586 5742
rect 12798 5730 12850 5742
rect 19182 5794 19234 5806
rect 19182 5730 19234 5742
rect 19630 5794 19682 5806
rect 19630 5730 19682 5742
rect 20078 5794 20130 5806
rect 20078 5730 20130 5742
rect 20526 5794 20578 5806
rect 20526 5730 20578 5742
rect 21198 5794 21250 5806
rect 21198 5730 21250 5742
rect 23214 5794 23266 5806
rect 26238 5794 26290 5806
rect 25442 5742 25454 5794
rect 25506 5742 25518 5794
rect 23214 5730 23266 5742
rect 26238 5730 26290 5742
rect 27246 5794 27298 5806
rect 33294 5794 33346 5806
rect 27570 5742 27582 5794
rect 27634 5742 27646 5794
rect 32498 5742 32510 5794
rect 32562 5742 32574 5794
rect 27246 5730 27298 5742
rect 33294 5730 33346 5742
rect 34302 5794 34354 5806
rect 34302 5730 34354 5742
rect 47294 5794 47346 5806
rect 47294 5730 47346 5742
rect 51214 5794 51266 5806
rect 51214 5730 51266 5742
rect 51662 5794 51714 5806
rect 51662 5730 51714 5742
rect 52558 5794 52610 5806
rect 70478 5794 70530 5806
rect 65538 5742 65550 5794
rect 65602 5742 65614 5794
rect 68898 5742 68910 5794
rect 68962 5742 68974 5794
rect 75618 5742 75630 5794
rect 75682 5742 75694 5794
rect 52558 5730 52610 5742
rect 70478 5730 70530 5742
rect 15486 5682 15538 5694
rect 7522 5630 7534 5682
rect 7586 5679 7598 5682
rect 8194 5679 8206 5682
rect 7586 5633 8206 5679
rect 7586 5630 7598 5633
rect 8194 5630 8206 5633
rect 8258 5630 8270 5682
rect 15486 5618 15538 5630
rect 17390 5682 17442 5694
rect 17390 5618 17442 5630
rect 21422 5682 21474 5694
rect 21422 5618 21474 5630
rect 25790 5682 25842 5694
rect 25790 5618 25842 5630
rect 33518 5682 33570 5694
rect 33518 5618 33570 5630
rect 33854 5682 33906 5694
rect 33854 5618 33906 5630
rect 41582 5682 41634 5694
rect 41582 5618 41634 5630
rect 42030 5682 42082 5694
rect 42030 5618 42082 5630
rect 57934 5682 57986 5694
rect 57934 5618 57986 5630
rect 60846 5682 60898 5694
rect 60846 5618 60898 5630
rect 73278 5682 73330 5694
rect 73278 5618 73330 5630
rect 1344 5514 78624 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 65918 5514
rect 65970 5462 66022 5514
rect 66074 5462 66126 5514
rect 66178 5462 78624 5514
rect 1344 5428 78624 5462
rect 8990 5346 9042 5358
rect 8990 5282 9042 5294
rect 10782 5346 10834 5358
rect 10782 5282 10834 5294
rect 12014 5346 12066 5358
rect 12014 5282 12066 5294
rect 20750 5346 20802 5358
rect 20750 5282 20802 5294
rect 21534 5346 21586 5358
rect 21534 5282 21586 5294
rect 26574 5346 26626 5358
rect 26574 5282 26626 5294
rect 28590 5346 28642 5358
rect 28590 5282 28642 5294
rect 30942 5346 30994 5358
rect 30942 5282 30994 5294
rect 69358 5346 69410 5358
rect 69358 5282 69410 5294
rect 10222 5234 10274 5246
rect 10222 5170 10274 5182
rect 10670 5234 10722 5246
rect 10670 5170 10722 5182
rect 11454 5234 11506 5246
rect 11454 5170 11506 5182
rect 12462 5234 12514 5246
rect 12462 5170 12514 5182
rect 13694 5234 13746 5246
rect 13694 5170 13746 5182
rect 14142 5234 14194 5246
rect 19518 5234 19570 5246
rect 14690 5182 14702 5234
rect 14754 5182 14766 5234
rect 16706 5182 16718 5234
rect 16770 5182 16782 5234
rect 18946 5182 18958 5234
rect 19010 5182 19022 5234
rect 14142 5170 14194 5182
rect 19518 5170 19570 5182
rect 20638 5234 20690 5246
rect 22430 5234 22482 5246
rect 26462 5234 26514 5246
rect 21746 5182 21758 5234
rect 21810 5182 21822 5234
rect 23650 5182 23662 5234
rect 23714 5182 23726 5234
rect 25778 5182 25790 5234
rect 25842 5182 25854 5234
rect 20638 5170 20690 5182
rect 22430 5170 22482 5182
rect 26462 5170 26514 5182
rect 27806 5234 27858 5246
rect 27806 5170 27858 5182
rect 27918 5234 27970 5246
rect 29598 5234 29650 5246
rect 28354 5182 28366 5234
rect 28418 5182 28430 5234
rect 27918 5170 27970 5182
rect 29598 5170 29650 5182
rect 30830 5234 30882 5246
rect 30830 5170 30882 5182
rect 31838 5234 31890 5246
rect 31838 5170 31890 5182
rect 49758 5234 49810 5246
rect 49758 5170 49810 5182
rect 50094 5234 50146 5246
rect 50094 5170 50146 5182
rect 55246 5234 55298 5246
rect 55246 5170 55298 5182
rect 58158 5234 58210 5246
rect 58158 5170 58210 5182
rect 64430 5234 64482 5246
rect 64430 5170 64482 5182
rect 66446 5234 66498 5246
rect 66446 5170 66498 5182
rect 67118 5234 67170 5246
rect 67118 5170 67170 5182
rect 67454 5234 67506 5246
rect 67454 5170 67506 5182
rect 72270 5234 72322 5246
rect 72270 5170 72322 5182
rect 74734 5234 74786 5246
rect 75506 5182 75518 5234
rect 75570 5182 75582 5234
rect 74734 5170 74786 5182
rect 1710 5122 1762 5134
rect 1710 5058 1762 5070
rect 2494 5122 2546 5134
rect 2494 5058 2546 5070
rect 6190 5122 6242 5134
rect 8878 5122 8930 5134
rect 6514 5070 6526 5122
rect 6578 5070 6590 5122
rect 7298 5070 7310 5122
rect 7362 5070 7374 5122
rect 8194 5070 8206 5122
rect 8258 5070 8270 5122
rect 8642 5070 8654 5122
rect 8706 5070 8718 5122
rect 6190 5058 6242 5070
rect 8878 5058 8930 5070
rect 9662 5122 9714 5134
rect 12350 5122 12402 5134
rect 15598 5122 15650 5134
rect 19406 5122 19458 5134
rect 27246 5122 27298 5134
rect 29486 5122 29538 5134
rect 32286 5122 32338 5134
rect 39566 5122 39618 5134
rect 11666 5070 11678 5122
rect 11730 5070 11742 5122
rect 12898 5070 12910 5122
rect 12962 5070 12974 5122
rect 15922 5070 15934 5122
rect 15986 5070 15998 5122
rect 19730 5070 19742 5122
rect 19794 5070 19806 5122
rect 20402 5070 20414 5122
rect 20466 5070 20478 5122
rect 21858 5070 21870 5122
rect 21922 5070 21934 5122
rect 22866 5070 22878 5122
rect 22930 5070 22942 5122
rect 27570 5070 27582 5122
rect 27634 5070 27646 5122
rect 28242 5070 28254 5122
rect 28306 5070 28318 5122
rect 29250 5070 29262 5122
rect 29314 5070 29326 5122
rect 30594 5070 30606 5122
rect 30658 5070 30670 5122
rect 31378 5070 31390 5122
rect 31442 5070 31454 5122
rect 32610 5070 32622 5122
rect 32674 5070 32686 5122
rect 36418 5070 36430 5122
rect 36482 5070 36494 5122
rect 37090 5070 37102 5122
rect 37154 5070 37166 5122
rect 37314 5070 37326 5122
rect 37378 5070 37390 5122
rect 37538 5070 37550 5122
rect 37602 5070 37614 5122
rect 9662 5058 9714 5070
rect 12350 5058 12402 5070
rect 15598 5058 15650 5070
rect 19406 5058 19458 5070
rect 27246 5058 27298 5070
rect 29486 5058 29538 5070
rect 32286 5058 32338 5070
rect 39566 5058 39618 5070
rect 40014 5122 40066 5134
rect 51102 5122 51154 5134
rect 40450 5070 40462 5122
rect 40514 5070 40526 5122
rect 42690 5070 42702 5122
rect 42754 5070 42766 5122
rect 44818 5070 44830 5122
rect 44882 5070 44894 5122
rect 46834 5070 46846 5122
rect 46898 5070 46910 5122
rect 49186 5070 49198 5122
rect 49250 5070 49262 5122
rect 50530 5070 50542 5122
rect 50594 5070 50606 5122
rect 40014 5058 40066 5070
rect 51102 5058 51154 5070
rect 51550 5122 51602 5134
rect 51550 5058 51602 5070
rect 53566 5122 53618 5134
rect 75070 5122 75122 5134
rect 54226 5070 54238 5122
rect 54290 5070 54302 5122
rect 57138 5070 57150 5122
rect 57202 5070 57214 5122
rect 60610 5070 60622 5122
rect 60674 5070 60686 5122
rect 63522 5070 63534 5122
rect 63586 5070 63598 5122
rect 68450 5070 68462 5122
rect 68514 5070 68526 5122
rect 71362 5070 71374 5122
rect 71426 5070 71438 5122
rect 53566 5058 53618 5070
rect 75070 5058 75122 5070
rect 76526 5122 76578 5134
rect 77870 5122 77922 5134
rect 77410 5070 77422 5122
rect 77474 5070 77486 5122
rect 76526 5058 76578 5070
rect 77870 5058 77922 5070
rect 6750 5010 6802 5022
rect 2034 4958 2046 5010
rect 2098 4958 2110 5010
rect 6750 4946 6802 4958
rect 7646 5010 7698 5022
rect 7646 4946 7698 4958
rect 7982 5010 8034 5022
rect 7982 4946 8034 4958
rect 9326 5010 9378 5022
rect 9326 4946 9378 4958
rect 10558 5010 10610 5022
rect 10558 4946 10610 4958
rect 12574 5010 12626 5022
rect 12574 4946 12626 4958
rect 14030 5010 14082 5022
rect 14030 4946 14082 4958
rect 14254 5010 14306 5022
rect 14254 4946 14306 4958
rect 14702 5010 14754 5022
rect 14702 4946 14754 4958
rect 14926 5010 14978 5022
rect 14926 4946 14978 4958
rect 22542 5010 22594 5022
rect 22542 4946 22594 4958
rect 26910 5010 26962 5022
rect 26910 4946 26962 4958
rect 29934 5010 29986 5022
rect 29934 4946 29986 4958
rect 30270 5010 30322 5022
rect 30270 4946 30322 4958
rect 33294 5010 33346 5022
rect 33294 4946 33346 4958
rect 35310 5010 35362 5022
rect 35310 4946 35362 4958
rect 38334 5010 38386 5022
rect 39790 5010 39842 5022
rect 38882 4958 38894 5010
rect 38946 4958 38958 5010
rect 39106 4958 39118 5010
rect 39170 4958 39182 5010
rect 38334 4946 38386 4958
rect 39790 4946 39842 4958
rect 40126 5010 40178 5022
rect 43150 5010 43202 5022
rect 40562 4958 40574 5010
rect 40626 4958 40638 5010
rect 40126 4946 40178 4958
rect 43150 4946 43202 4958
rect 45390 5010 45442 5022
rect 45390 4946 45442 4958
rect 47406 5010 47458 5022
rect 47406 4946 47458 4958
rect 48974 5010 49026 5022
rect 48974 4946 49026 4958
rect 76190 5010 76242 5022
rect 76190 4946 76242 4958
rect 77198 5010 77250 5022
rect 77198 4946 77250 4958
rect 78206 5010 78258 5022
rect 78206 4946 78258 4958
rect 4286 4898 4338 4910
rect 4286 4834 4338 4846
rect 4734 4898 4786 4910
rect 4734 4834 4786 4846
rect 5182 4898 5234 4910
rect 5182 4834 5234 4846
rect 7534 4898 7586 4910
rect 7534 4834 7586 4846
rect 11902 4898 11954 4910
rect 11902 4834 11954 4846
rect 15262 4898 15314 4910
rect 15262 4834 15314 4846
rect 22318 4898 22370 4910
rect 22318 4834 22370 4846
rect 26350 4898 26402 4910
rect 26350 4834 26402 4846
rect 33966 4898 34018 4910
rect 52110 4898 52162 4910
rect 42802 4846 42814 4898
rect 42866 4846 42878 4898
rect 45826 4846 45838 4898
rect 45890 4846 45902 4898
rect 33966 4834 34018 4846
rect 52110 4834 52162 4846
rect 53230 4898 53282 4910
rect 53230 4834 53282 4846
rect 61518 4898 61570 4910
rect 61518 4834 61570 4846
rect 1344 4730 78624 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 50558 4730
rect 50610 4678 50662 4730
rect 50714 4678 50766 4730
rect 50818 4678 78624 4730
rect 1344 4644 78624 4678
rect 4286 4562 4338 4574
rect 4286 4498 4338 4510
rect 4958 4562 5010 4574
rect 4958 4498 5010 4510
rect 5630 4562 5682 4574
rect 5630 4498 5682 4510
rect 6078 4562 6130 4574
rect 6078 4498 6130 4510
rect 6190 4562 6242 4574
rect 6190 4498 6242 4510
rect 8990 4562 9042 4574
rect 17838 4562 17890 4574
rect 16706 4510 16718 4562
rect 16770 4510 16782 4562
rect 8990 4498 9042 4510
rect 17838 4498 17890 4510
rect 18622 4562 18674 4574
rect 18622 4498 18674 4510
rect 19630 4562 19682 4574
rect 19630 4498 19682 4510
rect 20638 4562 20690 4574
rect 20638 4498 20690 4510
rect 21198 4562 21250 4574
rect 33182 4562 33234 4574
rect 42142 4562 42194 4574
rect 32386 4510 32398 4562
rect 32450 4510 32462 4562
rect 40226 4510 40238 4562
rect 40290 4510 40302 4562
rect 21198 4498 21250 4510
rect 33182 4498 33234 4510
rect 42142 4498 42194 4510
rect 48750 4562 48802 4574
rect 48750 4498 48802 4510
rect 55918 4562 55970 4574
rect 55918 4498 55970 4510
rect 63198 4562 63250 4574
rect 63198 4498 63250 4510
rect 71038 4562 71090 4574
rect 71038 4498 71090 4510
rect 71710 4562 71762 4574
rect 71710 4498 71762 4510
rect 78206 4562 78258 4574
rect 78206 4498 78258 4510
rect 7646 4450 7698 4462
rect 7646 4386 7698 4398
rect 8318 4450 8370 4462
rect 8318 4386 8370 4398
rect 9886 4450 9938 4462
rect 9886 4386 9938 4398
rect 17950 4450 18002 4462
rect 17950 4386 18002 4398
rect 18286 4450 18338 4462
rect 18286 4386 18338 4398
rect 19294 4450 19346 4462
rect 19294 4386 19346 4398
rect 19966 4450 20018 4462
rect 19966 4386 20018 4398
rect 20302 4450 20354 4462
rect 20302 4386 20354 4398
rect 21310 4450 21362 4462
rect 21310 4386 21362 4398
rect 21758 4450 21810 4462
rect 21758 4386 21810 4398
rect 21982 4450 22034 4462
rect 21982 4386 22034 4398
rect 22654 4450 22706 4462
rect 22654 4386 22706 4398
rect 22990 4450 23042 4462
rect 22990 4386 23042 4398
rect 23102 4450 23154 4462
rect 23102 4386 23154 4398
rect 23214 4450 23266 4462
rect 23214 4386 23266 4398
rect 23998 4450 24050 4462
rect 23998 4386 24050 4398
rect 24334 4450 24386 4462
rect 24334 4386 24386 4398
rect 24670 4450 24722 4462
rect 31390 4450 31442 4462
rect 28802 4398 28814 4450
rect 28866 4398 28878 4450
rect 24670 4386 24722 4398
rect 31390 4386 31442 4398
rect 33294 4450 33346 4462
rect 39118 4450 39170 4462
rect 41582 4450 41634 4462
rect 45614 4450 45666 4462
rect 62526 4450 62578 4462
rect 34178 4398 34190 4450
rect 34242 4398 34254 4450
rect 36642 4398 36654 4450
rect 36706 4398 36718 4450
rect 40898 4398 40910 4450
rect 40962 4398 40974 4450
rect 42578 4398 42590 4450
rect 42642 4398 42654 4450
rect 46610 4398 46622 4450
rect 46674 4398 46686 4450
rect 46946 4398 46958 4450
rect 47010 4398 47022 4450
rect 33294 4386 33346 4398
rect 39118 4386 39170 4398
rect 41582 4386 41634 4398
rect 45614 4386 45666 4398
rect 62526 4386 62578 4398
rect 4622 4338 4674 4350
rect 7310 4338 7362 4350
rect 30830 4338 30882 4350
rect 4050 4286 4062 4338
rect 4114 4286 4126 4338
rect 5394 4286 5406 4338
rect 5458 4286 5470 4338
rect 6626 4286 6638 4338
rect 6690 4286 6702 4338
rect 7970 4286 7982 4338
rect 8034 4286 8046 4338
rect 8754 4286 8766 4338
rect 8818 4286 8830 4338
rect 9650 4286 9662 4338
rect 9714 4286 9726 4338
rect 10210 4286 10222 4338
rect 10274 4286 10286 4338
rect 13682 4286 13694 4338
rect 13746 4286 13758 4338
rect 17602 4286 17614 4338
rect 17666 4286 17678 4338
rect 18946 4286 18958 4338
rect 19010 4286 19022 4338
rect 20962 4286 20974 4338
rect 21026 4286 21038 4338
rect 22418 4286 22430 4338
rect 22482 4286 22494 4338
rect 23762 4286 23774 4338
rect 23826 4286 23838 4338
rect 25218 4286 25230 4338
rect 25282 4286 25294 4338
rect 28690 4286 28702 4338
rect 28754 4286 28766 4338
rect 4622 4274 4674 4286
rect 7310 4274 7362 4286
rect 30830 4274 30882 4286
rect 32958 4338 33010 4350
rect 35982 4338 36034 4350
rect 38670 4338 38722 4350
rect 33954 4286 33966 4338
rect 34018 4286 34030 4338
rect 36530 4286 36542 4338
rect 36594 4286 36606 4338
rect 32958 4274 33010 4286
rect 35982 4274 36034 4286
rect 38670 4274 38722 4286
rect 44158 4338 44210 4350
rect 49086 4338 49138 4350
rect 52558 4338 52610 4350
rect 46274 4286 46286 4338
rect 46338 4286 46350 4338
rect 47282 4286 47294 4338
rect 47346 4286 47358 4338
rect 49522 4286 49534 4338
rect 49586 4286 49598 4338
rect 52882 4286 52894 4338
rect 52946 4286 52958 4338
rect 56578 4286 56590 4338
rect 56642 4286 56654 4338
rect 61618 4286 61630 4338
rect 61682 4286 61694 4338
rect 64530 4286 64542 4338
rect 64594 4286 64606 4338
rect 67442 4286 67454 4338
rect 67506 4286 67518 4338
rect 72258 4286 72270 4338
rect 72322 4286 72334 4338
rect 75170 4286 75182 4338
rect 75234 4286 75246 4338
rect 44158 4274 44210 4286
rect 49086 4274 49138 4286
rect 52558 4274 52610 4286
rect 2158 4226 2210 4238
rect 2158 4162 2210 4174
rect 2494 4226 2546 4238
rect 2494 4162 2546 4174
rect 3278 4226 3330 4238
rect 3278 4162 3330 4174
rect 3726 4226 3778 4238
rect 8206 4226 8258 4238
rect 13134 4226 13186 4238
rect 41246 4226 41298 4238
rect 63534 4226 63586 4238
rect 70478 4226 70530 4238
rect 6738 4174 6750 4226
rect 6802 4174 6814 4226
rect 10994 4174 11006 4226
rect 11058 4174 11070 4226
rect 14466 4174 14478 4226
rect 14530 4174 14542 4226
rect 19058 4174 19070 4226
rect 19122 4174 19134 4226
rect 21746 4174 21758 4226
rect 21810 4174 21822 4226
rect 26002 4174 26014 4226
rect 26066 4174 26078 4226
rect 28130 4174 28142 4226
rect 28194 4174 28206 4226
rect 35074 4174 35086 4226
rect 35138 4174 35150 4226
rect 45266 4174 45278 4226
rect 45330 4174 45342 4226
rect 65538 4174 65550 4226
rect 65602 4174 65614 4226
rect 3726 4162 3778 4174
rect 8206 4162 8258 4174
rect 13134 4162 13186 4174
rect 41246 4162 41298 4174
rect 63534 4162 63586 4174
rect 70478 4162 70530 4174
rect 6302 4114 6354 4126
rect 6302 4050 6354 4062
rect 6974 4114 7026 4126
rect 6974 4050 7026 4062
rect 50542 4114 50594 4126
rect 50542 4050 50594 4062
rect 53902 4114 53954 4126
rect 53902 4050 53954 4062
rect 57598 4114 57650 4126
rect 57598 4050 57650 4062
rect 59726 4114 59778 4126
rect 68350 4114 68402 4126
rect 62626 4062 62638 4114
rect 62690 4111 62702 4114
rect 63522 4111 63534 4114
rect 62690 4065 63534 4111
rect 62690 4062 62702 4065
rect 63522 4062 63534 4065
rect 63586 4062 63598 4114
rect 59726 4050 59778 4062
rect 68350 4050 68402 4062
rect 73278 4114 73330 4126
rect 73278 4050 73330 4062
rect 76190 4114 76242 4126
rect 76190 4050 76242 4062
rect 1344 3946 78624 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 65918 3946
rect 65970 3894 66022 3946
rect 66074 3894 66126 3946
rect 66178 3894 78624 3946
rect 1344 3860 78624 3894
rect 11230 3778 11282 3790
rect 11230 3714 11282 3726
rect 15710 3778 15762 3790
rect 15710 3714 15762 3726
rect 17502 3778 17554 3790
rect 17502 3714 17554 3726
rect 21646 3778 21698 3790
rect 21646 3714 21698 3726
rect 21982 3778 22034 3790
rect 21982 3714 22034 3726
rect 25118 3778 25170 3790
rect 25118 3714 25170 3726
rect 67454 3778 67506 3790
rect 67454 3714 67506 3726
rect 75070 3778 75122 3790
rect 75070 3714 75122 3726
rect 11118 3666 11170 3678
rect 11118 3602 11170 3614
rect 15598 3666 15650 3678
rect 25006 3666 25058 3678
rect 47406 3666 47458 3678
rect 17266 3614 17278 3666
rect 17330 3614 17342 3666
rect 23426 3614 23438 3666
rect 23490 3614 23502 3666
rect 39330 3614 39342 3666
rect 39394 3614 39406 3666
rect 41794 3614 41806 3666
rect 41858 3614 41870 3666
rect 45714 3614 45726 3666
rect 45778 3614 45790 3666
rect 15598 3602 15650 3614
rect 25006 3602 25058 3614
rect 47406 3602 47458 3614
rect 50654 3666 50706 3678
rect 50654 3602 50706 3614
rect 51774 3666 51826 3678
rect 51774 3602 51826 3614
rect 56030 3666 56082 3678
rect 56030 3602 56082 3614
rect 58046 3666 58098 3678
rect 58046 3602 58098 3614
rect 59054 3666 59106 3678
rect 59054 3602 59106 3614
rect 61854 3666 61906 3678
rect 65662 3666 65714 3678
rect 63858 3614 63870 3666
rect 63922 3614 63934 3666
rect 61854 3602 61906 3614
rect 65662 3602 65714 3614
rect 69806 3666 69858 3678
rect 69806 3602 69858 3614
rect 71262 3666 71314 3678
rect 71262 3602 71314 3614
rect 77198 3666 77250 3678
rect 77198 3602 77250 3614
rect 7086 3554 7138 3566
rect 1810 3502 1822 3554
rect 1874 3502 1886 3554
rect 3378 3502 3390 3554
rect 3442 3502 3454 3554
rect 4722 3502 4734 3554
rect 4786 3502 4798 3554
rect 5842 3502 5854 3554
rect 5906 3502 5918 3554
rect 6514 3502 6526 3554
rect 6578 3502 6590 3554
rect 7086 3490 7138 3502
rect 7758 3554 7810 3566
rect 10222 3554 10274 3566
rect 12238 3554 12290 3566
rect 16046 3554 16098 3566
rect 19182 3554 19234 3566
rect 22990 3554 23042 3566
rect 25454 3554 25506 3566
rect 8530 3502 8542 3554
rect 8594 3502 8606 3554
rect 9650 3502 9662 3554
rect 9714 3502 9726 3554
rect 10882 3502 10894 3554
rect 10946 3502 10958 3554
rect 11666 3502 11678 3554
rect 11730 3502 11742 3554
rect 13458 3502 13470 3554
rect 13522 3502 13534 3554
rect 14130 3502 14142 3554
rect 14194 3502 14206 3554
rect 14802 3502 14814 3554
rect 14866 3502 14878 3554
rect 15362 3502 15374 3554
rect 15426 3502 15438 3554
rect 18610 3502 18622 3554
rect 18674 3502 18686 3554
rect 19954 3502 19966 3554
rect 20018 3502 20030 3554
rect 21074 3502 21086 3554
rect 21138 3502 21150 3554
rect 21634 3502 21646 3554
rect 21698 3502 21710 3554
rect 24770 3502 24782 3554
rect 24834 3502 24846 3554
rect 7758 3490 7810 3502
rect 10222 3490 10274 3502
rect 12238 3490 12290 3502
rect 16046 3490 16098 3502
rect 19182 3490 19234 3502
rect 22990 3490 23042 3502
rect 25454 3490 25506 3502
rect 26126 3554 26178 3566
rect 28590 3554 28642 3566
rect 32398 3554 32450 3566
rect 26898 3502 26910 3554
rect 26962 3502 26974 3554
rect 27570 3502 27582 3554
rect 27634 3502 27646 3554
rect 29362 3502 29374 3554
rect 29426 3502 29438 3554
rect 30034 3502 30046 3554
rect 30098 3502 30110 3554
rect 31378 3502 31390 3554
rect 31442 3502 31454 3554
rect 26126 3490 26178 3502
rect 28590 3490 28642 3502
rect 32398 3490 32450 3502
rect 33070 3554 33122 3566
rect 33070 3490 33122 3502
rect 33742 3554 33794 3566
rect 35086 3554 35138 3566
rect 48190 3554 48242 3566
rect 54238 3554 54290 3566
rect 34514 3502 34526 3554
rect 34578 3502 34590 3554
rect 36866 3502 36878 3554
rect 36930 3502 36942 3554
rect 37650 3502 37662 3554
rect 37714 3502 37726 3554
rect 41346 3502 41358 3554
rect 41410 3502 41422 3554
rect 43026 3502 43038 3554
rect 43090 3502 43102 3554
rect 43698 3502 43710 3554
rect 43762 3502 43774 3554
rect 45266 3502 45278 3554
rect 45330 3502 45342 3554
rect 47954 3502 47966 3554
rect 48018 3502 48030 3554
rect 48738 3502 48750 3554
rect 48802 3502 48814 3554
rect 49410 3502 49422 3554
rect 49474 3502 49486 3554
rect 50082 3502 50094 3554
rect 50146 3502 50158 3554
rect 52322 3502 52334 3554
rect 52386 3502 52398 3554
rect 52994 3502 53006 3554
rect 53058 3502 53070 3554
rect 53666 3502 53678 3554
rect 53730 3502 53742 3554
rect 55010 3502 55022 3554
rect 55074 3502 55086 3554
rect 61394 3502 61406 3554
rect 61458 3502 61470 3554
rect 62626 3502 62638 3554
rect 62690 3502 62702 3554
rect 66434 3502 66446 3554
rect 66498 3502 66510 3554
rect 70242 3502 70254 3554
rect 70306 3502 70318 3554
rect 74050 3502 74062 3554
rect 74114 3502 74126 3554
rect 78082 3502 78094 3554
rect 78146 3502 78158 3554
rect 33742 3490 33794 3502
rect 35086 3490 35138 3502
rect 48190 3490 48242 3502
rect 54238 3490 54290 3502
rect 2382 3442 2434 3454
rect 3614 3442 3666 3454
rect 2034 3390 2046 3442
rect 2098 3390 2110 3442
rect 2706 3390 2718 3442
rect 2770 3390 2782 3442
rect 2382 3378 2434 3390
rect 3614 3378 3666 3390
rect 3950 3442 4002 3454
rect 3950 3378 4002 3390
rect 4286 3442 4338 3454
rect 4286 3378 4338 3390
rect 4958 3442 5010 3454
rect 4958 3378 5010 3390
rect 6078 3442 6130 3454
rect 6078 3378 6130 3390
rect 7422 3442 7474 3454
rect 7422 3378 7474 3390
rect 8766 3442 8818 3454
rect 8766 3378 8818 3390
rect 12574 3442 12626 3454
rect 12574 3378 12626 3390
rect 13694 3442 13746 3454
rect 13694 3378 13746 3390
rect 14366 3442 14418 3454
rect 14366 3378 14418 3390
rect 15038 3442 15090 3454
rect 15038 3378 15090 3390
rect 17838 3442 17890 3454
rect 17838 3378 17890 3390
rect 18174 3442 18226 3454
rect 18174 3378 18226 3390
rect 19518 3442 19570 3454
rect 19518 3378 19570 3390
rect 20190 3442 20242 3454
rect 20190 3378 20242 3390
rect 22318 3442 22370 3454
rect 22318 3378 22370 3390
rect 22654 3442 22706 3454
rect 22654 3378 22706 3390
rect 25790 3442 25842 3454
rect 25790 3378 25842 3390
rect 26462 3442 26514 3454
rect 26462 3378 26514 3390
rect 27134 3442 27186 3454
rect 27134 3378 27186 3390
rect 29598 3442 29650 3454
rect 29598 3378 29650 3390
rect 30270 3442 30322 3454
rect 30270 3378 30322 3390
rect 30606 3442 30658 3454
rect 30606 3378 30658 3390
rect 32734 3442 32786 3454
rect 32734 3378 32786 3390
rect 33406 3442 33458 3454
rect 33406 3378 33458 3390
rect 34078 3442 34130 3454
rect 34078 3378 34130 3390
rect 34750 3442 34802 3454
rect 34750 3378 34802 3390
rect 35422 3442 35474 3454
rect 48526 3442 48578 3454
rect 49870 3442 49922 3454
rect 36754 3390 36766 3442
rect 36818 3390 36830 3442
rect 37538 3390 37550 3442
rect 37602 3390 37614 3442
rect 41458 3390 41470 3442
rect 41522 3390 41534 3442
rect 42242 3390 42254 3442
rect 42306 3390 42318 3442
rect 44370 3390 44382 3442
rect 44434 3390 44446 3442
rect 45378 3390 45390 3442
rect 45442 3390 45454 3442
rect 49186 3390 49198 3442
rect 49250 3390 49262 3442
rect 35422 3378 35474 3390
rect 48526 3378 48578 3390
rect 49870 3378 49922 3390
rect 51214 3442 51266 3454
rect 73614 3442 73666 3454
rect 52770 3390 52782 3442
rect 52834 3390 52846 3442
rect 53442 3390 53454 3442
rect 53506 3390 53518 3442
rect 51214 3378 51266 3390
rect 73614 3378 73666 3390
rect 77870 3442 77922 3454
rect 77870 3378 77922 3390
rect 6750 3330 6802 3342
rect 6750 3266 6802 3278
rect 8094 3330 8146 3342
rect 8094 3266 8146 3278
rect 9886 3330 9938 3342
rect 9886 3266 9938 3278
rect 10558 3330 10610 3342
rect 10558 3266 10610 3278
rect 11902 3330 11954 3342
rect 11902 3266 11954 3278
rect 16382 3330 16434 3342
rect 16382 3266 16434 3278
rect 17278 3330 17330 3342
rect 17278 3266 17330 3278
rect 18846 3330 18898 3342
rect 24110 3330 24162 3342
rect 21298 3278 21310 3330
rect 21362 3278 21374 3330
rect 18846 3266 18898 3278
rect 24110 3266 24162 3278
rect 27806 3330 27858 3342
rect 30942 3330 30994 3342
rect 28914 3278 28926 3330
rect 28978 3278 28990 3330
rect 27806 3266 27858 3278
rect 30942 3266 30994 3278
rect 31614 3330 31666 3342
rect 52098 3278 52110 3330
rect 52162 3278 52174 3330
rect 31614 3266 31666 3278
rect 1344 3162 78624 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 50558 3162
rect 50610 3110 50662 3162
rect 50714 3110 50766 3162
rect 50818 3110 78624 3162
rect 1344 3076 78624 3110
rect 18610 2942 18622 2994
rect 18674 2991 18686 2994
rect 22418 2991 22430 2994
rect 18674 2945 22430 2991
rect 18674 2942 18686 2945
rect 22418 2942 22430 2945
rect 22482 2942 22494 2994
<< via1 >>
rect 69022 77198 69074 77250
rect 70254 77198 70306 77250
rect 75070 77198 75122 77250
rect 75854 77198 75906 77250
rect 76414 77198 76466 77250
rect 50878 77086 50930 77138
rect 51774 77086 51826 77138
rect 52110 77086 52162 77138
rect 66334 77086 66386 77138
rect 67118 77086 67170 77138
rect 67454 77086 67506 77138
rect 68686 77086 68738 77138
rect 42814 76974 42866 77026
rect 43598 76974 43650 77026
rect 45502 76974 45554 77026
rect 46286 76974 46338 77026
rect 47518 76974 47570 77026
rect 48302 76974 48354 77026
rect 48862 76974 48914 77026
rect 50094 76974 50146 77026
rect 51550 76974 51602 77026
rect 53006 76974 53058 77026
rect 60958 76974 61010 77026
rect 61854 76974 61906 77026
rect 62302 76974 62354 77026
rect 63310 76974 63362 77026
rect 64318 76974 64370 77026
rect 65326 76974 65378 77026
rect 65662 76974 65714 77026
rect 66446 76974 66498 77026
rect 67678 76974 67730 77026
rect 68462 76974 68514 77026
rect 71038 76974 71090 77026
rect 71934 76974 71986 77026
rect 72606 76974 72658 77026
rect 74398 76974 74450 77026
rect 75070 76974 75122 77026
rect 75742 76974 75794 77026
rect 76638 76974 76690 77026
rect 77198 76974 77250 77026
rect 19838 76806 19890 76858
rect 19942 76806 19994 76858
rect 20046 76806 20098 76858
rect 50558 76806 50610 76858
rect 50662 76806 50714 76858
rect 50766 76806 50818 76858
rect 4622 76638 4674 76690
rect 15374 76638 15426 76690
rect 19182 76638 19234 76690
rect 21086 76638 21138 76690
rect 24894 76638 24946 76690
rect 25566 76638 25618 76690
rect 26238 76638 26290 76690
rect 26910 76638 26962 76690
rect 27582 76638 27634 76690
rect 28366 76638 28418 76690
rect 28926 76638 28978 76690
rect 29598 76638 29650 76690
rect 30270 76638 30322 76690
rect 30942 76638 30994 76690
rect 31502 76638 31554 76690
rect 32286 76638 32338 76690
rect 36766 76638 36818 76690
rect 37662 76638 37714 76690
rect 39230 76638 39282 76690
rect 40126 76638 40178 76690
rect 41022 76638 41074 76690
rect 42030 76638 42082 76690
rect 42366 76638 42418 76690
rect 43598 76638 43650 76690
rect 44494 76638 44546 76690
rect 45390 76638 45442 76690
rect 46286 76638 46338 76690
rect 47406 76638 47458 76690
rect 48302 76638 48354 76690
rect 49198 76638 49250 76690
rect 50094 76638 50146 76690
rect 51214 76638 51266 76690
rect 52110 76638 52162 76690
rect 53006 76638 53058 76690
rect 53902 76638 53954 76690
rect 55134 76638 55186 76690
rect 59838 76638 59890 76690
rect 63310 76638 63362 76690
rect 63982 76638 64034 76690
rect 64654 76638 64706 76690
rect 65326 76638 65378 76690
rect 66446 76638 66498 76690
rect 67118 76638 67170 76690
rect 67790 76638 67842 76690
rect 68462 76638 68514 76690
rect 69134 76638 69186 76690
rect 72606 76638 72658 76690
rect 74062 76638 74114 76690
rect 75406 76638 75458 76690
rect 76414 76638 76466 76690
rect 4958 76526 5010 76578
rect 5518 76526 5570 76578
rect 36094 76526 36146 76578
rect 61742 76526 61794 76578
rect 62638 76526 62690 76578
rect 62974 76526 63026 76578
rect 63646 76526 63698 76578
rect 64318 76526 64370 76578
rect 64990 76526 65042 76578
rect 65662 76526 65714 76578
rect 66782 76526 66834 76578
rect 67454 76526 67506 76578
rect 68126 76526 68178 76578
rect 68798 76526 68850 76578
rect 69470 76526 69522 76578
rect 70254 76526 70306 76578
rect 70590 76526 70642 76578
rect 70926 76526 70978 76578
rect 71262 76526 71314 76578
rect 71598 76526 71650 76578
rect 72270 76526 72322 76578
rect 72942 76526 72994 76578
rect 74398 76526 74450 76578
rect 74734 76526 74786 76578
rect 75742 76526 75794 76578
rect 76078 76526 76130 76578
rect 78206 76526 78258 76578
rect 4286 76414 4338 76466
rect 5742 76414 5794 76466
rect 12126 76414 12178 76466
rect 16382 76414 16434 76466
rect 19742 76414 19794 76466
rect 23886 76414 23938 76466
rect 35086 76414 35138 76466
rect 36318 76414 36370 76466
rect 58270 76414 58322 76466
rect 58830 76414 58882 76466
rect 62078 76414 62130 76466
rect 71822 76414 71874 76466
rect 73166 76414 73218 76466
rect 74958 76414 75010 76466
rect 77198 76414 77250 76466
rect 77870 76414 77922 76466
rect 13358 76302 13410 76354
rect 17166 76302 17218 76354
rect 21646 76302 21698 76354
rect 33406 76302 33458 76354
rect 37326 76302 37378 76354
rect 38110 76302 38162 76354
rect 38670 76302 38722 76354
rect 40686 76302 40738 76354
rect 41582 76302 41634 76354
rect 42814 76302 42866 76354
rect 44158 76302 44210 76354
rect 45054 76302 45106 76354
rect 45950 76302 46002 76354
rect 46846 76302 46898 76354
rect 47854 76302 47906 76354
rect 48862 76302 48914 76354
rect 49758 76302 49810 76354
rect 50542 76302 50594 76354
rect 51662 76302 51714 76354
rect 52670 76302 52722 76354
rect 53454 76302 53506 76354
rect 54350 76302 54402 76354
rect 55918 76302 55970 76354
rect 76750 76302 76802 76354
rect 1934 76190 1986 76242
rect 11566 76190 11618 76242
rect 4478 76022 4530 76074
rect 4582 76022 4634 76074
rect 4686 76022 4738 76074
rect 35198 76022 35250 76074
rect 35302 76022 35354 76074
rect 35406 76022 35458 76074
rect 65918 76022 65970 76074
rect 66022 76022 66074 76074
rect 66126 76022 66178 76074
rect 11902 75854 11954 75906
rect 16830 75854 16882 75906
rect 21534 75854 21586 75906
rect 56702 75854 56754 75906
rect 62638 75854 62690 75906
rect 63086 75854 63138 75906
rect 71374 75854 71426 75906
rect 71822 75854 71874 75906
rect 1934 75742 1986 75794
rect 18622 75742 18674 75794
rect 24782 75742 24834 75794
rect 32734 75742 32786 75794
rect 34078 75742 34130 75794
rect 35422 75742 35474 75794
rect 36430 75742 36482 75794
rect 37326 75742 37378 75794
rect 37886 75742 37938 75794
rect 38558 75742 38610 75794
rect 40014 75742 40066 75794
rect 41470 75742 41522 75794
rect 42478 75742 42530 75794
rect 43374 75742 43426 75794
rect 43934 75742 43986 75794
rect 44382 75742 44434 75794
rect 46062 75742 46114 75794
rect 46510 75742 46562 75794
rect 48078 75742 48130 75794
rect 48526 75742 48578 75794
rect 49086 75742 49138 75794
rect 49534 75742 49586 75794
rect 50206 75742 50258 75794
rect 50766 75742 50818 75794
rect 51214 75742 51266 75794
rect 51774 75742 51826 75794
rect 52222 75742 52274 75794
rect 54238 75742 54290 75794
rect 55134 75742 55186 75794
rect 56030 75742 56082 75794
rect 63086 75742 63138 75794
rect 63534 75742 63586 75794
rect 63982 75742 64034 75794
rect 64542 75742 64594 75794
rect 64990 75742 65042 75794
rect 65998 75742 66050 75794
rect 66446 75742 66498 75794
rect 67006 75742 67058 75794
rect 67566 75742 67618 75794
rect 68462 75742 68514 75794
rect 69022 75742 69074 75794
rect 70030 75742 70082 75794
rect 70702 75742 70754 75794
rect 71374 75742 71426 75794
rect 71934 75742 71986 75794
rect 72382 75742 72434 75794
rect 73390 75742 73442 75794
rect 73950 75742 74002 75794
rect 74510 75742 74562 75794
rect 75070 75742 75122 75794
rect 4286 75630 4338 75682
rect 4958 75630 5010 75682
rect 12686 75630 12738 75682
rect 13582 75630 13634 75682
rect 17838 75630 17890 75682
rect 20302 75630 20354 75682
rect 23662 75630 23714 75682
rect 25230 75630 25282 75682
rect 32958 75630 33010 75682
rect 33518 75630 33570 75682
rect 34302 75630 34354 75682
rect 34862 75630 34914 75682
rect 35646 75630 35698 75682
rect 38222 75630 38274 75682
rect 39006 75630 39058 75682
rect 39566 75630 39618 75682
rect 40910 75630 40962 75682
rect 41694 75630 41746 75682
rect 45166 75630 45218 75682
rect 45614 75630 45666 75682
rect 47070 75630 47122 75682
rect 47630 75630 47682 75682
rect 49758 75630 49810 75682
rect 52670 75630 52722 75682
rect 53230 75630 53282 75682
rect 53790 75630 53842 75682
rect 54686 75630 54738 75682
rect 55582 75630 55634 75682
rect 59054 75630 59106 75682
rect 61854 75630 61906 75682
rect 62638 75630 62690 75682
rect 65214 75630 65266 75682
rect 72606 75630 72658 75682
rect 75406 75630 75458 75682
rect 76190 75630 76242 75682
rect 76862 75630 76914 75682
rect 78094 75630 78146 75682
rect 4622 75518 4674 75570
rect 24222 75518 24274 75570
rect 59390 75518 59442 75570
rect 61182 75518 61234 75570
rect 75630 75518 75682 75570
rect 76526 75518 76578 75570
rect 77870 75518 77922 75570
rect 14254 75406 14306 75458
rect 14702 75406 14754 75458
rect 35982 75406 36034 75458
rect 42030 75406 42082 75458
rect 59726 75406 59778 75458
rect 60510 75406 60562 75458
rect 60846 75406 60898 75458
rect 61518 75406 61570 75458
rect 62190 75406 62242 75458
rect 65550 75406 65602 75458
rect 72942 75406 72994 75458
rect 77198 75406 77250 75458
rect 19838 75238 19890 75290
rect 19942 75238 19994 75290
rect 20046 75238 20098 75290
rect 50558 75238 50610 75290
rect 50662 75238 50714 75290
rect 50766 75238 50818 75290
rect 4622 75070 4674 75122
rect 12910 75070 12962 75122
rect 15262 75070 15314 75122
rect 23102 75070 23154 75122
rect 23550 75070 23602 75122
rect 34750 75070 34802 75122
rect 37438 75070 37490 75122
rect 38894 75070 38946 75122
rect 46846 75070 46898 75122
rect 52782 75070 52834 75122
rect 53566 75070 53618 75122
rect 54462 75070 54514 75122
rect 55358 75070 55410 75122
rect 57486 75070 57538 75122
rect 61294 75070 61346 75122
rect 61742 75070 61794 75122
rect 62190 75070 62242 75122
rect 74062 75070 74114 75122
rect 74510 75070 74562 75122
rect 74958 75070 75010 75122
rect 75406 75070 75458 75122
rect 76862 75070 76914 75122
rect 34974 74958 35026 75010
rect 75630 74958 75682 75010
rect 75966 74958 76018 75010
rect 77534 74958 77586 75010
rect 77870 74958 77922 75010
rect 4174 74846 4226 74898
rect 4846 74846 4898 74898
rect 13470 74846 13522 74898
rect 14702 74846 14754 74898
rect 22766 74846 22818 74898
rect 35198 74846 35250 74898
rect 60398 74846 60450 74898
rect 60846 74846 60898 74898
rect 77310 74846 77362 74898
rect 78094 74846 78146 74898
rect 2158 74734 2210 74786
rect 17950 74734 18002 74786
rect 18286 74734 18338 74786
rect 19406 74734 19458 74786
rect 19854 74734 19906 74786
rect 20414 74734 20466 74786
rect 35758 74734 35810 74786
rect 58046 74734 58098 74786
rect 76302 74734 76354 74786
rect 4478 74454 4530 74506
rect 4582 74454 4634 74506
rect 4686 74454 4738 74506
rect 35198 74454 35250 74506
rect 35302 74454 35354 74506
rect 35406 74454 35458 74506
rect 65918 74454 65970 74506
rect 66022 74454 66074 74506
rect 66126 74454 66178 74506
rect 19182 74286 19234 74338
rect 77758 74286 77810 74338
rect 77982 74286 78034 74338
rect 1934 74174 1986 74226
rect 11230 74174 11282 74226
rect 16046 74174 16098 74226
rect 58494 74174 58546 74226
rect 59166 74174 59218 74226
rect 75294 74174 75346 74226
rect 75742 74174 75794 74226
rect 76414 74174 76466 74226
rect 77982 74174 78034 74226
rect 4286 74062 4338 74114
rect 4846 74062 4898 74114
rect 12910 74062 12962 74114
rect 14030 74062 14082 74114
rect 17838 74062 17890 74114
rect 18174 74062 18226 74114
rect 76974 74062 77026 74114
rect 77534 74062 77586 74114
rect 4622 73950 4674 74002
rect 14366 73950 14418 74002
rect 22990 73950 23042 74002
rect 59502 73838 59554 73890
rect 19838 73670 19890 73722
rect 19942 73670 19994 73722
rect 20046 73670 20098 73722
rect 50558 73670 50610 73722
rect 50662 73670 50714 73722
rect 50766 73670 50818 73722
rect 76078 73502 76130 73554
rect 76526 73502 76578 73554
rect 76974 73502 77026 73554
rect 77422 73502 77474 73554
rect 78206 73502 78258 73554
rect 4622 73390 4674 73442
rect 12126 73390 12178 73442
rect 4286 73278 4338 73330
rect 4846 73278 4898 73330
rect 13918 73278 13970 73330
rect 16382 73278 16434 73330
rect 14590 73166 14642 73218
rect 18062 73166 18114 73218
rect 77646 73166 77698 73218
rect 1934 73054 1986 73106
rect 76638 73054 76690 73106
rect 77198 73054 77250 73106
rect 4478 72886 4530 72938
rect 4582 72886 4634 72938
rect 4686 72886 4738 72938
rect 35198 72886 35250 72938
rect 35302 72886 35354 72938
rect 35406 72886 35458 72938
rect 65918 72886 65970 72938
rect 66022 72886 66074 72938
rect 66126 72886 66178 72938
rect 1934 72606 1986 72658
rect 77198 72606 77250 72658
rect 3838 72494 3890 72546
rect 4958 72494 5010 72546
rect 77646 72382 77698 72434
rect 78206 72382 78258 72434
rect 4622 72270 4674 72322
rect 14142 72270 14194 72322
rect 77870 72270 77922 72322
rect 19838 72102 19890 72154
rect 19942 72102 19994 72154
rect 20046 72102 20098 72154
rect 50558 72102 50610 72154
rect 50662 72102 50714 72154
rect 50766 72102 50818 72154
rect 2494 71934 2546 71986
rect 3166 71934 3218 71986
rect 3502 71934 3554 71986
rect 3838 71822 3890 71874
rect 77870 71822 77922 71874
rect 2158 71710 2210 71762
rect 2942 71710 2994 71762
rect 77646 71710 77698 71762
rect 78206 71710 78258 71762
rect 1934 71598 1986 71650
rect 4478 71318 4530 71370
rect 4582 71318 4634 71370
rect 4686 71318 4738 71370
rect 35198 71318 35250 71370
rect 35302 71318 35354 71370
rect 35406 71318 35458 71370
rect 65918 71318 65970 71370
rect 66022 71318 66074 71370
rect 66126 71318 66178 71370
rect 1934 71038 1986 71090
rect 77758 71038 77810 71090
rect 3950 70926 4002 70978
rect 77422 70702 77474 70754
rect 78206 70702 78258 70754
rect 19838 70534 19890 70586
rect 19942 70534 19994 70586
rect 20046 70534 20098 70586
rect 50558 70534 50610 70586
rect 50662 70534 50714 70586
rect 50766 70534 50818 70586
rect 3838 70142 3890 70194
rect 1934 69918 1986 69970
rect 4478 69750 4530 69802
rect 4582 69750 4634 69802
rect 4686 69750 4738 69802
rect 35198 69750 35250 69802
rect 35302 69750 35354 69802
rect 35406 69750 35458 69802
rect 65918 69750 65970 69802
rect 66022 69750 66074 69802
rect 66126 69750 66178 69802
rect 2942 69358 2994 69410
rect 2382 69246 2434 69298
rect 2718 69246 2770 69298
rect 2046 69134 2098 69186
rect 77646 69134 77698 69186
rect 77870 69134 77922 69186
rect 78206 69134 78258 69186
rect 19838 68966 19890 69018
rect 19942 68966 19994 69018
rect 20046 68966 20098 69018
rect 50558 68966 50610 69018
rect 50662 68966 50714 69018
rect 50766 68966 50818 69018
rect 2046 68574 2098 68626
rect 78206 68574 78258 68626
rect 77422 68462 77474 68514
rect 77646 68462 77698 68514
rect 2718 68350 2770 68402
rect 4478 68182 4530 68234
rect 4582 68182 4634 68234
rect 4686 68182 4738 68234
rect 35198 68182 35250 68234
rect 35302 68182 35354 68234
rect 35406 68182 35458 68234
rect 65918 68182 65970 68234
rect 66022 68182 66074 68234
rect 66126 68182 66178 68234
rect 1934 67902 1986 67954
rect 4062 67790 4114 67842
rect 19838 67398 19890 67450
rect 19942 67398 19994 67450
rect 20046 67398 20098 67450
rect 50558 67398 50610 67450
rect 50662 67398 50714 67450
rect 50766 67398 50818 67450
rect 4062 67230 4114 67282
rect 2046 67118 2098 67170
rect 2718 67118 2770 67170
rect 3054 67118 3106 67170
rect 3726 67118 3778 67170
rect 77870 67118 77922 67170
rect 2382 67006 2434 67058
rect 3390 67006 3442 67058
rect 4286 67006 4338 67058
rect 78206 67006 78258 67058
rect 77646 66894 77698 66946
rect 4478 66614 4530 66666
rect 4582 66614 4634 66666
rect 4686 66614 4738 66666
rect 35198 66614 35250 66666
rect 35302 66614 35354 66666
rect 35406 66614 35458 66666
rect 65918 66614 65970 66666
rect 66022 66614 66074 66666
rect 66126 66614 66178 66666
rect 1934 66334 1986 66386
rect 3838 66222 3890 66274
rect 77646 66222 77698 66274
rect 77422 65998 77474 66050
rect 78206 65998 78258 66050
rect 19838 65830 19890 65882
rect 19942 65830 19994 65882
rect 20046 65830 20098 65882
rect 50558 65830 50610 65882
rect 50662 65830 50714 65882
rect 50766 65830 50818 65882
rect 2046 65438 2098 65490
rect 2718 65214 2770 65266
rect 4478 65046 4530 65098
rect 4582 65046 4634 65098
rect 4686 65046 4738 65098
rect 35198 65046 35250 65098
rect 35302 65046 35354 65098
rect 35406 65046 35458 65098
rect 65918 65046 65970 65098
rect 66022 65046 66074 65098
rect 66126 65046 66178 65098
rect 1934 64766 1986 64818
rect 3838 64654 3890 64706
rect 77646 64654 77698 64706
rect 77422 64542 77474 64594
rect 78206 64542 78258 64594
rect 19838 64262 19890 64314
rect 19942 64262 19994 64314
rect 20046 64262 20098 64314
rect 50558 64262 50610 64314
rect 50662 64262 50714 64314
rect 50766 64262 50818 64314
rect 2494 64094 2546 64146
rect 3502 64094 3554 64146
rect 2830 63982 2882 64034
rect 3166 63982 3218 64034
rect 77870 63982 77922 64034
rect 2270 63870 2322 63922
rect 3726 63870 3778 63922
rect 77646 63870 77698 63922
rect 78206 63870 78258 63922
rect 4478 63478 4530 63530
rect 4582 63478 4634 63530
rect 4686 63478 4738 63530
rect 35198 63478 35250 63530
rect 35302 63478 35354 63530
rect 35406 63478 35458 63530
rect 65918 63478 65970 63530
rect 66022 63478 66074 63530
rect 66126 63478 66178 63530
rect 1934 63198 1986 63250
rect 3838 63086 3890 63138
rect 77646 63086 77698 63138
rect 77422 62862 77474 62914
rect 78206 62862 78258 62914
rect 19838 62694 19890 62746
rect 19942 62694 19994 62746
rect 20046 62694 20098 62746
rect 50558 62694 50610 62746
rect 50662 62694 50714 62746
rect 50766 62694 50818 62746
rect 3838 62302 3890 62354
rect 1934 62078 1986 62130
rect 4478 61910 4530 61962
rect 4582 61910 4634 61962
rect 4686 61910 4738 61962
rect 35198 61910 35250 61962
rect 35302 61910 35354 61962
rect 35406 61910 35458 61962
rect 65918 61910 65970 61962
rect 66022 61910 66074 61962
rect 66126 61910 66178 61962
rect 2270 61518 2322 61570
rect 3614 61518 3666 61570
rect 2718 61406 2770 61458
rect 3054 61406 3106 61458
rect 3390 61406 3442 61458
rect 2046 61294 2098 61346
rect 4286 61294 4338 61346
rect 77646 61294 77698 61346
rect 77870 61294 77922 61346
rect 78206 61294 78258 61346
rect 19838 61126 19890 61178
rect 19942 61126 19994 61178
rect 20046 61126 20098 61178
rect 50558 61126 50610 61178
rect 50662 61126 50714 61178
rect 50766 61126 50818 61178
rect 77870 60846 77922 60898
rect 2046 60734 2098 60786
rect 77646 60734 77698 60786
rect 78206 60734 78258 60786
rect 2718 60510 2770 60562
rect 4478 60342 4530 60394
rect 4582 60342 4634 60394
rect 4686 60342 4738 60394
rect 35198 60342 35250 60394
rect 35302 60342 35354 60394
rect 35406 60342 35458 60394
rect 65918 60342 65970 60394
rect 66022 60342 66074 60394
rect 66126 60342 66178 60394
rect 1934 60062 1986 60114
rect 3838 59950 3890 60002
rect 19838 59558 19890 59610
rect 19942 59558 19994 59610
rect 20046 59558 20098 59610
rect 50558 59558 50610 59610
rect 50662 59558 50714 59610
rect 50766 59558 50818 59610
rect 2718 59390 2770 59442
rect 2046 59278 2098 59330
rect 2382 59166 2434 59218
rect 2942 59166 2994 59218
rect 3502 59166 3554 59218
rect 78206 59166 78258 59218
rect 77422 59054 77474 59106
rect 77646 59054 77698 59106
rect 4478 58774 4530 58826
rect 4582 58774 4634 58826
rect 4686 58774 4738 58826
rect 35198 58774 35250 58826
rect 35302 58774 35354 58826
rect 35406 58774 35458 58826
rect 65918 58774 65970 58826
rect 66022 58774 66074 58826
rect 66126 58774 66178 58826
rect 2046 58382 2098 58434
rect 2718 58158 2770 58210
rect 77646 58158 77698 58210
rect 77870 58158 77922 58210
rect 78206 58158 78258 58210
rect 19838 57990 19890 58042
rect 19942 57990 19994 58042
rect 20046 57990 20098 58042
rect 50558 57990 50610 58042
rect 50662 57990 50714 58042
rect 50766 57990 50818 58042
rect 4286 57598 4338 57650
rect 1934 57374 1986 57426
rect 4478 57206 4530 57258
rect 4582 57206 4634 57258
rect 4686 57206 4738 57258
rect 35198 57206 35250 57258
rect 35302 57206 35354 57258
rect 35406 57206 35458 57258
rect 65918 57206 65970 57258
rect 66022 57206 66074 57258
rect 66126 57206 66178 57258
rect 1934 56926 1986 56978
rect 3838 56814 3890 56866
rect 4846 56814 4898 56866
rect 4622 56702 4674 56754
rect 77646 56702 77698 56754
rect 78206 56702 78258 56754
rect 77870 56590 77922 56642
rect 19838 56422 19890 56474
rect 19942 56422 19994 56474
rect 20046 56422 20098 56474
rect 50558 56422 50610 56474
rect 50662 56422 50714 56474
rect 50766 56422 50818 56474
rect 2718 56254 2770 56306
rect 3726 56254 3778 56306
rect 2046 56142 2098 56194
rect 2382 56142 2434 56194
rect 3390 56142 3442 56194
rect 2942 56030 2994 56082
rect 78206 56030 78258 56082
rect 77422 55918 77474 55970
rect 77646 55918 77698 55970
rect 4478 55638 4530 55690
rect 4582 55638 4634 55690
rect 4686 55638 4738 55690
rect 35198 55638 35250 55690
rect 35302 55638 35354 55690
rect 35406 55638 35458 55690
rect 65918 55638 65970 55690
rect 66022 55638 66074 55690
rect 66126 55638 66178 55690
rect 2046 55246 2098 55298
rect 77646 55134 77698 55186
rect 78206 55134 78258 55186
rect 2718 55022 2770 55074
rect 77870 55022 77922 55074
rect 19838 54854 19890 54906
rect 19942 54854 19994 54906
rect 20046 54854 20098 54906
rect 50558 54854 50610 54906
rect 50662 54854 50714 54906
rect 50766 54854 50818 54906
rect 3838 54462 3890 54514
rect 1934 54238 1986 54290
rect 4478 54070 4530 54122
rect 4582 54070 4634 54122
rect 4686 54070 4738 54122
rect 35198 54070 35250 54122
rect 35302 54070 35354 54122
rect 35406 54070 35458 54122
rect 65918 54070 65970 54122
rect 66022 54070 66074 54122
rect 66126 54070 66178 54122
rect 2270 53678 2322 53730
rect 2942 53678 2994 53730
rect 1934 53566 1986 53618
rect 3166 53566 3218 53618
rect 3502 53566 3554 53618
rect 3838 53566 3890 53618
rect 78206 53566 78258 53618
rect 2494 53454 2546 53506
rect 77646 53454 77698 53506
rect 77870 53454 77922 53506
rect 19838 53286 19890 53338
rect 19942 53286 19994 53338
rect 20046 53286 20098 53338
rect 50558 53286 50610 53338
rect 50662 53286 50714 53338
rect 50766 53286 50818 53338
rect 77870 53006 77922 53058
rect 3950 52894 4002 52946
rect 78206 52894 78258 52946
rect 77646 52782 77698 52834
rect 1934 52670 1986 52722
rect 4478 52502 4530 52554
rect 4582 52502 4634 52554
rect 4686 52502 4738 52554
rect 35198 52502 35250 52554
rect 35302 52502 35354 52554
rect 35406 52502 35458 52554
rect 65918 52502 65970 52554
rect 66022 52502 66074 52554
rect 66126 52502 66178 52554
rect 1934 52222 1986 52274
rect 3838 52110 3890 52162
rect 19838 51718 19890 51770
rect 19942 51718 19994 51770
rect 20046 51718 20098 51770
rect 50558 51718 50610 51770
rect 50662 51718 50714 51770
rect 50766 51718 50818 51770
rect 2494 51550 2546 51602
rect 3502 51550 3554 51602
rect 2830 51438 2882 51490
rect 3838 51438 3890 51490
rect 77870 51438 77922 51490
rect 2270 51326 2322 51378
rect 3166 51326 3218 51378
rect 78206 51326 78258 51378
rect 77646 51214 77698 51266
rect 4478 50934 4530 50986
rect 4582 50934 4634 50986
rect 4686 50934 4738 50986
rect 35198 50934 35250 50986
rect 35302 50934 35354 50986
rect 35406 50934 35458 50986
rect 65918 50934 65970 50986
rect 66022 50934 66074 50986
rect 66126 50934 66178 50986
rect 1934 50654 1986 50706
rect 3838 50542 3890 50594
rect 77646 50430 77698 50482
rect 78206 50430 78258 50482
rect 77870 50318 77922 50370
rect 19838 50150 19890 50202
rect 19942 50150 19994 50202
rect 20046 50150 20098 50202
rect 50558 50150 50610 50202
rect 50662 50150 50714 50202
rect 50766 50150 50818 50202
rect 3838 49758 3890 49810
rect 1934 49534 1986 49586
rect 4478 49366 4530 49418
rect 4582 49366 4634 49418
rect 4686 49366 4738 49418
rect 35198 49366 35250 49418
rect 35302 49366 35354 49418
rect 35406 49366 35458 49418
rect 65918 49366 65970 49418
rect 66022 49366 66074 49418
rect 66126 49366 66178 49418
rect 1934 49086 1986 49138
rect 3838 48974 3890 49026
rect 77646 48862 77698 48914
rect 78206 48862 78258 48914
rect 77870 48750 77922 48802
rect 19838 48582 19890 48634
rect 19942 48582 19994 48634
rect 20046 48582 20098 48634
rect 50558 48582 50610 48634
rect 50662 48582 50714 48634
rect 50766 48582 50818 48634
rect 2718 48414 2770 48466
rect 3390 48414 3442 48466
rect 2046 48302 2098 48354
rect 77870 48302 77922 48354
rect 2382 48190 2434 48242
rect 2942 48190 2994 48242
rect 3614 48190 3666 48242
rect 77646 48190 77698 48242
rect 78206 48190 78258 48242
rect 4478 47798 4530 47850
rect 4582 47798 4634 47850
rect 4686 47798 4738 47850
rect 35198 47798 35250 47850
rect 35302 47798 35354 47850
rect 35406 47798 35458 47850
rect 65918 47798 65970 47850
rect 66022 47798 66074 47850
rect 66126 47798 66178 47850
rect 2046 47406 2098 47458
rect 78206 47294 78258 47346
rect 2718 47182 2770 47234
rect 77646 47182 77698 47234
rect 77870 47182 77922 47234
rect 19838 47014 19890 47066
rect 19942 47014 19994 47066
rect 20046 47014 20098 47066
rect 50558 47014 50610 47066
rect 50662 47014 50714 47066
rect 50766 47014 50818 47066
rect 3838 46622 3890 46674
rect 1934 46398 1986 46450
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 65918 46230 65970 46282
rect 66022 46230 66074 46282
rect 66126 46230 66178 46282
rect 2382 45838 2434 45890
rect 2718 45838 2770 45890
rect 3614 45838 3666 45890
rect 4286 45838 4338 45890
rect 3054 45726 3106 45778
rect 3390 45726 3442 45778
rect 78206 45726 78258 45778
rect 2046 45614 2098 45666
rect 77646 45614 77698 45666
rect 77870 45614 77922 45666
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 50558 45446 50610 45498
rect 50662 45446 50714 45498
rect 50766 45446 50818 45498
rect 77870 45166 77922 45218
rect 2046 45054 2098 45106
rect 78206 45054 78258 45106
rect 77646 44942 77698 44994
rect 2718 44830 2770 44882
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 65918 44662 65970 44714
rect 66022 44662 66074 44714
rect 66126 44662 66178 44714
rect 2046 44270 2098 44322
rect 2718 44046 2770 44098
rect 78318 44046 78370 44098
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 50558 43878 50610 43930
rect 50662 43878 50714 43930
rect 50766 43878 50818 43930
rect 2046 43710 2098 43762
rect 2718 43598 2770 43650
rect 2270 43486 2322 43538
rect 3054 43486 3106 43538
rect 56590 43486 56642 43538
rect 77086 43486 77138 43538
rect 77422 43486 77474 43538
rect 77646 43486 77698 43538
rect 57038 43374 57090 43426
rect 76974 43374 77026 43426
rect 77310 43374 77362 43426
rect 78206 43374 78258 43426
rect 76638 43262 76690 43314
rect 76974 43262 77026 43314
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 65918 43094 65970 43146
rect 66022 43094 66074 43146
rect 66126 43094 66178 43146
rect 1934 42814 1986 42866
rect 56030 42814 56082 42866
rect 57262 42814 57314 42866
rect 58158 42814 58210 42866
rect 62302 42814 62354 42866
rect 75742 42814 75794 42866
rect 3838 42702 3890 42754
rect 55582 42702 55634 42754
rect 76526 42702 76578 42754
rect 77534 42702 77586 42754
rect 78094 42702 78146 42754
rect 76974 42590 77026 42642
rect 77310 42590 77362 42642
rect 56702 42478 56754 42530
rect 57598 42478 57650 42530
rect 76302 42478 76354 42530
rect 77198 42478 77250 42530
rect 77870 42478 77922 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 50558 42310 50610 42362
rect 50662 42310 50714 42362
rect 50766 42310 50818 42362
rect 55694 42142 55746 42194
rect 56590 42142 56642 42194
rect 57486 42142 57538 42194
rect 75294 42030 75346 42082
rect 3838 41918 3890 41970
rect 4734 41918 4786 41970
rect 60622 41918 60674 41970
rect 61070 41918 61122 41970
rect 61630 41918 61682 41970
rect 62526 41918 62578 41970
rect 62862 41918 62914 41970
rect 63198 41918 63250 41970
rect 64430 41918 64482 41970
rect 65438 41918 65490 41970
rect 65886 41918 65938 41970
rect 74062 41918 74114 41970
rect 74958 41918 75010 41970
rect 75630 41918 75682 41970
rect 54910 41806 54962 41858
rect 55134 41806 55186 41858
rect 57150 41806 57202 41858
rect 58046 41806 58098 41858
rect 60174 41806 60226 41858
rect 62078 41806 62130 41858
rect 62750 41806 62802 41858
rect 64990 41806 65042 41858
rect 69806 41806 69858 41858
rect 70254 41806 70306 41858
rect 70702 41806 70754 41858
rect 71150 41806 71202 41858
rect 74734 41806 74786 41858
rect 77982 41806 78034 41858
rect 1934 41694 1986 41746
rect 55358 41694 55410 41746
rect 56926 41694 56978 41746
rect 57822 41694 57874 41746
rect 69806 41694 69858 41746
rect 70142 41694 70194 41746
rect 71038 41694 71090 41746
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 65918 41526 65970 41578
rect 66022 41526 66074 41578
rect 66126 41526 66178 41578
rect 55582 41358 55634 41410
rect 55918 41358 55970 41410
rect 71150 41358 71202 41410
rect 71598 41358 71650 41410
rect 71710 41358 71762 41410
rect 74398 41358 74450 41410
rect 74734 41358 74786 41410
rect 1934 41246 1986 41298
rect 4734 41246 4786 41298
rect 56366 41246 56418 41298
rect 58942 41246 58994 41298
rect 60622 41246 60674 41298
rect 62414 41246 62466 41298
rect 64990 41246 65042 41298
rect 70478 41246 70530 41298
rect 71374 41246 71426 41298
rect 74174 41246 74226 41298
rect 75070 41246 75122 41298
rect 75294 41246 75346 41298
rect 78094 41246 78146 41298
rect 4174 41134 4226 41186
rect 55358 41134 55410 41186
rect 58494 41134 58546 41186
rect 59390 41134 59442 41186
rect 59950 41134 60002 41186
rect 60510 41134 60562 41186
rect 61630 41134 61682 41186
rect 62526 41134 62578 41186
rect 62862 41134 62914 41186
rect 63422 41134 63474 41186
rect 64318 41134 64370 41186
rect 65662 41134 65714 41186
rect 66782 41134 66834 41186
rect 70142 41134 70194 41186
rect 70926 41134 70978 41186
rect 73614 41134 73666 41186
rect 76078 41134 76130 41186
rect 76526 41134 76578 41186
rect 76974 41134 77026 41186
rect 77534 41134 77586 41186
rect 58158 41022 58210 41074
rect 59166 41022 59218 41074
rect 60958 41022 61010 41074
rect 61966 41022 62018 41074
rect 63534 41022 63586 41074
rect 65774 41022 65826 41074
rect 69582 41022 69634 41074
rect 73278 41022 73330 41074
rect 73838 41022 73890 41074
rect 76750 41022 76802 41074
rect 77422 41022 77474 41074
rect 55022 40910 55074 40962
rect 57150 40910 57202 40962
rect 64318 40910 64370 40962
rect 66558 40910 66610 40962
rect 69022 40910 69074 40962
rect 69246 40910 69298 40962
rect 73390 40910 73442 40962
rect 75630 40910 75682 40962
rect 76302 40910 76354 40962
rect 77198 40910 77250 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 50558 40742 50610 40794
rect 50662 40742 50714 40794
rect 50766 40742 50818 40794
rect 2270 40574 2322 40626
rect 5406 40574 5458 40626
rect 59950 40574 60002 40626
rect 61518 40574 61570 40626
rect 64654 40574 64706 40626
rect 66894 40574 66946 40626
rect 67454 40574 67506 40626
rect 67902 40574 67954 40626
rect 71374 40574 71426 40626
rect 72942 40574 72994 40626
rect 73950 40574 74002 40626
rect 74622 40574 74674 40626
rect 75182 40574 75234 40626
rect 4062 40462 4114 40514
rect 4510 40462 4562 40514
rect 60734 40462 60786 40514
rect 62974 40462 63026 40514
rect 63534 40462 63586 40514
rect 65102 40462 65154 40514
rect 66334 40462 66386 40514
rect 69358 40462 69410 40514
rect 70926 40462 70978 40514
rect 73614 40462 73666 40514
rect 74286 40462 74338 40514
rect 76638 40462 76690 40514
rect 1710 40350 1762 40402
rect 2606 40350 2658 40402
rect 3166 40350 3218 40402
rect 3502 40350 3554 40402
rect 4958 40350 5010 40402
rect 60062 40350 60114 40402
rect 60510 40350 60562 40402
rect 61742 40350 61794 40402
rect 62302 40350 62354 40402
rect 62638 40350 62690 40402
rect 63198 40350 63250 40402
rect 63758 40350 63810 40402
rect 64430 40350 64482 40402
rect 65550 40350 65602 40402
rect 65886 40350 65938 40402
rect 66782 40350 66834 40402
rect 68238 40350 68290 40402
rect 68574 40350 68626 40402
rect 69694 40350 69746 40402
rect 70142 40350 70194 40402
rect 70702 40350 70754 40402
rect 73390 40350 73442 40402
rect 77870 40350 77922 40402
rect 62750 40238 62802 40290
rect 69470 40238 69522 40290
rect 72494 40238 72546 40290
rect 74958 40126 75010 40178
rect 75294 40126 75346 40178
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 65918 39958 65970 40010
rect 66022 39958 66074 40010
rect 66126 39958 66178 40010
rect 1934 39678 1986 39730
rect 61294 39678 61346 39730
rect 61854 39678 61906 39730
rect 63422 39678 63474 39730
rect 67118 39678 67170 39730
rect 71934 39678 71986 39730
rect 72942 39678 72994 39730
rect 74622 39678 74674 39730
rect 76750 39678 76802 39730
rect 3838 39566 3890 39618
rect 4734 39566 4786 39618
rect 65214 39566 65266 39618
rect 65550 39566 65602 39618
rect 66670 39566 66722 39618
rect 68350 39566 68402 39618
rect 69246 39566 69298 39618
rect 70366 39566 70418 39618
rect 70590 39566 70642 39618
rect 71374 39566 71426 39618
rect 72382 39566 72434 39618
rect 73166 39566 73218 39618
rect 73614 39566 73666 39618
rect 74062 39566 74114 39618
rect 75070 39566 75122 39618
rect 75406 39566 75458 39618
rect 75518 39566 75570 39618
rect 76526 39566 76578 39618
rect 77310 39566 77362 39618
rect 78094 39566 78146 39618
rect 65774 39454 65826 39506
rect 68462 39454 68514 39506
rect 70030 39454 70082 39506
rect 70926 39454 70978 39506
rect 71262 39454 71314 39506
rect 76414 39454 76466 39506
rect 77870 39454 77922 39506
rect 64654 39342 64706 39394
rect 66446 39342 66498 39394
rect 67566 39342 67618 39394
rect 69358 39342 69410 39394
rect 70254 39342 70306 39394
rect 71150 39342 71202 39394
rect 75294 39342 75346 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 50558 39174 50610 39226
rect 50662 39174 50714 39226
rect 50766 39174 50818 39226
rect 42030 39006 42082 39058
rect 43598 39006 43650 39058
rect 62190 39006 62242 39058
rect 65326 39006 65378 39058
rect 69246 39006 69298 39058
rect 71374 39006 71426 39058
rect 73502 39006 73554 39058
rect 74398 39006 74450 39058
rect 41246 38894 41298 38946
rect 41470 38894 41522 38946
rect 42590 38894 42642 38946
rect 43038 38894 43090 38946
rect 43262 38894 43314 38946
rect 61854 38894 61906 38946
rect 67118 38894 67170 38946
rect 68014 38894 68066 38946
rect 69694 38894 69746 38946
rect 70926 38894 70978 38946
rect 72718 38894 72770 38946
rect 73054 38894 73106 38946
rect 73278 38894 73330 38946
rect 75182 38894 75234 38946
rect 76190 38894 76242 38946
rect 77646 38894 77698 38946
rect 2046 38782 2098 38834
rect 41582 38782 41634 38834
rect 42030 38782 42082 38834
rect 42926 38782 42978 38834
rect 44046 38782 44098 38834
rect 62526 38782 62578 38834
rect 65886 38782 65938 38834
rect 66334 38782 66386 38834
rect 67342 38782 67394 38834
rect 68238 38782 68290 38834
rect 68574 38782 68626 38834
rect 70366 38782 70418 38834
rect 70702 38782 70754 38834
rect 72494 38782 72546 38834
rect 73726 38782 73778 38834
rect 74174 38782 74226 38834
rect 74846 38782 74898 38834
rect 75630 38782 75682 38834
rect 75966 38782 76018 38834
rect 76638 38782 76690 38834
rect 77086 38782 77138 38834
rect 77534 38782 77586 38834
rect 78094 38782 78146 38834
rect 3390 38670 3442 38722
rect 41134 38670 41186 38722
rect 66670 38670 66722 38722
rect 67902 38670 67954 38722
rect 70478 38670 70530 38722
rect 76414 38670 76466 38722
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 65918 38390 65970 38442
rect 66022 38390 66074 38442
rect 66126 38390 66178 38442
rect 2046 38110 2098 38162
rect 2942 38110 2994 38162
rect 67230 38110 67282 38162
rect 70590 38110 70642 38162
rect 72942 38110 72994 38162
rect 75630 38110 75682 38162
rect 77534 38110 77586 38162
rect 78206 38110 78258 38162
rect 2494 37998 2546 38050
rect 68350 37998 68402 38050
rect 69246 37998 69298 38050
rect 69806 37998 69858 38050
rect 71038 37998 71090 38050
rect 71262 37998 71314 38050
rect 72158 37998 72210 38050
rect 73166 37998 73218 38050
rect 73278 37998 73330 38050
rect 74286 37998 74338 38050
rect 74622 37998 74674 38050
rect 75070 37998 75122 38050
rect 76190 37998 76242 38050
rect 76638 37998 76690 38050
rect 77086 37998 77138 38050
rect 68462 37886 68514 37938
rect 70142 37886 70194 37938
rect 71598 37886 71650 37938
rect 72830 37886 72882 37938
rect 73726 37886 73778 37938
rect 73950 37886 74002 37938
rect 74958 37886 75010 37938
rect 76526 37886 76578 37938
rect 77310 37886 77362 37938
rect 77646 37886 77698 37938
rect 67790 37774 67842 37826
rect 69246 37774 69298 37826
rect 71486 37774 71538 37826
rect 72494 37774 72546 37826
rect 74062 37774 74114 37826
rect 74734 37774 74786 37826
rect 76302 37774 76354 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 50558 37606 50610 37658
rect 50662 37606 50714 37658
rect 50766 37606 50818 37658
rect 68126 37438 68178 37490
rect 68686 37438 68738 37490
rect 69022 37438 69074 37490
rect 69694 37438 69746 37490
rect 70926 37438 70978 37490
rect 71598 37438 71650 37490
rect 75070 37438 75122 37490
rect 76414 37438 76466 37490
rect 2046 37326 2098 37378
rect 70590 37326 70642 37378
rect 71262 37326 71314 37378
rect 72270 37326 72322 37378
rect 74510 37326 74562 37378
rect 74846 37326 74898 37378
rect 75406 37326 75458 37378
rect 75966 37326 76018 37378
rect 1710 37214 1762 37266
rect 69358 37214 69410 37266
rect 72494 37214 72546 37266
rect 72718 37214 72770 37266
rect 73054 37214 73106 37266
rect 73390 37214 73442 37266
rect 73614 37214 73666 37266
rect 74286 37214 74338 37266
rect 75182 37214 75234 37266
rect 76190 37214 76242 37266
rect 76638 37214 76690 37266
rect 77198 37214 77250 37266
rect 77870 37214 77922 37266
rect 2494 37102 2546 37154
rect 72382 37102 72434 37154
rect 73278 37102 73330 37154
rect 77310 37102 77362 37154
rect 77422 36990 77474 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 65918 36822 65970 36874
rect 66022 36822 66074 36874
rect 66126 36822 66178 36874
rect 72494 36654 72546 36706
rect 73278 36654 73330 36706
rect 74958 36654 75010 36706
rect 77870 36654 77922 36706
rect 71262 36542 71314 36594
rect 71934 36542 71986 36594
rect 72942 36542 72994 36594
rect 73278 36542 73330 36594
rect 74846 36542 74898 36594
rect 76414 36542 76466 36594
rect 76750 36542 76802 36594
rect 77982 36542 78034 36594
rect 72494 36430 72546 36482
rect 74622 36430 74674 36482
rect 75406 36430 75458 36482
rect 76190 36430 76242 36482
rect 76862 36430 76914 36482
rect 78206 36430 78258 36482
rect 1710 36318 1762 36370
rect 44830 36318 44882 36370
rect 45390 36318 45442 36370
rect 73950 36318 74002 36370
rect 74398 36318 74450 36370
rect 2046 36206 2098 36258
rect 2494 36206 2546 36258
rect 44942 36206 44994 36258
rect 69022 36206 69074 36258
rect 75630 36206 75682 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 50558 36038 50610 36090
rect 50662 36038 50714 36090
rect 50766 36038 50818 36090
rect 44270 35870 44322 35922
rect 54350 35870 54402 35922
rect 72942 35870 72994 35922
rect 77646 35870 77698 35922
rect 78206 35870 78258 35922
rect 44606 35758 44658 35810
rect 45838 35758 45890 35810
rect 46622 35758 46674 35810
rect 46958 35758 47010 35810
rect 73278 35758 73330 35810
rect 73614 35758 73666 35810
rect 74174 35758 74226 35810
rect 74510 35758 74562 35810
rect 75182 35758 75234 35810
rect 76078 35758 76130 35810
rect 76526 35758 76578 35810
rect 76862 35758 76914 35810
rect 44718 35646 44770 35698
rect 45390 35646 45442 35698
rect 45950 35646 46002 35698
rect 46398 35646 46450 35698
rect 72606 35646 72658 35698
rect 73950 35646 74002 35698
rect 74734 35646 74786 35698
rect 75294 35646 75346 35698
rect 75742 35646 75794 35698
rect 76974 35646 77026 35698
rect 77870 35646 77922 35698
rect 45614 35534 45666 35586
rect 46846 35534 46898 35586
rect 71710 35534 71762 35586
rect 74398 35534 74450 35586
rect 74958 35534 75010 35586
rect 76638 35534 76690 35586
rect 54014 35422 54066 35474
rect 54350 35422 54402 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 65918 35254 65970 35306
rect 66022 35254 66074 35306
rect 66126 35254 66178 35306
rect 77870 35086 77922 35138
rect 55582 34974 55634 35026
rect 75406 34974 75458 35026
rect 76526 34974 76578 35026
rect 76750 34974 76802 35026
rect 78094 34974 78146 35026
rect 44942 34862 44994 34914
rect 45390 34862 45442 34914
rect 45614 34862 45666 34914
rect 45838 34862 45890 34914
rect 45950 34862 46002 34914
rect 53566 34862 53618 34914
rect 54462 34862 54514 34914
rect 71262 34862 71314 34914
rect 71598 34862 71650 34914
rect 71822 34862 71874 34914
rect 72158 34862 72210 34914
rect 72830 34862 72882 34914
rect 73054 34862 73106 34914
rect 73278 34862 73330 34914
rect 73502 34862 73554 34914
rect 73838 34862 73890 34914
rect 74062 34862 74114 34914
rect 74734 34862 74786 34914
rect 76078 34862 76130 34914
rect 76862 34862 76914 34914
rect 78206 34862 78258 34914
rect 1710 34750 1762 34802
rect 2494 34750 2546 34802
rect 44830 34750 44882 34802
rect 54014 34750 54066 34802
rect 54798 34750 54850 34802
rect 70926 34750 70978 34802
rect 72382 34750 72434 34802
rect 75294 34750 75346 34802
rect 2046 34638 2098 34690
rect 44382 34638 44434 34690
rect 53566 34638 53618 34690
rect 55022 34638 55074 34690
rect 71374 34638 71426 34690
rect 71934 34638 71986 34690
rect 73054 34638 73106 34690
rect 73726 34638 73778 34690
rect 74958 34638 75010 34690
rect 75518 34638 75570 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 50558 34470 50610 34522
rect 50662 34470 50714 34522
rect 50766 34470 50818 34522
rect 55470 34302 55522 34354
rect 71822 34302 71874 34354
rect 72494 34302 72546 34354
rect 73390 34302 73442 34354
rect 73838 34302 73890 34354
rect 75966 34302 76018 34354
rect 78206 34302 78258 34354
rect 2046 34190 2098 34242
rect 44158 34190 44210 34242
rect 44382 34190 44434 34242
rect 53342 34190 53394 34242
rect 54574 34190 54626 34242
rect 71374 34190 71426 34242
rect 76302 34190 76354 34242
rect 76638 34190 76690 34242
rect 77534 34190 77586 34242
rect 1710 34078 1762 34130
rect 53006 34078 53058 34130
rect 54238 34078 54290 34130
rect 72718 34078 72770 34130
rect 73054 34078 73106 34130
rect 74734 34078 74786 34130
rect 75070 34078 75122 34130
rect 76414 34078 76466 34130
rect 2494 33966 2546 34018
rect 54574 33966 54626 34018
rect 44494 33854 44546 33906
rect 53118 33854 53170 33906
rect 76862 34078 76914 34130
rect 77086 34078 77138 34130
rect 77646 34078 77698 34130
rect 74846 33966 74898 34018
rect 77310 33966 77362 34018
rect 73614 33854 73666 33906
rect 74734 33854 74786 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 65918 33686 65970 33738
rect 66022 33686 66074 33738
rect 66126 33686 66178 33738
rect 76750 33518 76802 33570
rect 54014 33406 54066 33458
rect 72718 33406 72770 33458
rect 73390 33406 73442 33458
rect 74398 33406 74450 33458
rect 74846 33406 74898 33458
rect 76526 33406 76578 33458
rect 78206 33406 78258 33458
rect 45390 33294 45442 33346
rect 45838 33294 45890 33346
rect 72046 33294 72098 33346
rect 72158 33294 72210 33346
rect 73614 33294 73666 33346
rect 74622 33294 74674 33346
rect 75294 33294 75346 33346
rect 77534 33294 77586 33346
rect 46062 33182 46114 33234
rect 46398 33182 46450 33234
rect 71710 33182 71762 33234
rect 76862 33182 76914 33234
rect 77086 33182 77138 33234
rect 77758 33182 77810 33234
rect 1710 33070 1762 33122
rect 2046 33070 2098 33122
rect 2494 33070 2546 33122
rect 45726 33070 45778 33122
rect 46734 33070 46786 33122
rect 71822 33070 71874 33122
rect 73950 33070 74002 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 50558 32902 50610 32954
rect 50662 32902 50714 32954
rect 50766 32902 50818 32954
rect 46062 32734 46114 32786
rect 74846 32734 74898 32786
rect 75630 32734 75682 32786
rect 76750 32734 76802 32786
rect 77870 32734 77922 32786
rect 45390 32622 45442 32674
rect 46734 32622 46786 32674
rect 71374 32622 71426 32674
rect 72606 32622 72658 32674
rect 73166 32622 73218 32674
rect 74286 32622 74338 32674
rect 74958 32622 75010 32674
rect 76862 32622 76914 32674
rect 45838 32510 45890 32562
rect 46510 32510 46562 32562
rect 71262 32510 71314 32562
rect 71710 32510 71762 32562
rect 72158 32510 72210 32562
rect 72830 32510 72882 32562
rect 73390 32510 73442 32562
rect 74062 32510 74114 32562
rect 74622 32510 74674 32562
rect 75294 32510 75346 32562
rect 76414 32510 76466 32562
rect 76974 32510 77026 32562
rect 77646 32510 77698 32562
rect 78206 32510 78258 32562
rect 45054 32398 45106 32450
rect 71598 32398 71650 32450
rect 72382 32398 72434 32450
rect 76078 32398 76130 32450
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 65918 32118 65970 32170
rect 66022 32118 66074 32170
rect 66126 32118 66178 32170
rect 72606 31950 72658 32002
rect 73166 31950 73218 32002
rect 76974 31950 77026 32002
rect 77198 31950 77250 32002
rect 77534 31950 77586 32002
rect 77870 31950 77922 32002
rect 45278 31838 45330 31890
rect 73166 31838 73218 31890
rect 74734 31838 74786 31890
rect 77310 31838 77362 31890
rect 44942 31726 44994 31778
rect 45726 31726 45778 31778
rect 45950 31726 46002 31778
rect 46286 31726 46338 31778
rect 51438 31726 51490 31778
rect 52782 31726 52834 31778
rect 72046 31726 72098 31778
rect 73278 31726 73330 31778
rect 75070 31726 75122 31778
rect 76190 31726 76242 31778
rect 76414 31726 76466 31778
rect 76638 31726 76690 31778
rect 1710 31614 1762 31666
rect 2046 31614 2098 31666
rect 44382 31614 44434 31666
rect 44830 31614 44882 31666
rect 45390 31614 45442 31666
rect 46174 31614 46226 31666
rect 51550 31614 51602 31666
rect 72718 31614 72770 31666
rect 2494 31502 2546 31554
rect 51774 31502 51826 31554
rect 73726 31502 73778 31554
rect 73838 31502 73890 31554
rect 73950 31502 74002 31554
rect 75406 31502 75458 31554
rect 76302 31502 76354 31554
rect 77758 31502 77810 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 50558 31334 50610 31386
rect 50662 31334 50714 31386
rect 50766 31334 50818 31386
rect 53678 31166 53730 31218
rect 73390 31166 73442 31218
rect 74062 31166 74114 31218
rect 74846 31166 74898 31218
rect 75182 31166 75234 31218
rect 77310 31166 77362 31218
rect 77534 31166 77586 31218
rect 2046 31054 2098 31106
rect 44158 31054 44210 31106
rect 44382 31054 44434 31106
rect 45502 31054 45554 31106
rect 46174 31054 46226 31106
rect 47070 31054 47122 31106
rect 51774 31054 51826 31106
rect 52558 31054 52610 31106
rect 72606 31054 72658 31106
rect 74174 31054 74226 31106
rect 75854 31054 75906 31106
rect 76414 31054 76466 31106
rect 77870 31054 77922 31106
rect 1710 30942 1762 30994
rect 45278 30942 45330 30994
rect 45726 30942 45778 30994
rect 46286 30942 46338 30994
rect 46846 30942 46898 30994
rect 51438 30942 51490 30994
rect 52446 30942 52498 30994
rect 72270 30942 72322 30994
rect 72718 30942 72770 30994
rect 73614 30942 73666 30994
rect 74286 30942 74338 30994
rect 75518 30942 75570 30994
rect 76078 30942 76130 30994
rect 76750 30942 76802 30994
rect 2494 30830 2546 30882
rect 45950 30830 46002 30882
rect 51998 30830 52050 30882
rect 52894 30830 52946 30882
rect 72382 30830 72434 30882
rect 75630 30830 75682 30882
rect 44494 30718 44546 30770
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 65918 30550 65970 30602
rect 66022 30550 66074 30602
rect 66126 30550 66178 30602
rect 72830 30382 72882 30434
rect 52894 30270 52946 30322
rect 71934 30270 71986 30322
rect 73614 30270 73666 30322
rect 74622 30270 74674 30322
rect 45726 30158 45778 30210
rect 46174 30158 46226 30210
rect 46286 30158 46338 30210
rect 46734 30158 46786 30210
rect 46958 30158 47010 30210
rect 47182 30158 47234 30210
rect 50878 30158 50930 30210
rect 72046 30158 72098 30210
rect 72494 30158 72546 30210
rect 72942 30158 72994 30210
rect 73726 30158 73778 30210
rect 75070 30158 75122 30210
rect 75406 30158 75458 30210
rect 76078 30158 76130 30210
rect 76638 30158 76690 30210
rect 77086 30158 77138 30210
rect 78206 30158 78258 30210
rect 47294 30046 47346 30098
rect 51214 30046 51266 30098
rect 51998 30046 52050 30098
rect 71486 30046 71538 30098
rect 76526 30046 76578 30098
rect 77422 30046 77474 30098
rect 77870 30046 77922 30098
rect 46062 29934 46114 29986
rect 51438 29934 51490 29986
rect 71150 29934 71202 29986
rect 71822 29934 71874 29986
rect 75630 29934 75682 29986
rect 76302 29934 76354 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 50558 29766 50610 29818
rect 50662 29766 50714 29818
rect 50766 29766 50818 29818
rect 44942 29598 44994 29650
rect 71374 29598 71426 29650
rect 71822 29598 71874 29650
rect 76302 29598 76354 29650
rect 77646 29598 77698 29650
rect 2046 29486 2098 29538
rect 44606 29486 44658 29538
rect 44830 29486 44882 29538
rect 73166 29486 73218 29538
rect 75854 29486 75906 29538
rect 76078 29486 76130 29538
rect 1710 29374 1762 29426
rect 72718 29374 72770 29426
rect 72830 29374 72882 29426
rect 73502 29374 73554 29426
rect 74398 29374 74450 29426
rect 74846 29374 74898 29426
rect 75518 29374 75570 29426
rect 75630 29374 75682 29426
rect 2494 29262 2546 29314
rect 70926 29262 70978 29314
rect 73054 29262 73106 29314
rect 77758 29598 77810 29650
rect 76638 29486 76690 29538
rect 76974 29486 77026 29538
rect 77086 29374 77138 29426
rect 76750 29262 76802 29314
rect 72158 29150 72210 29202
rect 72494 29150 72546 29202
rect 74062 29150 74114 29202
rect 76302 29150 76354 29202
rect 77534 29150 77586 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 65918 28982 65970 29034
rect 66022 28982 66074 29034
rect 66126 28982 66178 29034
rect 70814 28814 70866 28866
rect 37102 28702 37154 28754
rect 70590 28702 70642 28754
rect 73502 28702 73554 28754
rect 76302 28702 76354 28754
rect 78206 28702 78258 28754
rect 1710 28590 1762 28642
rect 2494 28590 2546 28642
rect 70366 28590 70418 28642
rect 70702 28590 70754 28642
rect 72494 28590 72546 28642
rect 73726 28590 73778 28642
rect 74398 28590 74450 28642
rect 75070 28590 75122 28642
rect 76078 28590 76130 28642
rect 76526 28590 76578 28642
rect 76974 28590 77026 28642
rect 77422 28590 77474 28642
rect 77646 28590 77698 28642
rect 2046 28478 2098 28530
rect 71822 28478 71874 28530
rect 72158 28478 72210 28530
rect 72830 28478 72882 28530
rect 74734 28478 74786 28530
rect 76750 28478 76802 28530
rect 74062 28366 74114 28418
rect 75406 28366 75458 28418
rect 77198 28366 77250 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 50558 28198 50610 28250
rect 50662 28198 50714 28250
rect 50766 28198 50818 28250
rect 36990 28030 37042 28082
rect 37438 28030 37490 28082
rect 38670 28030 38722 28082
rect 39342 28030 39394 28082
rect 41022 28030 41074 28082
rect 42478 28030 42530 28082
rect 44718 28030 44770 28082
rect 72606 28030 72658 28082
rect 77646 28030 77698 28082
rect 35086 27918 35138 27970
rect 36430 27918 36482 27970
rect 38222 27918 38274 27970
rect 41582 27918 41634 27970
rect 45054 27918 45106 27970
rect 72830 27918 72882 27970
rect 73726 27918 73778 27970
rect 75182 27918 75234 27970
rect 75854 27918 75906 27970
rect 76414 27918 76466 27970
rect 76638 27918 76690 27970
rect 76750 27918 76802 27970
rect 77534 27918 77586 27970
rect 77758 27918 77810 27970
rect 35534 27806 35586 27858
rect 35982 27806 36034 27858
rect 37774 27806 37826 27858
rect 38782 27806 38834 27858
rect 40350 27806 40402 27858
rect 41022 27806 41074 27858
rect 41470 27806 41522 27858
rect 70254 27806 70306 27858
rect 70702 27806 70754 27858
rect 70926 27806 70978 27858
rect 73166 27806 73218 27858
rect 73390 27806 73442 27858
rect 73950 27806 74002 27858
rect 74286 27806 74338 27858
rect 74734 27806 74786 27858
rect 74958 27806 75010 27858
rect 75630 27806 75682 27858
rect 76862 27806 76914 27858
rect 77086 27806 77138 27858
rect 36094 27694 36146 27746
rect 70142 27694 70194 27746
rect 70814 27694 70866 27746
rect 71486 27694 71538 27746
rect 72942 27694 72994 27746
rect 73838 27694 73890 27746
rect 75070 27694 75122 27746
rect 45166 27582 45218 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 65918 27414 65970 27466
rect 66022 27414 66074 27466
rect 66126 27414 66178 27466
rect 45166 27246 45218 27298
rect 46286 27246 46338 27298
rect 49646 27246 49698 27298
rect 76862 27246 76914 27298
rect 77198 27246 77250 27298
rect 35870 27134 35922 27186
rect 38558 27134 38610 27186
rect 39678 27134 39730 27186
rect 42590 27134 42642 27186
rect 43038 27134 43090 27186
rect 44830 27134 44882 27186
rect 45390 27134 45442 27186
rect 45838 27134 45890 27186
rect 46622 27134 46674 27186
rect 50206 27134 50258 27186
rect 71822 27134 71874 27186
rect 72270 27134 72322 27186
rect 72718 27134 72770 27186
rect 75406 27134 75458 27186
rect 33854 27022 33906 27074
rect 34862 27022 34914 27074
rect 35534 27022 35586 27074
rect 36206 27022 36258 27074
rect 37550 27022 37602 27074
rect 38110 27022 38162 27074
rect 38782 27022 38834 27074
rect 39790 27022 39842 27074
rect 40686 27022 40738 27074
rect 41022 27022 41074 27074
rect 42142 27022 42194 27074
rect 46398 27022 46450 27074
rect 47294 27022 47346 27074
rect 47518 27022 47570 27074
rect 47854 27022 47906 27074
rect 48974 27022 49026 27074
rect 49534 27022 49586 27074
rect 70702 27022 70754 27074
rect 71038 27022 71090 27074
rect 73166 27022 73218 27074
rect 73502 27022 73554 27074
rect 74062 27022 74114 27074
rect 75294 27022 75346 27074
rect 76414 27022 76466 27074
rect 77870 27022 77922 27074
rect 1710 26910 1762 26962
rect 2046 26910 2098 26962
rect 2494 26910 2546 26962
rect 34302 26910 34354 26962
rect 36430 26910 36482 26962
rect 36990 26910 37042 26962
rect 38222 26910 38274 26962
rect 40014 26910 40066 26962
rect 42030 26910 42082 26962
rect 44942 26910 44994 26962
rect 46846 26910 46898 26962
rect 47070 26910 47122 26962
rect 47742 26910 47794 26962
rect 49086 26910 49138 26962
rect 49646 26910 49698 26962
rect 50654 26910 50706 26962
rect 70590 26910 70642 26962
rect 72942 26910 72994 26962
rect 74622 26910 74674 26962
rect 74958 26910 75010 26962
rect 75630 26910 75682 26962
rect 76190 26910 76242 26962
rect 77534 26910 77586 26962
rect 34862 26798 34914 26850
rect 41134 26798 41186 26850
rect 49310 26798 49362 26850
rect 70478 26798 70530 26850
rect 73166 26798 73218 26850
rect 76974 26798 77026 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 50558 26630 50610 26682
rect 50662 26630 50714 26682
rect 50766 26630 50818 26682
rect 36654 26462 36706 26514
rect 42366 26462 42418 26514
rect 44494 26462 44546 26514
rect 48862 26462 48914 26514
rect 50094 26462 50146 26514
rect 50542 26462 50594 26514
rect 72494 26462 72546 26514
rect 76190 26462 76242 26514
rect 76750 26462 76802 26514
rect 77310 26462 77362 26514
rect 77758 26462 77810 26514
rect 2046 26350 2098 26402
rect 35534 26350 35586 26402
rect 37998 26350 38050 26402
rect 39118 26350 39170 26402
rect 42030 26350 42082 26402
rect 43486 26350 43538 26402
rect 46174 26350 46226 26402
rect 46846 26350 46898 26402
rect 47742 26350 47794 26402
rect 49422 26350 49474 26402
rect 74622 26350 74674 26402
rect 75518 26350 75570 26402
rect 1710 26238 1762 26290
rect 33742 26238 33794 26290
rect 34302 26238 34354 26290
rect 35198 26238 35250 26290
rect 36094 26238 36146 26290
rect 37662 26238 37714 26290
rect 39678 26238 39730 26290
rect 40014 26238 40066 26290
rect 40910 26238 40962 26290
rect 41918 26238 41970 26290
rect 42926 26238 42978 26290
rect 44046 26238 44098 26290
rect 44382 26238 44434 26290
rect 45054 26238 45106 26290
rect 45950 26238 46002 26290
rect 46398 26238 46450 26290
rect 46622 26238 46674 26290
rect 46958 26238 47010 26290
rect 47294 26238 47346 26290
rect 47854 26238 47906 26290
rect 48750 26238 48802 26290
rect 49310 26238 49362 26290
rect 49646 26238 49698 26290
rect 73390 26238 73442 26290
rect 74174 26238 74226 26290
rect 74734 26238 74786 26290
rect 75294 26238 75346 26290
rect 76526 26238 76578 26290
rect 77534 26238 77586 26290
rect 77646 26238 77698 26290
rect 2494 26126 2546 26178
rect 34750 26126 34802 26178
rect 39790 26126 39842 26178
rect 41470 26126 41522 26178
rect 44942 26126 44994 26178
rect 45502 26126 45554 26178
rect 47518 26126 47570 26178
rect 71374 26126 71426 26178
rect 71822 26126 71874 26178
rect 73166 26126 73218 26178
rect 48862 26014 48914 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 65918 25846 65970 25898
rect 66022 25846 66074 25898
rect 66126 25846 66178 25898
rect 39678 25678 39730 25730
rect 40126 25678 40178 25730
rect 47070 25678 47122 25730
rect 71262 25678 71314 25730
rect 74398 25678 74450 25730
rect 74734 25678 74786 25730
rect 35982 25566 36034 25618
rect 40126 25566 40178 25618
rect 40910 25566 40962 25618
rect 41918 25566 41970 25618
rect 44270 25566 44322 25618
rect 45278 25566 45330 25618
rect 72046 25566 72098 25618
rect 72942 25566 72994 25618
rect 73726 25566 73778 25618
rect 74734 25566 74786 25618
rect 34974 25454 35026 25506
rect 35534 25454 35586 25506
rect 37214 25454 37266 25506
rect 37774 25454 37826 25506
rect 38334 25454 38386 25506
rect 38670 25454 38722 25506
rect 40462 25454 40514 25506
rect 41358 25454 41410 25506
rect 42814 25454 42866 25506
rect 43374 25454 43426 25506
rect 43710 25454 43762 25506
rect 44942 25454 44994 25506
rect 45838 25454 45890 25506
rect 46286 25454 46338 25506
rect 70926 25454 70978 25506
rect 71038 25454 71090 25506
rect 71822 25454 71874 25506
rect 72718 25454 72770 25506
rect 73502 25454 73554 25506
rect 75406 25454 75458 25506
rect 77422 25454 77474 25506
rect 78206 25454 78258 25506
rect 2046 25342 2098 25394
rect 35758 25342 35810 25394
rect 39118 25342 39170 25394
rect 42702 25342 42754 25394
rect 45502 25342 45554 25394
rect 46622 25342 46674 25394
rect 46958 25342 47010 25394
rect 47518 25342 47570 25394
rect 70478 25342 70530 25394
rect 76190 25342 76242 25394
rect 76526 25342 76578 25394
rect 77870 25342 77922 25394
rect 1710 25230 1762 25282
rect 2494 25230 2546 25282
rect 34750 25230 34802 25282
rect 38222 25230 38274 25282
rect 39678 25230 39730 25282
rect 43262 25230 43314 25282
rect 75630 25230 75682 25282
rect 77086 25230 77138 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 50558 25062 50610 25114
rect 50662 25062 50714 25114
rect 50766 25062 50818 25114
rect 25566 24894 25618 24946
rect 26574 24894 26626 24946
rect 36878 24894 36930 24946
rect 40910 24894 40962 24946
rect 42030 24894 42082 24946
rect 44046 24894 44098 24946
rect 44606 24894 44658 24946
rect 45502 24894 45554 24946
rect 46622 24894 46674 24946
rect 63086 24894 63138 24946
rect 63310 24894 63362 24946
rect 64654 24894 64706 24946
rect 71710 24894 71762 24946
rect 75854 24894 75906 24946
rect 76526 24894 76578 24946
rect 77646 24894 77698 24946
rect 17502 24782 17554 24834
rect 19742 24782 19794 24834
rect 20974 24782 21026 24834
rect 35310 24782 35362 24834
rect 35534 24782 35586 24834
rect 36206 24782 36258 24834
rect 37998 24782 38050 24834
rect 39342 24782 39394 24834
rect 40350 24782 40402 24834
rect 41246 24782 41298 24834
rect 43038 24782 43090 24834
rect 45166 24782 45218 24834
rect 46174 24782 46226 24834
rect 75742 24782 75794 24834
rect 77198 24782 77250 24834
rect 77534 24782 77586 24834
rect 17390 24670 17442 24722
rect 17726 24670 17778 24722
rect 19630 24670 19682 24722
rect 20302 24670 20354 24722
rect 25118 24670 25170 24722
rect 25790 24670 25842 24722
rect 26686 24670 26738 24722
rect 27134 24670 27186 24722
rect 30270 24670 30322 24722
rect 34974 24670 35026 24722
rect 35198 24670 35250 24722
rect 35982 24670 36034 24722
rect 37886 24670 37938 24722
rect 39678 24670 39730 24722
rect 40126 24670 40178 24722
rect 42366 24670 42418 24722
rect 43598 24670 43650 24722
rect 44158 24670 44210 24722
rect 45950 24670 46002 24722
rect 63534 24670 63586 24722
rect 72158 24670 72210 24722
rect 72942 24670 72994 24722
rect 73502 24670 73554 24722
rect 73838 24670 73890 24722
rect 74622 24670 74674 24722
rect 75182 24670 75234 24722
rect 76862 24670 76914 24722
rect 77870 24670 77922 24722
rect 18062 24558 18114 24610
rect 19294 24558 19346 24610
rect 23102 24558 23154 24610
rect 23438 24558 23490 24610
rect 23774 24558 23826 24610
rect 25678 24558 25730 24610
rect 27806 24558 27858 24610
rect 29934 24558 29986 24610
rect 30382 24558 30434 24610
rect 41694 24558 41746 24610
rect 47070 24558 47122 24610
rect 63422 24558 63474 24610
rect 71374 24558 71426 24610
rect 74062 24558 74114 24610
rect 19742 24446 19794 24498
rect 72382 24446 72434 24498
rect 75966 24446 76018 24498
rect 76862 24446 76914 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 65918 24278 65970 24330
rect 66022 24278 66074 24330
rect 66126 24278 66178 24330
rect 42590 24110 42642 24162
rect 43374 24110 43426 24162
rect 74062 24110 74114 24162
rect 77534 24110 77586 24162
rect 19630 23998 19682 24050
rect 19966 23998 20018 24050
rect 21422 23998 21474 24050
rect 23102 23998 23154 24050
rect 24782 23998 24834 24050
rect 26910 23998 26962 24050
rect 27918 23998 27970 24050
rect 34078 23998 34130 24050
rect 41806 23998 41858 24050
rect 44942 23998 44994 24050
rect 48078 23998 48130 24050
rect 62862 23998 62914 24050
rect 63534 23998 63586 24050
rect 64094 23998 64146 24050
rect 73166 23998 73218 24050
rect 74510 23998 74562 24050
rect 75294 23998 75346 24050
rect 76414 23998 76466 24050
rect 16830 23886 16882 23938
rect 21870 23886 21922 23938
rect 23998 23886 24050 23938
rect 34526 23886 34578 23938
rect 35646 23886 35698 23938
rect 35982 23886 36034 23938
rect 37662 23886 37714 23938
rect 38446 23886 38498 23938
rect 40350 23886 40402 23938
rect 45726 23886 45778 23938
rect 46062 23886 46114 23938
rect 46734 23886 46786 23938
rect 48526 23886 48578 23938
rect 62974 23886 63026 23938
rect 63422 23886 63474 23938
rect 72158 23886 72210 23938
rect 72718 23886 72770 23938
rect 73278 23886 73330 23938
rect 74398 23886 74450 23938
rect 77086 23886 77138 23938
rect 2046 23774 2098 23826
rect 17502 23774 17554 23826
rect 20302 23774 20354 23826
rect 23550 23774 23602 23826
rect 23662 23774 23714 23826
rect 27806 23774 27858 23826
rect 35758 23774 35810 23826
rect 36206 23774 36258 23826
rect 36318 23774 36370 23826
rect 37102 23774 37154 23826
rect 37214 23774 37266 23826
rect 37774 23774 37826 23826
rect 37998 23774 38050 23826
rect 38558 23774 38610 23826
rect 40462 23774 40514 23826
rect 46398 23774 46450 23826
rect 47406 23774 47458 23826
rect 47518 23774 47570 23826
rect 75630 23774 75682 23826
rect 76190 23774 76242 23826
rect 77758 23774 77810 23826
rect 1710 23662 1762 23714
rect 2494 23662 2546 23714
rect 21310 23662 21362 23714
rect 21534 23662 21586 23714
rect 22318 23662 22370 23714
rect 23326 23662 23378 23714
rect 27582 23662 27634 23714
rect 28030 23662 28082 23714
rect 34862 23662 34914 23714
rect 35422 23662 35474 23714
rect 36542 23662 36594 23714
rect 37438 23662 37490 23714
rect 40238 23662 40290 23714
rect 42366 23662 42418 23714
rect 42814 23662 42866 23714
rect 43262 23662 43314 23714
rect 44270 23662 44322 23714
rect 45390 23662 45442 23714
rect 46062 23662 46114 23714
rect 47070 23662 47122 23714
rect 47742 23662 47794 23714
rect 48974 23662 49026 23714
rect 49534 23662 49586 23714
rect 63646 23662 63698 23714
rect 75406 23662 75458 23714
rect 76414 23662 76466 23714
rect 76862 23662 76914 23714
rect 77646 23662 77698 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 50558 23494 50610 23546
rect 50662 23494 50714 23546
rect 50766 23494 50818 23546
rect 17502 23326 17554 23378
rect 17614 23326 17666 23378
rect 17838 23326 17890 23378
rect 18398 23326 18450 23378
rect 19294 23326 19346 23378
rect 21870 23326 21922 23378
rect 24670 23326 24722 23378
rect 26126 23326 26178 23378
rect 28030 23326 28082 23378
rect 38222 23326 38274 23378
rect 45166 23326 45218 23378
rect 46286 23326 46338 23378
rect 46846 23326 46898 23378
rect 47406 23326 47458 23378
rect 48974 23326 49026 23378
rect 50318 23326 50370 23378
rect 50766 23326 50818 23378
rect 71710 23326 71762 23378
rect 75742 23326 75794 23378
rect 76526 23326 76578 23378
rect 77646 23326 77698 23378
rect 2046 23214 2098 23266
rect 19966 23214 20018 23266
rect 20078 23214 20130 23266
rect 24334 23214 24386 23266
rect 24446 23214 24498 23266
rect 25230 23214 25282 23266
rect 25342 23214 25394 23266
rect 36430 23214 36482 23266
rect 37550 23214 37602 23266
rect 39678 23214 39730 23266
rect 41694 23214 41746 23266
rect 45054 23214 45106 23266
rect 46734 23214 46786 23266
rect 47966 23214 48018 23266
rect 49422 23214 49474 23266
rect 75630 23214 75682 23266
rect 76750 23214 76802 23266
rect 77086 23214 77138 23266
rect 77534 23214 77586 23266
rect 1710 23102 1762 23154
rect 17390 23102 17442 23154
rect 19518 23102 19570 23154
rect 20302 23102 20354 23154
rect 21198 23102 21250 23154
rect 21646 23102 21698 23154
rect 23550 23102 23602 23154
rect 25566 23102 25618 23154
rect 25902 23102 25954 23154
rect 27358 23102 27410 23154
rect 27806 23102 27858 23154
rect 28366 23102 28418 23154
rect 31614 23102 31666 23154
rect 31726 23102 31778 23154
rect 34078 23102 34130 23154
rect 34974 23102 35026 23154
rect 36542 23102 36594 23154
rect 37326 23102 37378 23154
rect 39230 23102 39282 23154
rect 41022 23102 41074 23154
rect 44270 23102 44322 23154
rect 45950 23102 46002 23154
rect 46174 23102 46226 23154
rect 46510 23102 46562 23154
rect 47294 23102 47346 23154
rect 47854 23102 47906 23154
rect 72158 23102 72210 23154
rect 72942 23102 72994 23154
rect 73950 23102 74002 23154
rect 74958 23102 75010 23154
rect 75966 23102 76018 23154
rect 77870 23102 77922 23154
rect 2494 22990 2546 23042
rect 20638 22990 20690 23042
rect 21198 22990 21250 23042
rect 21758 22990 21810 23042
rect 20414 22878 20466 22930
rect 23998 22990 24050 23042
rect 27918 22990 27970 23042
rect 29150 22990 29202 23042
rect 31278 22990 31330 23042
rect 33854 22990 33906 23042
rect 43822 22990 43874 23042
rect 44718 22990 44770 23042
rect 49758 22990 49810 23042
rect 72382 22990 72434 23042
rect 73278 22990 73330 23042
rect 74734 22990 74786 23042
rect 46846 22878 46898 22930
rect 47406 22878 47458 22930
rect 47966 22878 48018 22930
rect 49870 22878 49922 22930
rect 50206 22878 50258 22930
rect 74062 22878 74114 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 65918 22710 65970 22762
rect 66022 22710 66074 22762
rect 66126 22710 66178 22762
rect 35758 22542 35810 22594
rect 46734 22542 46786 22594
rect 74286 22542 74338 22594
rect 76862 22542 76914 22594
rect 77198 22542 77250 22594
rect 77534 22542 77586 22594
rect 15598 22430 15650 22482
rect 19406 22430 19458 22482
rect 19742 22430 19794 22482
rect 20078 22430 20130 22482
rect 22094 22430 22146 22482
rect 24222 22430 24274 22482
rect 24558 22430 24610 22482
rect 28366 22430 28418 22482
rect 29150 22430 29202 22482
rect 34414 22430 34466 22482
rect 37326 22430 37378 22482
rect 42142 22430 42194 22482
rect 46286 22430 46338 22482
rect 51774 22430 51826 22482
rect 52782 22430 52834 22482
rect 71934 22430 71986 22482
rect 72270 22430 72322 22482
rect 77646 22430 77698 22482
rect 16158 22318 16210 22370
rect 16606 22318 16658 22370
rect 21310 22318 21362 22370
rect 25566 22318 25618 22370
rect 38334 22318 38386 22370
rect 40350 22318 40402 22370
rect 42478 22318 42530 22370
rect 43374 22318 43426 22370
rect 45166 22318 45218 22370
rect 45950 22318 46002 22370
rect 46174 22318 46226 22370
rect 47182 22318 47234 22370
rect 48078 22318 48130 22370
rect 48638 22318 48690 22370
rect 48974 22318 49026 22370
rect 50094 22318 50146 22370
rect 50878 22318 50930 22370
rect 51326 22318 51378 22370
rect 72046 22318 72098 22370
rect 72830 22318 72882 22370
rect 73390 22318 73442 22370
rect 74062 22318 74114 22370
rect 74846 22318 74898 22370
rect 75406 22318 75458 22370
rect 76190 22318 76242 22370
rect 16046 22206 16098 22258
rect 17278 22206 17330 22258
rect 20414 22206 20466 22258
rect 26238 22206 26290 22258
rect 35198 22206 35250 22258
rect 35310 22206 35362 22258
rect 35870 22206 35922 22258
rect 36206 22206 36258 22258
rect 36318 22206 36370 22258
rect 38446 22206 38498 22258
rect 40462 22206 40514 22258
rect 42366 22206 42418 22258
rect 43710 22206 43762 22258
rect 43822 22206 43874 22258
rect 46398 22206 46450 22258
rect 46846 22206 46898 22258
rect 49870 22206 49922 22258
rect 76526 22206 76578 22258
rect 15822 22094 15874 22146
rect 20750 22094 20802 22146
rect 24670 22094 24722 22146
rect 29262 22094 29314 22146
rect 33966 22094 34018 22146
rect 34750 22094 34802 22146
rect 34974 22094 35026 22146
rect 35758 22094 35810 22146
rect 36542 22094 36594 22146
rect 37774 22094 37826 22146
rect 40014 22094 40066 22146
rect 43038 22094 43090 22146
rect 44046 22094 44098 22146
rect 45502 22094 45554 22146
rect 47742 22094 47794 22146
rect 49086 22094 49138 22146
rect 76974 22094 77026 22146
rect 77758 22094 77810 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 50558 21926 50610 21978
rect 50662 21926 50714 21978
rect 50766 21926 50818 21978
rect 17502 21758 17554 21810
rect 17726 21758 17778 21810
rect 17838 21758 17890 21810
rect 17950 21758 18002 21810
rect 18510 21758 18562 21810
rect 23886 21758 23938 21810
rect 26462 21758 26514 21810
rect 26574 21758 26626 21810
rect 39230 21758 39282 21810
rect 45726 21758 45778 21810
rect 48078 21758 48130 21810
rect 53790 21758 53842 21810
rect 55358 21758 55410 21810
rect 55918 21758 55970 21810
rect 2046 21646 2098 21698
rect 25230 21646 25282 21698
rect 25342 21646 25394 21698
rect 35198 21646 35250 21698
rect 35982 21646 36034 21698
rect 36878 21646 36930 21698
rect 39902 21646 39954 21698
rect 43262 21646 43314 21698
rect 44270 21646 44322 21698
rect 46398 21646 46450 21698
rect 47182 21646 47234 21698
rect 47406 21646 47458 21698
rect 47630 21646 47682 21698
rect 48190 21646 48242 21698
rect 49870 21646 49922 21698
rect 51326 21646 51378 21698
rect 54350 21646 54402 21698
rect 71710 21646 71762 21698
rect 73950 21646 74002 21698
rect 76078 21646 76130 21698
rect 76638 21646 76690 21698
rect 76974 21646 77026 21698
rect 77534 21646 77586 21698
rect 77758 21646 77810 21698
rect 1710 21534 1762 21586
rect 18846 21534 18898 21586
rect 24222 21534 24274 21586
rect 25566 21534 25618 21586
rect 25902 21534 25954 21586
rect 26350 21534 26402 21586
rect 29150 21534 29202 21586
rect 32398 21534 32450 21586
rect 34974 21534 35026 21586
rect 35422 21534 35474 21586
rect 35646 21534 35698 21586
rect 36318 21534 36370 21586
rect 37662 21534 37714 21586
rect 38558 21534 38610 21586
rect 39118 21534 39170 21586
rect 41358 21534 41410 21586
rect 42478 21534 42530 21586
rect 44158 21534 44210 21586
rect 45614 21534 45666 21586
rect 47854 21534 47906 21586
rect 48974 21534 49026 21586
rect 49534 21534 49586 21586
rect 50206 21534 50258 21586
rect 51886 21534 51938 21586
rect 52446 21534 52498 21586
rect 52782 21534 52834 21586
rect 53342 21534 53394 21586
rect 54910 21534 54962 21586
rect 55470 21534 55522 21586
rect 72158 21534 72210 21586
rect 72942 21534 72994 21586
rect 73502 21534 73554 21586
rect 74286 21534 74338 21586
rect 74958 21534 75010 21586
rect 75742 21534 75794 21586
rect 2494 21422 2546 21474
rect 19630 21422 19682 21474
rect 21758 21422 21810 21474
rect 24670 21422 24722 21474
rect 29934 21422 29986 21474
rect 32062 21422 32114 21474
rect 34862 21422 34914 21474
rect 41022 21422 41074 21474
rect 49198 21422 49250 21474
rect 50654 21422 50706 21474
rect 51998 21422 52050 21474
rect 74622 21422 74674 21474
rect 77870 21422 77922 21474
rect 32510 21310 32562 21362
rect 42142 21310 42194 21362
rect 72382 21310 72434 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 65918 21142 65970 21194
rect 66022 21142 66074 21194
rect 66126 21142 66178 21194
rect 32510 20974 32562 21026
rect 32958 20974 33010 21026
rect 38782 20974 38834 21026
rect 75294 20974 75346 21026
rect 76526 20974 76578 21026
rect 76862 20974 76914 21026
rect 77198 20974 77250 21026
rect 19518 20862 19570 20914
rect 29822 20862 29874 20914
rect 33182 20862 33234 20914
rect 35310 20862 35362 20914
rect 37214 20862 37266 20914
rect 51886 20862 51938 20914
rect 54126 20862 54178 20914
rect 55022 20862 55074 20914
rect 56926 20862 56978 20914
rect 71262 20862 71314 20914
rect 74286 20862 74338 20914
rect 75070 20862 75122 20914
rect 77310 20862 77362 20914
rect 20078 20750 20130 20802
rect 26574 20750 26626 20802
rect 35086 20750 35138 20802
rect 35534 20750 35586 20802
rect 35646 20750 35698 20802
rect 36430 20750 36482 20802
rect 38110 20750 38162 20802
rect 39454 20750 39506 20802
rect 40126 20750 40178 20802
rect 41246 20750 41298 20802
rect 43150 20750 43202 20802
rect 45054 20750 45106 20802
rect 45502 20750 45554 20802
rect 45950 20750 46002 20802
rect 47070 20750 47122 20802
rect 47630 20750 47682 20802
rect 48414 20750 48466 20802
rect 48974 20750 49026 20802
rect 49534 20750 49586 20802
rect 50318 20750 50370 20802
rect 51438 20750 51490 20802
rect 53566 20750 53618 20802
rect 54014 20750 54066 20802
rect 55134 20750 55186 20802
rect 55806 20750 55858 20802
rect 56478 20750 56530 20802
rect 71374 20750 71426 20802
rect 72494 20750 72546 20802
rect 72718 20750 72770 20802
rect 73054 20750 73106 20802
rect 73950 20750 74002 20802
rect 75294 20750 75346 20802
rect 77534 20750 77586 20802
rect 78206 20750 78258 20802
rect 2046 20638 2098 20690
rect 24446 20638 24498 20690
rect 24782 20638 24834 20690
rect 25230 20638 25282 20690
rect 25790 20638 25842 20690
rect 33518 20638 33570 20690
rect 34302 20638 34354 20690
rect 34638 20638 34690 20690
rect 34862 20638 34914 20690
rect 36094 20638 36146 20690
rect 41134 20638 41186 20690
rect 42926 20638 42978 20690
rect 46398 20638 46450 20690
rect 48526 20638 48578 20690
rect 49982 20638 50034 20690
rect 50990 20638 51042 20690
rect 54350 20638 54402 20690
rect 55022 20638 55074 20690
rect 72270 20638 72322 20690
rect 74062 20638 74114 20690
rect 75630 20638 75682 20690
rect 77870 20638 77922 20690
rect 1710 20526 1762 20578
rect 2494 20526 2546 20578
rect 19406 20526 19458 20578
rect 19630 20526 19682 20578
rect 20526 20526 20578 20578
rect 22990 20526 23042 20578
rect 23662 20526 23714 20578
rect 24110 20526 24162 20578
rect 25342 20526 25394 20578
rect 25566 20526 25618 20578
rect 25902 20526 25954 20578
rect 26126 20526 26178 20578
rect 26910 20526 26962 20578
rect 29486 20526 29538 20578
rect 29710 20526 29762 20578
rect 29934 20526 29986 20578
rect 30494 20526 30546 20578
rect 32398 20526 32450 20578
rect 32958 20526 33010 20578
rect 34078 20526 34130 20578
rect 34526 20526 34578 20578
rect 37438 20526 37490 20578
rect 37774 20526 37826 20578
rect 38446 20526 38498 20578
rect 39902 20526 39954 20578
rect 40686 20526 40738 20578
rect 42142 20526 42194 20578
rect 46846 20526 46898 20578
rect 47630 20526 47682 20578
rect 48974 20526 49026 20578
rect 50430 20526 50482 20578
rect 52782 20526 52834 20578
rect 76638 20526 76690 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 50558 20358 50610 20410
rect 50662 20358 50714 20410
rect 50766 20358 50818 20410
rect 19070 20190 19122 20242
rect 19854 20190 19906 20242
rect 33406 20190 33458 20242
rect 33854 20190 33906 20242
rect 34302 20190 34354 20242
rect 37550 20190 37602 20242
rect 39902 20190 39954 20242
rect 42814 20190 42866 20242
rect 48078 20190 48130 20242
rect 51550 20190 51602 20242
rect 52334 20190 52386 20242
rect 72942 20190 72994 20242
rect 73950 20190 74002 20242
rect 18622 20078 18674 20130
rect 19630 20078 19682 20130
rect 21310 20078 21362 20130
rect 25566 20078 25618 20130
rect 35086 20078 35138 20130
rect 35534 20078 35586 20130
rect 35870 20078 35922 20130
rect 40910 20078 40962 20130
rect 42926 20078 42978 20130
rect 44494 20078 44546 20130
rect 47406 20078 47458 20130
rect 48190 20078 48242 20130
rect 49422 20078 49474 20130
rect 51102 20078 51154 20130
rect 53230 20078 53282 20130
rect 54350 20078 54402 20130
rect 57598 20078 57650 20130
rect 75070 20078 75122 20130
rect 75630 20078 75682 20130
rect 76078 20078 76130 20130
rect 76750 20078 76802 20130
rect 77646 20078 77698 20130
rect 78318 20078 78370 20130
rect 18958 19966 19010 20018
rect 19518 19966 19570 20018
rect 20190 19966 20242 20018
rect 21646 19966 21698 20018
rect 25230 19966 25282 20018
rect 26462 19966 26514 20018
rect 29598 19966 29650 20018
rect 33742 19966 33794 20018
rect 34862 19966 34914 20018
rect 35198 19966 35250 20018
rect 36318 19966 36370 20018
rect 37662 19966 37714 20018
rect 37998 19966 38050 20018
rect 39454 19966 39506 20018
rect 39678 19966 39730 20018
rect 40014 19966 40066 20018
rect 41134 19966 41186 20018
rect 43038 19966 43090 20018
rect 44718 19966 44770 20018
rect 46286 19966 46338 20018
rect 46734 19966 46786 20018
rect 48750 19966 48802 20018
rect 49310 19966 49362 20018
rect 50878 19966 50930 20018
rect 51774 19966 51826 20018
rect 52110 19966 52162 20018
rect 52894 19966 52946 20018
rect 53566 19966 53618 20018
rect 54238 19966 54290 20018
rect 55022 19966 55074 20018
rect 56702 19966 56754 20018
rect 74846 19966 74898 20018
rect 76302 19966 76354 20018
rect 77086 19966 77138 20018
rect 77422 19966 77474 20018
rect 20974 19854 21026 19906
rect 22430 19854 22482 19906
rect 24558 19854 24610 19906
rect 26014 19854 26066 19906
rect 27134 19854 27186 19906
rect 29262 19854 29314 19906
rect 30382 19854 30434 19906
rect 32510 19854 32562 19906
rect 33294 19854 33346 19906
rect 34190 19854 34242 19906
rect 49534 19854 49586 19906
rect 50318 19854 50370 19906
rect 54014 19854 54066 19906
rect 55470 19854 55522 19906
rect 56030 19854 56082 19906
rect 57150 19854 57202 19906
rect 75406 19854 75458 19906
rect 75742 19854 75794 19906
rect 76974 19854 77026 19906
rect 77646 19854 77698 19906
rect 19070 19742 19122 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 65918 19574 65970 19626
rect 66022 19574 66074 19626
rect 66126 19574 66178 19626
rect 32174 19406 32226 19458
rect 32846 19406 32898 19458
rect 33966 19406 34018 19458
rect 22654 19294 22706 19346
rect 27470 19294 27522 19346
rect 28590 19294 28642 19346
rect 29038 19294 29090 19346
rect 29262 19294 29314 19346
rect 30382 19294 30434 19346
rect 31278 19294 31330 19346
rect 33070 19294 33122 19346
rect 35422 19294 35474 19346
rect 38110 19294 38162 19346
rect 48526 19294 48578 19346
rect 53678 19294 53730 19346
rect 75070 19294 75122 19346
rect 19294 19182 19346 19234
rect 21758 19182 21810 19234
rect 22094 19182 22146 19234
rect 22542 19182 22594 19234
rect 26910 19182 26962 19234
rect 27582 19182 27634 19234
rect 29934 19182 29986 19234
rect 30270 19182 30322 19234
rect 30494 19182 30546 19234
rect 34638 19182 34690 19234
rect 35646 19182 35698 19234
rect 36430 19182 36482 19234
rect 37326 19182 37378 19234
rect 37998 19182 38050 19234
rect 38334 19182 38386 19234
rect 38446 19182 38498 19234
rect 39118 19182 39170 19234
rect 39342 19182 39394 19234
rect 40238 19182 40290 19234
rect 40798 19182 40850 19234
rect 41022 19182 41074 19234
rect 41694 19182 41746 19234
rect 43374 19182 43426 19234
rect 44830 19182 44882 19234
rect 45390 19182 45442 19234
rect 46622 19182 46674 19234
rect 47182 19182 47234 19234
rect 49758 19182 49810 19234
rect 50990 19182 51042 19234
rect 52670 19182 52722 19234
rect 53342 19182 53394 19234
rect 54574 19182 54626 19234
rect 56142 19182 56194 19234
rect 57038 19182 57090 19234
rect 76862 19182 76914 19234
rect 78206 19182 78258 19234
rect 1710 19070 1762 19122
rect 2046 19070 2098 19122
rect 2494 19070 2546 19122
rect 19070 19070 19122 19122
rect 21534 19070 21586 19122
rect 22766 19070 22818 19122
rect 23102 19070 23154 19122
rect 23326 19070 23378 19122
rect 24446 19070 24498 19122
rect 24782 19070 24834 19122
rect 25118 19070 25170 19122
rect 25566 19070 25618 19122
rect 25902 19070 25954 19122
rect 26238 19070 26290 19122
rect 29710 19070 29762 19122
rect 33406 19070 33458 19122
rect 33854 19070 33906 19122
rect 34974 19070 35026 19122
rect 35310 19070 35362 19122
rect 35870 19070 35922 19122
rect 36318 19070 36370 19122
rect 37102 19070 37154 19122
rect 38894 19070 38946 19122
rect 39902 19070 39954 19122
rect 40462 19070 40514 19122
rect 40574 19070 40626 19122
rect 42926 19070 42978 19122
rect 49310 19070 49362 19122
rect 51102 19070 51154 19122
rect 53454 19070 53506 19122
rect 54798 19070 54850 19122
rect 76526 19070 76578 19122
rect 77198 19070 77250 19122
rect 77534 19070 77586 19122
rect 23214 18958 23266 19010
rect 23550 18958 23602 19010
rect 24110 18958 24162 19010
rect 24334 18958 24386 19010
rect 26350 18958 26402 19010
rect 26574 18958 26626 19010
rect 27358 18958 27410 19010
rect 28478 18958 28530 19010
rect 29486 18958 29538 19010
rect 29822 18958 29874 19010
rect 30718 18958 30770 19010
rect 31950 18958 32002 19010
rect 32286 18958 32338 19010
rect 32734 18958 32786 19010
rect 39118 18958 39170 19010
rect 40014 18958 40066 19010
rect 43038 18958 43090 19010
rect 46622 18958 46674 19010
rect 49982 18958 50034 19010
rect 56366 18958 56418 19010
rect 75406 18958 75458 19010
rect 76638 18958 76690 19010
rect 77870 18958 77922 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 50558 18790 50610 18842
rect 50662 18790 50714 18842
rect 50766 18790 50818 18842
rect 17838 18622 17890 18674
rect 41358 18622 41410 18674
rect 41918 18622 41970 18674
rect 42366 18622 42418 18674
rect 49870 18622 49922 18674
rect 54798 18622 54850 18674
rect 71262 18622 71314 18674
rect 76750 18622 76802 18674
rect 2046 18510 2098 18562
rect 17950 18510 18002 18562
rect 24334 18510 24386 18562
rect 30046 18510 30098 18562
rect 41806 18510 41858 18562
rect 44046 18510 44098 18562
rect 48862 18510 48914 18562
rect 51102 18510 51154 18562
rect 53230 18510 53282 18562
rect 55134 18510 55186 18562
rect 77422 18510 77474 18562
rect 1710 18398 1762 18450
rect 23438 18398 23490 18450
rect 24670 18398 24722 18450
rect 25342 18398 25394 18450
rect 25790 18398 25842 18450
rect 29374 18398 29426 18450
rect 33630 18398 33682 18450
rect 39230 18398 39282 18450
rect 39342 18398 39394 18450
rect 39790 18398 39842 18450
rect 40014 18398 40066 18450
rect 41246 18398 41298 18450
rect 42702 18398 42754 18450
rect 44270 18398 44322 18450
rect 45614 18398 45666 18450
rect 47854 18398 47906 18450
rect 49982 18398 50034 18450
rect 50878 18398 50930 18450
rect 53006 18398 53058 18450
rect 54910 18398 54962 18450
rect 56702 18398 56754 18450
rect 70926 18398 70978 18450
rect 77198 18398 77250 18450
rect 77758 18398 77810 18450
rect 78318 18398 78370 18450
rect 2494 18286 2546 18338
rect 18846 18286 18898 18338
rect 23998 18286 24050 18338
rect 26462 18286 26514 18338
rect 28590 18286 28642 18338
rect 32174 18286 32226 18338
rect 38222 18286 38274 18338
rect 39566 18286 39618 18338
rect 43038 18286 43090 18338
rect 43150 18286 43202 18338
rect 45502 18286 45554 18338
rect 52558 18286 52610 18338
rect 57150 18286 57202 18338
rect 70590 18286 70642 18338
rect 17838 18174 17890 18226
rect 41358 18174 41410 18226
rect 41918 18174 41970 18226
rect 44046 18174 44098 18226
rect 47182 18174 47234 18226
rect 77758 18174 77810 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 65918 18006 65970 18058
rect 66022 18006 66074 18058
rect 66126 18006 66178 18058
rect 17726 17726 17778 17778
rect 18174 17726 18226 17778
rect 22318 17726 22370 17778
rect 27918 17726 27970 17778
rect 28590 17726 28642 17778
rect 36318 17726 36370 17778
rect 37102 17726 37154 17778
rect 39118 17726 39170 17778
rect 47742 17726 47794 17778
rect 48526 17726 48578 17778
rect 18846 17614 18898 17666
rect 19182 17614 19234 17666
rect 19854 17614 19906 17666
rect 19966 17614 20018 17666
rect 27246 17614 27298 17666
rect 33630 17614 33682 17666
rect 35646 17614 35698 17666
rect 35870 17614 35922 17666
rect 37214 17614 37266 17666
rect 37998 17614 38050 17666
rect 38446 17614 38498 17666
rect 38670 17614 38722 17666
rect 39342 17614 39394 17666
rect 39790 17614 39842 17666
rect 40014 17614 40066 17666
rect 40686 17614 40738 17666
rect 41358 17614 41410 17666
rect 42926 17614 42978 17666
rect 43150 17614 43202 17666
rect 44830 17614 44882 17666
rect 45390 17614 45442 17666
rect 46958 17614 47010 17666
rect 49646 17614 49698 17666
rect 51326 17614 51378 17666
rect 53230 17614 53282 17666
rect 55470 17614 55522 17666
rect 56590 17614 56642 17666
rect 56814 17614 56866 17666
rect 58718 17614 58770 17666
rect 78206 17614 78258 17666
rect 1710 17502 1762 17554
rect 2046 17502 2098 17554
rect 19518 17502 19570 17554
rect 21310 17502 21362 17554
rect 21646 17502 21698 17554
rect 29598 17502 29650 17554
rect 35310 17502 35362 17554
rect 36990 17502 37042 17554
rect 37550 17502 37602 17554
rect 40350 17502 40402 17554
rect 41470 17502 41522 17554
rect 47070 17502 47122 17554
rect 49198 17502 49250 17554
rect 51102 17502 51154 17554
rect 51774 17502 51826 17554
rect 53454 17502 53506 17554
rect 55134 17502 55186 17554
rect 58830 17502 58882 17554
rect 76974 17502 77026 17554
rect 77198 17502 77250 17554
rect 77534 17502 77586 17554
rect 77870 17502 77922 17554
rect 2494 17390 2546 17442
rect 18958 17390 19010 17442
rect 19742 17390 19794 17442
rect 20414 17390 20466 17442
rect 28478 17390 28530 17442
rect 35534 17390 35586 17442
rect 38222 17390 38274 17442
rect 39678 17390 39730 17442
rect 43038 17390 43090 17442
rect 54126 17390 54178 17442
rect 57710 17390 57762 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 50558 17222 50610 17274
rect 50662 17222 50714 17274
rect 50766 17222 50818 17274
rect 26350 17054 26402 17106
rect 26686 17054 26738 17106
rect 26798 17054 26850 17106
rect 27582 17054 27634 17106
rect 28142 17054 28194 17106
rect 32510 17054 32562 17106
rect 33854 17054 33906 17106
rect 34302 17054 34354 17106
rect 35198 17054 35250 17106
rect 35982 17054 36034 17106
rect 37102 17054 37154 17106
rect 37550 17054 37602 17106
rect 37998 17054 38050 17106
rect 39006 17054 39058 17106
rect 39790 17054 39842 17106
rect 41134 17054 41186 17106
rect 41694 17054 41746 17106
rect 42142 17054 42194 17106
rect 42590 17054 42642 17106
rect 44270 17054 44322 17106
rect 48078 17054 48130 17106
rect 49982 17054 50034 17106
rect 57150 17054 57202 17106
rect 77646 17054 77698 17106
rect 77870 17054 77922 17106
rect 19294 16942 19346 16994
rect 22542 16942 22594 16994
rect 27022 16942 27074 16994
rect 32062 16942 32114 16994
rect 36094 16942 36146 16994
rect 39902 16942 39954 16994
rect 41358 16942 41410 16994
rect 41470 16942 41522 16994
rect 42926 16942 42978 16994
rect 45614 16942 45666 16994
rect 47406 16942 47458 16994
rect 49310 16942 49362 16994
rect 51102 16942 51154 16994
rect 52446 16942 52498 16994
rect 18622 16830 18674 16882
rect 21870 16830 21922 16882
rect 26574 16830 26626 16882
rect 28590 16830 28642 16882
rect 33518 16830 33570 16882
rect 34638 16830 34690 16882
rect 34750 16830 34802 16882
rect 35646 16830 35698 16882
rect 36206 16830 36258 16882
rect 37438 16830 37490 16882
rect 38670 16830 38722 16882
rect 38894 16830 38946 16882
rect 39230 16830 39282 16882
rect 39454 16830 39506 16882
rect 40126 16830 40178 16882
rect 44606 16830 44658 16882
rect 46734 16830 46786 16882
rect 47070 16830 47122 16882
rect 48190 16830 48242 16882
rect 49086 16830 49138 16882
rect 50990 16830 51042 16882
rect 52670 16830 52722 16882
rect 54350 16830 54402 16882
rect 54574 16830 54626 16882
rect 56702 16830 56754 16882
rect 77198 16830 77250 16882
rect 78094 16830 78146 16882
rect 21422 16718 21474 16770
rect 24670 16718 24722 16770
rect 29262 16718 29314 16770
rect 31390 16718 31442 16770
rect 31726 16718 31778 16770
rect 33742 16718 33794 16770
rect 34190 16718 34242 16770
rect 37886 16718 37938 16770
rect 55358 16718 55410 16770
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 65918 16438 65970 16490
rect 66022 16438 66074 16490
rect 66126 16438 66178 16490
rect 37102 16270 37154 16322
rect 37998 16270 38050 16322
rect 38446 16270 38498 16322
rect 44046 16270 44098 16322
rect 51102 16270 51154 16322
rect 23774 16158 23826 16210
rect 27918 16158 27970 16210
rect 28254 16158 28306 16210
rect 29262 16158 29314 16210
rect 30158 16158 30210 16210
rect 34974 16158 35026 16210
rect 36094 16158 36146 16210
rect 36542 16158 36594 16210
rect 36990 16158 37042 16210
rect 39678 16158 39730 16210
rect 40462 16158 40514 16210
rect 40910 16158 40962 16210
rect 41470 16158 41522 16210
rect 41918 16158 41970 16210
rect 44942 16158 44994 16210
rect 51998 16158 52050 16210
rect 56478 16158 56530 16210
rect 25006 16046 25058 16098
rect 29374 16046 29426 16098
rect 32174 16046 32226 16098
rect 35310 16046 35362 16098
rect 38894 16046 38946 16098
rect 43038 16046 43090 16098
rect 43374 16046 43426 16098
rect 43710 16046 43762 16098
rect 43934 16046 43986 16098
rect 45502 16046 45554 16098
rect 46062 16046 46114 16098
rect 47294 16046 47346 16098
rect 48974 16046 49026 16098
rect 50430 16046 50482 16098
rect 52670 16046 52722 16098
rect 52894 16046 52946 16098
rect 54462 16046 54514 16098
rect 54798 16046 54850 16098
rect 1710 15934 1762 15986
rect 2046 15934 2098 15986
rect 25790 15934 25842 15986
rect 32846 15934 32898 15986
rect 37550 15934 37602 15986
rect 37886 15934 37938 15986
rect 38334 15934 38386 15986
rect 39230 15934 39282 15986
rect 42142 15934 42194 15986
rect 43486 15934 43538 15986
rect 47742 15934 47794 15986
rect 49534 15934 49586 15986
rect 77870 15934 77922 15986
rect 78206 15934 78258 15986
rect 2494 15822 2546 15874
rect 28366 15822 28418 15874
rect 29150 15822 29202 15874
rect 29598 15822 29650 15874
rect 35422 15822 35474 15874
rect 37438 15822 37490 15874
rect 42254 15822 42306 15874
rect 44046 15822 44098 15874
rect 45726 15822 45778 15874
rect 46398 15822 46450 15874
rect 47966 15822 48018 15874
rect 51438 15822 51490 15874
rect 53790 15822 53842 15874
rect 77646 15822 77698 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 50558 15654 50610 15706
rect 50662 15654 50714 15706
rect 50766 15654 50818 15706
rect 33518 15486 33570 15538
rect 34078 15486 34130 15538
rect 34526 15486 34578 15538
rect 38558 15486 38610 15538
rect 39006 15486 39058 15538
rect 39454 15486 39506 15538
rect 40126 15486 40178 15538
rect 46510 15486 46562 15538
rect 2046 15374 2098 15426
rect 27246 15374 27298 15426
rect 33406 15374 33458 15426
rect 38894 15374 38946 15426
rect 47742 15374 47794 15426
rect 48862 15374 48914 15426
rect 50654 15374 50706 15426
rect 52334 15374 52386 15426
rect 1710 15262 1762 15314
rect 30830 15262 30882 15314
rect 32958 15262 33010 15314
rect 33630 15262 33682 15314
rect 35198 15262 35250 15314
rect 39678 15262 39730 15314
rect 40350 15262 40402 15314
rect 41694 15262 41746 15314
rect 45502 15262 45554 15314
rect 46398 15262 46450 15314
rect 47182 15262 47234 15314
rect 48974 15262 49026 15314
rect 50878 15262 50930 15314
rect 52558 15262 52610 15314
rect 54238 15262 54290 15314
rect 54462 15262 54514 15314
rect 2494 15150 2546 15202
rect 31390 15150 31442 15202
rect 32510 15150 32562 15202
rect 35982 15150 36034 15202
rect 38110 15150 38162 15202
rect 40238 15150 40290 15202
rect 42478 15150 42530 15202
rect 44606 15150 44658 15202
rect 51662 15150 51714 15202
rect 55246 15150 55298 15202
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 65918 14870 65970 14922
rect 66022 14870 66074 14922
rect 66126 14870 66178 14922
rect 43934 14702 43986 14754
rect 44270 14702 44322 14754
rect 45166 14702 45218 14754
rect 53454 14702 53506 14754
rect 26686 14590 26738 14642
rect 34190 14590 34242 14642
rect 34526 14590 34578 14642
rect 34862 14590 34914 14642
rect 35982 14590 36034 14642
rect 40014 14590 40066 14642
rect 42142 14590 42194 14642
rect 42590 14590 42642 14642
rect 43934 14590 43986 14642
rect 44382 14590 44434 14642
rect 45726 14590 45778 14642
rect 50094 14590 50146 14642
rect 50654 14590 50706 14642
rect 26126 14478 26178 14530
rect 31390 14478 31442 14530
rect 35422 14478 35474 14530
rect 35870 14478 35922 14530
rect 39230 14478 39282 14530
rect 42702 14478 42754 14530
rect 45054 14478 45106 14530
rect 47518 14478 47570 14530
rect 48190 14478 48242 14530
rect 48750 14478 48802 14530
rect 51326 14478 51378 14530
rect 52670 14478 52722 14530
rect 26798 14366 26850 14418
rect 28254 14366 28306 14418
rect 29150 14366 29202 14418
rect 30942 14366 30994 14418
rect 32062 14366 32114 14418
rect 42926 14366 42978 14418
rect 46846 14366 46898 14418
rect 77870 14366 77922 14418
rect 78206 14366 78258 14418
rect 26574 14254 26626 14306
rect 27246 14254 27298 14306
rect 28590 14254 28642 14306
rect 29262 14254 29314 14306
rect 29374 14254 29426 14306
rect 29598 14254 29650 14306
rect 30158 14254 30210 14306
rect 30830 14254 30882 14306
rect 36094 14254 36146 14306
rect 42478 14254 42530 14306
rect 48414 14254 48466 14306
rect 51998 14254 52050 14306
rect 77646 14254 77698 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 50558 14086 50610 14138
rect 50662 14086 50714 14138
rect 50766 14086 50818 14138
rect 2046 13918 2098 13970
rect 25902 13918 25954 13970
rect 27022 13918 27074 13970
rect 28142 13918 28194 13970
rect 33406 13918 33458 13970
rect 33518 13918 33570 13970
rect 33630 13918 33682 13970
rect 34190 13918 34242 13970
rect 34414 13918 34466 13970
rect 39342 13918 39394 13970
rect 40238 13918 40290 13970
rect 41582 13918 41634 13970
rect 48302 13918 48354 13970
rect 48974 13918 49026 13970
rect 49422 13918 49474 13970
rect 52222 13918 52274 13970
rect 77870 13918 77922 13970
rect 26126 13806 26178 13858
rect 26686 13806 26738 13858
rect 27246 13806 27298 13858
rect 27918 13806 27970 13858
rect 29150 13806 29202 13858
rect 34750 13806 34802 13858
rect 40014 13806 40066 13858
rect 51998 13806 52050 13858
rect 53902 13806 53954 13858
rect 1710 13694 1762 13746
rect 19630 13694 19682 13746
rect 23438 13694 23490 13746
rect 26238 13694 26290 13746
rect 26574 13694 26626 13746
rect 27358 13694 27410 13746
rect 27806 13694 27858 13746
rect 28478 13694 28530 13746
rect 33070 13694 33122 13746
rect 35086 13694 35138 13746
rect 38334 13694 38386 13746
rect 39006 13694 39058 13746
rect 39566 13694 39618 13746
rect 42030 13694 42082 13746
rect 45278 13694 45330 13746
rect 45390 13694 45442 13746
rect 51326 13694 51378 13746
rect 53566 13694 53618 13746
rect 78094 13694 78146 13746
rect 2494 13582 2546 13634
rect 20414 13582 20466 13634
rect 22542 13582 22594 13634
rect 23662 13582 23714 13634
rect 31278 13582 31330 13634
rect 35870 13582 35922 13634
rect 37998 13582 38050 13634
rect 40126 13582 40178 13634
rect 41694 13582 41746 13634
rect 42814 13582 42866 13634
rect 44942 13582 44994 13634
rect 46958 13582 47010 13634
rect 77646 13582 77698 13634
rect 23774 13470 23826 13522
rect 26686 13470 26738 13522
rect 38446 13470 38498 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 65918 13302 65970 13354
rect 66022 13302 66074 13354
rect 66126 13302 66178 13354
rect 32510 13134 32562 13186
rect 33070 13134 33122 13186
rect 33966 13134 34018 13186
rect 19518 13022 19570 13074
rect 21422 13022 21474 13074
rect 23662 13022 23714 13074
rect 25790 13022 25842 13074
rect 26574 13022 26626 13074
rect 35870 13022 35922 13074
rect 39902 13022 39954 13074
rect 42030 13022 42082 13074
rect 42926 13022 42978 13074
rect 16606 12910 16658 12962
rect 19966 12910 20018 12962
rect 20078 12910 20130 12962
rect 22990 12910 23042 12962
rect 26462 12910 26514 12962
rect 32622 12910 32674 12962
rect 33182 12910 33234 12962
rect 33854 12910 33906 12962
rect 34414 12910 34466 12962
rect 34750 12910 34802 12962
rect 35422 12910 35474 12962
rect 35758 12910 35810 12962
rect 35982 12910 36034 12962
rect 37662 12910 37714 12962
rect 38446 12910 38498 12962
rect 39230 12910 39282 12962
rect 42366 12910 42418 12962
rect 43038 12910 43090 12962
rect 1710 12798 1762 12850
rect 2046 12798 2098 12850
rect 17278 12798 17330 12850
rect 27806 12798 27858 12850
rect 28142 12798 28194 12850
rect 29150 12798 29202 12850
rect 29486 12798 29538 12850
rect 37326 12798 37378 12850
rect 42814 12798 42866 12850
rect 2494 12686 2546 12738
rect 20190 12686 20242 12738
rect 20414 12686 20466 12738
rect 26238 12686 26290 12738
rect 26686 12686 26738 12738
rect 32510 12686 32562 12738
rect 33070 12686 33122 12738
rect 33966 12686 34018 12738
rect 34526 12686 34578 12738
rect 37438 12686 37490 12738
rect 38782 12686 38834 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 50558 12518 50610 12570
rect 50662 12518 50714 12570
rect 50766 12518 50818 12570
rect 12574 12350 12626 12402
rect 19182 12350 19234 12402
rect 19406 12350 19458 12402
rect 20974 12350 21026 12402
rect 25454 12350 25506 12402
rect 28254 12350 28306 12402
rect 33742 12350 33794 12402
rect 36206 12350 36258 12402
rect 37214 12350 37266 12402
rect 41694 12350 41746 12402
rect 42366 12350 42418 12402
rect 74622 12350 74674 12402
rect 75966 12350 76018 12402
rect 77870 12350 77922 12402
rect 17726 12238 17778 12290
rect 20078 12238 20130 12290
rect 20302 12238 20354 12290
rect 36430 12238 36482 12290
rect 36990 12238 37042 12290
rect 9662 12126 9714 12178
rect 19854 12126 19906 12178
rect 21758 12126 21810 12178
rect 25230 12126 25282 12178
rect 25902 12126 25954 12178
rect 27918 12126 27970 12178
rect 29262 12126 29314 12178
rect 33966 12126 34018 12178
rect 36542 12126 36594 12178
rect 36878 12126 36930 12178
rect 37550 12126 37602 12178
rect 41582 12126 41634 12178
rect 74958 12126 75010 12178
rect 75182 12126 75234 12178
rect 78206 12126 78258 12178
rect 10334 12014 10386 12066
rect 17614 12014 17666 12066
rect 17950 12014 18002 12066
rect 19294 12014 19346 12066
rect 20414 12014 20466 12066
rect 22430 12014 22482 12066
rect 24558 12014 24610 12066
rect 25342 12014 25394 12066
rect 29934 12014 29986 12066
rect 32062 12014 32114 12066
rect 38222 12014 38274 12066
rect 40350 12014 40402 12066
rect 41022 12014 41074 12066
rect 77646 12014 77698 12066
rect 40910 11902 40962 11954
rect 75518 11902 75570 11954
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 65918 11734 65970 11786
rect 66022 11734 66074 11786
rect 66126 11734 66178 11786
rect 22430 11566 22482 11618
rect 37998 11566 38050 11618
rect 9438 11454 9490 11506
rect 12462 11454 12514 11506
rect 13470 11454 13522 11506
rect 18398 11454 18450 11506
rect 20638 11454 20690 11506
rect 22318 11454 22370 11506
rect 28254 11454 28306 11506
rect 29934 11454 29986 11506
rect 35982 11454 36034 11506
rect 9214 11342 9266 11394
rect 11678 11342 11730 11394
rect 15374 11342 15426 11394
rect 19630 11342 19682 11394
rect 19854 11342 19906 11394
rect 20190 11342 20242 11394
rect 22094 11342 22146 11394
rect 25342 11342 25394 11394
rect 31502 11342 31554 11394
rect 31950 11342 32002 11394
rect 32398 11342 32450 11394
rect 33182 11342 33234 11394
rect 36990 11342 37042 11394
rect 38782 11342 38834 11394
rect 76414 11342 76466 11394
rect 1710 11230 1762 11282
rect 2046 11230 2098 11282
rect 9550 11230 9602 11282
rect 11566 11230 11618 11282
rect 13806 11230 13858 11282
rect 16158 11230 16210 11282
rect 24894 11230 24946 11282
rect 25006 11230 25058 11282
rect 26126 11230 26178 11282
rect 30046 11230 30098 11282
rect 31390 11230 31442 11282
rect 32622 11230 32674 11282
rect 33854 11230 33906 11282
rect 37326 11230 37378 11282
rect 37886 11230 37938 11282
rect 41470 11230 41522 11282
rect 44830 11230 44882 11282
rect 45166 11230 45218 11282
rect 77870 11230 77922 11282
rect 78206 11230 78258 11282
rect 2494 11118 2546 11170
rect 11454 11118 11506 11170
rect 11902 11118 11954 11170
rect 13582 11118 13634 11170
rect 19742 11118 19794 11170
rect 24782 11118 24834 11170
rect 29822 11118 29874 11170
rect 31278 11118 31330 11170
rect 32174 11118 32226 11170
rect 32286 11118 32338 11170
rect 36430 11118 36482 11170
rect 37998 11118 38050 11170
rect 76190 11118 76242 11170
rect 77198 11118 77250 11170
rect 77646 11118 77698 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 50558 10950 50610 11002
rect 50662 10950 50714 11002
rect 50766 10950 50818 11002
rect 11118 10782 11170 10834
rect 11566 10782 11618 10834
rect 21758 10782 21810 10834
rect 24110 10782 24162 10834
rect 24334 10782 24386 10834
rect 25678 10782 25730 10834
rect 25790 10782 25842 10834
rect 25902 10782 25954 10834
rect 26798 10782 26850 10834
rect 31502 10782 31554 10834
rect 32510 10782 32562 10834
rect 39566 10782 39618 10834
rect 39678 10782 39730 10834
rect 39790 10782 39842 10834
rect 40350 10782 40402 10834
rect 2046 10670 2098 10722
rect 13358 10670 13410 10722
rect 18174 10670 18226 10722
rect 18398 10670 18450 10722
rect 33294 10670 33346 10722
rect 38782 10670 38834 10722
rect 39006 10670 39058 10722
rect 1710 10558 1762 10610
rect 11342 10558 11394 10610
rect 11902 10558 11954 10610
rect 12686 10558 12738 10610
rect 18846 10558 18898 10610
rect 22206 10558 22258 10610
rect 24782 10558 24834 10610
rect 26238 10558 26290 10610
rect 28142 10558 28194 10610
rect 31278 10558 31330 10610
rect 31950 10558 32002 10610
rect 38334 10558 38386 10610
rect 38670 10558 38722 10610
rect 39118 10558 39170 10610
rect 41470 10558 41522 10610
rect 78206 10558 78258 10610
rect 2494 10446 2546 10498
rect 11454 10446 11506 10498
rect 15486 10446 15538 10498
rect 18286 10446 18338 10498
rect 19518 10446 19570 10498
rect 22318 10446 22370 10498
rect 22542 10446 22594 10498
rect 24222 10446 24274 10498
rect 27806 10446 27858 10498
rect 28814 10446 28866 10498
rect 30942 10446 30994 10498
rect 31390 10446 31442 10498
rect 42142 10446 42194 10498
rect 44270 10446 44322 10498
rect 75854 10334 75906 10386
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 65918 10166 65970 10218
rect 66022 10166 66074 10218
rect 66126 10166 66178 10218
rect 8206 9998 8258 10050
rect 29150 9998 29202 10050
rect 29486 9998 29538 10050
rect 30270 9998 30322 10050
rect 31390 9998 31442 10050
rect 32398 9998 32450 10050
rect 32846 9998 32898 10050
rect 33070 9998 33122 10050
rect 35198 9998 35250 10050
rect 11566 9886 11618 9938
rect 13582 9886 13634 9938
rect 14478 9886 14530 9938
rect 15374 9886 15426 9938
rect 20750 9886 20802 9938
rect 31726 9886 31778 9938
rect 33182 9886 33234 9938
rect 34862 9886 34914 9938
rect 41806 9886 41858 9938
rect 42478 9886 42530 9938
rect 76302 9886 76354 9938
rect 8654 9774 8706 9826
rect 12238 9774 12290 9826
rect 12574 9774 12626 9826
rect 14030 9774 14082 9826
rect 20190 9774 20242 9826
rect 22766 9774 22818 9826
rect 31838 9774 31890 9826
rect 32286 9774 32338 9826
rect 35086 9774 35138 9826
rect 36990 9774 37042 9826
rect 37662 9774 37714 9826
rect 38222 9774 38274 9826
rect 38782 9774 38834 9826
rect 42366 9774 42418 9826
rect 42590 9774 42642 9826
rect 42926 9774 42978 9826
rect 1710 9662 1762 9714
rect 2046 9662 2098 9714
rect 8094 9662 8146 9714
rect 9326 9662 9378 9714
rect 13694 9662 13746 9714
rect 23550 9662 23602 9714
rect 26910 9662 26962 9714
rect 33742 9662 33794 9714
rect 37326 9662 37378 9714
rect 39454 9662 39506 9714
rect 40798 9662 40850 9714
rect 77646 9662 77698 9714
rect 77870 9662 77922 9714
rect 78206 9662 78258 9714
rect 2494 9550 2546 9602
rect 7982 9550 8034 9602
rect 12014 9550 12066 9602
rect 12126 9550 12178 9602
rect 13470 9550 13522 9602
rect 27246 9550 27298 9602
rect 27806 9550 27858 9602
rect 28254 9550 28306 9602
rect 28702 9550 28754 9602
rect 29262 9550 29314 9602
rect 30046 9550 30098 9602
rect 30494 9550 30546 9602
rect 30942 9550 30994 9602
rect 31278 9550 31330 9602
rect 31614 9550 31666 9602
rect 32846 9550 32898 9602
rect 33294 9550 33346 9602
rect 34078 9550 34130 9602
rect 37774 9550 37826 9602
rect 37998 9550 38050 9602
rect 38334 9550 38386 9602
rect 38558 9550 38610 9602
rect 38894 9550 38946 9602
rect 39118 9550 39170 9602
rect 40014 9550 40066 9602
rect 40910 9550 40962 9602
rect 42142 9550 42194 9602
rect 43038 9550 43090 9602
rect 43150 9550 43202 9602
rect 43374 9550 43426 9602
rect 43934 9550 43986 9602
rect 74846 9550 74898 9602
rect 75294 9550 75346 9602
rect 75630 9550 75682 9602
rect 77198 9550 77250 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 50558 9382 50610 9434
rect 50662 9382 50714 9434
rect 50766 9382 50818 9434
rect 13470 9214 13522 9266
rect 13806 9214 13858 9266
rect 14142 9214 14194 9266
rect 14478 9214 14530 9266
rect 14926 9214 14978 9266
rect 16158 9214 16210 9266
rect 18286 9214 18338 9266
rect 19182 9214 19234 9266
rect 22542 9214 22594 9266
rect 24670 9214 24722 9266
rect 25230 9214 25282 9266
rect 8766 9102 8818 9154
rect 15374 9102 15426 9154
rect 42590 9102 42642 9154
rect 9662 8990 9714 9042
rect 15934 8990 15986 9042
rect 18062 8990 18114 9042
rect 18734 8990 18786 9042
rect 19518 8990 19570 9042
rect 25454 8990 25506 9042
rect 26126 8990 26178 9042
rect 29374 8990 29426 9042
rect 33294 8990 33346 9042
rect 33966 8990 34018 9042
rect 37550 8990 37602 9042
rect 41470 8990 41522 9042
rect 41806 8990 41858 9042
rect 75182 8990 75234 9042
rect 76078 8990 76130 9042
rect 8878 8878 8930 8930
rect 10334 8878 10386 8930
rect 12462 8878 12514 8930
rect 13246 8878 13298 8930
rect 15374 8878 15426 8930
rect 16270 8878 16322 8930
rect 17726 8878 17778 8930
rect 18174 8878 18226 8930
rect 20302 8878 20354 8930
rect 23438 8878 23490 8930
rect 23886 8878 23938 8930
rect 24334 8878 24386 8930
rect 26910 8878 26962 8930
rect 29038 8878 29090 8930
rect 30158 8878 30210 8930
rect 32286 8878 32338 8930
rect 33518 8878 33570 8930
rect 34750 8878 34802 8930
rect 36878 8878 36930 8930
rect 38222 8878 38274 8930
rect 40350 8878 40402 8930
rect 41022 8878 41074 8930
rect 44718 8878 44770 8930
rect 45054 8878 45106 8930
rect 45278 8878 45330 8930
rect 77870 8878 77922 8930
rect 8990 8766 9042 8818
rect 15598 8766 15650 8818
rect 33630 8766 33682 8818
rect 73838 8766 73890 8818
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 65918 8598 65970 8650
rect 66022 8598 66074 8650
rect 66126 8598 66178 8650
rect 19294 8430 19346 8482
rect 28142 8430 28194 8482
rect 30270 8430 30322 8482
rect 41694 8430 41746 8482
rect 15374 8318 15426 8370
rect 17614 8318 17666 8370
rect 18174 8318 18226 8370
rect 19070 8318 19122 8370
rect 19854 8318 19906 8370
rect 20750 8318 20802 8370
rect 22430 8318 22482 8370
rect 24558 8318 24610 8370
rect 26910 8318 26962 8370
rect 27358 8318 27410 8370
rect 27582 8318 27634 8370
rect 30158 8318 30210 8370
rect 32286 8318 32338 8370
rect 34190 8318 34242 8370
rect 9774 8206 9826 8258
rect 14030 8206 14082 8258
rect 14702 8206 14754 8258
rect 18286 8206 18338 8258
rect 18734 8206 18786 8258
rect 19966 8206 20018 8258
rect 20414 8206 20466 8258
rect 21646 8206 21698 8258
rect 26350 8206 26402 8258
rect 26798 8206 26850 8258
rect 29038 8206 29090 8258
rect 32622 8206 32674 8258
rect 34302 8206 34354 8258
rect 34638 8206 34690 8258
rect 35310 8206 35362 8258
rect 38110 8206 38162 8258
rect 38670 8206 38722 8258
rect 39566 8206 39618 8258
rect 39902 8206 39954 8258
rect 40798 8206 40850 8258
rect 41358 8206 41410 8258
rect 42478 8206 42530 8258
rect 43038 8206 43090 8258
rect 44718 8206 44770 8258
rect 75294 8206 75346 8258
rect 78206 8206 78258 8258
rect 1710 8094 1762 8146
rect 2046 8094 2098 8146
rect 10558 8094 10610 8146
rect 14254 8094 14306 8146
rect 19742 8094 19794 8146
rect 28254 8094 28306 8146
rect 29262 8094 29314 8146
rect 29374 8094 29426 8146
rect 31502 8094 31554 8146
rect 34974 8094 35026 8146
rect 39118 8094 39170 8146
rect 40910 8094 40962 8146
rect 41022 8094 41074 8146
rect 42366 8094 42418 8146
rect 43710 8094 43762 8146
rect 44046 8094 44098 8146
rect 45054 8094 45106 8146
rect 76862 8094 76914 8146
rect 77198 8094 77250 8146
rect 77534 8094 77586 8146
rect 77870 8094 77922 8146
rect 2494 7982 2546 8034
rect 12798 7982 12850 8034
rect 13694 7982 13746 8034
rect 18062 7982 18114 8034
rect 19070 7982 19122 8034
rect 25342 7982 25394 8034
rect 25790 7982 25842 8034
rect 26238 7982 26290 8034
rect 27022 7982 27074 8034
rect 27582 7982 27634 8034
rect 28142 7982 28194 8034
rect 30046 7982 30098 8034
rect 30830 7982 30882 8034
rect 31278 7982 31330 8034
rect 31838 7982 31890 8034
rect 32958 7982 33010 8034
rect 33518 7982 33570 8034
rect 34078 7982 34130 8034
rect 35086 7982 35138 8034
rect 35870 7982 35922 8034
rect 37102 7982 37154 8034
rect 37662 7982 37714 8034
rect 37886 7982 37938 8034
rect 38782 7982 38834 8034
rect 38894 7982 38946 8034
rect 39678 7982 39730 8034
rect 42926 7982 42978 8034
rect 44942 7982 44994 8034
rect 45502 7982 45554 8034
rect 45950 7982 46002 8034
rect 74622 7982 74674 8034
rect 76526 7982 76578 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 50558 7814 50610 7866
rect 50662 7814 50714 7866
rect 50766 7814 50818 7866
rect 2046 7646 2098 7698
rect 8542 7646 8594 7698
rect 13134 7646 13186 7698
rect 13582 7646 13634 7698
rect 16942 7646 16994 7698
rect 18622 7646 18674 7698
rect 18846 7646 18898 7698
rect 19294 7646 19346 7698
rect 20078 7646 20130 7698
rect 20414 7646 20466 7698
rect 20862 7646 20914 7698
rect 23102 7646 23154 7698
rect 24782 7646 24834 7698
rect 25678 7646 25730 7698
rect 25902 7646 25954 7698
rect 27806 7646 27858 7698
rect 28366 7646 28418 7698
rect 29262 7646 29314 7698
rect 30046 7646 30098 7698
rect 30270 7646 30322 7698
rect 31726 7646 31778 7698
rect 33966 7646 34018 7698
rect 38110 7646 38162 7698
rect 39678 7646 39730 7698
rect 42030 7646 42082 7698
rect 71710 7646 71762 7698
rect 11006 7534 11058 7586
rect 14254 7534 14306 7586
rect 15598 7534 15650 7586
rect 18062 7534 18114 7586
rect 18398 7534 18450 7586
rect 26574 7534 26626 7586
rect 30382 7534 30434 7586
rect 31054 7534 31106 7586
rect 32510 7534 32562 7586
rect 33854 7534 33906 7586
rect 35198 7534 35250 7586
rect 38670 7534 38722 7586
rect 39230 7534 39282 7586
rect 40910 7534 40962 7586
rect 43038 7534 43090 7586
rect 44494 7534 44546 7586
rect 66670 7534 66722 7586
rect 1710 7422 1762 7474
rect 8318 7422 8370 7474
rect 13358 7422 13410 7474
rect 13918 7422 13970 7474
rect 14478 7422 14530 7474
rect 17726 7422 17778 7474
rect 19630 7422 19682 7474
rect 23438 7422 23490 7474
rect 25342 7422 25394 7474
rect 26350 7422 26402 7474
rect 26910 7422 26962 7474
rect 28926 7422 28978 7474
rect 29822 7422 29874 7474
rect 30718 7422 30770 7474
rect 32174 7422 32226 7474
rect 33406 7422 33458 7474
rect 34078 7422 34130 7474
rect 34414 7422 34466 7474
rect 40014 7422 40066 7474
rect 41246 7422 41298 7474
rect 41918 7422 41970 7474
rect 43934 7422 43986 7474
rect 46510 7422 46562 7474
rect 67006 7422 67058 7474
rect 72382 7422 72434 7474
rect 75294 7422 75346 7474
rect 2494 7310 2546 7362
rect 10222 7310 10274 7362
rect 10894 7310 10946 7362
rect 11230 7310 11282 7362
rect 11790 7310 11842 7362
rect 12686 7310 12738 7362
rect 13470 7310 13522 7362
rect 15262 7310 15314 7362
rect 15710 7310 15762 7362
rect 15822 7310 15874 7362
rect 16494 7310 16546 7362
rect 18510 7310 18562 7362
rect 21422 7310 21474 7362
rect 21870 7310 21922 7362
rect 22318 7310 22370 7362
rect 22766 7310 22818 7362
rect 23774 7310 23826 7362
rect 24334 7310 24386 7362
rect 25790 7310 25842 7362
rect 27470 7310 27522 7362
rect 31838 7310 31890 7362
rect 33294 7310 33346 7362
rect 37326 7310 37378 7362
rect 41582 7310 41634 7362
rect 46174 7310 46226 7362
rect 47070 7310 47122 7362
rect 47630 7310 47682 7362
rect 60174 7310 60226 7362
rect 73950 7310 74002 7362
rect 8654 7198 8706 7250
rect 21870 7198 21922 7250
rect 22094 7198 22146 7250
rect 22430 7198 22482 7250
rect 23214 7198 23266 7250
rect 23438 7198 23490 7250
rect 28702 7198 28754 7250
rect 29598 7198 29650 7250
rect 31502 7198 31554 7250
rect 38446 7198 38498 7250
rect 68014 7198 68066 7250
rect 76302 7198 76354 7250
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 65918 7030 65970 7082
rect 66022 7030 66074 7082
rect 66126 7030 66178 7082
rect 8206 6862 8258 6914
rect 8878 6862 8930 6914
rect 9214 6862 9266 6914
rect 7982 6750 8034 6802
rect 8766 6750 8818 6802
rect 9326 6750 9378 6802
rect 13582 6750 13634 6802
rect 15710 6750 15762 6802
rect 17838 6750 17890 6802
rect 25566 6750 25618 6802
rect 26238 6750 26290 6802
rect 28478 6750 28530 6802
rect 31502 6750 31554 6802
rect 31838 6750 31890 6802
rect 32734 6750 32786 6802
rect 36430 6750 36482 6802
rect 37998 6750 38050 6802
rect 40126 6750 40178 6802
rect 74734 6750 74786 6802
rect 76414 6750 76466 6802
rect 78094 6750 78146 6802
rect 12126 6638 12178 6690
rect 13694 6638 13746 6690
rect 14926 6638 14978 6690
rect 19966 6638 20018 6690
rect 21870 6638 21922 6690
rect 22654 6638 22706 6690
rect 23438 6638 23490 6690
rect 26126 6638 26178 6690
rect 26350 6638 26402 6690
rect 26798 6638 26850 6690
rect 27246 6638 27298 6690
rect 27918 6638 27970 6690
rect 28254 6638 28306 6690
rect 29374 6638 29426 6690
rect 30046 6638 30098 6690
rect 30606 6638 30658 6690
rect 30830 6638 30882 6690
rect 32622 6638 32674 6690
rect 32846 6638 32898 6690
rect 33294 6638 33346 6690
rect 33630 6638 33682 6690
rect 37326 6638 37378 6690
rect 40462 6638 40514 6690
rect 44270 6638 44322 6690
rect 46622 6638 46674 6690
rect 47070 6638 47122 6690
rect 49982 6638 50034 6690
rect 50990 6638 51042 6690
rect 51438 6638 51490 6690
rect 59502 6638 59554 6690
rect 60062 6638 60114 6690
rect 60510 6638 60562 6690
rect 63422 6638 63474 6690
rect 67902 6638 67954 6690
rect 68350 6638 68402 6690
rect 71262 6638 71314 6690
rect 74958 6638 75010 6690
rect 75182 6638 75234 6690
rect 76190 6638 76242 6690
rect 77086 6638 77138 6690
rect 77310 6638 77362 6690
rect 9438 6526 9490 6578
rect 19630 6526 19682 6578
rect 21534 6526 21586 6578
rect 22206 6526 22258 6578
rect 27022 6526 27074 6578
rect 30270 6526 30322 6578
rect 31166 6526 31218 6578
rect 34302 6526 34354 6578
rect 41582 6526 41634 6578
rect 43598 6526 43650 6578
rect 46062 6526 46114 6578
rect 48638 6526 48690 6578
rect 50542 6526 50594 6578
rect 6638 6414 6690 6466
rect 7086 6414 7138 6466
rect 7646 6414 7698 6466
rect 7982 6414 8034 6466
rect 8654 6414 8706 6466
rect 10222 6414 10274 6466
rect 10894 6414 10946 6466
rect 11678 6414 11730 6466
rect 12574 6414 12626 6466
rect 13022 6414 13074 6466
rect 13470 6414 13522 6466
rect 13918 6414 13970 6466
rect 14702 6414 14754 6466
rect 18958 6414 19010 6466
rect 19406 6414 19458 6466
rect 20862 6414 20914 6466
rect 29598 6414 29650 6466
rect 31614 6414 31666 6466
rect 32398 6414 32450 6466
rect 40686 6414 40738 6466
rect 47070 6414 47122 6466
rect 49086 6414 49138 6466
rect 49646 6414 49698 6466
rect 51886 6414 51938 6466
rect 56814 6414 56866 6466
rect 61518 6414 61570 6466
rect 64430 6414 64482 6466
rect 67342 6414 67394 6466
rect 69358 6414 69410 6466
rect 72270 6414 72322 6466
rect 75518 6414 75570 6466
rect 76750 6414 76802 6466
rect 77646 6414 77698 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 50558 6246 50610 6298
rect 50662 6246 50714 6298
rect 50766 6246 50818 6298
rect 2046 6078 2098 6130
rect 8318 6078 8370 6130
rect 8654 6078 8706 6130
rect 13918 6078 13970 6130
rect 14366 6078 14418 6130
rect 14814 6078 14866 6130
rect 15150 6078 15202 6130
rect 15598 6078 15650 6130
rect 18062 6078 18114 6130
rect 18286 6078 18338 6130
rect 21534 6078 21586 6130
rect 26350 6078 26402 6130
rect 27918 6078 27970 6130
rect 28926 6078 28978 6130
rect 34190 6078 34242 6130
rect 34414 6078 34466 6130
rect 34638 6078 34690 6130
rect 36094 6078 36146 6130
rect 40238 6078 40290 6130
rect 41134 6078 41186 6130
rect 44046 6078 44098 6130
rect 46734 6078 46786 6130
rect 47966 6078 48018 6130
rect 49646 6078 49698 6130
rect 50766 6078 50818 6130
rect 53902 6078 53954 6130
rect 56030 6078 56082 6130
rect 63870 6078 63922 6130
rect 71038 6078 71090 6130
rect 78206 6078 78258 6130
rect 6638 5966 6690 6018
rect 8990 5966 9042 6018
rect 13694 5966 13746 6018
rect 14142 5966 14194 6018
rect 15710 5966 15762 6018
rect 16494 5966 16546 6018
rect 16830 5966 16882 6018
rect 22654 5966 22706 6018
rect 23326 5966 23378 6018
rect 23662 5966 23714 6018
rect 23998 5966 24050 6018
rect 24334 5966 24386 6018
rect 24670 5966 24722 6018
rect 25566 5966 25618 6018
rect 26126 5966 26178 6018
rect 27470 5966 27522 6018
rect 30382 5966 30434 6018
rect 35646 5966 35698 6018
rect 37662 5966 37714 6018
rect 39566 5966 39618 6018
rect 40014 5966 40066 6018
rect 42254 5966 42306 6018
rect 43150 5966 43202 6018
rect 45166 5966 45218 6018
rect 48750 5966 48802 6018
rect 63198 5966 63250 6018
rect 1710 5854 1762 5906
rect 7982 5854 8034 5906
rect 9886 5854 9938 5906
rect 14030 5854 14082 5906
rect 17390 5854 17442 5906
rect 17726 5854 17778 5906
rect 18174 5854 18226 5906
rect 18734 5854 18786 5906
rect 21758 5854 21810 5906
rect 22318 5854 22370 5906
rect 22990 5854 23042 5906
rect 26798 5854 26850 5906
rect 28254 5854 28306 5906
rect 28478 5854 28530 5906
rect 29262 5854 29314 5906
rect 29710 5854 29762 5906
rect 33854 5854 33906 5906
rect 35086 5854 35138 5906
rect 37102 5854 37154 5906
rect 39342 5854 39394 5906
rect 41806 5854 41858 5906
rect 44270 5854 44322 5906
rect 46398 5854 46450 5906
rect 47070 5854 47122 5906
rect 47630 5854 47682 5906
rect 49086 5854 49138 5906
rect 49870 5854 49922 5906
rect 56926 5854 56978 5906
rect 59838 5854 59890 5906
rect 64430 5854 64482 5906
rect 67342 5854 67394 5906
rect 71710 5854 71762 5906
rect 72270 5854 72322 5906
rect 77310 5854 77362 5906
rect 2494 5742 2546 5794
rect 5294 5742 5346 5794
rect 5742 5742 5794 5794
rect 6190 5742 6242 5794
rect 7086 5742 7138 5794
rect 7534 5742 7586 5794
rect 10670 5742 10722 5794
rect 12798 5742 12850 5794
rect 19182 5742 19234 5794
rect 19630 5742 19682 5794
rect 20078 5742 20130 5794
rect 20526 5742 20578 5794
rect 21198 5742 21250 5794
rect 23214 5742 23266 5794
rect 25454 5742 25506 5794
rect 26238 5742 26290 5794
rect 27246 5742 27298 5794
rect 27582 5742 27634 5794
rect 32510 5742 32562 5794
rect 33294 5742 33346 5794
rect 34302 5742 34354 5794
rect 47294 5742 47346 5794
rect 51214 5742 51266 5794
rect 51662 5742 51714 5794
rect 52558 5742 52610 5794
rect 65550 5742 65602 5794
rect 68910 5742 68962 5794
rect 70478 5742 70530 5794
rect 75630 5742 75682 5794
rect 7534 5630 7586 5682
rect 8206 5630 8258 5682
rect 15486 5630 15538 5682
rect 17390 5630 17442 5682
rect 21422 5630 21474 5682
rect 25790 5630 25842 5682
rect 33518 5630 33570 5682
rect 33854 5630 33906 5682
rect 41582 5630 41634 5682
rect 42030 5630 42082 5682
rect 57934 5630 57986 5682
rect 60846 5630 60898 5682
rect 73278 5630 73330 5682
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 65918 5462 65970 5514
rect 66022 5462 66074 5514
rect 66126 5462 66178 5514
rect 8990 5294 9042 5346
rect 10782 5294 10834 5346
rect 12014 5294 12066 5346
rect 20750 5294 20802 5346
rect 21534 5294 21586 5346
rect 26574 5294 26626 5346
rect 28590 5294 28642 5346
rect 30942 5294 30994 5346
rect 69358 5294 69410 5346
rect 10222 5182 10274 5234
rect 10670 5182 10722 5234
rect 11454 5182 11506 5234
rect 12462 5182 12514 5234
rect 13694 5182 13746 5234
rect 14142 5182 14194 5234
rect 14702 5182 14754 5234
rect 16718 5182 16770 5234
rect 18958 5182 19010 5234
rect 19518 5182 19570 5234
rect 20638 5182 20690 5234
rect 21758 5182 21810 5234
rect 22430 5182 22482 5234
rect 23662 5182 23714 5234
rect 25790 5182 25842 5234
rect 26462 5182 26514 5234
rect 27806 5182 27858 5234
rect 27918 5182 27970 5234
rect 28366 5182 28418 5234
rect 29598 5182 29650 5234
rect 30830 5182 30882 5234
rect 31838 5182 31890 5234
rect 49758 5182 49810 5234
rect 50094 5182 50146 5234
rect 55246 5182 55298 5234
rect 58158 5182 58210 5234
rect 64430 5182 64482 5234
rect 66446 5182 66498 5234
rect 67118 5182 67170 5234
rect 67454 5182 67506 5234
rect 72270 5182 72322 5234
rect 74734 5182 74786 5234
rect 75518 5182 75570 5234
rect 1710 5070 1762 5122
rect 2494 5070 2546 5122
rect 6190 5070 6242 5122
rect 6526 5070 6578 5122
rect 7310 5070 7362 5122
rect 8206 5070 8258 5122
rect 8654 5070 8706 5122
rect 8878 5070 8930 5122
rect 9662 5070 9714 5122
rect 11678 5070 11730 5122
rect 12350 5070 12402 5122
rect 12910 5070 12962 5122
rect 15598 5070 15650 5122
rect 15934 5070 15986 5122
rect 19406 5070 19458 5122
rect 19742 5070 19794 5122
rect 20414 5070 20466 5122
rect 21870 5070 21922 5122
rect 22878 5070 22930 5122
rect 27246 5070 27298 5122
rect 27582 5070 27634 5122
rect 28254 5070 28306 5122
rect 29262 5070 29314 5122
rect 29486 5070 29538 5122
rect 30606 5070 30658 5122
rect 31390 5070 31442 5122
rect 32286 5070 32338 5122
rect 32622 5070 32674 5122
rect 36430 5070 36482 5122
rect 37102 5070 37154 5122
rect 37326 5070 37378 5122
rect 37550 5070 37602 5122
rect 39566 5070 39618 5122
rect 40014 5070 40066 5122
rect 40462 5070 40514 5122
rect 42702 5070 42754 5122
rect 44830 5070 44882 5122
rect 46846 5070 46898 5122
rect 49198 5070 49250 5122
rect 50542 5070 50594 5122
rect 51102 5070 51154 5122
rect 51550 5070 51602 5122
rect 53566 5070 53618 5122
rect 54238 5070 54290 5122
rect 57150 5070 57202 5122
rect 60622 5070 60674 5122
rect 63534 5070 63586 5122
rect 68462 5070 68514 5122
rect 71374 5070 71426 5122
rect 75070 5070 75122 5122
rect 76526 5070 76578 5122
rect 77422 5070 77474 5122
rect 77870 5070 77922 5122
rect 2046 4958 2098 5010
rect 6750 4958 6802 5010
rect 7646 4958 7698 5010
rect 7982 4958 8034 5010
rect 9326 4958 9378 5010
rect 10558 4958 10610 5010
rect 12574 4958 12626 5010
rect 14030 4958 14082 5010
rect 14254 4958 14306 5010
rect 14702 4958 14754 5010
rect 14926 4958 14978 5010
rect 22542 4958 22594 5010
rect 26910 4958 26962 5010
rect 29934 4958 29986 5010
rect 30270 4958 30322 5010
rect 33294 4958 33346 5010
rect 35310 4958 35362 5010
rect 38334 4958 38386 5010
rect 38894 4958 38946 5010
rect 39118 4958 39170 5010
rect 39790 4958 39842 5010
rect 40126 4958 40178 5010
rect 40574 4958 40626 5010
rect 43150 4958 43202 5010
rect 45390 4958 45442 5010
rect 47406 4958 47458 5010
rect 48974 4958 49026 5010
rect 76190 4958 76242 5010
rect 77198 4958 77250 5010
rect 78206 4958 78258 5010
rect 4286 4846 4338 4898
rect 4734 4846 4786 4898
rect 5182 4846 5234 4898
rect 7534 4846 7586 4898
rect 11902 4846 11954 4898
rect 15262 4846 15314 4898
rect 22318 4846 22370 4898
rect 26350 4846 26402 4898
rect 33966 4846 34018 4898
rect 42814 4846 42866 4898
rect 45838 4846 45890 4898
rect 52110 4846 52162 4898
rect 53230 4846 53282 4898
rect 61518 4846 61570 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 50558 4678 50610 4730
rect 50662 4678 50714 4730
rect 50766 4678 50818 4730
rect 4286 4510 4338 4562
rect 4958 4510 5010 4562
rect 5630 4510 5682 4562
rect 6078 4510 6130 4562
rect 6190 4510 6242 4562
rect 8990 4510 9042 4562
rect 16718 4510 16770 4562
rect 17838 4510 17890 4562
rect 18622 4510 18674 4562
rect 19630 4510 19682 4562
rect 20638 4510 20690 4562
rect 21198 4510 21250 4562
rect 32398 4510 32450 4562
rect 33182 4510 33234 4562
rect 40238 4510 40290 4562
rect 42142 4510 42194 4562
rect 48750 4510 48802 4562
rect 55918 4510 55970 4562
rect 63198 4510 63250 4562
rect 71038 4510 71090 4562
rect 71710 4510 71762 4562
rect 78206 4510 78258 4562
rect 7646 4398 7698 4450
rect 8318 4398 8370 4450
rect 9886 4398 9938 4450
rect 17950 4398 18002 4450
rect 18286 4398 18338 4450
rect 19294 4398 19346 4450
rect 19966 4398 20018 4450
rect 20302 4398 20354 4450
rect 21310 4398 21362 4450
rect 21758 4398 21810 4450
rect 21982 4398 22034 4450
rect 22654 4398 22706 4450
rect 22990 4398 23042 4450
rect 23102 4398 23154 4450
rect 23214 4398 23266 4450
rect 23998 4398 24050 4450
rect 24334 4398 24386 4450
rect 24670 4398 24722 4450
rect 28814 4398 28866 4450
rect 31390 4398 31442 4450
rect 33294 4398 33346 4450
rect 34190 4398 34242 4450
rect 36654 4398 36706 4450
rect 39118 4398 39170 4450
rect 40910 4398 40962 4450
rect 41582 4398 41634 4450
rect 42590 4398 42642 4450
rect 45614 4398 45666 4450
rect 46622 4398 46674 4450
rect 46958 4398 47010 4450
rect 62526 4398 62578 4450
rect 4062 4286 4114 4338
rect 4622 4286 4674 4338
rect 5406 4286 5458 4338
rect 6638 4286 6690 4338
rect 7310 4286 7362 4338
rect 7982 4286 8034 4338
rect 8766 4286 8818 4338
rect 9662 4286 9714 4338
rect 10222 4286 10274 4338
rect 13694 4286 13746 4338
rect 17614 4286 17666 4338
rect 18958 4286 19010 4338
rect 20974 4286 21026 4338
rect 22430 4286 22482 4338
rect 23774 4286 23826 4338
rect 25230 4286 25282 4338
rect 28702 4286 28754 4338
rect 30830 4286 30882 4338
rect 32958 4286 33010 4338
rect 33966 4286 34018 4338
rect 35982 4286 36034 4338
rect 36542 4286 36594 4338
rect 38670 4286 38722 4338
rect 44158 4286 44210 4338
rect 46286 4286 46338 4338
rect 47294 4286 47346 4338
rect 49086 4286 49138 4338
rect 49534 4286 49586 4338
rect 52558 4286 52610 4338
rect 52894 4286 52946 4338
rect 56590 4286 56642 4338
rect 61630 4286 61682 4338
rect 64542 4286 64594 4338
rect 67454 4286 67506 4338
rect 72270 4286 72322 4338
rect 75182 4286 75234 4338
rect 2158 4174 2210 4226
rect 2494 4174 2546 4226
rect 3278 4174 3330 4226
rect 3726 4174 3778 4226
rect 6750 4174 6802 4226
rect 8206 4174 8258 4226
rect 11006 4174 11058 4226
rect 13134 4174 13186 4226
rect 14478 4174 14530 4226
rect 19070 4174 19122 4226
rect 21758 4174 21810 4226
rect 26014 4174 26066 4226
rect 28142 4174 28194 4226
rect 35086 4174 35138 4226
rect 41246 4174 41298 4226
rect 45278 4174 45330 4226
rect 63534 4174 63586 4226
rect 65550 4174 65602 4226
rect 70478 4174 70530 4226
rect 6302 4062 6354 4114
rect 6974 4062 7026 4114
rect 50542 4062 50594 4114
rect 53902 4062 53954 4114
rect 57598 4062 57650 4114
rect 59726 4062 59778 4114
rect 62638 4062 62690 4114
rect 63534 4062 63586 4114
rect 68350 4062 68402 4114
rect 73278 4062 73330 4114
rect 76190 4062 76242 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 65918 3894 65970 3946
rect 66022 3894 66074 3946
rect 66126 3894 66178 3946
rect 11230 3726 11282 3778
rect 15710 3726 15762 3778
rect 17502 3726 17554 3778
rect 21646 3726 21698 3778
rect 21982 3726 22034 3778
rect 25118 3726 25170 3778
rect 67454 3726 67506 3778
rect 75070 3726 75122 3778
rect 11118 3614 11170 3666
rect 15598 3614 15650 3666
rect 17278 3614 17330 3666
rect 23438 3614 23490 3666
rect 25006 3614 25058 3666
rect 39342 3614 39394 3666
rect 41806 3614 41858 3666
rect 45726 3614 45778 3666
rect 47406 3614 47458 3666
rect 50654 3614 50706 3666
rect 51774 3614 51826 3666
rect 56030 3614 56082 3666
rect 58046 3614 58098 3666
rect 59054 3614 59106 3666
rect 61854 3614 61906 3666
rect 63870 3614 63922 3666
rect 65662 3614 65714 3666
rect 69806 3614 69858 3666
rect 71262 3614 71314 3666
rect 77198 3614 77250 3666
rect 1822 3502 1874 3554
rect 3390 3502 3442 3554
rect 4734 3502 4786 3554
rect 5854 3502 5906 3554
rect 6526 3502 6578 3554
rect 7086 3502 7138 3554
rect 7758 3502 7810 3554
rect 8542 3502 8594 3554
rect 9662 3502 9714 3554
rect 10222 3502 10274 3554
rect 10894 3502 10946 3554
rect 11678 3502 11730 3554
rect 12238 3502 12290 3554
rect 13470 3502 13522 3554
rect 14142 3502 14194 3554
rect 14814 3502 14866 3554
rect 15374 3502 15426 3554
rect 16046 3502 16098 3554
rect 18622 3502 18674 3554
rect 19182 3502 19234 3554
rect 19966 3502 20018 3554
rect 21086 3502 21138 3554
rect 21646 3502 21698 3554
rect 22990 3502 23042 3554
rect 24782 3502 24834 3554
rect 25454 3502 25506 3554
rect 26126 3502 26178 3554
rect 26910 3502 26962 3554
rect 27582 3502 27634 3554
rect 28590 3502 28642 3554
rect 29374 3502 29426 3554
rect 30046 3502 30098 3554
rect 31390 3502 31442 3554
rect 32398 3502 32450 3554
rect 33070 3502 33122 3554
rect 33742 3502 33794 3554
rect 34526 3502 34578 3554
rect 35086 3502 35138 3554
rect 36878 3502 36930 3554
rect 37662 3502 37714 3554
rect 41358 3502 41410 3554
rect 43038 3502 43090 3554
rect 43710 3502 43762 3554
rect 45278 3502 45330 3554
rect 47966 3502 48018 3554
rect 48190 3502 48242 3554
rect 48750 3502 48802 3554
rect 49422 3502 49474 3554
rect 50094 3502 50146 3554
rect 52334 3502 52386 3554
rect 53006 3502 53058 3554
rect 53678 3502 53730 3554
rect 54238 3502 54290 3554
rect 55022 3502 55074 3554
rect 61406 3502 61458 3554
rect 62638 3502 62690 3554
rect 66446 3502 66498 3554
rect 70254 3502 70306 3554
rect 74062 3502 74114 3554
rect 78094 3502 78146 3554
rect 2046 3390 2098 3442
rect 2382 3390 2434 3442
rect 2718 3390 2770 3442
rect 3614 3390 3666 3442
rect 3950 3390 4002 3442
rect 4286 3390 4338 3442
rect 4958 3390 5010 3442
rect 6078 3390 6130 3442
rect 7422 3390 7474 3442
rect 8766 3390 8818 3442
rect 12574 3390 12626 3442
rect 13694 3390 13746 3442
rect 14366 3390 14418 3442
rect 15038 3390 15090 3442
rect 17838 3390 17890 3442
rect 18174 3390 18226 3442
rect 19518 3390 19570 3442
rect 20190 3390 20242 3442
rect 22318 3390 22370 3442
rect 22654 3390 22706 3442
rect 25790 3390 25842 3442
rect 26462 3390 26514 3442
rect 27134 3390 27186 3442
rect 29598 3390 29650 3442
rect 30270 3390 30322 3442
rect 30606 3390 30658 3442
rect 32734 3390 32786 3442
rect 33406 3390 33458 3442
rect 34078 3390 34130 3442
rect 34750 3390 34802 3442
rect 35422 3390 35474 3442
rect 36766 3390 36818 3442
rect 37550 3390 37602 3442
rect 41470 3390 41522 3442
rect 42254 3390 42306 3442
rect 44382 3390 44434 3442
rect 45390 3390 45442 3442
rect 48526 3390 48578 3442
rect 49198 3390 49250 3442
rect 49870 3390 49922 3442
rect 51214 3390 51266 3442
rect 52782 3390 52834 3442
rect 53454 3390 53506 3442
rect 73614 3390 73666 3442
rect 77870 3390 77922 3442
rect 6750 3278 6802 3330
rect 8094 3278 8146 3330
rect 9886 3278 9938 3330
rect 10558 3278 10610 3330
rect 11902 3278 11954 3330
rect 16382 3278 16434 3330
rect 17278 3278 17330 3330
rect 18846 3278 18898 3330
rect 21310 3278 21362 3330
rect 24110 3278 24162 3330
rect 27806 3278 27858 3330
rect 28926 3278 28978 3330
rect 30942 3278 30994 3330
rect 31614 3278 31666 3330
rect 52110 3278 52162 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
rect 50558 3110 50610 3162
rect 50662 3110 50714 3162
rect 50766 3110 50818 3162
rect 18622 2942 18674 2994
rect 22430 2942 22482 2994
<< metal2 >>
rect 448 79200 560 80000
rect 1120 79200 1232 80000
rect 1792 79200 1904 80000
rect 2464 79200 2576 80000
rect 3136 79200 3248 80000
rect 3808 79200 3920 80000
rect 4480 79200 4592 80000
rect 5152 79200 5264 80000
rect 5824 79200 5936 80000
rect 6496 79200 6608 80000
rect 7168 79200 7280 80000
rect 7840 79200 7952 80000
rect 8512 79200 8624 80000
rect 9184 79200 9296 80000
rect 9856 79200 9968 80000
rect 10528 79200 10640 80000
rect 11200 79200 11312 80000
rect 11872 79200 11984 80000
rect 12544 79200 12656 80000
rect 13216 79200 13328 80000
rect 13888 79200 14000 80000
rect 14560 79200 14672 80000
rect 15232 79200 15344 80000
rect 15904 79200 16016 80000
rect 16576 79200 16688 80000
rect 17248 79200 17360 80000
rect 17920 79200 18032 80000
rect 18592 79200 18704 80000
rect 19264 79200 19376 80000
rect 19936 79200 20048 80000
rect 20608 79200 20720 80000
rect 21280 79200 21392 80000
rect 21952 79200 22064 80000
rect 22624 79200 22736 80000
rect 23296 79200 23408 80000
rect 23968 79200 24080 80000
rect 24640 79200 24752 80000
rect 25312 79200 25424 80000
rect 25984 79200 26096 80000
rect 26656 79200 26768 80000
rect 27328 79200 27440 80000
rect 28000 79200 28112 80000
rect 28672 79200 28784 80000
rect 29344 79200 29456 80000
rect 30016 79200 30128 80000
rect 30688 79200 30800 80000
rect 31360 79200 31472 80000
rect 32032 79200 32144 80000
rect 32704 79200 32816 80000
rect 33376 79200 33488 80000
rect 34048 79200 34160 80000
rect 34720 79200 34832 80000
rect 35392 79200 35504 80000
rect 36064 79200 36176 80000
rect 36736 79200 36848 80000
rect 37408 79200 37520 80000
rect 38080 79200 38192 80000
rect 38752 79200 38864 80000
rect 39424 79200 39536 80000
rect 40096 79200 40208 80000
rect 40768 79200 40880 80000
rect 41440 79200 41552 80000
rect 42112 79200 42224 80000
rect 42784 79200 42896 80000
rect 43456 79200 43568 80000
rect 44128 79200 44240 80000
rect 44800 79200 44912 80000
rect 45472 79200 45584 80000
rect 46144 79200 46256 80000
rect 46816 79200 46928 80000
rect 47488 79200 47600 80000
rect 48160 79200 48272 80000
rect 48832 79200 48944 80000
rect 49504 79200 49616 80000
rect 50176 79200 50288 80000
rect 50848 79200 50960 80000
rect 51520 79200 51632 80000
rect 52192 79200 52304 80000
rect 52864 79200 52976 80000
rect 53536 79200 53648 80000
rect 54208 79200 54320 80000
rect 54880 79200 54992 80000
rect 55552 79200 55664 80000
rect 56224 79200 56336 80000
rect 56896 79200 57008 80000
rect 57568 79200 57680 80000
rect 58240 79200 58352 80000
rect 58912 79200 59024 80000
rect 59584 79200 59696 80000
rect 60256 79200 60368 80000
rect 60928 79200 61040 80000
rect 61600 79200 61712 80000
rect 62272 79200 62384 80000
rect 62944 79200 63056 80000
rect 63616 79200 63728 80000
rect 64288 79200 64400 80000
rect 64960 79200 65072 80000
rect 65632 79200 65744 80000
rect 66304 79200 66416 80000
rect 66976 79200 67088 80000
rect 67648 79200 67760 80000
rect 68320 79200 68432 80000
rect 68992 79200 69104 80000
rect 69664 79200 69776 80000
rect 70336 79200 70448 80000
rect 71008 79200 71120 80000
rect 71680 79200 71792 80000
rect 72352 79200 72464 80000
rect 73024 79200 73136 80000
rect 73696 79200 73808 80000
rect 74368 79200 74480 80000
rect 75040 79200 75152 80000
rect 75712 79200 75824 80000
rect 76384 79200 76496 80000
rect 77056 79200 77168 80000
rect 77728 79200 77840 80000
rect 78400 79200 78512 80000
rect 79072 79200 79184 80000
rect 2156 77364 2212 77374
rect 1932 76244 1988 76254
rect 1932 76150 1988 76188
rect 1932 75794 1988 75806
rect 1932 75742 1934 75794
rect 1986 75742 1988 75794
rect 1932 75348 1988 75742
rect 1932 75282 1988 75292
rect 2156 74786 2212 77308
rect 4620 76692 4676 76702
rect 4172 76690 4676 76692
rect 4172 76638 4622 76690
rect 4674 76638 4676 76690
rect 4172 76636 4676 76638
rect 4172 74898 4228 76636
rect 4620 76626 4676 76636
rect 4956 76580 5012 76590
rect 5516 76580 5572 76590
rect 4956 76578 5572 76580
rect 4956 76526 4958 76578
rect 5010 76526 5518 76578
rect 5570 76526 5572 76578
rect 4956 76524 5572 76526
rect 4284 76466 4340 76478
rect 4284 76414 4286 76466
rect 4338 76414 4340 76466
rect 4284 75908 4340 76414
rect 4476 76076 4740 76086
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4476 76010 4740 76020
rect 4284 75852 4676 75908
rect 4284 75684 4340 75694
rect 4284 75682 4564 75684
rect 4284 75630 4286 75682
rect 4338 75630 4564 75682
rect 4284 75628 4564 75630
rect 4284 75618 4340 75628
rect 4508 75124 4564 75628
rect 4620 75570 4676 75852
rect 4956 75682 5012 76524
rect 5516 76514 5572 76524
rect 4956 75630 4958 75682
rect 5010 75630 5012 75682
rect 4956 75618 5012 75630
rect 5740 76466 5796 76478
rect 5740 76414 5742 76466
rect 5794 76414 5796 76466
rect 4620 75518 4622 75570
rect 4674 75518 4676 75570
rect 4620 75506 4676 75518
rect 4620 75124 4676 75134
rect 4508 75122 4676 75124
rect 4508 75070 4622 75122
rect 4674 75070 4676 75122
rect 4508 75068 4676 75070
rect 4620 75058 4676 75068
rect 4172 74846 4174 74898
rect 4226 74846 4228 74898
rect 4172 74834 4228 74846
rect 4844 74898 4900 74910
rect 4844 74846 4846 74898
rect 4898 74846 4900 74898
rect 2156 74734 2158 74786
rect 2210 74734 2212 74786
rect 2156 74722 2212 74734
rect 4476 74508 4740 74518
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4476 74442 4740 74452
rect 1932 74228 1988 74238
rect 1932 74134 1988 74172
rect 4284 74116 4340 74126
rect 4284 74114 4676 74116
rect 4284 74062 4286 74114
rect 4338 74062 4676 74114
rect 4284 74060 4676 74062
rect 4284 74050 4340 74060
rect 4620 74002 4676 74060
rect 4620 73950 4622 74002
rect 4674 73950 4676 74002
rect 4620 73938 4676 73950
rect 4844 74114 4900 74846
rect 4844 74062 4846 74114
rect 4898 74062 4900 74114
rect 4620 73444 4676 73454
rect 4284 73442 4676 73444
rect 4284 73390 4622 73442
rect 4674 73390 4676 73442
rect 4284 73388 4676 73390
rect 4284 73330 4340 73388
rect 4620 73378 4676 73388
rect 4284 73278 4286 73330
rect 4338 73278 4340 73330
rect 4284 73266 4340 73278
rect 4844 73330 4900 74062
rect 4844 73278 4846 73330
rect 4898 73278 4900 73330
rect 1932 73108 1988 73118
rect 1932 73014 1988 73052
rect 4476 72940 4740 72950
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4476 72874 4740 72884
rect 1932 72658 1988 72670
rect 1932 72606 1934 72658
rect 1986 72606 1988 72658
rect 1932 71988 1988 72606
rect 2940 72548 2996 72558
rect 3836 72548 3892 72558
rect 1932 71922 1988 71932
rect 2492 71988 2548 71998
rect 2940 71988 2996 72492
rect 3500 72546 3892 72548
rect 3500 72494 3838 72546
rect 3890 72494 3892 72546
rect 3500 72492 3892 72494
rect 2492 71986 2996 71988
rect 2492 71934 2494 71986
rect 2546 71934 2996 71986
rect 2492 71932 2996 71934
rect 2492 71922 2548 71932
rect 2156 71762 2212 71774
rect 2156 71710 2158 71762
rect 2210 71710 2212 71762
rect 1932 71652 1988 71662
rect 2156 71652 2212 71710
rect 1820 71650 2212 71652
rect 1820 71598 1934 71650
rect 1986 71598 2212 71650
rect 1820 71596 2212 71598
rect 2940 71762 2996 71932
rect 3164 71988 3220 71998
rect 3164 71894 3220 71932
rect 3500 71986 3556 72492
rect 3836 72482 3892 72492
rect 4620 72324 4676 72334
rect 4844 72324 4900 73278
rect 4956 72548 5012 72558
rect 4956 72454 5012 72492
rect 5740 72548 5796 76414
rect 5740 72482 5796 72492
rect 8316 76356 8372 76366
rect 4620 72322 4900 72324
rect 4620 72270 4622 72322
rect 4674 72270 4900 72322
rect 4620 72268 4900 72270
rect 4620 72212 4676 72268
rect 3500 71934 3502 71986
rect 3554 71934 3556 71986
rect 3500 71922 3556 71934
rect 3836 72156 4676 72212
rect 3836 71874 3892 72156
rect 3836 71822 3838 71874
rect 3890 71822 3892 71874
rect 3836 71810 3892 71822
rect 3948 71988 4004 71998
rect 2940 71710 2942 71762
rect 2994 71710 2996 71762
rect 1820 43708 1876 71596
rect 1932 71586 1988 71596
rect 1932 71090 1988 71102
rect 1932 71038 1934 71090
rect 1986 71038 1988 71090
rect 1932 70644 1988 71038
rect 1932 70578 1988 70588
rect 2716 70196 2772 70206
rect 1932 69970 1988 69982
rect 1932 69918 1934 69970
rect 1986 69918 1988 69970
rect 1932 69524 1988 69918
rect 1932 69458 1988 69468
rect 2380 69298 2436 69310
rect 2380 69246 2382 69298
rect 2434 69246 2436 69298
rect 2044 69186 2100 69198
rect 2044 69134 2046 69186
rect 2098 69134 2100 69186
rect 2044 68626 2100 69134
rect 2044 68574 2046 68626
rect 2098 68574 2100 68626
rect 2044 68562 2100 68574
rect 1932 67954 1988 67966
rect 1932 67902 1934 67954
rect 1986 67902 1988 67954
rect 1932 67284 1988 67902
rect 1932 67218 1988 67228
rect 2380 67228 2436 69246
rect 2716 69298 2772 70140
rect 2940 69410 2996 71710
rect 3948 70978 4004 71932
rect 4476 71372 4740 71382
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4476 71306 4740 71316
rect 3948 70926 3950 70978
rect 4002 70926 4004 70978
rect 3948 70914 4004 70926
rect 3836 70196 3892 70206
rect 3836 70102 3892 70140
rect 4476 69804 4740 69814
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4476 69738 4740 69748
rect 2940 69358 2942 69410
rect 2994 69358 2996 69410
rect 2940 69346 2996 69358
rect 2716 69246 2718 69298
rect 2770 69246 2772 69298
rect 2716 69234 2772 69246
rect 2716 68404 2772 68414
rect 2716 68310 2772 68348
rect 4476 68236 4740 68246
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4476 68170 4740 68180
rect 4060 67842 4116 67854
rect 4060 67790 4062 67842
rect 4114 67790 4116 67842
rect 4060 67282 4116 67790
rect 4060 67230 4062 67282
rect 4114 67230 4116 67282
rect 2044 67170 2100 67182
rect 2380 67172 2772 67228
rect 4060 67218 4116 67230
rect 2044 67118 2046 67170
rect 2098 67118 2100 67170
rect 1932 66388 1988 66398
rect 1932 66294 1988 66332
rect 2044 65490 2100 67118
rect 2716 67078 2772 67116
rect 3052 67170 3108 67182
rect 3052 67118 3054 67170
rect 3106 67118 3108 67170
rect 2044 65438 2046 65490
rect 2098 65438 2100 65490
rect 2044 65426 2100 65438
rect 2268 67060 2324 67070
rect 1932 64818 1988 64830
rect 1932 64766 1934 64818
rect 1986 64766 1988 64818
rect 1932 63924 1988 64766
rect 1932 63858 1988 63868
rect 2268 63922 2324 67004
rect 2380 67058 2436 67070
rect 2380 67006 2382 67058
rect 2434 67006 2436 67058
rect 2380 64148 2436 67006
rect 3052 66276 3108 67118
rect 3724 67172 3780 67182
rect 3724 67078 3780 67116
rect 4284 67172 4340 67182
rect 3388 67060 3444 67070
rect 3388 66966 3444 67004
rect 4284 67058 4340 67116
rect 4284 67006 4286 67058
rect 4338 67006 4340 67058
rect 4284 66994 4340 67006
rect 4476 66668 4740 66678
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4476 66602 4740 66612
rect 3052 66210 3108 66220
rect 3836 66276 3892 66286
rect 3836 66182 3892 66220
rect 2716 65268 2772 65278
rect 2716 65174 2772 65212
rect 4476 65100 4740 65110
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4476 65034 4740 65044
rect 3836 64708 3892 64718
rect 3500 64706 3892 64708
rect 3500 64654 3838 64706
rect 3890 64654 3892 64706
rect 3500 64652 3892 64654
rect 2492 64148 2548 64158
rect 2380 64146 2884 64148
rect 2380 64094 2494 64146
rect 2546 64094 2884 64146
rect 2380 64092 2884 64094
rect 2492 64082 2548 64092
rect 2268 63870 2270 63922
rect 2322 63870 2324 63922
rect 1932 63250 1988 63262
rect 1932 63198 1934 63250
rect 1986 63198 1988 63250
rect 1932 62804 1988 63198
rect 1932 62738 1988 62748
rect 1932 62130 1988 62142
rect 1932 62078 1934 62130
rect 1986 62078 1988 62130
rect 1932 61684 1988 62078
rect 1932 61618 1988 61628
rect 2268 61684 2324 63870
rect 2828 64036 2884 64092
rect 3500 64146 3556 64652
rect 3836 64642 3892 64652
rect 3500 64094 3502 64146
rect 3554 64094 3556 64146
rect 3500 64082 3556 64094
rect 2828 62132 2884 63980
rect 3164 64034 3220 64046
rect 3164 63982 3166 64034
rect 3218 63982 3220 64034
rect 3164 63140 3220 63982
rect 3724 64036 3780 64046
rect 3724 63922 3780 63980
rect 3724 63870 3726 63922
rect 3778 63870 3780 63922
rect 3724 63858 3780 63870
rect 4476 63532 4740 63542
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4476 63466 4740 63476
rect 3836 63140 3892 63150
rect 3164 63138 3892 63140
rect 3164 63086 3838 63138
rect 3890 63086 3892 63138
rect 3164 63084 3892 63086
rect 3836 63074 3892 63084
rect 3836 62356 3892 62366
rect 2828 62066 2884 62076
rect 3388 62354 3892 62356
rect 3388 62302 3838 62354
rect 3890 62302 3892 62354
rect 3388 62300 3892 62302
rect 2268 61628 3108 61684
rect 2268 61570 2324 61628
rect 2268 61518 2270 61570
rect 2322 61518 2324 61570
rect 2268 61506 2324 61518
rect 2716 61460 2772 61470
rect 2716 61458 2884 61460
rect 2716 61406 2718 61458
rect 2770 61406 2884 61458
rect 2716 61404 2884 61406
rect 2716 61394 2772 61404
rect 2044 61346 2100 61358
rect 2044 61294 2046 61346
rect 2098 61294 2100 61346
rect 2044 60786 2100 61294
rect 2828 61348 2884 61404
rect 3052 61458 3108 61628
rect 3052 61406 3054 61458
rect 3106 61406 3108 61458
rect 3052 61394 3108 61406
rect 3388 61458 3444 62300
rect 3836 62290 3892 62300
rect 3612 62132 3668 62142
rect 3612 61570 3668 62076
rect 4476 61964 4740 61974
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4476 61898 4740 61908
rect 3612 61518 3614 61570
rect 3666 61518 3668 61570
rect 3612 61506 3668 61518
rect 3388 61406 3390 61458
rect 3442 61406 3444 61458
rect 3388 61394 3444 61406
rect 2828 61282 2884 61292
rect 4172 61348 4228 61358
rect 4284 61348 4340 61358
rect 4228 61346 4340 61348
rect 4228 61294 4286 61346
rect 4338 61294 4340 61346
rect 4228 61292 4340 61294
rect 2044 60734 2046 60786
rect 2098 60734 2100 60786
rect 2044 60722 2100 60734
rect 2716 60564 2772 60574
rect 2716 60470 2772 60508
rect 1932 60114 1988 60126
rect 1932 60062 1934 60114
rect 1986 60062 1988 60114
rect 1932 59444 1988 60062
rect 1932 59378 1988 59388
rect 2716 60004 2772 60014
rect 2716 59442 2772 59948
rect 3836 60004 3892 60014
rect 3836 59910 3892 59948
rect 2716 59390 2718 59442
rect 2770 59390 2772 59442
rect 2716 59378 2772 59390
rect 2044 59330 2100 59342
rect 2044 59278 2046 59330
rect 2098 59278 2100 59330
rect 2044 58434 2100 59278
rect 2044 58382 2046 58434
rect 2098 58382 2100 58434
rect 2044 58370 2100 58382
rect 2156 59220 2212 59230
rect 1932 57428 1988 57438
rect 1932 57334 1988 57372
rect 1932 56978 1988 56990
rect 1932 56926 1934 56978
rect 1986 56926 1988 56978
rect 1932 56084 1988 56926
rect 1932 56018 1988 56028
rect 2044 56194 2100 56206
rect 2044 56142 2046 56194
rect 2098 56142 2100 56194
rect 2044 55298 2100 56142
rect 2044 55246 2046 55298
rect 2098 55246 2100 55298
rect 2044 55234 2100 55246
rect 1932 54290 1988 54302
rect 1932 54238 1934 54290
rect 1986 54238 1988 54290
rect 1932 53844 1988 54238
rect 1932 53778 1988 53788
rect 2156 53732 2212 59164
rect 2380 59218 2436 59230
rect 2380 59166 2382 59218
rect 2434 59166 2436 59218
rect 2380 56308 2436 59166
rect 2940 59220 2996 59230
rect 2940 59126 2996 59164
rect 3500 59220 3556 59230
rect 3500 59126 3556 59164
rect 2716 58212 2772 58222
rect 2716 58118 2772 58156
rect 3836 56868 3892 56878
rect 3724 56866 3892 56868
rect 3724 56814 3838 56866
rect 3890 56814 3892 56866
rect 3724 56812 3892 56814
rect 2716 56308 2772 56318
rect 2380 56306 2772 56308
rect 2380 56254 2718 56306
rect 2770 56254 2772 56306
rect 2380 56252 2772 56254
rect 2380 56194 2436 56252
rect 2380 56142 2382 56194
rect 2434 56142 2436 56194
rect 2380 56130 2436 56142
rect 2716 56196 2772 56252
rect 3724 56306 3780 56812
rect 3836 56802 3892 56812
rect 3724 56254 3726 56306
rect 3778 56254 3780 56306
rect 3724 56242 3780 56254
rect 2716 56130 2772 56140
rect 3388 56196 3444 56206
rect 3388 56102 3444 56140
rect 2940 56082 2996 56094
rect 2940 56030 2942 56082
rect 2994 56030 2996 56082
rect 2716 55076 2772 55086
rect 2716 54982 2772 55020
rect 2268 53732 2324 53742
rect 2044 53730 2436 53732
rect 2044 53678 2270 53730
rect 2322 53678 2436 53730
rect 2044 53676 2436 53678
rect 1932 53620 1988 53630
rect 2044 53620 2100 53676
rect 2268 53666 2324 53676
rect 1932 53618 2100 53620
rect 1932 53566 1934 53618
rect 1986 53566 2100 53618
rect 1932 53564 2100 53566
rect 1932 53554 1988 53564
rect 1932 52724 1988 52734
rect 1932 52630 1988 52668
rect 1932 52274 1988 52286
rect 1932 52222 1934 52274
rect 1986 52222 1988 52274
rect 1932 51604 1988 52222
rect 1932 51538 1988 51548
rect 2268 51378 2324 51390
rect 2268 51326 2270 51378
rect 2322 51326 2324 51378
rect 1932 50708 1988 50718
rect 1932 50614 1988 50652
rect 1932 49588 1988 49598
rect 1932 49494 1988 49532
rect 1932 49138 1988 49150
rect 1932 49086 1934 49138
rect 1986 49086 1988 49138
rect 1932 48244 1988 49086
rect 1932 48178 1988 48188
rect 2044 48354 2100 48366
rect 2044 48302 2046 48354
rect 2098 48302 2100 48354
rect 2044 47458 2100 48302
rect 2044 47406 2046 47458
rect 2098 47406 2100 47458
rect 2044 47394 2100 47406
rect 1932 46450 1988 46462
rect 1932 46398 1934 46450
rect 1986 46398 1988 46450
rect 1932 46004 1988 46398
rect 1932 45938 1988 45948
rect 2044 45666 2100 45678
rect 2044 45614 2046 45666
rect 2098 45614 2100 45666
rect 2044 45106 2100 45614
rect 2044 45054 2046 45106
rect 2098 45054 2100 45106
rect 2044 45042 2100 45054
rect 1708 43652 1876 43708
rect 2044 44322 2100 44334
rect 2044 44270 2046 44322
rect 2098 44270 2100 44322
rect 2044 43762 2100 44270
rect 2044 43710 2046 43762
rect 2098 43710 2100 43762
rect 2044 43698 2100 43710
rect 2268 43652 2324 51326
rect 2380 51380 2436 53676
rect 2940 53730 2996 56030
rect 3836 54516 3892 54526
rect 2940 53678 2942 53730
rect 2994 53678 2996 53730
rect 2492 53508 2548 53518
rect 2492 53414 2548 53452
rect 2940 53508 2996 53678
rect 3500 54514 3892 54516
rect 3500 54462 3838 54514
rect 3890 54462 3892 54514
rect 3500 54460 3892 54462
rect 3164 53620 3220 53630
rect 3164 53526 3220 53564
rect 3500 53618 3556 54460
rect 3836 54450 3892 54460
rect 3500 53566 3502 53618
rect 3554 53566 3556 53618
rect 3500 53554 3556 53566
rect 3836 53618 3892 53630
rect 3836 53566 3838 53618
rect 3890 53566 3892 53618
rect 2940 53442 2996 53452
rect 3836 53508 3892 53566
rect 3836 52724 3892 53452
rect 3948 53620 4004 53630
rect 3948 52946 4004 53564
rect 3948 52894 3950 52946
rect 4002 52894 4004 52946
rect 3948 52882 4004 52894
rect 3836 52668 4004 52724
rect 3836 52164 3892 52174
rect 3500 52162 3892 52164
rect 3500 52110 3838 52162
rect 3890 52110 3892 52162
rect 3500 52108 3892 52110
rect 2492 51660 2996 51716
rect 2492 51602 2548 51660
rect 2492 51550 2494 51602
rect 2546 51550 2548 51602
rect 2492 51538 2548 51550
rect 2828 51490 2884 51502
rect 2828 51438 2830 51490
rect 2882 51438 2884 51490
rect 2380 51324 2548 51380
rect 2380 48244 2436 48254
rect 2380 45890 2436 48188
rect 2380 45838 2382 45890
rect 2434 45838 2436 45890
rect 2380 45780 2436 45838
rect 2380 45714 2436 45724
rect 2492 43708 2548 51324
rect 2828 50596 2884 51438
rect 2940 51380 2996 51660
rect 3500 51602 3556 52108
rect 3836 52098 3892 52108
rect 3500 51550 3502 51602
rect 3554 51550 3556 51602
rect 3500 51538 3556 51550
rect 3836 51492 3892 51502
rect 3948 51492 4004 52668
rect 3836 51490 4004 51492
rect 3836 51438 3838 51490
rect 3890 51438 4004 51490
rect 3836 51436 4004 51438
rect 3836 51426 3892 51436
rect 3164 51380 3220 51390
rect 2940 51378 3220 51380
rect 2940 51326 3166 51378
rect 3218 51326 3220 51378
rect 2940 51324 3220 51326
rect 2828 50530 2884 50540
rect 3164 49588 3220 51324
rect 3836 50596 3892 50606
rect 3836 50502 3892 50540
rect 3836 49812 3892 49822
rect 3164 49522 3220 49532
rect 3388 49810 3892 49812
rect 3388 49758 3838 49810
rect 3890 49758 3892 49810
rect 3388 49756 3892 49758
rect 2716 49028 2772 49038
rect 2716 48466 2772 48972
rect 2716 48414 2718 48466
rect 2770 48414 2772 48466
rect 2716 48402 2772 48414
rect 3388 48466 3444 49756
rect 3836 49746 3892 49756
rect 3388 48414 3390 48466
rect 3442 48414 3444 48466
rect 3388 48402 3444 48414
rect 3612 49588 3668 49598
rect 2940 48244 2996 48254
rect 2940 48150 2996 48188
rect 3612 48242 3668 49532
rect 3836 49028 3892 49038
rect 3836 48934 3892 48972
rect 3612 48190 3614 48242
rect 3666 48190 3668 48242
rect 3612 48178 3668 48190
rect 2716 47236 2772 47246
rect 2716 47142 2772 47180
rect 3836 46676 3892 46686
rect 3388 46674 3892 46676
rect 3388 46622 3838 46674
rect 3890 46622 3892 46674
rect 3388 46620 3892 46622
rect 2716 45892 2772 45902
rect 2716 45798 2772 45836
rect 3276 45892 3332 45902
rect 3052 45780 3108 45790
rect 3052 45686 3108 45724
rect 2716 44884 2772 44894
rect 2716 44790 2772 44828
rect 2716 44100 2772 44110
rect 2716 44006 2772 44044
rect 2492 43652 2660 43708
rect 1708 41972 1764 43652
rect 2156 43596 2324 43652
rect 1932 42868 1988 42878
rect 1932 42774 1988 42812
rect 1708 40402 1764 41916
rect 1932 41748 1988 41758
rect 1932 41654 1988 41692
rect 1708 40350 1710 40402
rect 1762 40350 1764 40402
rect 1708 40338 1764 40350
rect 1932 41298 1988 41310
rect 1932 41246 1934 41298
rect 1986 41246 1988 41298
rect 1932 40404 1988 41246
rect 1932 40338 1988 40348
rect 1932 39730 1988 39742
rect 1932 39678 1934 39730
rect 1986 39678 1988 39730
rect 1932 39284 1988 39678
rect 1932 39218 1988 39228
rect 2044 38836 2100 38846
rect 2156 38836 2212 43596
rect 2268 43540 2324 43596
rect 2268 43446 2324 43484
rect 2268 40628 2324 40638
rect 2268 40534 2324 40572
rect 2604 40402 2660 43652
rect 2716 43650 2772 43662
rect 2716 43598 2718 43650
rect 2770 43598 2772 43650
rect 2716 42756 2772 43598
rect 2828 43540 2884 43550
rect 3052 43540 3108 43550
rect 2884 43538 3108 43540
rect 2884 43486 3054 43538
rect 3106 43486 3108 43538
rect 2884 43484 3108 43486
rect 2828 43474 2884 43484
rect 3052 43474 3108 43484
rect 2716 42690 2772 42700
rect 2604 40350 2606 40402
rect 2658 40350 2660 40402
rect 2604 39620 2660 40350
rect 3164 40404 3220 40414
rect 3164 40310 3220 40348
rect 2604 39554 2660 39564
rect 2044 38834 2212 38836
rect 2044 38782 2046 38834
rect 2098 38782 2212 38834
rect 2044 38780 2212 38782
rect 2940 39060 2996 39070
rect 2044 38162 2100 38780
rect 2940 38164 2996 39004
rect 3276 39060 3332 45836
rect 3388 45778 3444 46620
rect 3836 46610 3892 46620
rect 3388 45726 3390 45778
rect 3442 45726 3444 45778
rect 3388 45714 3444 45726
rect 3612 45890 3668 45902
rect 3612 45838 3614 45890
rect 3666 45838 3668 45890
rect 3612 45780 3668 45838
rect 3612 45714 3668 45724
rect 3836 42756 3892 42766
rect 3836 42662 3892 42700
rect 3836 41972 3892 41982
rect 3836 41878 3892 41916
rect 4172 41300 4228 61292
rect 4284 61282 4340 61292
rect 4476 60396 4740 60406
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4476 60330 4740 60340
rect 4476 58828 4740 58838
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4476 58762 4740 58772
rect 4284 57650 4340 57662
rect 4284 57598 4286 57650
rect 4338 57598 4340 57650
rect 4284 56756 4340 57598
rect 4476 57260 4740 57270
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4476 57194 4740 57204
rect 4844 56866 4900 56878
rect 4844 56814 4846 56866
rect 4898 56814 4900 56866
rect 4620 56756 4676 56766
rect 4284 56754 4676 56756
rect 4284 56702 4622 56754
rect 4674 56702 4676 56754
rect 4284 56700 4676 56702
rect 4620 56690 4676 56700
rect 4844 56196 4900 56814
rect 4844 56130 4900 56140
rect 4476 55692 4740 55702
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4476 55626 4740 55636
rect 4476 54124 4740 54134
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4476 54058 4740 54068
rect 4476 52556 4740 52566
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4476 52490 4740 52500
rect 4476 50988 4740 50998
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4476 50922 4740 50932
rect 4476 49420 4740 49430
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4476 49354 4740 49364
rect 4476 47852 4740 47862
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4476 47786 4740 47796
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 4284 45892 4340 45902
rect 4284 45798 4340 45836
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 4732 41972 4788 41982
rect 4732 41878 4788 41916
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 4732 41300 4788 41310
rect 4172 41298 4788 41300
rect 4172 41246 4734 41298
rect 4786 41246 4788 41298
rect 4172 41244 4788 41246
rect 4172 41188 4228 41244
rect 4732 41234 4788 41244
rect 3500 41186 4228 41188
rect 3500 41134 4174 41186
rect 4226 41134 4228 41186
rect 3500 41132 4228 41134
rect 3500 40402 3556 41132
rect 4172 41122 4228 41132
rect 5404 40628 5460 40638
rect 5404 40534 5460 40572
rect 4060 40516 4116 40526
rect 4060 40422 4116 40460
rect 4508 40516 4564 40526
rect 4508 40422 4564 40460
rect 5180 40516 5236 40526
rect 3500 40350 3502 40402
rect 3554 40350 3556 40402
rect 3500 40338 3556 40350
rect 4956 40404 5012 40414
rect 4956 40310 5012 40348
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 3836 39620 3892 39630
rect 3836 39526 3892 39564
rect 4732 39620 4788 39630
rect 4732 39526 4788 39564
rect 5180 39396 5236 40460
rect 5180 39330 5236 39340
rect 3276 38994 3332 39004
rect 2044 38110 2046 38162
rect 2098 38110 2100 38162
rect 2044 38098 2100 38110
rect 2492 38162 2996 38164
rect 2492 38110 2942 38162
rect 2994 38110 2996 38162
rect 2492 38108 2996 38110
rect 2492 38050 2548 38108
rect 2940 38098 2996 38108
rect 3388 38722 3444 38734
rect 3388 38670 3390 38722
rect 3442 38670 3444 38722
rect 3388 38164 3444 38670
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 3388 38098 3444 38108
rect 2492 37998 2494 38050
rect 2546 37998 2548 38050
rect 2492 37986 2548 37998
rect 2044 37380 2100 37390
rect 2044 37286 2100 37324
rect 1708 37266 1764 37278
rect 1708 37214 1710 37266
rect 1762 37214 1764 37266
rect 1708 37044 1764 37214
rect 1708 36978 1764 36988
rect 2492 37154 2548 37166
rect 2492 37102 2494 37154
rect 2546 37102 2548 37154
rect 2492 37044 2548 37102
rect 2492 36978 2548 36988
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 1708 36370 1764 36382
rect 1708 36318 1710 36370
rect 1762 36318 1764 36370
rect 1708 35924 1764 36318
rect 2044 36260 2100 36270
rect 2044 36166 2100 36204
rect 2492 36258 2548 36270
rect 2492 36206 2494 36258
rect 2546 36206 2548 36258
rect 1708 35858 1764 35868
rect 2492 35924 2548 36206
rect 2492 35858 2548 35868
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 1708 34804 1764 34814
rect 1708 34710 1764 34748
rect 2492 34804 2548 34814
rect 2492 34710 2548 34748
rect 2044 34692 2100 34702
rect 2044 34598 2100 34636
rect 2044 34244 2100 34254
rect 2044 34150 2100 34188
rect 1708 34130 1764 34142
rect 1708 34078 1710 34130
rect 1762 34078 1764 34130
rect 1708 33684 1764 34078
rect 1708 33618 1764 33628
rect 2492 34018 2548 34030
rect 2492 33966 2494 34018
rect 2546 33966 2548 34018
rect 2492 33684 2548 33966
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 2492 33618 2548 33628
rect 1708 33122 1764 33134
rect 1708 33070 1710 33122
rect 1762 33070 1764 33122
rect 1708 32564 1764 33070
rect 2044 33124 2100 33134
rect 2044 33030 2100 33068
rect 2492 33122 2548 33134
rect 2492 33070 2494 33122
rect 2546 33070 2548 33122
rect 1708 32498 1764 32508
rect 2492 32564 2548 33070
rect 2492 32498 2548 32508
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 2044 31780 2100 31790
rect 1708 31666 1764 31678
rect 1708 31614 1710 31666
rect 1762 31614 1764 31666
rect 1708 31444 1764 31614
rect 2044 31666 2100 31724
rect 2044 31614 2046 31666
rect 2098 31614 2100 31666
rect 2044 31602 2100 31614
rect 1708 31378 1764 31388
rect 2492 31554 2548 31566
rect 2492 31502 2494 31554
rect 2546 31502 2548 31554
rect 2492 31444 2548 31502
rect 2492 31378 2548 31388
rect 2044 31108 2100 31118
rect 2044 31014 2100 31052
rect 1708 30994 1764 31006
rect 1708 30942 1710 30994
rect 1762 30942 1764 30994
rect 1708 30884 1764 30942
rect 1708 30324 1764 30828
rect 2492 30884 2548 30894
rect 2492 30790 2548 30828
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 1708 30258 1764 30268
rect 2044 29540 2100 29550
rect 2044 29446 2100 29484
rect 1708 29426 1764 29438
rect 1708 29374 1710 29426
rect 1762 29374 1764 29426
rect 1708 29204 1764 29374
rect 1708 29138 1764 29148
rect 2492 29314 2548 29326
rect 2492 29262 2494 29314
rect 2546 29262 2548 29314
rect 2492 29204 2548 29262
rect 2492 29138 2548 29148
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 2044 28756 2100 28766
rect 1708 28642 1764 28654
rect 1708 28590 1710 28642
rect 1762 28590 1764 28642
rect 1708 28084 1764 28590
rect 2044 28530 2100 28700
rect 2044 28478 2046 28530
rect 2098 28478 2100 28530
rect 2044 28466 2100 28478
rect 2492 28642 2548 28654
rect 2492 28590 2494 28642
rect 2546 28590 2548 28642
rect 1708 28018 1764 28028
rect 2492 28084 2548 28590
rect 2492 28018 2548 28028
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 2044 27300 2100 27310
rect 1708 26964 1764 26974
rect 1708 26870 1764 26908
rect 2044 26962 2100 27244
rect 2044 26910 2046 26962
rect 2098 26910 2100 26962
rect 2044 26898 2100 26910
rect 2492 26964 2548 26974
rect 2492 26870 2548 26908
rect 2044 26402 2100 26414
rect 2044 26350 2046 26402
rect 2098 26350 2100 26402
rect 1708 26290 1764 26302
rect 1708 26238 1710 26290
rect 1762 26238 1764 26290
rect 1708 25844 1764 26238
rect 2044 26068 2100 26350
rect 2044 26002 2100 26012
rect 2492 26178 2548 26190
rect 2492 26126 2494 26178
rect 2546 26126 2548 26178
rect 1708 25778 1764 25788
rect 2492 25844 2548 26126
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 2492 25778 2548 25788
rect 2044 25620 2100 25630
rect 2044 25394 2100 25564
rect 2044 25342 2046 25394
rect 2098 25342 2100 25394
rect 2044 25330 2100 25342
rect 1708 25282 1764 25294
rect 1708 25230 1710 25282
rect 1762 25230 1764 25282
rect 1708 24724 1764 25230
rect 1708 24658 1764 24668
rect 2492 25282 2548 25294
rect 2492 25230 2494 25282
rect 2546 25230 2548 25282
rect 2492 24724 2548 25230
rect 2492 24658 2548 24668
rect 8316 24388 8372 76300
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 8316 24322 8372 24332
rect 9996 74900 10052 74910
rect 4476 24266 4740 24276
rect 2044 23940 2100 23950
rect 2044 23826 2100 23884
rect 2044 23774 2046 23826
rect 2098 23774 2100 23826
rect 2044 23762 2100 23774
rect 1708 23714 1764 23726
rect 1708 23662 1710 23714
rect 1762 23662 1764 23714
rect 1708 23604 1764 23662
rect 1708 23538 1764 23548
rect 2492 23714 2548 23726
rect 2492 23662 2494 23714
rect 2546 23662 2548 23714
rect 2492 23604 2548 23662
rect 2492 23538 2548 23548
rect 2044 23266 2100 23278
rect 2044 23214 2046 23266
rect 2098 23214 2100 23266
rect 1708 23154 1764 23166
rect 1708 23102 1710 23154
rect 1762 23102 1764 23154
rect 1708 23044 1764 23102
rect 1708 22484 1764 22988
rect 2044 22596 2100 23214
rect 2492 23044 2548 23054
rect 2492 22950 2548 22988
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 2044 22530 2100 22540
rect 1708 22418 1764 22428
rect 9996 21812 10052 74844
rect 11228 74226 11284 79200
rect 11900 77924 11956 79200
rect 11900 77868 12068 77924
rect 11564 76242 11620 76254
rect 11564 76190 11566 76242
rect 11618 76190 11620 76242
rect 11564 75572 11620 76190
rect 11900 75908 11956 75918
rect 11900 75814 11956 75852
rect 11564 75506 11620 75516
rect 11228 74174 11230 74226
rect 11282 74174 11284 74226
rect 11228 74162 11284 74174
rect 11676 74788 11732 74798
rect 9996 21746 10052 21756
rect 11452 22932 11508 22942
rect 2044 21700 2100 21710
rect 2044 21606 2100 21644
rect 1708 21586 1764 21598
rect 1708 21534 1710 21586
rect 1762 21534 1764 21586
rect 1708 21364 1764 21534
rect 1708 21298 1764 21308
rect 2492 21474 2548 21486
rect 2492 21422 2494 21474
rect 2546 21422 2548 21474
rect 2492 21364 2548 21422
rect 2492 21298 2548 21308
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 2044 20916 2100 20926
rect 2044 20690 2100 20860
rect 2044 20638 2046 20690
rect 2098 20638 2100 20690
rect 2044 20626 2100 20638
rect 1708 20578 1764 20590
rect 1708 20526 1710 20578
rect 1762 20526 1764 20578
rect 1708 20244 1764 20526
rect 2492 20578 2548 20590
rect 2492 20526 2494 20578
rect 2546 20526 2548 20578
rect 1708 20178 1764 20188
rect 2044 20356 2100 20366
rect 1708 19124 1764 19134
rect 1708 19030 1764 19068
rect 2044 19122 2100 20300
rect 2492 20244 2548 20526
rect 11452 20188 11508 22876
rect 2492 20178 2548 20188
rect 11228 20132 11508 20188
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 7532 19348 7588 19358
rect 2044 19070 2046 19122
rect 2098 19070 2100 19122
rect 2044 19058 2100 19070
rect 2492 19124 2548 19134
rect 2492 19030 2548 19068
rect 6300 18676 6356 18686
rect 2044 18562 2100 18574
rect 2044 18510 2046 18562
rect 2098 18510 2100 18562
rect 1708 18450 1764 18462
rect 1708 18398 1710 18450
rect 1762 18398 1764 18450
rect 1708 18004 1764 18398
rect 2044 18340 2100 18510
rect 2044 18274 2100 18284
rect 2492 18338 2548 18350
rect 2492 18286 2494 18338
rect 2546 18286 2548 18338
rect 1708 17938 1764 17948
rect 2492 18004 2548 18286
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 2492 17938 2548 17948
rect 2044 17892 2100 17902
rect 1708 17554 1764 17566
rect 1708 17502 1710 17554
rect 1762 17502 1764 17554
rect 1708 17444 1764 17502
rect 2044 17554 2100 17836
rect 2044 17502 2046 17554
rect 2098 17502 2100 17554
rect 2044 17490 2100 17502
rect 1708 16884 1764 17388
rect 2492 17444 2548 17454
rect 2492 17350 2548 17388
rect 1708 16818 1764 16828
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 2044 16324 2100 16334
rect 1708 15986 1764 15998
rect 1708 15934 1710 15986
rect 1762 15934 1764 15986
rect 1708 15764 1764 15934
rect 2044 15986 2100 16268
rect 2044 15934 2046 15986
rect 2098 15934 2100 15986
rect 2044 15922 2100 15934
rect 2156 16100 2212 16110
rect 1708 15698 1764 15708
rect 2044 15428 2100 15438
rect 2044 15334 2100 15372
rect 1708 15314 1764 15326
rect 1708 15262 1710 15314
rect 1762 15262 1764 15314
rect 1708 14644 1764 15262
rect 1708 14578 1764 14588
rect 1596 14420 1652 14430
rect 1596 5012 1652 14364
rect 2044 13972 2100 13982
rect 2044 13878 2100 13916
rect 1708 13746 1764 13758
rect 1708 13694 1710 13746
rect 1762 13694 1764 13746
rect 1708 13524 1764 13694
rect 1708 13458 1764 13468
rect 1932 13076 1988 13086
rect 1708 12850 1764 12862
rect 1708 12798 1710 12850
rect 1762 12798 1764 12850
rect 1708 12404 1764 12798
rect 1708 12338 1764 12348
rect 1708 11284 1764 11294
rect 1708 11190 1764 11228
rect 1708 10610 1764 10622
rect 1708 10558 1710 10610
rect 1762 10558 1764 10610
rect 1708 10164 1764 10558
rect 1708 10098 1764 10108
rect 1708 9714 1764 9726
rect 1708 9662 1710 9714
rect 1762 9662 1764 9714
rect 1708 9604 1764 9662
rect 1708 9044 1764 9548
rect 1708 8978 1764 8988
rect 1708 8146 1764 8158
rect 1708 8094 1710 8146
rect 1762 8094 1764 8146
rect 1708 7924 1764 8094
rect 1708 7858 1764 7868
rect 1708 7474 1764 7486
rect 1708 7422 1710 7474
rect 1762 7422 1764 7474
rect 1708 7364 1764 7422
rect 1708 6804 1764 7308
rect 1708 6738 1764 6748
rect 1932 6132 1988 13020
rect 2044 12852 2100 12862
rect 2044 12758 2100 12796
rect 2044 11284 2100 11294
rect 2044 11190 2100 11228
rect 2044 10724 2100 10734
rect 2044 10630 2100 10668
rect 2156 10500 2212 16044
rect 2492 15874 2548 15886
rect 2492 15822 2494 15874
rect 2546 15822 2548 15874
rect 2492 15764 2548 15822
rect 2492 15698 2548 15708
rect 2492 15202 2548 15214
rect 2492 15150 2494 15202
rect 2546 15150 2548 15202
rect 2492 14644 2548 15150
rect 5852 15204 5908 15214
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 2492 14578 2548 14588
rect 2492 13634 2548 13646
rect 2492 13582 2494 13634
rect 2546 13582 2548 13634
rect 2492 13524 2548 13582
rect 2492 13458 2548 13468
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 2492 12738 2548 12750
rect 2492 12686 2494 12738
rect 2546 12686 2548 12738
rect 2492 12404 2548 12686
rect 2492 12338 2548 12348
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 2492 11172 2548 11182
rect 2492 11078 2548 11116
rect 2044 10444 2212 10500
rect 2492 10498 2548 10510
rect 2492 10446 2494 10498
rect 2546 10446 2548 10498
rect 2044 9714 2100 10444
rect 2044 9662 2046 9714
rect 2098 9662 2100 9714
rect 2044 9650 2100 9662
rect 2380 10388 2436 10398
rect 2380 8428 2436 10332
rect 2492 10164 2548 10446
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 2492 10098 2548 10108
rect 2492 9604 2548 9614
rect 2492 9510 2548 9548
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 2044 8372 2436 8428
rect 2044 8146 2100 8372
rect 2044 8094 2046 8146
rect 2098 8094 2100 8146
rect 2044 8082 2100 8094
rect 2492 8034 2548 8046
rect 2492 7982 2494 8034
rect 2546 7982 2548 8034
rect 2492 7924 2548 7982
rect 2492 7858 2548 7868
rect 2044 7700 2100 7710
rect 2044 7606 2100 7644
rect 5852 7700 5908 15148
rect 5852 7634 5908 7644
rect 2492 7364 2548 7374
rect 2492 7270 2548 7308
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 6076 7028 6132 7038
rect 4476 7018 4740 7028
rect 5964 6972 6076 7028
rect 2156 6804 2212 6814
rect 2044 6132 2100 6142
rect 1932 6130 2100 6132
rect 1932 6078 2046 6130
rect 2098 6078 2100 6130
rect 1932 6076 2100 6078
rect 2044 6066 2100 6076
rect 1708 5906 1764 5918
rect 2156 5908 2212 6748
rect 4284 6580 4340 6590
rect 3612 6132 3668 6142
rect 2380 6020 2436 6030
rect 1708 5854 1710 5906
rect 1762 5854 1764 5906
rect 1708 5684 1764 5854
rect 1708 5618 1764 5628
rect 2044 5852 2212 5908
rect 2268 5964 2380 6020
rect 1596 4946 1652 4956
rect 1708 5122 1764 5134
rect 1708 5070 1710 5122
rect 1762 5070 1764 5122
rect 1708 4564 1764 5070
rect 2044 5010 2100 5852
rect 2044 4958 2046 5010
rect 2098 4958 2100 5010
rect 2044 4946 2100 4958
rect 2268 4788 2324 5964
rect 2380 5954 2436 5964
rect 2492 5794 2548 5806
rect 2492 5742 2494 5794
rect 2546 5742 2548 5794
rect 2492 5684 2548 5742
rect 2492 5618 2548 5628
rect 1708 4498 1764 4508
rect 2044 4732 2324 4788
rect 2492 5122 2548 5134
rect 2492 5070 2494 5122
rect 2546 5070 2548 5122
rect 1820 4228 1876 4238
rect 1820 3556 1876 4172
rect 1820 3462 1876 3500
rect 2044 3442 2100 4732
rect 2492 4564 2548 5070
rect 2492 4498 2548 4508
rect 2716 5012 2772 5022
rect 2044 3390 2046 3442
rect 2098 3390 2100 3442
rect 2044 3378 2100 3390
rect 2156 4226 2212 4238
rect 2156 4174 2158 4226
rect 2210 4174 2212 4226
rect 2156 3444 2212 4174
rect 2492 4228 2548 4238
rect 2492 4134 2548 4172
rect 2380 3444 2436 3454
rect 2156 3442 2436 3444
rect 2156 3390 2382 3442
rect 2434 3390 2436 3442
rect 2156 3388 2436 3390
rect 2380 2324 2436 3388
rect 2716 3442 2772 4956
rect 3276 4228 3332 4238
rect 3276 4226 3444 4228
rect 3276 4174 3278 4226
rect 3330 4174 3444 4226
rect 3276 4172 3444 4174
rect 3276 4162 3332 4172
rect 3388 3556 3444 4172
rect 3388 3462 3444 3500
rect 2716 3390 2718 3442
rect 2770 3390 2772 3442
rect 2716 3378 2772 3390
rect 3612 3442 3668 6076
rect 4284 5124 4340 6524
rect 4956 6468 5012 6478
rect 4844 5572 4900 5582
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 4284 5068 4452 5124
rect 4284 4900 4340 4910
rect 4172 4898 4340 4900
rect 4172 4846 4286 4898
rect 4338 4846 4340 4898
rect 4172 4844 4340 4846
rect 4060 4338 4116 4350
rect 4060 4286 4062 4338
rect 4114 4286 4116 4338
rect 3724 4228 3780 4238
rect 4060 4228 4116 4286
rect 3724 4226 4116 4228
rect 3724 4174 3726 4226
rect 3778 4174 4116 4226
rect 3724 4172 4116 4174
rect 3724 4162 3780 4172
rect 3612 3390 3614 3442
rect 3666 3390 3668 3442
rect 3612 3378 3668 3390
rect 3948 3444 4004 3482
rect 3948 3378 4004 3388
rect 2380 2258 2436 2268
rect 4060 756 4116 4172
rect 4172 3444 4228 4844
rect 4284 4834 4340 4844
rect 4284 4564 4340 4574
rect 4396 4564 4452 5068
rect 4284 4562 4452 4564
rect 4284 4510 4286 4562
rect 4338 4510 4452 4562
rect 4284 4508 4452 4510
rect 4732 4898 4788 4910
rect 4732 4846 4734 4898
rect 4786 4846 4788 4898
rect 4284 4498 4340 4508
rect 4508 4340 4564 4350
rect 4396 4284 4508 4340
rect 4396 4116 4452 4284
rect 4508 4274 4564 4284
rect 4620 4340 4676 4350
rect 4732 4340 4788 4846
rect 4620 4338 4788 4340
rect 4620 4286 4622 4338
rect 4674 4286 4788 4338
rect 4620 4284 4788 4286
rect 4620 4228 4676 4284
rect 4620 4162 4676 4172
rect 4172 3378 4228 3388
rect 4284 4060 4452 4116
rect 4284 3442 4340 4060
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 4732 3780 4788 3790
rect 4732 3554 4788 3724
rect 4732 3502 4734 3554
rect 4786 3502 4788 3554
rect 4732 3490 4788 3502
rect 4284 3390 4286 3442
rect 4338 3390 4340 3442
rect 4284 3378 4340 3390
rect 4844 3444 4900 5516
rect 4956 4562 5012 6412
rect 5628 5908 5684 5918
rect 5292 5796 5348 5806
rect 4956 4510 4958 4562
rect 5010 4510 5012 4562
rect 4956 4498 5012 4510
rect 5068 5794 5348 5796
rect 5068 5742 5294 5794
rect 5346 5742 5348 5794
rect 5068 5740 5348 5742
rect 5068 3780 5124 5740
rect 5292 5730 5348 5740
rect 5180 4898 5236 4910
rect 5180 4846 5182 4898
rect 5234 4846 5236 4898
rect 5180 4340 5236 4846
rect 5628 4562 5684 5852
rect 5628 4510 5630 4562
rect 5682 4510 5684 4562
rect 5628 4498 5684 4510
rect 5740 5794 5796 5806
rect 5740 5742 5742 5794
rect 5794 5742 5796 5794
rect 5404 4340 5460 4350
rect 5180 4338 5460 4340
rect 5180 4286 5406 4338
rect 5458 4286 5460 4338
rect 5180 4284 5460 4286
rect 5404 3892 5460 4284
rect 5404 3826 5460 3836
rect 5068 3714 5124 3724
rect 5740 3668 5796 5742
rect 5852 3668 5908 3678
rect 5740 3612 5852 3668
rect 5628 3556 5684 3566
rect 4956 3444 5012 3454
rect 4844 3442 5012 3444
rect 4844 3390 4958 3442
rect 5010 3390 5012 3442
rect 4844 3388 5012 3390
rect 4956 3378 5012 3388
rect 4620 924 5012 980
rect 4620 756 4676 924
rect 4956 800 5012 924
rect 5628 800 5684 3500
rect 5852 3554 5908 3612
rect 5852 3502 5854 3554
rect 5906 3502 5908 3554
rect 5852 3490 5908 3502
rect 5964 3444 6020 6972
rect 6076 6962 6132 6972
rect 6300 6020 6356 18620
rect 7532 6804 7588 19292
rect 9996 15316 10052 15326
rect 8316 14644 8372 14654
rect 8316 12852 8372 14588
rect 8316 12786 8372 12796
rect 8316 12404 8372 12414
rect 8316 11284 8372 12348
rect 9660 12178 9716 12190
rect 9660 12126 9662 12178
rect 9714 12126 9716 12178
rect 9436 12068 9492 12078
rect 9436 11506 9492 12012
rect 9436 11454 9438 11506
rect 9490 11454 9492 11506
rect 9436 11442 9492 11454
rect 9212 11396 9268 11406
rect 8316 11218 8372 11228
rect 8540 11394 9268 11396
rect 8540 11342 9214 11394
rect 9266 11342 9268 11394
rect 8540 11340 9268 11342
rect 8204 10500 8260 10510
rect 8204 10050 8260 10444
rect 8204 9998 8206 10050
rect 8258 9998 8260 10050
rect 8204 9986 8260 9998
rect 8428 9940 8484 9950
rect 8092 9716 8148 9726
rect 8092 9622 8148 9660
rect 7532 6738 7588 6748
rect 7980 9602 8036 9614
rect 7980 9550 7982 9602
rect 8034 9550 8036 9602
rect 7980 6802 8036 9550
rect 8428 7700 8484 9884
rect 8540 8820 8596 11340
rect 9212 11330 9268 11340
rect 9548 11284 9604 11294
rect 9548 11190 9604 11228
rect 9660 9940 9716 12126
rect 9996 10388 10052 15260
rect 10332 12068 10388 12078
rect 10332 11974 10388 12012
rect 11116 10836 11172 10846
rect 11116 10742 11172 10780
rect 9996 10322 10052 10332
rect 11228 10052 11284 20132
rect 11676 13076 11732 74732
rect 12012 73444 12068 77868
rect 12124 76466 12180 76478
rect 12124 76414 12126 76466
rect 12178 76414 12180 76466
rect 12124 76356 12180 76414
rect 12124 76290 12180 76300
rect 12572 75908 12628 79200
rect 13244 76132 13300 79200
rect 13356 76356 13412 76366
rect 13356 76262 13412 76300
rect 12572 75842 12628 75852
rect 12908 76076 13300 76132
rect 12684 75684 12740 75694
rect 12124 73444 12180 73454
rect 12012 73442 12180 73444
rect 12012 73390 12126 73442
rect 12178 73390 12180 73442
rect 12012 73388 12180 73390
rect 12124 73378 12180 73388
rect 12684 24052 12740 75628
rect 12908 75122 12964 76076
rect 13580 75684 13636 75694
rect 13580 75590 13636 75628
rect 13916 75572 13972 79200
rect 13916 75506 13972 75516
rect 12908 75070 12910 75122
rect 12962 75070 12964 75122
rect 12908 75058 12964 75070
rect 14252 75458 14308 75470
rect 14252 75406 14254 75458
rect 14306 75406 14308 75458
rect 13468 74900 13524 74910
rect 13468 74806 13524 74844
rect 14252 74900 14308 75406
rect 14252 74834 14308 74844
rect 12908 74114 12964 74126
rect 12908 74062 12910 74114
rect 12962 74062 12964 74114
rect 12908 74004 12964 74062
rect 14028 74116 14084 74126
rect 14028 74022 14084 74060
rect 12908 73938 12964 73948
rect 14364 74004 14420 74014
rect 13916 73330 13972 73342
rect 13916 73278 13918 73330
rect 13970 73278 13972 73330
rect 13916 72324 13972 73278
rect 14140 72324 14196 72334
rect 13916 72322 14196 72324
rect 13916 72270 14142 72322
rect 14194 72270 14196 72322
rect 13916 72268 14196 72270
rect 14140 55468 14196 72268
rect 12684 20188 12740 23996
rect 13468 55412 14196 55468
rect 13468 23492 13524 55412
rect 13468 23426 13524 23436
rect 14252 24388 14308 24398
rect 11676 13010 11732 13020
rect 12572 20132 12740 20188
rect 12908 22484 12964 22494
rect 12572 12402 12628 20132
rect 12908 15148 12964 22428
rect 12572 12350 12574 12402
rect 12626 12350 12628 12402
rect 11676 11508 11732 11518
rect 11676 11394 11732 11452
rect 12460 11508 12516 11518
rect 12572 11508 12628 12350
rect 12516 11452 12628 11508
rect 12796 15092 12964 15148
rect 14252 15148 14308 24332
rect 14364 22932 14420 73948
rect 14588 73218 14644 79200
rect 14588 73166 14590 73218
rect 14642 73166 14644 73218
rect 14588 73154 14644 73166
rect 14700 75458 14756 75470
rect 14700 75406 14702 75458
rect 14754 75406 14756 75458
rect 14700 74898 14756 75406
rect 15260 75122 15316 79200
rect 15372 76692 15428 76702
rect 15932 76692 15988 79200
rect 16604 76692 16660 79200
rect 17276 77252 17332 79200
rect 15932 76636 16100 76692
rect 15372 76598 15428 76636
rect 15260 75070 15262 75122
rect 15314 75070 15316 75122
rect 15260 75058 15316 75070
rect 14700 74846 14702 74898
rect 14754 74846 14756 74898
rect 14364 22866 14420 22876
rect 14700 22484 14756 74846
rect 16044 74226 16100 76636
rect 16604 76626 16660 76636
rect 17052 77196 17332 77252
rect 16380 76466 16436 76478
rect 16380 76414 16382 76466
rect 16434 76414 16436 76466
rect 16380 76356 16436 76414
rect 16380 76290 16436 76300
rect 16828 75908 16884 75918
rect 17052 75908 17108 77196
rect 16828 75906 17108 75908
rect 16828 75854 16830 75906
rect 16882 75854 17108 75906
rect 16828 75852 17108 75854
rect 17164 76356 17220 76366
rect 16828 75842 16884 75852
rect 16044 74174 16046 74226
rect 16098 74174 16100 74226
rect 16044 74162 16100 74174
rect 16380 74116 16436 74126
rect 16380 73330 16436 74060
rect 16380 73278 16382 73330
rect 16434 73278 16436 73330
rect 16380 24612 16436 73278
rect 17164 31948 17220 76300
rect 17836 75682 17892 75694
rect 17836 75630 17838 75682
rect 17890 75630 17892 75682
rect 17836 75012 17892 75630
rect 17948 75572 18004 79200
rect 18620 75794 18676 79200
rect 19180 76692 19236 76702
rect 19292 76692 19348 79200
rect 19964 77028 20020 79200
rect 19964 76972 20244 77028
rect 19836 76860 20100 76870
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 19836 76794 20100 76804
rect 20188 76692 20244 76972
rect 19180 76690 19348 76692
rect 19180 76638 19182 76690
rect 19234 76638 19348 76690
rect 19180 76636 19348 76638
rect 20076 76636 20244 76692
rect 19180 76626 19236 76636
rect 19740 76468 19796 76478
rect 18620 75742 18622 75794
rect 18674 75742 18676 75794
rect 18620 75730 18676 75742
rect 19404 76466 19796 76468
rect 19404 76414 19742 76466
rect 19794 76414 19796 76466
rect 19404 76412 19796 76414
rect 17948 75506 18004 75516
rect 19180 75572 19236 75582
rect 17836 74956 18116 75012
rect 17948 74786 18004 74798
rect 17948 74734 17950 74786
rect 18002 74734 18004 74786
rect 17948 74340 18004 74734
rect 18060 74788 18116 74956
rect 18284 74788 18340 74798
rect 18060 74786 18340 74788
rect 18060 74734 18286 74786
rect 18338 74734 18340 74786
rect 18060 74732 18340 74734
rect 17612 74284 18228 74340
rect 17612 31948 17668 74284
rect 17836 74114 17892 74126
rect 17836 74062 17838 74114
rect 17890 74062 17892 74114
rect 17836 73220 17892 74062
rect 18172 74114 18228 74284
rect 18172 74062 18174 74114
rect 18226 74062 18228 74114
rect 18172 74050 18228 74062
rect 18060 73220 18116 73230
rect 17836 73218 18116 73220
rect 17836 73166 18062 73218
rect 18114 73166 18116 73218
rect 17836 73164 18116 73166
rect 18060 43708 18116 73164
rect 18060 43652 18228 43708
rect 14700 22418 14756 22428
rect 14924 23492 14980 23502
rect 14924 23156 14980 23436
rect 14252 15092 14420 15148
rect 12460 11414 12516 11452
rect 11676 11342 11678 11394
rect 11730 11342 11732 11394
rect 11676 11330 11732 11342
rect 11564 11284 11620 11294
rect 11564 11190 11620 11228
rect 11452 11172 11508 11182
rect 11228 9986 11284 9996
rect 11340 11170 11508 11172
rect 11340 11118 11454 11170
rect 11506 11118 11508 11170
rect 11340 11116 11508 11118
rect 11340 10610 11396 11116
rect 11452 11106 11508 11116
rect 11900 11170 11956 11182
rect 11900 11118 11902 11170
rect 11954 11118 11956 11170
rect 11340 10558 11342 10610
rect 11394 10558 11396 10610
rect 8652 9884 9716 9940
rect 8652 9826 8708 9884
rect 8652 9774 8654 9826
rect 8706 9774 8708 9826
rect 8652 9762 8708 9774
rect 9324 9716 9380 9726
rect 9324 9622 9380 9660
rect 8764 9156 8820 9166
rect 8764 9154 9380 9156
rect 8764 9102 8766 9154
rect 8818 9102 9380 9154
rect 8764 9100 9380 9102
rect 8764 9090 8820 9100
rect 8876 8932 8932 8942
rect 8876 8838 8932 8876
rect 8988 8820 9044 8830
rect 8540 8764 8820 8820
rect 8540 7700 8596 7710
rect 8428 7698 8596 7700
rect 8428 7646 8542 7698
rect 8594 7646 8596 7698
rect 8428 7644 8596 7646
rect 8540 7634 8596 7644
rect 8316 7476 8372 7486
rect 7980 6750 7982 6802
rect 8034 6750 8036 6802
rect 7980 6738 8036 6750
rect 8092 7474 8372 7476
rect 8092 7422 8318 7474
rect 8370 7422 8372 7474
rect 8092 7420 8372 7422
rect 6636 6468 6692 6478
rect 7084 6468 7140 6478
rect 7644 6468 7700 6478
rect 6636 6466 7028 6468
rect 6636 6414 6638 6466
rect 6690 6414 7028 6466
rect 6636 6412 7028 6414
rect 6636 6402 6692 6412
rect 6300 5954 6356 5964
rect 6636 6020 6692 6030
rect 6636 5926 6692 5964
rect 6188 5794 6244 5806
rect 6188 5742 6190 5794
rect 6242 5742 6244 5794
rect 6188 5684 6244 5742
rect 6860 5796 6916 5806
rect 6188 5628 6580 5684
rect 6300 5460 6356 5470
rect 6076 5124 6132 5134
rect 6076 4562 6132 5068
rect 6188 5122 6244 5134
rect 6188 5070 6190 5122
rect 6242 5070 6244 5122
rect 6188 4900 6244 5070
rect 6188 4834 6244 4844
rect 6076 4510 6078 4562
rect 6130 4510 6132 4562
rect 6076 4498 6132 4510
rect 6188 4564 6244 4574
rect 6300 4564 6356 5404
rect 6524 5348 6580 5628
rect 6188 4562 6356 4564
rect 6188 4510 6190 4562
rect 6242 4510 6356 4562
rect 6188 4508 6356 4510
rect 6412 5292 6580 5348
rect 6188 4498 6244 4508
rect 6188 4228 6244 4238
rect 6076 3444 6132 3454
rect 5964 3442 6132 3444
rect 5964 3390 6078 3442
rect 6130 3390 6132 3442
rect 5964 3388 6132 3390
rect 6076 3378 6132 3388
rect 6188 3388 6244 4172
rect 6412 4228 6468 5292
rect 6860 5236 6916 5740
rect 6636 5180 6916 5236
rect 6412 4162 6468 4172
rect 6524 5122 6580 5134
rect 6524 5070 6526 5122
rect 6578 5070 6580 5122
rect 6524 4900 6580 5070
rect 6300 4116 6356 4126
rect 6300 4022 6356 4060
rect 6524 4004 6580 4844
rect 6636 4788 6692 5180
rect 6748 5012 6804 5022
rect 6748 4918 6804 4956
rect 6860 4900 6916 4910
rect 6636 4732 6804 4788
rect 6636 4340 6692 4350
rect 6636 4246 6692 4284
rect 6748 4226 6804 4732
rect 6748 4174 6750 4226
rect 6802 4174 6804 4226
rect 6748 4162 6804 4174
rect 6860 4116 6916 4844
rect 6972 4452 7028 6412
rect 7084 6466 7252 6468
rect 7084 6414 7086 6466
rect 7138 6414 7252 6466
rect 7084 6412 7252 6414
rect 7084 6402 7140 6412
rect 7084 5794 7140 5806
rect 7084 5742 7086 5794
rect 7138 5742 7140 5794
rect 7084 4676 7140 5742
rect 7084 4610 7140 4620
rect 6972 4396 7140 4452
rect 6972 4116 7028 4154
rect 6860 4060 6972 4116
rect 6972 4050 7028 4060
rect 6524 3938 6580 3948
rect 6972 3892 7028 3902
rect 6524 3556 6580 3566
rect 6524 3462 6580 3500
rect 6188 3332 6356 3388
rect 6300 800 6356 3332
rect 6748 3332 6804 3342
rect 6748 3238 6804 3276
rect 6972 800 7028 3836
rect 7084 3554 7140 4396
rect 7084 3502 7086 3554
rect 7138 3502 7140 3554
rect 7084 2660 7140 3502
rect 7196 3556 7252 6412
rect 7420 6466 7700 6468
rect 7420 6414 7646 6466
rect 7698 6414 7700 6466
rect 7420 6412 7700 6414
rect 7308 5122 7364 5134
rect 7308 5070 7310 5122
rect 7362 5070 7364 5122
rect 7308 5012 7364 5070
rect 7308 4946 7364 4956
rect 7308 4338 7364 4350
rect 7308 4286 7310 4338
rect 7362 4286 7364 4338
rect 7308 4116 7364 4286
rect 7420 4228 7476 6412
rect 7644 6402 7700 6412
rect 7980 6466 8036 6478
rect 7980 6414 7982 6466
rect 8034 6414 8036 6466
rect 7868 6244 7924 6254
rect 7868 5908 7924 6188
rect 7980 6132 8036 6414
rect 7980 6066 8036 6076
rect 7980 5908 8036 5918
rect 7868 5906 8036 5908
rect 7868 5854 7982 5906
rect 8034 5854 8036 5906
rect 7868 5852 8036 5854
rect 7980 5842 8036 5852
rect 8092 5908 8148 7420
rect 8316 7410 8372 7420
rect 8652 7250 8708 7262
rect 8652 7198 8654 7250
rect 8706 7198 8708 7250
rect 8204 6916 8260 6926
rect 8204 6822 8260 6860
rect 8652 6916 8708 7198
rect 8652 6850 8708 6860
rect 8764 6802 8820 8764
rect 8988 8726 9044 8764
rect 8764 6750 8766 6802
rect 8818 6750 8820 6802
rect 8764 6738 8820 6750
rect 8876 6916 8932 6926
rect 9212 6916 9268 6926
rect 8932 6914 9268 6916
rect 8932 6862 9214 6914
rect 9266 6862 9268 6914
rect 8932 6860 9268 6862
rect 8652 6468 8708 6478
rect 8652 6374 8708 6412
rect 8876 6244 8932 6860
rect 9212 6850 9268 6860
rect 9324 6802 9380 9100
rect 9660 9042 9716 9884
rect 9660 8990 9662 9042
rect 9714 8990 9716 9042
rect 9660 8260 9716 8990
rect 9996 9716 10052 9726
rect 9772 8260 9828 8270
rect 9660 8258 9940 8260
rect 9660 8206 9774 8258
rect 9826 8206 9940 8258
rect 9660 8204 9940 8206
rect 9772 8194 9828 8204
rect 9324 6750 9326 6802
rect 9378 6750 9380 6802
rect 9324 6738 9380 6750
rect 9548 7140 9604 7150
rect 9436 6580 9492 6590
rect 9436 6486 9492 6524
rect 8652 6188 8932 6244
rect 8988 6468 9044 6478
rect 8316 6132 8372 6142
rect 8316 6038 8372 6076
rect 8652 6130 8708 6188
rect 8652 6078 8654 6130
rect 8706 6078 8708 6130
rect 8652 6066 8708 6078
rect 8988 6132 9044 6412
rect 8092 5842 8148 5852
rect 8428 6020 8484 6030
rect 7532 5794 7588 5806
rect 7532 5742 7534 5794
rect 7586 5742 7588 5794
rect 7532 5682 7588 5742
rect 7532 5630 7534 5682
rect 7586 5630 7588 5682
rect 7532 5618 7588 5630
rect 8204 5682 8260 5694
rect 8204 5630 8206 5682
rect 8258 5630 8260 5682
rect 7644 5348 7700 5358
rect 7644 5010 7700 5292
rect 7644 4958 7646 5010
rect 7698 4958 7700 5010
rect 7532 4898 7588 4910
rect 7532 4846 7534 4898
rect 7586 4846 7588 4898
rect 7532 4676 7588 4846
rect 7644 4900 7700 4958
rect 7980 5124 8036 5134
rect 8204 5124 8260 5630
rect 7980 5010 8036 5068
rect 7980 4958 7982 5010
rect 8034 4958 8036 5010
rect 7980 4946 8036 4958
rect 8092 5122 8260 5124
rect 8092 5070 8206 5122
rect 8258 5070 8260 5122
rect 8092 5068 8260 5070
rect 7644 4834 7700 4844
rect 7532 4620 8036 4676
rect 7644 4452 7700 4462
rect 7644 4358 7700 4396
rect 7980 4338 8036 4620
rect 7980 4286 7982 4338
rect 8034 4286 8036 4338
rect 7980 4274 8036 4286
rect 7420 4172 7812 4228
rect 7308 4050 7364 4060
rect 7196 3490 7252 3500
rect 7420 3892 7476 3902
rect 7420 3442 7476 3836
rect 7756 3554 7812 4172
rect 8092 3892 8148 5068
rect 8204 5058 8260 5068
rect 8316 5236 8372 5246
rect 8316 4450 8372 5180
rect 8428 4676 8484 5964
rect 8988 6018 9044 6076
rect 8988 5966 8990 6018
rect 9042 5966 9044 6018
rect 8988 5954 9044 5966
rect 8652 5572 8708 5582
rect 8652 5122 8708 5516
rect 8988 5348 9044 5358
rect 9044 5292 9380 5348
rect 8988 5254 9044 5292
rect 8652 5070 8654 5122
rect 8706 5070 8708 5122
rect 8652 5058 8708 5070
rect 8876 5124 8932 5134
rect 8876 5030 8932 5068
rect 9324 5010 9380 5292
rect 9324 4958 9326 5010
rect 9378 4958 9380 5010
rect 9324 4946 9380 4958
rect 9548 4788 9604 7084
rect 9660 6468 9716 6478
rect 9660 5122 9716 6412
rect 9884 5908 9940 8204
rect 9996 6468 10052 9660
rect 11340 9604 11396 10558
rect 11564 10836 11620 10846
rect 11452 10500 11508 10510
rect 11452 10406 11508 10444
rect 11564 9938 11620 10780
rect 11564 9886 11566 9938
rect 11618 9886 11620 9938
rect 11564 9874 11620 9886
rect 11900 10610 11956 11118
rect 11900 10558 11902 10610
rect 11954 10558 11956 10610
rect 11900 9828 11956 10558
rect 12684 10612 12740 10622
rect 12684 10518 12740 10556
rect 11900 9762 11956 9772
rect 12236 10052 12292 10062
rect 12236 9826 12292 9996
rect 12236 9774 12238 9826
rect 12290 9774 12292 9826
rect 11340 9538 11396 9548
rect 12012 9604 12068 9614
rect 12012 9510 12068 9548
rect 12124 9602 12180 9614
rect 12124 9550 12126 9602
rect 12178 9550 12180 9602
rect 10332 8932 10388 8942
rect 10332 8838 10388 8876
rect 12124 8820 12180 9550
rect 12236 8932 12292 9774
rect 12572 9828 12628 9838
rect 12572 9734 12628 9772
rect 12460 8932 12516 8942
rect 12236 8876 12460 8932
rect 12460 8838 12516 8876
rect 12124 8754 12180 8764
rect 12796 8260 12852 15092
rect 13468 11508 13524 11518
rect 13356 11506 13524 11508
rect 13356 11454 13470 11506
rect 13522 11454 13524 11506
rect 13356 11452 13524 11454
rect 13356 10722 13412 11452
rect 13468 11442 13524 11452
rect 13804 11284 13860 11294
rect 13692 11282 13860 11284
rect 13692 11230 13806 11282
rect 13858 11230 13860 11282
rect 13692 11228 13860 11230
rect 13580 11172 13636 11182
rect 13356 10670 13358 10722
rect 13410 10670 13412 10722
rect 13356 10658 13412 10670
rect 13468 11170 13636 11172
rect 13468 11118 13582 11170
rect 13634 11118 13636 11170
rect 13468 11116 13636 11118
rect 13468 9940 13524 11116
rect 13580 11106 13636 11116
rect 13468 9874 13524 9884
rect 13580 9940 13636 9950
rect 13692 9940 13748 11228
rect 13804 11218 13860 11228
rect 13916 9940 13972 9950
rect 13580 9938 13748 9940
rect 13580 9886 13582 9938
rect 13634 9886 13748 9938
rect 13580 9884 13748 9886
rect 13804 9884 13916 9940
rect 13580 9874 13636 9884
rect 13244 9828 13300 9838
rect 13300 9772 13412 9828
rect 13244 9762 13300 9772
rect 13356 9268 13412 9772
rect 13692 9716 13748 9726
rect 13804 9716 13860 9884
rect 13916 9874 13972 9884
rect 14028 9828 14084 9838
rect 14028 9734 14084 9772
rect 13692 9714 13860 9716
rect 13692 9662 13694 9714
rect 13746 9662 13860 9714
rect 13692 9660 13860 9662
rect 13692 9650 13748 9660
rect 13468 9604 13524 9614
rect 13468 9510 13524 9548
rect 14140 9604 14196 9614
rect 13468 9268 13524 9278
rect 13356 9266 13524 9268
rect 13356 9214 13470 9266
rect 13522 9214 13524 9266
rect 13356 9212 13524 9214
rect 13468 9202 13524 9212
rect 13804 9268 13860 9278
rect 13804 9174 13860 9212
rect 14140 9266 14196 9548
rect 14140 9214 14142 9266
rect 14194 9214 14196 9266
rect 14140 9202 14196 9214
rect 14252 9268 14308 9278
rect 13244 8932 13300 8942
rect 13244 8838 13300 8876
rect 12460 8204 12852 8260
rect 14028 8258 14084 8270
rect 14028 8206 14030 8258
rect 14082 8206 14084 8258
rect 10556 8148 10612 8158
rect 10556 8146 10948 8148
rect 10556 8094 10558 8146
rect 10610 8094 10948 8146
rect 10556 8092 10948 8094
rect 10556 8082 10612 8092
rect 10220 7364 10276 7374
rect 9996 6402 10052 6412
rect 10108 7362 10276 7364
rect 10108 7310 10222 7362
rect 10274 7310 10276 7362
rect 10108 7308 10276 7310
rect 10108 6244 10164 7308
rect 10220 7298 10276 7308
rect 10892 7362 10948 8092
rect 10892 7310 10894 7362
rect 10946 7310 10948 7362
rect 10892 7298 10948 7310
rect 11004 7586 11060 7598
rect 11004 7534 11006 7586
rect 11058 7534 11060 7586
rect 10780 6804 10836 6814
rect 10220 6468 10276 6478
rect 10220 6466 10500 6468
rect 10220 6414 10222 6466
rect 10274 6414 10500 6466
rect 10220 6412 10500 6414
rect 10220 6402 10276 6412
rect 10108 6188 10388 6244
rect 10220 5908 10276 5918
rect 9884 5906 10052 5908
rect 9884 5854 9886 5906
rect 9938 5854 10052 5906
rect 9884 5852 10052 5854
rect 9884 5842 9940 5852
rect 9660 5070 9662 5122
rect 9714 5070 9716 5122
rect 9660 5058 9716 5070
rect 9996 5012 10052 5852
rect 10220 5234 10276 5852
rect 10220 5182 10222 5234
rect 10274 5182 10276 5234
rect 10220 5170 10276 5182
rect 9996 4956 10164 5012
rect 8988 4732 9604 4788
rect 8540 4676 8596 4686
rect 8428 4620 8540 4676
rect 8316 4398 8318 4450
rect 8370 4398 8372 4450
rect 8316 4386 8372 4398
rect 8204 4228 8260 4238
rect 8204 4134 8260 4172
rect 8092 3836 8372 3892
rect 7756 3502 7758 3554
rect 7810 3502 7812 3554
rect 7420 3390 7422 3442
rect 7474 3390 7476 3442
rect 7420 3378 7476 3390
rect 7532 3444 7588 3454
rect 7532 3220 7588 3388
rect 7532 3164 7700 3220
rect 7084 2594 7140 2604
rect 7644 800 7700 3164
rect 7756 2548 7812 3502
rect 7756 2482 7812 2492
rect 8092 3330 8148 3342
rect 8092 3278 8094 3330
rect 8146 3278 8148 3330
rect 8092 2324 8148 3278
rect 8092 2258 8148 2268
rect 8316 800 8372 3836
rect 8540 3554 8596 4620
rect 8764 4564 8820 4574
rect 8764 4338 8820 4508
rect 8988 4562 9044 4732
rect 8988 4510 8990 4562
rect 9042 4510 9044 4562
rect 8988 4498 9044 4510
rect 9884 4452 9940 4462
rect 9884 4450 10052 4452
rect 9884 4398 9886 4450
rect 9938 4398 10052 4450
rect 9884 4396 10052 4398
rect 9884 4386 9940 4396
rect 8764 4286 8766 4338
rect 8818 4286 8820 4338
rect 8764 4274 8820 4286
rect 9660 4338 9716 4350
rect 9660 4286 9662 4338
rect 9714 4286 9716 4338
rect 9660 4116 9716 4286
rect 9660 4050 9716 4060
rect 8540 3502 8542 3554
rect 8594 3502 8596 3554
rect 8540 3490 8596 3502
rect 8988 4004 9044 4014
rect 8764 3442 8820 3454
rect 8764 3390 8766 3442
rect 8818 3390 8820 3442
rect 8764 3220 8820 3390
rect 8764 3154 8820 3164
rect 8988 800 9044 3948
rect 9548 3780 9604 3790
rect 9548 3388 9604 3724
rect 9660 3556 9716 3594
rect 9660 3490 9716 3500
rect 9548 3332 9716 3388
rect 9660 800 9716 3332
rect 9884 3330 9940 3342
rect 9884 3278 9886 3330
rect 9938 3278 9940 3330
rect 9884 2884 9940 3278
rect 9996 3332 10052 4396
rect 10108 4340 10164 4956
rect 10220 4340 10276 4350
rect 10108 4284 10220 4340
rect 10220 4246 10276 4284
rect 10220 4116 10276 4126
rect 10332 4116 10388 6188
rect 10276 4060 10388 4116
rect 10220 4050 10276 4060
rect 10332 3892 10388 3902
rect 10220 3836 10332 3892
rect 10220 3554 10276 3836
rect 10332 3826 10388 3836
rect 10220 3502 10222 3554
rect 10274 3502 10276 3554
rect 10220 3490 10276 3502
rect 10332 3668 10388 3678
rect 9996 3266 10052 3276
rect 9884 2818 9940 2828
rect 10332 800 10388 3612
rect 10444 3556 10500 6412
rect 10668 5794 10724 5806
rect 10668 5742 10670 5794
rect 10722 5742 10724 5794
rect 10556 5460 10612 5470
rect 10556 5010 10612 5404
rect 10668 5234 10724 5742
rect 10780 5346 10836 6748
rect 10780 5294 10782 5346
rect 10834 5294 10836 5346
rect 10780 5282 10836 5294
rect 10892 6466 10948 6478
rect 10892 6414 10894 6466
rect 10946 6414 10948 6466
rect 10668 5182 10670 5234
rect 10722 5182 10724 5234
rect 10668 5170 10724 5182
rect 10556 4958 10558 5010
rect 10610 4958 10612 5010
rect 10556 4946 10612 4958
rect 10892 4676 10948 6414
rect 11004 5796 11060 7534
rect 11004 5730 11060 5740
rect 11116 7476 11172 7486
rect 10780 4620 10948 4676
rect 10780 3892 10836 4620
rect 10780 3826 10836 3836
rect 10892 4452 10948 4462
rect 10444 3108 10500 3500
rect 10892 3554 10948 4396
rect 11004 4228 11060 4238
rect 11004 4134 11060 4172
rect 11116 3666 11172 7420
rect 11228 7364 11284 7374
rect 11228 7270 11284 7308
rect 11788 7364 11844 7374
rect 11788 7362 12292 7364
rect 11788 7310 11790 7362
rect 11842 7310 12292 7362
rect 11788 7308 12292 7310
rect 11788 7298 11844 7308
rect 12124 6692 12180 6702
rect 12124 6598 12180 6636
rect 11676 6468 11732 6478
rect 11564 6466 11732 6468
rect 11564 6414 11678 6466
rect 11730 6414 11732 6466
rect 11564 6412 11732 6414
rect 11228 5684 11284 5694
rect 11228 3778 11284 5628
rect 11452 5348 11508 5358
rect 11452 5234 11508 5292
rect 11452 5182 11454 5234
rect 11506 5182 11508 5234
rect 11452 5170 11508 5182
rect 11228 3726 11230 3778
rect 11282 3726 11284 3778
rect 11228 3714 11284 3726
rect 11452 4004 11508 4014
rect 11116 3614 11118 3666
rect 11170 3614 11172 3666
rect 11116 3602 11172 3614
rect 10892 3502 10894 3554
rect 10946 3502 10948 3554
rect 10892 3490 10948 3502
rect 11004 3444 11060 3454
rect 10444 3042 10500 3052
rect 10556 3330 10612 3342
rect 10556 3278 10558 3330
rect 10610 3278 10612 3330
rect 10556 2436 10612 3278
rect 10556 2370 10612 2380
rect 11004 800 11060 3388
rect 11452 3388 11508 3948
rect 11564 3556 11620 6412
rect 11676 6402 11732 6412
rect 12012 5796 12068 5806
rect 12012 5346 12068 5740
rect 12012 5294 12014 5346
rect 12066 5294 12068 5346
rect 12012 5282 12068 5294
rect 11676 5124 11732 5134
rect 11676 5030 11732 5068
rect 11900 4898 11956 4910
rect 11900 4846 11902 4898
rect 11954 4846 11956 4898
rect 11900 4228 11956 4846
rect 11900 4162 11956 4172
rect 12236 4452 12292 7308
rect 12348 6916 12404 6926
rect 12348 5122 12404 6860
rect 12460 6244 12516 8204
rect 12796 8034 12852 8046
rect 12796 7982 12798 8034
rect 12850 7982 12852 8034
rect 12796 7700 12852 7982
rect 13692 8036 13748 8046
rect 14028 8036 14084 8206
rect 14252 8146 14308 9212
rect 14252 8094 14254 8146
rect 14306 8094 14308 8146
rect 14252 8082 14308 8094
rect 13692 8034 14084 8036
rect 13692 7982 13694 8034
rect 13746 7982 14084 8034
rect 13692 7980 14084 7982
rect 13692 7970 13748 7980
rect 13132 7700 13188 7710
rect 12796 7644 13132 7700
rect 13132 7606 13188 7644
rect 13580 7700 13636 7710
rect 13580 7606 13636 7644
rect 13804 7588 13860 7598
rect 13692 7532 13804 7588
rect 13356 7474 13412 7486
rect 13356 7422 13358 7474
rect 13410 7422 13412 7474
rect 12684 7364 12740 7374
rect 12684 7362 13300 7364
rect 12684 7310 12686 7362
rect 12738 7310 13300 7362
rect 12684 7308 13300 7310
rect 12684 7298 12740 7308
rect 12796 6692 12852 6702
rect 12572 6468 12628 6478
rect 12572 6466 12740 6468
rect 12572 6414 12574 6466
rect 12626 6414 12740 6466
rect 12572 6412 12740 6414
rect 12572 6402 12628 6412
rect 12684 6244 12740 6412
rect 12460 6188 12628 6244
rect 12572 5908 12628 6188
rect 12684 6178 12740 6188
rect 12460 5236 12516 5246
rect 12460 5142 12516 5180
rect 12348 5070 12350 5122
rect 12402 5070 12404 5122
rect 12348 5058 12404 5070
rect 11676 3556 11732 3594
rect 11564 3500 11676 3556
rect 11676 3490 11732 3500
rect 12236 3554 12292 4396
rect 12572 5010 12628 5852
rect 12796 5794 12852 6636
rect 12796 5742 12798 5794
rect 12850 5742 12852 5794
rect 12796 5730 12852 5742
rect 12908 6468 12964 6478
rect 12908 5122 12964 6412
rect 12908 5070 12910 5122
rect 12962 5070 12964 5122
rect 12908 5058 12964 5070
rect 13020 6466 13076 6478
rect 13020 6414 13022 6466
rect 13074 6414 13076 6466
rect 13020 5124 13076 6414
rect 13244 5236 13300 7308
rect 13356 6916 13412 7422
rect 13468 7364 13524 7374
rect 13468 7270 13524 7308
rect 13468 6916 13524 6926
rect 13356 6860 13468 6916
rect 13468 6468 13524 6860
rect 13580 6804 13636 6814
rect 13580 6710 13636 6748
rect 13692 6804 13748 7532
rect 13804 7522 13860 7532
rect 13916 7474 13972 7486
rect 13916 7422 13918 7474
rect 13970 7422 13972 7474
rect 13804 6804 13860 6814
rect 13692 6748 13804 6804
rect 13692 6690 13748 6748
rect 13804 6738 13860 6748
rect 13692 6638 13694 6690
rect 13746 6638 13748 6690
rect 13692 6626 13748 6638
rect 13916 6468 13972 7422
rect 14028 6580 14084 7980
rect 14364 7700 14420 15092
rect 14588 11732 14644 11742
rect 14476 9940 14532 9950
rect 14476 9846 14532 9884
rect 14364 7634 14420 7644
rect 14476 9716 14532 9726
rect 14476 9266 14532 9660
rect 14476 9214 14478 9266
rect 14530 9214 14532 9266
rect 14252 7586 14308 7598
rect 14252 7534 14254 7586
rect 14306 7534 14308 7586
rect 14252 6916 14308 7534
rect 14476 7474 14532 9214
rect 14588 7588 14644 11676
rect 14924 10836 14980 23100
rect 16156 23492 16212 23502
rect 15596 22484 15652 22494
rect 15652 22428 16100 22484
rect 15596 22390 15652 22428
rect 16044 22258 16100 22428
rect 16156 22370 16212 23436
rect 16156 22318 16158 22370
rect 16210 22318 16212 22370
rect 16156 22306 16212 22318
rect 16044 22206 16046 22258
rect 16098 22206 16100 22258
rect 16044 22194 16100 22206
rect 15820 22146 15876 22158
rect 15820 22094 15822 22146
rect 15874 22094 15876 22146
rect 15484 21812 15540 21822
rect 15484 21476 15540 21756
rect 15820 21812 15876 22094
rect 15820 21746 15876 21756
rect 14924 10770 14980 10780
rect 15372 11394 15428 11406
rect 15372 11342 15374 11394
rect 15426 11342 15428 11394
rect 15372 10612 15428 11342
rect 14924 10052 14980 10062
rect 14924 9268 14980 9996
rect 15372 9940 15428 10556
rect 14924 9174 14980 9212
rect 15148 9938 15428 9940
rect 15148 9886 15374 9938
rect 15426 9886 15428 9938
rect 15148 9884 15428 9886
rect 15148 8428 15204 9884
rect 15372 9874 15428 9884
rect 15484 10498 15540 21420
rect 15484 10446 15486 10498
rect 15538 10446 15540 10498
rect 15484 9940 15540 10446
rect 15484 9874 15540 9884
rect 16044 11844 16100 11854
rect 15372 9156 15428 9166
rect 15372 9154 15540 9156
rect 15372 9102 15374 9154
rect 15426 9102 15540 9154
rect 15372 9100 15540 9102
rect 15372 9090 15428 9100
rect 14924 8372 15204 8428
rect 15372 8930 15428 8942
rect 15372 8878 15374 8930
rect 15426 8878 15428 8930
rect 14588 7522 14644 7532
rect 14700 8260 14756 8270
rect 14924 8260 14980 8372
rect 15372 8370 15428 8878
rect 15372 8318 15374 8370
rect 15426 8318 15428 8370
rect 15372 8306 15428 8318
rect 14700 8258 14980 8260
rect 14700 8206 14702 8258
rect 14754 8206 14980 8258
rect 14700 8204 14980 8206
rect 14476 7422 14478 7474
rect 14530 7422 14532 7474
rect 14476 7410 14532 7422
rect 14700 7252 14756 8204
rect 14252 6850 14308 6860
rect 14588 7196 14756 7252
rect 15260 7362 15316 7374
rect 15260 7310 15262 7362
rect 15314 7310 15316 7362
rect 14028 6514 14084 6524
rect 14252 6692 14308 6702
rect 13468 6466 13636 6468
rect 13468 6414 13470 6466
rect 13522 6414 13636 6466
rect 13468 6412 13636 6414
rect 13468 6402 13524 6412
rect 13580 6244 13636 6412
rect 13916 6374 13972 6412
rect 14140 6244 14196 6254
rect 13580 6188 13972 6244
rect 13468 6132 13524 6142
rect 13524 6076 13636 6132
rect 13468 6066 13524 6076
rect 13468 5572 13524 5582
rect 13580 5572 13636 6076
rect 13916 6130 13972 6188
rect 13916 6078 13918 6130
rect 13970 6078 13972 6130
rect 13916 6066 13972 6078
rect 13692 6020 13748 6030
rect 13692 5926 13748 5964
rect 14140 6018 14196 6188
rect 14140 5966 14142 6018
rect 14194 5966 14196 6018
rect 14140 5954 14196 5966
rect 14028 5908 14084 5946
rect 14028 5842 14084 5852
rect 13804 5684 13860 5694
rect 13580 5516 13748 5572
rect 13468 5236 13524 5516
rect 13244 5180 13412 5236
rect 13020 5058 13076 5068
rect 12572 4958 12574 5010
rect 12626 4958 12628 5010
rect 12572 4228 12628 4958
rect 13356 5012 13412 5180
rect 13468 5170 13524 5180
rect 13692 5234 13748 5516
rect 13692 5182 13694 5234
rect 13746 5182 13748 5234
rect 13692 5170 13748 5182
rect 13356 4956 13524 5012
rect 13132 4228 13188 4238
rect 12572 4226 13188 4228
rect 12572 4174 13134 4226
rect 13186 4174 13188 4226
rect 12572 4172 13188 4174
rect 13132 4162 13188 4172
rect 12236 3502 12238 3554
rect 12290 3502 12292 3554
rect 12236 3490 12292 3502
rect 13468 3780 13524 4956
rect 13804 4900 13860 5628
rect 14028 5572 14084 5582
rect 13804 4834 13860 4844
rect 13916 5460 13972 5470
rect 13692 4340 13748 4350
rect 13692 4246 13748 4284
rect 13468 3554 13524 3724
rect 13468 3502 13470 3554
rect 13522 3502 13524 3554
rect 13468 3490 13524 3502
rect 13580 4116 13636 4126
rect 12572 3444 12628 3482
rect 11452 3332 11732 3388
rect 12572 3378 12628 3388
rect 11676 800 11732 3332
rect 11900 3330 11956 3342
rect 11900 3278 11902 3330
rect 11954 3278 11956 3330
rect 11900 2996 11956 3278
rect 13580 3220 13636 4060
rect 13692 3444 13748 3454
rect 13916 3444 13972 5404
rect 14028 5010 14084 5516
rect 14252 5348 14308 6636
rect 14588 6692 14644 7196
rect 14924 6692 14980 6702
rect 14588 6690 14980 6692
rect 14588 6638 14926 6690
rect 14978 6638 14980 6690
rect 14588 6636 14980 6638
rect 14364 6468 14420 6478
rect 14364 6130 14420 6412
rect 14364 6078 14366 6130
rect 14418 6078 14420 6130
rect 14364 6066 14420 6078
rect 14140 5292 14308 5348
rect 14140 5234 14196 5292
rect 14140 5182 14142 5234
rect 14194 5182 14196 5234
rect 14140 5170 14196 5182
rect 14588 5124 14644 6636
rect 14924 6626 14980 6636
rect 14700 6468 14756 6478
rect 14700 6374 14756 6412
rect 14812 6356 14868 6366
rect 14812 6130 14868 6300
rect 14812 6078 14814 6130
rect 14866 6078 14868 6130
rect 14812 6066 14868 6078
rect 15148 6132 15204 6142
rect 15148 6038 15204 6076
rect 14700 5908 14756 5918
rect 14700 5234 14756 5852
rect 15260 5460 15316 7310
rect 15484 6132 15540 9100
rect 15932 9042 15988 9054
rect 15932 8990 15934 9042
rect 15986 8990 15988 9042
rect 15596 8818 15652 8830
rect 15596 8766 15598 8818
rect 15650 8766 15652 8818
rect 15596 8372 15652 8766
rect 15596 8306 15652 8316
rect 15596 7588 15652 7598
rect 15596 7494 15652 7532
rect 15708 7362 15764 7374
rect 15708 7310 15710 7362
rect 15762 7310 15764 7362
rect 15708 6802 15764 7310
rect 15820 7364 15876 7374
rect 15820 7270 15876 7308
rect 15708 6750 15710 6802
rect 15762 6750 15764 6802
rect 15708 6738 15764 6750
rect 15932 6692 15988 8990
rect 15932 6626 15988 6636
rect 15596 6132 15652 6142
rect 15484 6130 15652 6132
rect 15484 6078 15598 6130
rect 15650 6078 15652 6130
rect 15484 6076 15652 6078
rect 15596 6066 15652 6076
rect 15708 6018 15764 6030
rect 15708 5966 15710 6018
rect 15762 5966 15764 6018
rect 15596 5796 15652 5806
rect 15148 5404 15316 5460
rect 15484 5682 15540 5694
rect 15484 5630 15486 5682
rect 15538 5630 15540 5682
rect 14700 5182 14702 5234
rect 14754 5182 14756 5234
rect 14700 5170 14756 5182
rect 14812 5348 14868 5358
rect 14028 4958 14030 5010
rect 14082 4958 14084 5010
rect 14028 4946 14084 4958
rect 14140 5012 14196 5022
rect 14140 3892 14196 4956
rect 14252 5010 14308 5022
rect 14252 4958 14254 5010
rect 14306 4958 14308 5010
rect 14252 4900 14308 4958
rect 14252 4834 14308 4844
rect 14364 4788 14420 4798
rect 14140 3554 14196 3836
rect 14140 3502 14142 3554
rect 14194 3502 14196 3554
rect 14140 3490 14196 3502
rect 14252 4564 14308 4574
rect 13692 3442 13972 3444
rect 13692 3390 13694 3442
rect 13746 3390 13972 3442
rect 13692 3388 13972 3390
rect 13692 3378 13748 3388
rect 13580 3164 13748 3220
rect 11900 2930 11956 2940
rect 12348 2660 12404 2670
rect 12348 800 12404 2604
rect 13020 2548 13076 2558
rect 13020 800 13076 2492
rect 13692 800 13748 3164
rect 14252 3108 14308 4508
rect 14364 3442 14420 4732
rect 14588 4340 14644 5068
rect 14700 5012 14756 5022
rect 14700 4918 14756 4956
rect 14588 4274 14644 4284
rect 14476 4228 14532 4238
rect 14476 4134 14532 4172
rect 14812 3668 14868 5292
rect 14924 5010 14980 5022
rect 14924 4958 14926 5010
rect 14978 4958 14980 5010
rect 14924 4900 14980 4958
rect 14924 4834 14980 4844
rect 14812 3554 14868 3612
rect 14812 3502 14814 3554
rect 14866 3502 14868 3554
rect 14812 3490 14868 3502
rect 14924 4676 14980 4686
rect 14364 3390 14366 3442
rect 14418 3390 14420 3442
rect 14364 3378 14420 3390
rect 14924 3220 14980 4620
rect 15148 4676 15204 5404
rect 15260 4900 15316 4910
rect 15484 4900 15540 5630
rect 15596 5122 15652 5740
rect 15596 5070 15598 5122
rect 15650 5070 15652 5122
rect 15596 5058 15652 5070
rect 15316 4844 15540 4900
rect 15260 4806 15316 4844
rect 15708 4676 15764 5966
rect 16044 5460 16100 11788
rect 16380 11732 16436 24556
rect 17052 31892 17220 31948
rect 17276 31892 17668 31948
rect 16828 23938 16884 23950
rect 16828 23886 16830 23938
rect 16882 23886 16884 23938
rect 16604 22372 16660 22382
rect 16828 22372 16884 23886
rect 16604 22370 16828 22372
rect 16604 22318 16606 22370
rect 16658 22318 16828 22370
rect 16604 22316 16828 22318
rect 16604 22306 16660 22316
rect 16828 22278 16884 22316
rect 16716 22148 16772 22158
rect 16604 13636 16660 13646
rect 16604 12962 16660 13580
rect 16604 12910 16606 12962
rect 16658 12910 16660 12962
rect 16604 12898 16660 12910
rect 16380 11666 16436 11676
rect 16156 11282 16212 11294
rect 16156 11230 16158 11282
rect 16210 11230 16212 11282
rect 16156 9266 16212 11230
rect 16156 9214 16158 9266
rect 16210 9214 16212 9266
rect 16156 9202 16212 9214
rect 16268 8932 16324 8942
rect 16268 8838 16324 8876
rect 16492 7364 16548 7374
rect 16492 7362 16660 7364
rect 16492 7310 16494 7362
rect 16546 7310 16660 7362
rect 16492 7308 16660 7310
rect 16492 7298 16548 7308
rect 15148 4610 15204 4620
rect 15260 4620 15764 4676
rect 15820 5404 16100 5460
rect 16492 6018 16548 6030
rect 16492 5966 16494 6018
rect 16546 5966 16548 6018
rect 15036 4340 15092 4350
rect 15036 3442 15092 4284
rect 15036 3390 15038 3442
rect 15090 3390 15092 3442
rect 15036 3378 15092 3390
rect 14924 3164 15092 3220
rect 14252 3052 14420 3108
rect 14364 800 14420 3052
rect 15036 800 15092 3164
rect 15260 2772 15316 4620
rect 15820 4564 15876 5404
rect 15932 5124 15988 5134
rect 15932 5030 15988 5068
rect 16492 5124 16548 5966
rect 16604 5348 16660 7308
rect 16716 6244 16772 22092
rect 17052 20132 17108 31892
rect 17276 26908 17332 31892
rect 17052 20066 17108 20076
rect 17164 26852 17332 26908
rect 17164 19236 17220 26852
rect 17500 24834 17556 24846
rect 17500 24782 17502 24834
rect 17554 24782 17556 24834
rect 17388 24722 17444 24734
rect 17388 24670 17390 24722
rect 17442 24670 17444 24722
rect 17388 23604 17444 24670
rect 17500 24388 17556 24782
rect 17500 24322 17556 24332
rect 17724 24722 17780 24734
rect 17724 24670 17726 24722
rect 17778 24670 17780 24722
rect 17388 23538 17444 23548
rect 17500 23826 17556 23838
rect 17500 23774 17502 23826
rect 17554 23774 17556 23826
rect 17500 23378 17556 23774
rect 17500 23326 17502 23378
rect 17554 23326 17556 23378
rect 17500 23314 17556 23326
rect 17612 23380 17668 23390
rect 17724 23380 17780 24670
rect 18060 24610 18116 24622
rect 18060 24558 18062 24610
rect 18114 24558 18116 24610
rect 18060 24388 18116 24558
rect 18060 24322 18116 24332
rect 17836 23380 17892 23390
rect 17724 23378 17892 23380
rect 17724 23326 17838 23378
rect 17890 23326 17892 23378
rect 17724 23324 17892 23326
rect 17612 23286 17668 23324
rect 17836 23314 17892 23324
rect 17388 23156 17444 23166
rect 17388 23154 17556 23156
rect 17388 23102 17390 23154
rect 17442 23102 17556 23154
rect 17388 23100 17556 23102
rect 17388 23090 17444 23100
rect 17500 22820 17556 23100
rect 17500 22764 18004 22820
rect 17276 22260 17332 22270
rect 17948 22260 18004 22764
rect 17276 22258 17892 22260
rect 17276 22206 17278 22258
rect 17330 22206 17892 22258
rect 17276 22204 17892 22206
rect 17276 22194 17332 22204
rect 17500 21812 17556 21822
rect 17500 21718 17556 21756
rect 17724 21812 17780 21822
rect 17724 21718 17780 21756
rect 17836 21810 17892 22204
rect 17836 21758 17838 21810
rect 17890 21758 17892 21810
rect 17836 21746 17892 21758
rect 17948 21810 18004 22204
rect 18172 22148 18228 43652
rect 18172 22082 18228 22092
rect 17948 21758 17950 21810
rect 18002 21758 18004 21810
rect 17948 21746 18004 21758
rect 18284 19572 18340 74732
rect 19180 74338 19236 75516
rect 19404 74788 19460 76412
rect 19740 76402 19796 76412
rect 19628 75684 19684 75694
rect 19628 74788 19684 75628
rect 20076 75572 20132 76636
rect 20636 75908 20692 79200
rect 21084 76692 21140 76702
rect 21084 76598 21140 76636
rect 21308 76356 21364 79200
rect 21980 76692 22036 79200
rect 22652 77252 22708 79200
rect 22652 77196 23156 77252
rect 21980 76626 22036 76636
rect 21644 76356 21700 76366
rect 21308 76354 21700 76356
rect 21308 76302 21646 76354
rect 21698 76302 21700 76354
rect 21308 76300 21700 76302
rect 21644 76290 21700 76300
rect 20636 75842 20692 75852
rect 21532 75908 21588 75918
rect 21532 75814 21588 75852
rect 20300 75684 20356 75694
rect 20300 75590 20356 75628
rect 20076 75516 20244 75572
rect 19836 75292 20100 75302
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 19836 75226 20100 75236
rect 19852 74788 19908 74798
rect 19628 74786 19908 74788
rect 19628 74734 19854 74786
rect 19906 74734 19908 74786
rect 19628 74732 19908 74734
rect 20188 74788 20244 75516
rect 23100 75122 23156 77196
rect 23100 75070 23102 75122
rect 23154 75070 23156 75122
rect 23100 75058 23156 75070
rect 23324 75124 23380 79200
rect 23884 76466 23940 76478
rect 23884 76414 23886 76466
rect 23938 76414 23940 76466
rect 23660 75796 23716 75806
rect 23660 75682 23716 75740
rect 23660 75630 23662 75682
rect 23714 75630 23716 75682
rect 23548 75124 23604 75134
rect 23324 75122 23604 75124
rect 23324 75070 23550 75122
rect 23602 75070 23604 75122
rect 23324 75068 23604 75070
rect 23548 75058 23604 75068
rect 22764 74898 22820 74910
rect 22764 74846 22766 74898
rect 22818 74846 22820 74898
rect 20412 74788 20468 74798
rect 20188 74786 20468 74788
rect 20188 74734 20414 74786
rect 20466 74734 20468 74786
rect 20188 74732 20468 74734
rect 19404 74694 19460 74732
rect 19180 74286 19182 74338
rect 19234 74286 19236 74338
rect 19180 74274 19236 74286
rect 19852 73892 19908 74732
rect 20412 74722 20468 74732
rect 22764 74004 22820 74846
rect 22988 74004 23044 74014
rect 22764 74002 23044 74004
rect 22764 73950 22990 74002
rect 23042 73950 23044 74002
rect 22764 73948 23044 73950
rect 19628 73836 19908 73892
rect 19628 55468 19684 73836
rect 19836 73724 20100 73734
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 19836 73658 20100 73668
rect 19836 72156 20100 72166
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 19836 72090 20100 72100
rect 19836 70588 20100 70598
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 19836 70522 20100 70532
rect 19836 69020 20100 69030
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 19836 68954 20100 68964
rect 19836 67452 20100 67462
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 19836 67386 20100 67396
rect 19836 65884 20100 65894
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 19836 65818 20100 65828
rect 19836 64316 20100 64326
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 19836 64250 20100 64260
rect 19836 62748 20100 62758
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 19836 62682 20100 62692
rect 19836 61180 20100 61190
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 19836 61114 20100 61124
rect 19836 59612 20100 59622
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 19836 59546 20100 59556
rect 19836 58044 20100 58054
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 19836 57978 20100 57988
rect 19836 56476 20100 56486
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 19836 56410 20100 56420
rect 22988 55468 23044 73948
rect 19068 55412 19684 55468
rect 22428 55412 23044 55468
rect 18396 23380 18452 23390
rect 18396 23286 18452 23324
rect 18508 22820 18564 22830
rect 18508 21812 18564 22764
rect 18508 21718 18564 21756
rect 18844 22372 18900 22382
rect 18844 21586 18900 22316
rect 18844 21534 18846 21586
rect 18898 21534 18900 21586
rect 18620 20132 18676 20142
rect 17836 19516 18340 19572
rect 18396 20076 18620 20132
rect 17164 19180 17780 19236
rect 16940 17780 16996 17790
rect 16716 5572 16772 6188
rect 16828 8596 16884 8606
rect 16828 6018 16884 8540
rect 16940 7700 16996 17724
rect 17724 17780 17780 19180
rect 17836 18674 17892 19516
rect 17836 18622 17838 18674
rect 17890 18622 17892 18674
rect 17836 18610 17892 18622
rect 17948 19124 18004 19134
rect 17948 18562 18004 19068
rect 17948 18510 17950 18562
rect 18002 18510 18004 18562
rect 17948 18498 18004 18510
rect 17724 17686 17780 17724
rect 17836 18226 17892 18238
rect 17836 18174 17838 18226
rect 17890 18174 17892 18226
rect 17836 17444 17892 18174
rect 17836 17378 17892 17388
rect 18172 17778 18228 19516
rect 18172 17726 18174 17778
rect 18226 17726 18228 17778
rect 18172 15148 18228 17726
rect 17836 15092 18228 15148
rect 17276 12852 17332 12862
rect 17276 12850 17668 12852
rect 17276 12798 17278 12850
rect 17330 12798 17668 12850
rect 17276 12796 17668 12798
rect 17276 12786 17332 12796
rect 17612 12066 17668 12796
rect 17612 12014 17614 12066
rect 17666 12014 17668 12066
rect 17612 12002 17668 12014
rect 17724 12290 17780 12302
rect 17724 12238 17726 12290
rect 17778 12238 17780 12290
rect 17724 9156 17780 12238
rect 16940 7606 16996 7644
rect 17276 9100 17780 9156
rect 16828 5966 16830 6018
rect 16882 5966 16884 6018
rect 16828 5796 16884 5966
rect 16828 5730 16884 5740
rect 16716 5516 16884 5572
rect 16604 5282 16660 5292
rect 16716 5236 16772 5246
rect 16716 5142 16772 5180
rect 16492 5058 16548 5068
rect 15596 4508 15876 4564
rect 16044 4676 16100 4686
rect 15596 3666 15652 4508
rect 16044 4228 16100 4620
rect 16716 4564 16772 4574
rect 16828 4564 16884 5516
rect 16716 4562 16884 4564
rect 16716 4510 16718 4562
rect 16770 4510 16884 4562
rect 16716 4508 16884 4510
rect 16716 4498 16772 4508
rect 15708 4004 15764 4014
rect 15708 3778 15764 3948
rect 15708 3726 15710 3778
rect 15762 3726 15764 3778
rect 15708 3714 15764 3726
rect 15596 3614 15598 3666
rect 15650 3614 15652 3666
rect 15596 3602 15652 3614
rect 15372 3554 15428 3566
rect 15372 3502 15374 3554
rect 15426 3502 15428 3554
rect 15372 3332 15428 3502
rect 16044 3554 16100 4172
rect 16044 3502 16046 3554
rect 16098 3502 16100 3554
rect 16044 3490 16100 3502
rect 16268 4116 16324 4126
rect 15372 3266 15428 3276
rect 15260 2706 15316 2716
rect 15708 3108 15764 3118
rect 15708 800 15764 3052
rect 16268 1764 16324 4060
rect 17276 3666 17332 9100
rect 17724 8932 17780 8942
rect 17836 8932 17892 15092
rect 17948 12068 18004 12078
rect 17948 11974 18004 12012
rect 18396 11508 18452 20076
rect 18620 20038 18676 20076
rect 18844 18340 18900 21534
rect 19068 20242 19124 55412
rect 19836 54908 20100 54918
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 19836 54842 20100 54852
rect 19836 53340 20100 53350
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 19836 53274 20100 53284
rect 19836 51772 20100 51782
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 19836 51706 20100 51716
rect 19836 50204 20100 50214
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 19836 50138 20100 50148
rect 19836 48636 20100 48646
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 19836 48570 20100 48580
rect 19836 47068 20100 47078
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 19836 47002 20100 47012
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 20972 40516 21028 40526
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 20972 27972 21028 40460
rect 20972 27906 21028 27916
rect 22428 26908 22484 55412
rect 22204 26852 22484 26908
rect 23660 26908 23716 75630
rect 23884 75684 23940 76414
rect 23884 75236 23940 75628
rect 23996 75572 24052 79200
rect 24668 76692 24724 79200
rect 24892 76692 24948 76702
rect 24668 76690 24948 76692
rect 24668 76638 24894 76690
rect 24946 76638 24948 76690
rect 24668 76636 24948 76638
rect 25340 76692 25396 79200
rect 25564 76692 25620 76702
rect 25340 76690 25620 76692
rect 25340 76638 25566 76690
rect 25618 76638 25620 76690
rect 25340 76636 25620 76638
rect 26012 76692 26068 79200
rect 26236 76692 26292 76702
rect 26012 76690 26292 76692
rect 26012 76638 26238 76690
rect 26290 76638 26292 76690
rect 26012 76636 26292 76638
rect 26684 76692 26740 79200
rect 26908 76692 26964 76702
rect 26684 76690 26964 76692
rect 26684 76638 26910 76690
rect 26962 76638 26964 76690
rect 26684 76636 26964 76638
rect 27356 76692 27412 79200
rect 28028 77924 28084 79200
rect 28028 77868 28420 77924
rect 27580 76692 27636 76702
rect 27356 76690 27636 76692
rect 27356 76638 27582 76690
rect 27634 76638 27636 76690
rect 27356 76636 27636 76638
rect 24892 76626 24948 76636
rect 25564 76626 25620 76636
rect 26236 76626 26292 76636
rect 26908 76626 26964 76636
rect 27580 76626 27636 76636
rect 28364 76690 28420 77868
rect 28364 76638 28366 76690
rect 28418 76638 28420 76690
rect 28364 76626 28420 76638
rect 28700 76692 28756 79200
rect 28924 76692 28980 76702
rect 28700 76690 28980 76692
rect 28700 76638 28926 76690
rect 28978 76638 28980 76690
rect 28700 76636 28980 76638
rect 29372 76692 29428 79200
rect 29596 76692 29652 76702
rect 29372 76690 29652 76692
rect 29372 76638 29598 76690
rect 29650 76638 29652 76690
rect 29372 76636 29652 76638
rect 30044 76692 30100 79200
rect 30268 76692 30324 76702
rect 30044 76690 30324 76692
rect 30044 76638 30270 76690
rect 30322 76638 30324 76690
rect 30044 76636 30324 76638
rect 30716 76692 30772 79200
rect 30940 76692 30996 76702
rect 30716 76690 30996 76692
rect 30716 76638 30942 76690
rect 30994 76638 30996 76690
rect 30716 76636 30996 76638
rect 31388 76692 31444 79200
rect 31500 76692 31556 76702
rect 31388 76690 31556 76692
rect 31388 76638 31502 76690
rect 31554 76638 31556 76690
rect 31388 76636 31556 76638
rect 32060 76692 32116 79200
rect 32284 76692 32340 76702
rect 32060 76690 32340 76692
rect 32060 76638 32286 76690
rect 32338 76638 32340 76690
rect 32060 76636 32340 76638
rect 28924 76626 28980 76636
rect 29596 76626 29652 76636
rect 30268 76626 30324 76636
rect 30940 76626 30996 76636
rect 31500 76626 31556 76636
rect 32284 76626 32340 76636
rect 31836 76356 31892 76366
rect 24780 75796 24836 75806
rect 24780 75702 24836 75740
rect 25228 75684 25284 75694
rect 25228 75590 25284 75628
rect 30156 75684 30212 75694
rect 24220 75572 24276 75582
rect 23996 75570 24276 75572
rect 23996 75518 24222 75570
rect 24274 75518 24276 75570
rect 23996 75516 24276 75518
rect 24220 75506 24276 75516
rect 23884 75180 24164 75236
rect 23660 26852 23940 26908
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 21084 24892 21476 24948
rect 19740 24834 19796 24846
rect 19740 24782 19742 24834
rect 19794 24782 19796 24834
rect 19628 24724 19684 24734
rect 19516 24722 19684 24724
rect 19516 24670 19630 24722
rect 19682 24670 19684 24722
rect 19516 24668 19684 24670
rect 19292 24612 19348 24622
rect 19292 24518 19348 24556
rect 19292 23492 19348 23502
rect 19516 23492 19572 24668
rect 19628 24658 19684 24668
rect 19740 24724 19796 24782
rect 20972 24836 21028 24846
rect 21084 24836 21140 24892
rect 20972 24834 21140 24836
rect 20972 24782 20974 24834
rect 21026 24782 21140 24834
rect 20972 24780 21140 24782
rect 20972 24770 21028 24780
rect 19740 24658 19796 24668
rect 20300 24724 20356 24734
rect 20300 24630 20356 24668
rect 21196 24724 21252 24734
rect 19740 24500 19796 24510
rect 19740 24406 19796 24444
rect 19628 24052 19684 24062
rect 19964 24052 20020 24062
rect 19628 24050 20020 24052
rect 19628 23998 19630 24050
rect 19682 23998 19966 24050
rect 20018 23998 20020 24050
rect 19628 23996 20020 23998
rect 19628 23986 19684 23996
rect 19964 23986 20020 23996
rect 21196 23940 21252 24668
rect 21420 24050 21476 24892
rect 21420 23998 21422 24050
rect 21474 23998 21476 24050
rect 21420 23986 21476 23998
rect 21868 24500 21924 24510
rect 20300 23826 20356 23838
rect 20300 23774 20302 23826
rect 20354 23774 20356 23826
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19348 23436 19684 23492
rect 19836 23482 20100 23492
rect 20300 23492 20356 23774
rect 19292 23378 19348 23436
rect 19292 23326 19294 23378
rect 19346 23326 19348 23378
rect 19292 23314 19348 23326
rect 19628 23380 19684 23436
rect 20300 23426 20356 23436
rect 21196 23380 21252 23884
rect 21868 23938 21924 24444
rect 21868 23886 21870 23938
rect 21922 23886 21924 23938
rect 21868 23874 21924 23886
rect 21308 23716 21364 23726
rect 21308 23714 21476 23716
rect 21308 23662 21310 23714
rect 21362 23662 21476 23714
rect 21308 23660 21476 23662
rect 21308 23650 21364 23660
rect 21420 23380 21476 23660
rect 21532 23714 21588 23726
rect 21532 23662 21534 23714
rect 21586 23662 21588 23714
rect 21532 23604 21588 23662
rect 21532 23538 21588 23548
rect 21868 23380 21924 23390
rect 19628 23324 20020 23380
rect 21196 23324 21364 23380
rect 19964 23266 20020 23324
rect 19964 23214 19966 23266
rect 20018 23214 20020 23266
rect 19964 23202 20020 23214
rect 20076 23266 20132 23278
rect 20076 23214 20078 23266
rect 20130 23214 20132 23266
rect 19516 23156 19572 23166
rect 19068 20190 19070 20242
rect 19122 20190 19124 20242
rect 19068 20132 19124 20190
rect 18620 18338 18900 18340
rect 18620 18286 18846 18338
rect 18898 18286 18900 18338
rect 18620 18284 18900 18286
rect 18620 16882 18676 18284
rect 18844 18274 18900 18284
rect 18956 20020 19012 20030
rect 19068 20020 19124 20076
rect 19292 23154 19572 23156
rect 19292 23102 19518 23154
rect 19570 23102 19572 23154
rect 19292 23100 19572 23102
rect 19068 19964 19236 20020
rect 18956 19124 19012 19964
rect 19068 19796 19124 19806
rect 19068 19702 19124 19740
rect 19068 19124 19124 19134
rect 19012 19122 19124 19124
rect 19012 19070 19070 19122
rect 19122 19070 19124 19122
rect 19012 19068 19124 19070
rect 18732 17780 18788 17790
rect 18732 17444 18788 17724
rect 18844 17668 18900 17678
rect 18956 17668 19012 19068
rect 19068 19058 19124 19068
rect 19180 18900 19236 19964
rect 19292 19684 19348 23100
rect 19516 23090 19572 23100
rect 20076 23044 20132 23214
rect 20300 23156 20356 23166
rect 20300 23154 20468 23156
rect 20300 23102 20302 23154
rect 20354 23102 20468 23154
rect 20300 23100 20468 23102
rect 20300 23090 20356 23100
rect 19852 22988 20076 23044
rect 19404 22484 19460 22494
rect 19740 22484 19796 22494
rect 19404 22482 19796 22484
rect 19404 22430 19406 22482
rect 19458 22430 19742 22482
rect 19794 22430 19796 22482
rect 19404 22428 19796 22430
rect 19404 22418 19460 22428
rect 19740 22418 19796 22428
rect 19852 22148 19908 22988
rect 20076 22950 20132 22988
rect 20412 22930 20468 23100
rect 21196 23154 21252 23166
rect 21196 23102 21198 23154
rect 21250 23102 21252 23154
rect 20636 23044 20692 23054
rect 20636 22950 20692 22988
rect 21196 23042 21252 23102
rect 21196 22990 21198 23042
rect 21250 22990 21252 23042
rect 21196 22978 21252 22990
rect 20412 22878 20414 22930
rect 20466 22878 20468 22930
rect 20412 22866 20468 22878
rect 20076 22820 20132 22830
rect 20076 22482 20132 22764
rect 20076 22430 20078 22482
rect 20130 22430 20132 22482
rect 20076 22418 20132 22430
rect 20412 22708 20468 22718
rect 20412 22260 20468 22652
rect 21308 22372 21364 23324
rect 21420 23378 21924 23380
rect 21420 23326 21870 23378
rect 21922 23326 21924 23378
rect 21420 23324 21924 23326
rect 21420 22708 21476 23324
rect 21868 23314 21924 23324
rect 21420 22642 21476 22652
rect 21644 23154 21700 23166
rect 21644 23102 21646 23154
rect 21698 23102 21700 23154
rect 21644 22708 21700 23102
rect 21644 22642 21700 22652
rect 21756 23042 21812 23054
rect 21756 22990 21758 23042
rect 21810 22990 21812 23042
rect 21756 22484 21812 22990
rect 22092 22484 22148 22494
rect 21756 22482 22148 22484
rect 21756 22430 22094 22482
rect 22146 22430 22148 22482
rect 21756 22428 22148 22430
rect 22092 22418 22148 22428
rect 20412 22166 20468 22204
rect 21196 22370 21364 22372
rect 21196 22318 21310 22370
rect 21362 22318 21364 22370
rect 21196 22316 21364 22318
rect 19852 22082 19908 22092
rect 20748 22146 20804 22158
rect 20748 22094 20750 22146
rect 20802 22094 20804 22146
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 19628 21476 19684 21486
rect 19516 21474 19684 21476
rect 19516 21422 19630 21474
rect 19682 21422 19684 21474
rect 19516 21420 19684 21422
rect 19516 20914 19572 21420
rect 19628 21410 19684 21420
rect 19516 20862 19518 20914
rect 19570 20862 19572 20914
rect 19516 20850 19572 20862
rect 20076 20802 20132 20814
rect 20076 20750 20078 20802
rect 20130 20750 20132 20802
rect 19292 19234 19348 19628
rect 19404 20578 19460 20590
rect 19404 20526 19406 20578
rect 19458 20526 19460 20578
rect 19404 19348 19460 20526
rect 19628 20580 19684 20590
rect 20076 20580 20132 20750
rect 20524 20580 20580 20590
rect 20076 20524 20244 20580
rect 19628 20486 19684 20524
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 19852 20244 19908 20254
rect 20188 20244 20244 20524
rect 19852 20242 20244 20244
rect 19852 20190 19854 20242
rect 19906 20190 20244 20242
rect 19852 20188 20244 20190
rect 19852 20178 19908 20188
rect 19628 20130 19684 20142
rect 19628 20078 19630 20130
rect 19682 20078 19684 20130
rect 19516 20020 19572 20030
rect 19516 19926 19572 19964
rect 19628 19908 19684 20078
rect 20300 20132 20356 20142
rect 20188 20020 20244 20030
rect 20300 20020 20356 20076
rect 20188 20018 20356 20020
rect 20188 19966 20190 20018
rect 20242 19966 20356 20018
rect 20188 19964 20356 19966
rect 20188 19954 20244 19964
rect 20524 19908 20580 20524
rect 20748 20132 20804 22094
rect 20748 20066 20804 20076
rect 20972 19908 21028 19918
rect 20524 19852 20972 19908
rect 21196 19908 21252 22316
rect 21308 22306 21364 22316
rect 21756 21476 21812 21486
rect 21308 21474 21812 21476
rect 21308 21422 21758 21474
rect 21810 21422 21812 21474
rect 21308 21420 21812 21422
rect 21308 20130 21364 21420
rect 21756 21410 21812 21420
rect 21308 20078 21310 20130
rect 21362 20078 21364 20130
rect 21308 20066 21364 20078
rect 21756 20132 21812 20142
rect 21644 20018 21700 20030
rect 21644 19966 21646 20018
rect 21698 19966 21700 20018
rect 21644 19908 21700 19966
rect 21196 19852 21700 19908
rect 19628 19842 19684 19852
rect 20972 19814 21028 19852
rect 19404 19292 19684 19348
rect 19292 19182 19294 19234
rect 19346 19182 19348 19234
rect 19292 19170 19348 19182
rect 19628 19124 19684 19292
rect 18844 17666 19012 17668
rect 18844 17614 18846 17666
rect 18898 17614 19012 17666
rect 18844 17612 19012 17614
rect 19068 18844 19236 18900
rect 19516 19012 19572 19022
rect 18844 17602 18900 17612
rect 18956 17444 19012 17454
rect 18732 17442 19012 17444
rect 18732 17390 18958 17442
rect 19010 17390 19012 17442
rect 18732 17388 19012 17390
rect 18956 17378 19012 17388
rect 18620 16830 18622 16882
rect 18674 16830 18676 16882
rect 18620 13636 18676 16830
rect 19068 15148 19124 18844
rect 19516 18228 19572 18956
rect 19628 18676 19684 19068
rect 21532 19124 21588 19134
rect 21532 19030 21588 19068
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 21532 18788 21588 18798
rect 19628 18620 20020 18676
rect 19180 18172 19572 18228
rect 19180 17666 19236 18172
rect 19852 17668 19908 17678
rect 19180 17614 19182 17666
rect 19234 17614 19236 17666
rect 19180 17602 19236 17614
rect 19628 17666 19908 17668
rect 19628 17614 19854 17666
rect 19906 17614 19908 17666
rect 19628 17612 19908 17614
rect 19516 17554 19572 17566
rect 19516 17502 19518 17554
rect 19570 17502 19572 17554
rect 19404 17444 19460 17454
rect 19516 17444 19572 17502
rect 19460 17388 19572 17444
rect 19404 17378 19460 17388
rect 19628 17108 19684 17612
rect 19852 17602 19908 17612
rect 19964 17666 20020 18620
rect 19964 17614 19966 17666
rect 20018 17614 20020 17666
rect 19964 17602 20020 17614
rect 21308 17554 21364 17566
rect 21308 17502 21310 17554
rect 21362 17502 21364 17554
rect 19740 17444 19796 17482
rect 19740 17378 19796 17388
rect 20412 17444 20468 17454
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 20412 17220 20468 17388
rect 20412 17154 20468 17164
rect 19292 17052 19684 17108
rect 19292 16994 19348 17052
rect 19292 16942 19294 16994
rect 19346 16942 19348 16994
rect 19292 16930 19348 16942
rect 21308 16772 21364 17502
rect 21420 16772 21476 16782
rect 21308 16770 21476 16772
rect 21308 16718 21422 16770
rect 21474 16718 21476 16770
rect 21308 16716 21476 16718
rect 21420 16706 21476 16716
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 18620 13570 18676 13580
rect 18732 15092 19124 15148
rect 18060 11506 18452 11508
rect 18060 11454 18398 11506
rect 18450 11454 18452 11506
rect 18060 11452 18452 11454
rect 18060 9268 18116 11452
rect 18396 11442 18452 11452
rect 18620 11172 18676 11182
rect 18508 11116 18620 11172
rect 18172 10722 18228 10734
rect 18172 10670 18174 10722
rect 18226 10670 18228 10722
rect 18172 9492 18228 10670
rect 18396 10724 18452 10734
rect 18508 10724 18564 11116
rect 18620 11106 18676 11116
rect 18396 10722 18564 10724
rect 18396 10670 18398 10722
rect 18450 10670 18564 10722
rect 18396 10668 18564 10670
rect 18396 10658 18452 10668
rect 18284 10500 18340 10510
rect 18284 10406 18340 10444
rect 18172 9436 18452 9492
rect 18284 9268 18340 9278
rect 18060 9212 18284 9268
rect 18284 9174 18340 9212
rect 17724 8930 17892 8932
rect 17724 8878 17726 8930
rect 17778 8878 17892 8930
rect 17724 8876 17892 8878
rect 18060 9042 18116 9054
rect 18060 8990 18062 9042
rect 18114 8990 18116 9042
rect 17612 8372 17668 8382
rect 17724 8372 17780 8876
rect 17612 8370 17780 8372
rect 17612 8318 17614 8370
rect 17666 8318 17780 8370
rect 17612 8316 17780 8318
rect 17612 8306 17668 8316
rect 17724 8260 17780 8316
rect 17724 8194 17780 8204
rect 18060 8034 18116 8990
rect 18172 8932 18228 8942
rect 18172 8838 18228 8876
rect 18172 8372 18228 8382
rect 18172 8278 18228 8316
rect 18284 8260 18340 8270
rect 18284 8166 18340 8204
rect 18060 7982 18062 8034
rect 18114 7982 18116 8034
rect 17836 7700 17892 7710
rect 17724 7476 17780 7486
rect 17724 7382 17780 7420
rect 17724 7028 17780 7038
rect 17612 6972 17724 7028
rect 17388 5908 17444 5946
rect 17388 5842 17444 5852
rect 17388 5682 17444 5694
rect 17388 5630 17390 5682
rect 17442 5630 17444 5682
rect 17388 5236 17444 5630
rect 17612 5684 17668 6972
rect 17724 6962 17780 6972
rect 17836 6802 17892 7644
rect 17836 6750 17838 6802
rect 17890 6750 17892 6802
rect 17836 6738 17892 6750
rect 18060 7588 18116 7982
rect 18396 7812 18452 9436
rect 18732 9380 18788 15092
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 19628 13746 19684 13758
rect 21420 13748 21476 13758
rect 19628 13694 19630 13746
rect 19682 13694 19684 13746
rect 19628 13636 19684 13694
rect 21308 13692 21420 13748
rect 19628 13570 19684 13580
rect 20412 13636 20468 13646
rect 20412 13634 20580 13636
rect 20412 13582 20414 13634
rect 20466 13582 20580 13634
rect 20412 13580 20580 13582
rect 20412 13570 20468 13580
rect 19180 13244 20020 13300
rect 19180 12402 19236 13244
rect 19516 13074 19572 13086
rect 19516 13022 19518 13074
rect 19570 13022 19572 13074
rect 19516 12964 19572 13022
rect 19516 12898 19572 12908
rect 19964 12962 20020 13244
rect 19964 12910 19966 12962
rect 20018 12910 20020 12962
rect 19964 12898 20020 12910
rect 20076 12964 20132 12974
rect 20076 12962 20356 12964
rect 20076 12910 20078 12962
rect 20130 12910 20356 12962
rect 20076 12908 20356 12910
rect 20076 12898 20132 12908
rect 20188 12740 20244 12750
rect 20188 12646 20244 12684
rect 19836 12572 20100 12582
rect 19516 12516 19572 12526
rect 19180 12350 19182 12402
rect 19234 12350 19236 12402
rect 19180 11788 19236 12350
rect 19404 12460 19516 12516
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20300 12516 20356 12908
rect 19836 12506 20100 12516
rect 19404 12402 19460 12460
rect 19516 12450 19572 12460
rect 20188 12460 20356 12516
rect 20412 12738 20468 12750
rect 20412 12686 20414 12738
rect 20466 12686 20468 12738
rect 19404 12350 19406 12402
rect 19458 12350 19460 12402
rect 19404 12338 19460 12350
rect 19852 12292 19908 12302
rect 19852 12180 19908 12236
rect 20076 12292 20132 12302
rect 20188 12292 20244 12460
rect 20076 12290 20244 12292
rect 20076 12238 20078 12290
rect 20130 12238 20244 12290
rect 20076 12236 20244 12238
rect 20300 12290 20356 12302
rect 20300 12238 20302 12290
rect 20354 12238 20356 12290
rect 20076 12226 20132 12236
rect 19852 12178 20020 12180
rect 19852 12126 19854 12178
rect 19906 12126 20020 12178
rect 19852 12124 20020 12126
rect 19852 12114 19908 12124
rect 19292 12068 19348 12078
rect 19292 11974 19348 12012
rect 19964 11844 20020 12124
rect 20300 11844 20356 12238
rect 20412 12292 20468 12686
rect 20412 12226 20468 12236
rect 20412 12068 20468 12078
rect 20524 12068 20580 13580
rect 20972 12964 21028 12974
rect 20972 12402 21028 12908
rect 20972 12350 20974 12402
rect 21026 12350 21028 12402
rect 20972 12338 21028 12350
rect 20412 12066 20580 12068
rect 20412 12014 20414 12066
rect 20466 12014 20580 12066
rect 20412 12012 20580 12014
rect 20412 12002 20468 12012
rect 19964 11788 20244 11844
rect 19180 11732 19684 11788
rect 19068 11396 19124 11406
rect 18956 11340 19068 11396
rect 18732 9314 18788 9324
rect 18844 10610 18900 10622
rect 18844 10558 18846 10610
rect 18898 10558 18900 10610
rect 18396 7746 18452 7756
rect 18732 9042 18788 9054
rect 18732 8990 18734 9042
rect 18786 8990 18788 9042
rect 18732 8258 18788 8990
rect 18844 9044 18900 10558
rect 18844 8978 18900 8988
rect 18732 8206 18734 8258
rect 18786 8206 18788 8258
rect 18620 7700 18676 7710
rect 18508 7698 18676 7700
rect 18508 7646 18622 7698
rect 18674 7646 18676 7698
rect 18508 7644 18676 7646
rect 18732 7700 18788 8206
rect 18844 7700 18900 7710
rect 18732 7698 18900 7700
rect 18732 7646 18846 7698
rect 18898 7646 18900 7698
rect 18732 7644 18900 7646
rect 18396 7588 18452 7598
rect 18060 7586 18452 7588
rect 18060 7534 18062 7586
rect 18114 7534 18398 7586
rect 18450 7534 18452 7586
rect 18060 7532 18452 7534
rect 18060 6130 18116 7532
rect 18396 7522 18452 7532
rect 18508 7588 18564 7644
rect 18620 7634 18676 7644
rect 18508 7522 18564 7532
rect 18508 7364 18564 7374
rect 18508 7270 18564 7308
rect 18844 6692 18900 7644
rect 18956 6804 19012 11340
rect 19068 11330 19124 11340
rect 19628 11394 19684 11732
rect 19628 11342 19630 11394
rect 19682 11342 19684 11394
rect 19516 10500 19572 10510
rect 19516 10406 19572 10444
rect 19180 9268 19236 9278
rect 19180 9174 19236 9212
rect 19628 9268 19684 11342
rect 19852 11508 19908 11518
rect 19852 11394 19908 11452
rect 19852 11342 19854 11394
rect 19906 11342 19908 11394
rect 19852 11330 19908 11342
rect 20188 11396 20244 11788
rect 20300 11778 20356 11788
rect 20636 11508 20692 11518
rect 20636 11414 20692 11452
rect 20188 11394 20468 11396
rect 20188 11342 20190 11394
rect 20242 11342 20468 11394
rect 20188 11340 20468 11342
rect 20188 11330 20244 11340
rect 19740 11172 19796 11210
rect 19740 11106 19796 11116
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 20188 9940 20244 9950
rect 20188 9826 20244 9884
rect 20188 9774 20190 9826
rect 20242 9774 20244 9826
rect 20188 9762 20244 9774
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 19628 9202 19684 9212
rect 19516 9044 19572 9054
rect 19516 8950 19572 8988
rect 19180 8932 19236 8942
rect 19068 8372 19124 8382
rect 19180 8372 19236 8876
rect 20300 8932 20356 8942
rect 20300 8838 20356 8876
rect 19292 8484 19348 8494
rect 19292 8482 19908 8484
rect 19292 8430 19294 8482
rect 19346 8430 19908 8482
rect 19292 8428 19908 8430
rect 19292 8418 19348 8428
rect 19068 8370 19236 8372
rect 19068 8318 19070 8370
rect 19122 8318 19236 8370
rect 19068 8316 19236 8318
rect 19852 8370 19908 8428
rect 19852 8318 19854 8370
rect 19906 8318 19908 8370
rect 19068 8306 19124 8316
rect 19852 8306 19908 8318
rect 19964 8372 20020 8382
rect 19964 8258 20020 8316
rect 20412 8260 20468 11340
rect 20972 10276 21028 10286
rect 20748 9940 20804 9950
rect 20748 9846 20804 9884
rect 20636 8820 20692 8830
rect 19964 8206 19966 8258
rect 20018 8206 20020 8258
rect 19964 8194 20020 8206
rect 20188 8258 20468 8260
rect 20188 8206 20414 8258
rect 20466 8206 20468 8258
rect 20188 8204 20468 8206
rect 19292 8148 19348 8158
rect 19068 8034 19124 8046
rect 19068 7982 19070 8034
rect 19122 7982 19124 8034
rect 19068 7028 19124 7982
rect 19068 6962 19124 6972
rect 19180 7812 19236 7822
rect 18956 6748 19124 6804
rect 18508 6356 18564 6366
rect 18060 6078 18062 6130
rect 18114 6078 18116 6130
rect 18060 6066 18116 6078
rect 18284 6132 18340 6142
rect 18284 6038 18340 6076
rect 18396 6020 18452 6030
rect 17724 5908 17780 5918
rect 18172 5908 18228 5918
rect 17724 5906 18228 5908
rect 17724 5854 17726 5906
rect 17778 5854 18174 5906
rect 18226 5854 18228 5906
rect 17724 5852 18228 5854
rect 17724 5842 17780 5852
rect 18172 5842 18228 5852
rect 17612 5628 17892 5684
rect 17388 5170 17444 5180
rect 17836 4562 17892 5628
rect 18284 5348 18340 5358
rect 17836 4510 17838 4562
rect 17890 4510 17892 4562
rect 17836 4498 17892 4510
rect 17948 5012 18004 5022
rect 17724 4452 17780 4462
rect 17612 4340 17668 4350
rect 17276 3614 17278 3666
rect 17330 3614 17332 3666
rect 17276 3602 17332 3614
rect 17388 4338 17668 4340
rect 17388 4286 17614 4338
rect 17666 4286 17668 4338
rect 17388 4284 17668 4286
rect 17052 3556 17108 3566
rect 16380 3330 16436 3342
rect 16380 3278 16382 3330
rect 16434 3278 16436 3330
rect 16380 2772 16436 3278
rect 16380 2706 16436 2716
rect 16268 1708 16436 1764
rect 16380 800 16436 1708
rect 17052 800 17108 3500
rect 17276 3330 17332 3342
rect 17276 3278 17278 3330
rect 17330 3278 17332 3330
rect 17276 2324 17332 3278
rect 17388 3220 17444 4284
rect 17612 4274 17668 4284
rect 17500 4116 17556 4126
rect 17500 3778 17556 4060
rect 17500 3726 17502 3778
rect 17554 3726 17556 3778
rect 17500 3714 17556 3726
rect 17388 3154 17444 3164
rect 17276 2258 17332 2268
rect 17724 800 17780 4396
rect 17948 4450 18004 4956
rect 17948 4398 17950 4450
rect 18002 4398 18004 4450
rect 17948 4116 18004 4398
rect 18284 4452 18340 5292
rect 18284 4358 18340 4396
rect 18396 4228 18452 5964
rect 17948 4050 18004 4060
rect 18172 4172 18452 4228
rect 17836 4004 17892 4014
rect 17836 3442 17892 3948
rect 17836 3390 17838 3442
rect 17890 3390 17892 3442
rect 17836 3378 17892 3390
rect 18172 3442 18228 4172
rect 18172 3390 18174 3442
rect 18226 3390 18228 3442
rect 18172 3378 18228 3390
rect 18396 3780 18452 3790
rect 18396 800 18452 3724
rect 18508 3556 18564 6300
rect 18620 5908 18676 5918
rect 18620 4562 18676 5852
rect 18732 5908 18788 5918
rect 18844 5908 18900 6636
rect 18956 6468 19012 6478
rect 18956 6374 19012 6412
rect 18732 5906 18900 5908
rect 18732 5854 18734 5906
rect 18786 5854 18900 5906
rect 18732 5852 18900 5854
rect 18732 5842 18788 5852
rect 18732 5236 18788 5246
rect 18956 5236 19012 5246
rect 18788 5234 19012 5236
rect 18788 5182 18958 5234
rect 19010 5182 19012 5234
rect 18788 5180 19012 5182
rect 18732 5170 18788 5180
rect 18956 5170 19012 5180
rect 18620 4510 18622 4562
rect 18674 4510 18676 4562
rect 18620 4498 18676 4510
rect 18956 4340 19012 4350
rect 18956 4246 19012 4284
rect 19068 4226 19124 6748
rect 19180 6020 19236 7756
rect 19292 7698 19348 8092
rect 19740 8148 19796 8158
rect 19740 8054 19796 8092
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19292 7646 19294 7698
rect 19346 7646 19348 7698
rect 19292 7634 19348 7646
rect 19964 7700 20020 7710
rect 19628 7476 19684 7486
rect 19684 7420 19796 7476
rect 19628 7382 19684 7420
rect 19516 7140 19572 7150
rect 19404 6468 19460 6478
rect 19404 6374 19460 6412
rect 19516 6020 19572 7084
rect 19628 6692 19684 6702
rect 19740 6692 19796 7420
rect 19852 6692 19908 6702
rect 19740 6636 19852 6692
rect 19628 6578 19684 6636
rect 19852 6626 19908 6636
rect 19964 6690 20020 7644
rect 20076 7700 20132 7710
rect 20188 7700 20244 8204
rect 20412 8194 20468 8204
rect 20524 8764 20636 8820
rect 20076 7698 20244 7700
rect 20076 7646 20078 7698
rect 20130 7646 20244 7698
rect 20076 7644 20244 7646
rect 20412 7700 20468 7710
rect 20076 7634 20132 7644
rect 20412 7606 20468 7644
rect 19964 6638 19966 6690
rect 20018 6638 20020 6690
rect 19628 6526 19630 6578
rect 19682 6526 19684 6578
rect 19628 6514 19684 6526
rect 19964 6468 20020 6638
rect 19964 6402 20020 6412
rect 20188 6916 20244 6926
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 19180 5964 19460 6020
rect 19516 5964 19796 6020
rect 19404 5908 19460 5964
rect 19404 5852 19572 5908
rect 19068 4174 19070 4226
rect 19122 4174 19124 4226
rect 19068 4162 19124 4174
rect 19180 5794 19236 5806
rect 19180 5742 19182 5794
rect 19234 5742 19236 5794
rect 18508 3490 18564 3500
rect 18620 4116 18676 4126
rect 18620 3554 18676 4060
rect 19180 4116 19236 5742
rect 19404 5348 19460 5358
rect 19292 5292 19404 5348
rect 19292 4564 19348 5292
rect 19404 5282 19460 5292
rect 19516 5234 19572 5852
rect 19628 5796 19684 5806
rect 19628 5702 19684 5740
rect 19516 5182 19518 5234
rect 19570 5182 19572 5234
rect 19516 5170 19572 5182
rect 19404 5124 19460 5134
rect 19404 5030 19460 5068
rect 19740 5122 19796 5964
rect 19740 5070 19742 5122
rect 19794 5070 19796 5122
rect 19740 5058 19796 5070
rect 20076 5794 20132 5806
rect 20076 5742 20078 5794
rect 20130 5742 20132 5794
rect 20076 5124 20132 5742
rect 20076 5058 20132 5068
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 19628 4564 19684 4574
rect 19292 4562 19684 4564
rect 19292 4510 19630 4562
rect 19682 4510 19684 4562
rect 19292 4508 19684 4510
rect 19292 4450 19348 4508
rect 19628 4498 19684 4508
rect 19964 4564 20020 4574
rect 19292 4398 19294 4450
rect 19346 4398 19348 4450
rect 19292 4386 19348 4398
rect 19964 4450 20020 4508
rect 19964 4398 19966 4450
rect 20018 4398 20020 4450
rect 19964 4386 20020 4398
rect 19404 4340 19460 4350
rect 19404 4228 19460 4284
rect 19180 4050 19236 4060
rect 19292 4172 19460 4228
rect 18620 3502 18622 3554
rect 18674 3502 18676 3554
rect 18620 2994 18676 3502
rect 19068 3892 19124 3902
rect 18844 3332 18900 3342
rect 18844 3238 18900 3276
rect 18620 2942 18622 2994
rect 18674 2942 18676 2994
rect 18620 2930 18676 2942
rect 19068 800 19124 3836
rect 19180 3556 19236 3566
rect 19292 3556 19348 4172
rect 19964 4116 20020 4126
rect 19236 3500 19348 3556
rect 19404 3668 19460 3678
rect 19180 3462 19236 3500
rect 19404 980 19460 3612
rect 19964 3668 20020 4060
rect 19516 3556 19572 3566
rect 19516 3442 19572 3500
rect 19964 3554 20020 3612
rect 19964 3502 19966 3554
rect 20018 3502 20020 3554
rect 19964 3490 20020 3502
rect 19516 3390 19518 3442
rect 19570 3390 19572 3442
rect 19516 3378 19572 3390
rect 20188 3442 20244 6860
rect 20524 6020 20580 8764
rect 20636 8754 20692 8764
rect 20300 5964 20580 6020
rect 20636 8484 20692 8494
rect 20300 4564 20356 5964
rect 20524 5794 20580 5806
rect 20524 5742 20526 5794
rect 20578 5742 20580 5794
rect 20412 5460 20468 5470
rect 20412 5122 20468 5404
rect 20412 5070 20414 5122
rect 20466 5070 20468 5122
rect 20412 5058 20468 5070
rect 20300 4450 20356 4508
rect 20300 4398 20302 4450
rect 20354 4398 20356 4450
rect 20300 4386 20356 4398
rect 20412 4452 20468 4462
rect 20188 3390 20190 3442
rect 20242 3390 20244 3442
rect 20188 3378 20244 3390
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 19404 924 19796 980
rect 19740 800 19796 924
rect 20412 800 20468 4396
rect 20524 4004 20580 5742
rect 20636 5234 20692 8428
rect 20748 8372 20804 8382
rect 20748 8278 20804 8316
rect 20860 7700 20916 7710
rect 20860 7606 20916 7644
rect 20972 6916 21028 10220
rect 20972 6850 21028 6860
rect 20860 6466 20916 6478
rect 20860 6414 20862 6466
rect 20914 6414 20916 6466
rect 20748 5348 20804 5358
rect 20748 5254 20804 5292
rect 20636 5182 20638 5234
rect 20690 5182 20692 5234
rect 20636 5170 20692 5182
rect 20636 4564 20692 4574
rect 20636 4470 20692 4508
rect 20860 4452 20916 6414
rect 21308 6244 21364 13692
rect 21420 13682 21476 13692
rect 21420 13076 21476 13086
rect 21420 12740 21476 13020
rect 21420 12674 21476 12684
rect 21532 11508 21588 18732
rect 21644 17780 21700 19852
rect 21756 19236 21812 20076
rect 21756 19142 21812 19180
rect 22092 19796 22148 19806
rect 22092 19234 22148 19740
rect 22092 19182 22094 19234
rect 22146 19182 22148 19234
rect 22092 19170 22148 19182
rect 22204 18452 22260 26852
rect 23100 24612 23156 24622
rect 23436 24612 23492 24622
rect 23100 24610 23492 24612
rect 23100 24558 23102 24610
rect 23154 24558 23438 24610
rect 23490 24558 23492 24610
rect 23100 24556 23492 24558
rect 23100 24546 23156 24556
rect 23436 24546 23492 24556
rect 23772 24610 23828 24622
rect 23772 24558 23774 24610
rect 23826 24558 23828 24610
rect 23100 24052 23156 24062
rect 23156 23996 23604 24052
rect 23100 23958 23156 23996
rect 23548 23826 23604 23996
rect 23548 23774 23550 23826
rect 23602 23774 23604 23826
rect 23548 23762 23604 23774
rect 23660 23826 23716 23838
rect 23660 23774 23662 23826
rect 23714 23774 23716 23826
rect 22316 23714 22372 23726
rect 22316 23662 22318 23714
rect 22370 23662 22372 23714
rect 22316 23604 22372 23662
rect 23324 23716 23380 23726
rect 23324 23622 23380 23660
rect 22316 23538 22372 23548
rect 23660 23380 23716 23774
rect 23772 23604 23828 24558
rect 23772 23538 23828 23548
rect 23884 23380 23940 26852
rect 23996 23940 24052 23950
rect 23996 23846 24052 23884
rect 23660 23314 23716 23324
rect 23772 23324 23940 23380
rect 23996 23380 24052 23390
rect 23548 23156 23604 23166
rect 23548 23062 23604 23100
rect 22988 20578 23044 20590
rect 22988 20526 22990 20578
rect 23042 20526 23044 20578
rect 22428 20468 22484 20478
rect 22316 20412 22428 20468
rect 22316 19236 22372 20412
rect 22428 20402 22484 20412
rect 22988 20468 23044 20526
rect 22988 20402 23044 20412
rect 23436 20580 23492 20590
rect 22428 19908 22484 19918
rect 22428 19906 22708 19908
rect 22428 19854 22430 19906
rect 22482 19854 22708 19906
rect 22428 19852 22708 19854
rect 22428 19842 22484 19852
rect 22652 19346 22708 19852
rect 22652 19294 22654 19346
rect 22706 19294 22708 19346
rect 22652 19282 22708 19294
rect 22540 19236 22596 19246
rect 22316 19234 22596 19236
rect 22316 19182 22542 19234
rect 22594 19182 22596 19234
rect 22316 19180 22596 19182
rect 22540 19170 22596 19180
rect 22764 19124 22820 19134
rect 23100 19124 23156 19134
rect 22820 19122 23156 19124
rect 22820 19070 23102 19122
rect 23154 19070 23156 19122
rect 22820 19068 23156 19070
rect 22764 19030 22820 19068
rect 23100 19058 23156 19068
rect 23324 19124 23380 19134
rect 23324 19030 23380 19068
rect 21700 17724 21924 17780
rect 21644 17714 21700 17724
rect 21644 17554 21700 17566
rect 21644 17502 21646 17554
rect 21698 17502 21700 17554
rect 21644 17220 21700 17502
rect 21644 17154 21700 17164
rect 21868 16882 21924 17724
rect 21868 16830 21870 16882
rect 21922 16830 21924 16882
rect 21868 16818 21924 16830
rect 22204 15148 22260 18396
rect 23212 19010 23268 19022
rect 23212 18958 23214 19010
rect 23266 18958 23268 19010
rect 23212 18004 23268 18958
rect 23436 18676 23492 20524
rect 23660 20580 23716 20590
rect 23772 20580 23828 23324
rect 23996 23268 24052 23324
rect 23884 23212 24052 23268
rect 23884 21810 23940 23212
rect 23996 23042 24052 23054
rect 23996 22990 23998 23042
rect 24050 22990 24052 23042
rect 23996 22932 24052 22990
rect 23996 22866 24052 22876
rect 23884 21758 23886 21810
rect 23938 21758 23940 21810
rect 23884 21746 23940 21758
rect 23660 20578 23828 20580
rect 23660 20526 23662 20578
rect 23714 20526 23828 20578
rect 23660 20524 23828 20526
rect 24108 20580 24164 75180
rect 26908 40404 26964 40414
rect 26908 38948 26964 40348
rect 26908 38882 26964 38892
rect 26908 37380 26964 37390
rect 26908 36372 26964 37324
rect 26908 36306 26964 36316
rect 28476 33124 28532 33134
rect 28476 31668 28532 33068
rect 28476 31602 28532 31612
rect 30156 28084 30212 75628
rect 30156 28018 30212 28028
rect 31836 27748 31892 76300
rect 32732 75794 32788 79200
rect 33404 76354 33460 79200
rect 33404 76302 33406 76354
rect 33458 76302 33460 76354
rect 33404 76290 33460 76302
rect 33516 75908 33572 75918
rect 32732 75742 32734 75794
rect 32786 75742 32788 75794
rect 32732 75684 32788 75742
rect 33404 75852 33516 75908
rect 32956 75684 33012 75694
rect 32732 75682 33012 75684
rect 32732 75630 32958 75682
rect 33010 75630 33012 75682
rect 32732 75628 33012 75630
rect 32956 75618 33012 75628
rect 33404 67228 33460 75852
rect 33516 75842 33572 75852
rect 34076 75796 34132 79200
rect 34748 75908 34804 79200
rect 35084 76468 35140 76478
rect 35084 76374 35140 76412
rect 35420 76244 35476 79200
rect 36092 77028 36148 79200
rect 36092 76972 36372 77028
rect 36092 76578 36148 76590
rect 36092 76526 36094 76578
rect 36146 76526 36148 76578
rect 35756 76468 35812 76478
rect 35420 76188 35588 76244
rect 35196 76076 35460 76086
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35196 76010 35460 76020
rect 34748 75852 35252 75908
rect 34076 75794 34356 75796
rect 34076 75742 34078 75794
rect 34130 75742 34356 75794
rect 34076 75740 34356 75742
rect 34076 75730 34132 75740
rect 33516 75684 33572 75694
rect 33516 75590 33572 75628
rect 34300 75682 34356 75740
rect 34300 75630 34302 75682
rect 34354 75630 34356 75682
rect 34300 75618 34356 75630
rect 34748 75122 34804 75852
rect 34748 75070 34750 75122
rect 34802 75070 34804 75122
rect 34748 75058 34804 75070
rect 34860 75682 34916 75694
rect 34860 75630 34862 75682
rect 34914 75630 34916 75682
rect 33964 75012 34020 75022
rect 33404 67172 33572 67228
rect 31836 27682 31892 27692
rect 33516 27636 33572 67172
rect 33964 55468 34020 74956
rect 34860 55468 34916 75630
rect 34972 75012 35028 75022
rect 34972 74918 35028 74956
rect 35196 74898 35252 75852
rect 35420 75796 35476 75806
rect 35532 75796 35588 76188
rect 35420 75794 35700 75796
rect 35420 75742 35422 75794
rect 35474 75742 35700 75794
rect 35420 75740 35700 75742
rect 35420 75730 35476 75740
rect 35644 75682 35700 75740
rect 35644 75630 35646 75682
rect 35698 75630 35700 75682
rect 35644 75618 35700 75630
rect 35196 74846 35198 74898
rect 35250 74846 35252 74898
rect 35196 74834 35252 74846
rect 35756 74788 35812 76412
rect 35756 74694 35812 74732
rect 35980 75458 36036 75470
rect 35980 75406 35982 75458
rect 36034 75406 36036 75458
rect 35196 74508 35460 74518
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35196 74442 35460 74452
rect 35196 72940 35460 72950
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35196 72874 35460 72884
rect 35196 71372 35460 71382
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35196 71306 35460 71316
rect 35196 69804 35460 69814
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35196 69738 35460 69748
rect 35196 68236 35460 68246
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35196 68170 35460 68180
rect 35196 66668 35460 66678
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35196 66602 35460 66612
rect 35196 65100 35460 65110
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35196 65034 35460 65044
rect 35196 63532 35460 63542
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35196 63466 35460 63476
rect 35196 61964 35460 61974
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35196 61898 35460 61908
rect 35196 60396 35460 60406
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35196 60330 35460 60340
rect 35196 58828 35460 58838
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35196 58762 35460 58772
rect 35196 57260 35460 57270
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35196 57194 35460 57204
rect 35196 55692 35460 55702
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35196 55626 35460 55636
rect 33516 27570 33572 27580
rect 33852 55412 34020 55468
rect 34748 55412 34916 55468
rect 33852 27972 33908 55412
rect 33852 27074 33908 27916
rect 34748 27188 34804 55412
rect 35196 54124 35460 54134
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35196 54058 35460 54068
rect 35196 52556 35460 52566
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35196 52490 35460 52500
rect 35196 50988 35460 50998
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35196 50922 35460 50932
rect 35196 49420 35460 49430
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35196 49354 35460 49364
rect 35196 47852 35460 47862
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35196 47786 35460 47796
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35980 28084 36036 75406
rect 36092 29092 36148 76526
rect 36316 76466 36372 76972
rect 36316 76414 36318 76466
rect 36370 76414 36372 76466
rect 36316 75796 36372 76414
rect 36764 76690 36820 79200
rect 36764 76638 36766 76690
rect 36818 76638 36820 76690
rect 36428 75796 36484 75806
rect 36316 75794 36484 75796
rect 36316 75742 36430 75794
rect 36482 75742 36484 75794
rect 36316 75740 36484 75742
rect 36428 75730 36484 75740
rect 36764 75796 36820 76638
rect 37436 76692 37492 79200
rect 37660 76692 37716 76702
rect 37436 76690 37716 76692
rect 37436 76638 37662 76690
rect 37714 76638 37716 76690
rect 37436 76636 37716 76638
rect 37324 76356 37380 76366
rect 36764 75730 36820 75740
rect 37212 76354 37380 76356
rect 37212 76302 37326 76354
rect 37378 76302 37380 76354
rect 37212 76300 37380 76302
rect 37212 67228 37268 76300
rect 37324 76290 37380 76300
rect 37324 75796 37380 75806
rect 37324 75702 37380 75740
rect 37436 75122 37492 76636
rect 37660 76626 37716 76636
rect 38108 76580 38164 79200
rect 38780 76692 38836 79200
rect 39228 76692 39284 76702
rect 39452 76692 39508 79200
rect 38780 76636 39060 76692
rect 38108 76524 38276 76580
rect 38108 76356 38164 76366
rect 37996 76354 38164 76356
rect 37996 76302 38110 76354
rect 38162 76302 38164 76354
rect 37996 76300 38164 76302
rect 37884 75796 37940 75806
rect 37884 75702 37940 75740
rect 37436 75070 37438 75122
rect 37490 75070 37492 75122
rect 37436 75058 37492 75070
rect 37212 67172 37492 67228
rect 37100 29092 37156 29102
rect 36148 29036 36260 29092
rect 36092 29026 36148 29036
rect 34860 27972 34916 27982
rect 35084 27972 35140 27982
rect 34916 27970 35140 27972
rect 34916 27918 35086 27970
rect 35138 27918 35140 27970
rect 34916 27916 35140 27918
rect 34860 27906 34916 27916
rect 35084 27906 35140 27916
rect 35532 27858 35588 27870
rect 35532 27806 35534 27858
rect 35586 27806 35588 27858
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 33852 27022 33854 27074
rect 33906 27022 33908 27074
rect 33852 27010 33908 27022
rect 34636 27132 34804 27188
rect 34300 26962 34356 26974
rect 34300 26910 34302 26962
rect 34354 26910 34356 26962
rect 33740 26516 33796 26526
rect 33740 26290 33796 26460
rect 34300 26516 34356 26910
rect 34300 26450 34356 26460
rect 33740 26238 33742 26290
rect 33794 26238 33796 26290
rect 33740 26226 33796 26238
rect 34300 26290 34356 26302
rect 34300 26238 34302 26290
rect 34354 26238 34356 26290
rect 34300 26180 34356 26238
rect 34300 26114 34356 26124
rect 25564 25732 25620 25742
rect 25564 24946 25620 25676
rect 25564 24894 25566 24946
rect 25618 24894 25620 24946
rect 25564 24882 25620 24894
rect 26572 25732 26628 25742
rect 26572 24946 26628 25676
rect 26572 24894 26574 24946
rect 26626 24894 26628 24946
rect 26572 24882 26628 24894
rect 31836 25508 31892 25518
rect 25116 24724 25172 24734
rect 24892 24722 25172 24724
rect 24892 24670 25118 24722
rect 25170 24670 25172 24722
rect 24892 24668 25172 24670
rect 24780 24612 24836 24622
rect 24780 24050 24836 24556
rect 24780 23998 24782 24050
rect 24834 23998 24836 24050
rect 24780 23986 24836 23998
rect 24892 23828 24948 24668
rect 25116 24658 25172 24668
rect 25788 24724 25844 24734
rect 26684 24724 26740 24734
rect 25788 24722 26180 24724
rect 25788 24670 25790 24722
rect 25842 24670 26180 24722
rect 25788 24668 26180 24670
rect 25788 24658 25844 24668
rect 25676 24612 25732 24622
rect 25676 24518 25732 24556
rect 24668 23772 24948 23828
rect 24332 23380 24388 23390
rect 24332 23266 24388 23324
rect 24668 23378 24724 23772
rect 24668 23326 24670 23378
rect 24722 23326 24724 23378
rect 24668 23314 24724 23326
rect 25228 23380 25284 23390
rect 24332 23214 24334 23266
rect 24386 23214 24388 23266
rect 24332 23202 24388 23214
rect 24444 23266 24500 23278
rect 24444 23214 24446 23266
rect 24498 23214 24500 23266
rect 24444 23156 24500 23214
rect 24444 23090 24500 23100
rect 25228 23266 25284 23324
rect 26124 23380 26180 24668
rect 26684 24722 26964 24724
rect 26684 24670 26686 24722
rect 26738 24670 26964 24722
rect 26684 24668 26964 24670
rect 26684 24658 26740 24668
rect 26908 24050 26964 24668
rect 26908 23998 26910 24050
rect 26962 23998 26964 24050
rect 26908 23986 26964 23998
rect 27132 24722 27188 24734
rect 30268 24724 30324 24734
rect 27132 24670 27134 24722
rect 27186 24670 27188 24722
rect 26124 23286 26180 23324
rect 26572 23380 26628 23390
rect 25228 23214 25230 23266
rect 25282 23214 25284 23266
rect 24668 22708 24724 22718
rect 24220 22484 24276 22494
rect 24556 22484 24612 22494
rect 24220 22482 24612 22484
rect 24220 22430 24222 22482
rect 24274 22430 24558 22482
rect 24610 22430 24612 22482
rect 24220 22428 24612 22430
rect 24220 22418 24276 22428
rect 24556 22418 24612 22428
rect 24668 22146 24724 22652
rect 24668 22094 24670 22146
rect 24722 22094 24724 22146
rect 24668 21812 24724 22094
rect 24668 21746 24724 21756
rect 25228 21698 25284 23214
rect 25340 23266 25396 23278
rect 25340 23214 25342 23266
rect 25394 23214 25396 23266
rect 25340 22932 25396 23214
rect 25564 23156 25620 23166
rect 25564 23062 25620 23100
rect 25900 23156 25956 23166
rect 25900 23154 26068 23156
rect 25900 23102 25902 23154
rect 25954 23102 26068 23154
rect 25900 23100 26068 23102
rect 25900 23090 25956 23100
rect 25340 22866 25396 22876
rect 25564 22708 25620 22718
rect 25564 22370 25620 22652
rect 25564 22318 25566 22370
rect 25618 22318 25620 22370
rect 25564 22306 25620 22318
rect 25228 21646 25230 21698
rect 25282 21646 25284 21698
rect 25228 21634 25284 21646
rect 25340 21698 25396 21710
rect 25340 21646 25342 21698
rect 25394 21646 25396 21698
rect 23548 19012 23604 19022
rect 23548 18918 23604 18956
rect 23660 18788 23716 20524
rect 24108 20486 24164 20524
rect 24220 21586 24276 21598
rect 24220 21534 24222 21586
rect 24274 21534 24276 21586
rect 24220 20020 24276 21534
rect 24668 21476 24724 21486
rect 24668 21382 24724 21420
rect 25340 21476 25396 21646
rect 25564 21588 25620 21598
rect 25900 21588 25956 21598
rect 25564 21586 25956 21588
rect 25564 21534 25566 21586
rect 25618 21534 25902 21586
rect 25954 21534 25956 21586
rect 25564 21532 25956 21534
rect 25564 21522 25620 21532
rect 25900 21522 25956 21532
rect 25340 21410 25396 21420
rect 26012 20804 26068 23100
rect 26236 22260 26292 22270
rect 26236 22258 26516 22260
rect 26236 22206 26238 22258
rect 26290 22206 26516 22258
rect 26236 22204 26516 22206
rect 26236 22194 26292 22204
rect 26460 21810 26516 22204
rect 26460 21758 26462 21810
rect 26514 21758 26516 21810
rect 26460 21746 26516 21758
rect 26572 21810 26628 23324
rect 27132 22708 27188 24670
rect 29932 24722 30324 24724
rect 29932 24670 30270 24722
rect 30322 24670 30324 24722
rect 29932 24668 30324 24670
rect 27692 24612 27748 24622
rect 27692 23828 27748 24556
rect 27804 24610 27860 24622
rect 27804 24558 27806 24610
rect 27858 24558 27860 24610
rect 27804 24052 27860 24558
rect 29932 24610 29988 24668
rect 30268 24658 30324 24668
rect 29932 24558 29934 24610
rect 29986 24558 29988 24610
rect 29932 24546 29988 24558
rect 30380 24612 30436 24622
rect 30380 24518 30436 24556
rect 27916 24052 27972 24062
rect 27804 24050 27972 24052
rect 27804 23998 27918 24050
rect 27970 23998 27972 24050
rect 27804 23996 27972 23998
rect 27916 23986 27972 23996
rect 27804 23828 27860 23838
rect 27692 23826 27860 23828
rect 27692 23774 27806 23826
rect 27858 23774 27860 23826
rect 27692 23772 27860 23774
rect 27804 23762 27860 23772
rect 27580 23716 27636 23726
rect 27580 23622 27636 23660
rect 28028 23714 28084 23726
rect 28028 23662 28030 23714
rect 28082 23662 28084 23714
rect 28028 23380 28084 23662
rect 28028 23286 28084 23324
rect 27356 23156 27412 23166
rect 27356 23062 27412 23100
rect 27804 23156 27860 23166
rect 27804 23062 27860 23100
rect 28364 23154 28420 23166
rect 31612 23156 31668 23166
rect 28364 23102 28366 23154
rect 28418 23102 28420 23154
rect 27916 23044 27972 23054
rect 27916 22950 27972 22988
rect 27132 22642 27188 22652
rect 28364 22708 28420 23102
rect 31276 23154 31668 23156
rect 31276 23102 31614 23154
rect 31666 23102 31668 23154
rect 31276 23100 31668 23102
rect 29148 23044 29204 23054
rect 29148 22950 29204 22988
rect 31276 23042 31332 23100
rect 31612 23090 31668 23100
rect 31724 23156 31780 23166
rect 31724 23062 31780 23100
rect 31276 22990 31278 23042
rect 31330 22990 31332 23042
rect 31276 22978 31332 22990
rect 28364 22642 28420 22652
rect 29036 22708 29092 22718
rect 28364 22484 28420 22494
rect 28364 22390 28420 22428
rect 26572 21758 26574 21810
rect 26626 21758 26628 21810
rect 26572 21746 26628 21758
rect 26348 21588 26404 21598
rect 29036 21588 29092 22652
rect 29148 22484 29204 22494
rect 29148 22390 29204 22428
rect 29260 22146 29316 22158
rect 29260 22094 29262 22146
rect 29314 22094 29316 22146
rect 29148 21588 29204 21598
rect 26348 21586 26740 21588
rect 26348 21534 26350 21586
rect 26402 21534 26740 21586
rect 26348 21532 26740 21534
rect 29036 21586 29204 21588
rect 29036 21534 29150 21586
rect 29202 21534 29204 21586
rect 29036 21532 29204 21534
rect 26348 21522 26404 21532
rect 26572 20804 26628 20814
rect 26012 20802 26628 20804
rect 26012 20750 26574 20802
rect 26626 20750 26628 20802
rect 26012 20748 26628 20750
rect 24108 19684 24164 19694
rect 24220 19684 24276 19964
rect 24444 20690 24500 20702
rect 24444 20638 24446 20690
rect 24498 20638 24500 20690
rect 24444 19908 24500 20638
rect 24780 20690 24836 20702
rect 24780 20638 24782 20690
rect 24834 20638 24836 20690
rect 24780 20468 24836 20638
rect 24780 20402 24836 20412
rect 25228 20690 25284 20702
rect 25228 20638 25230 20690
rect 25282 20638 25284 20690
rect 25228 20188 25284 20638
rect 25788 20690 25844 20702
rect 25788 20638 25790 20690
rect 25842 20638 25844 20690
rect 25340 20580 25396 20590
rect 25340 20486 25396 20524
rect 25564 20580 25620 20590
rect 25564 20486 25620 20524
rect 25228 20132 25396 20188
rect 25564 20132 25620 20142
rect 25788 20132 25844 20638
rect 25340 20130 25844 20132
rect 25340 20078 25566 20130
rect 25618 20078 25844 20130
rect 25340 20076 25844 20078
rect 25900 20578 25956 20590
rect 25900 20526 25902 20578
rect 25954 20526 25956 20578
rect 25228 20020 25284 20030
rect 25228 19926 25284 19964
rect 24556 19908 24612 19918
rect 24444 19906 24612 19908
rect 24444 19854 24558 19906
rect 24610 19854 24612 19906
rect 24444 19852 24612 19854
rect 24556 19842 24612 19852
rect 24164 19628 24276 19684
rect 24108 19618 24164 19628
rect 23660 18722 23716 18732
rect 23996 19124 24052 19134
rect 22540 17948 23268 18004
rect 23324 18620 23492 18676
rect 22316 17780 22372 17790
rect 22316 17686 22372 17724
rect 22540 16994 22596 17948
rect 22540 16942 22542 16994
rect 22594 16942 22596 16994
rect 22540 16930 22596 16942
rect 23324 15148 23380 18620
rect 23436 18450 23492 18462
rect 23436 18398 23438 18450
rect 23490 18398 23492 18450
rect 23436 16772 23492 18398
rect 23996 18338 24052 19068
rect 24108 19012 24164 19022
rect 24108 18918 24164 18956
rect 24220 18564 24276 19628
rect 24444 19124 24500 19134
rect 24444 19030 24500 19068
rect 24780 19122 24836 19134
rect 24780 19070 24782 19122
rect 24834 19070 24836 19122
rect 24332 19010 24388 19022
rect 24332 18958 24334 19010
rect 24386 18958 24388 19010
rect 24332 18788 24388 18958
rect 24332 18722 24388 18732
rect 24332 18564 24388 18574
rect 24220 18562 24388 18564
rect 24220 18510 24334 18562
rect 24386 18510 24388 18562
rect 24220 18508 24388 18510
rect 24332 18498 24388 18508
rect 23996 18286 23998 18338
rect 24050 18286 24052 18338
rect 23996 18004 24052 18286
rect 24668 18450 24724 18462
rect 24668 18398 24670 18450
rect 24722 18398 24724 18450
rect 24668 18340 24724 18398
rect 24668 18274 24724 18284
rect 23996 17938 24052 17948
rect 24668 16772 24724 16782
rect 24780 16772 24836 19070
rect 25116 19122 25172 19134
rect 25116 19070 25118 19122
rect 25170 19070 25172 19122
rect 25116 18004 25172 19070
rect 25452 19124 25508 20076
rect 25564 20066 25620 20076
rect 25900 19908 25956 20526
rect 26124 20578 26180 20590
rect 26124 20526 26126 20578
rect 26178 20526 26180 20578
rect 26012 19908 26068 19918
rect 25676 19906 26068 19908
rect 25676 19854 26014 19906
rect 26066 19854 26068 19906
rect 25676 19852 26068 19854
rect 25452 19058 25508 19068
rect 25564 19236 25620 19246
rect 25564 19122 25620 19180
rect 25564 19070 25566 19122
rect 25618 19070 25620 19122
rect 25564 19058 25620 19070
rect 25340 18452 25396 18462
rect 25340 18358 25396 18396
rect 25116 17938 25172 17948
rect 23436 16716 23828 16772
rect 23772 16210 23828 16716
rect 24668 16770 24836 16772
rect 24668 16718 24670 16770
rect 24722 16718 24836 16770
rect 24668 16716 24836 16718
rect 25004 17780 25060 17790
rect 24668 16706 24724 16716
rect 23772 16158 23774 16210
rect 23826 16158 23828 16210
rect 23772 15876 23828 16158
rect 23772 15810 23828 15820
rect 25004 16098 25060 17724
rect 25004 16046 25006 16098
rect 25058 16046 25060 16098
rect 22204 15092 22596 15148
rect 22540 13634 22596 15092
rect 22540 13582 22542 13634
rect 22594 13582 22596 13634
rect 21756 13412 21812 13422
rect 21756 12178 21812 13356
rect 22540 13076 22596 13582
rect 22540 13010 22596 13020
rect 22652 15092 23380 15148
rect 21756 12126 21758 12178
rect 21810 12126 21812 12178
rect 21756 12114 21812 12126
rect 22428 12068 22484 12078
rect 22316 12066 22484 12068
rect 22316 12014 22430 12066
rect 22482 12014 22484 12066
rect 22316 12012 22484 12014
rect 21588 11452 21812 11508
rect 21532 11442 21588 11452
rect 21756 10834 21812 11452
rect 22316 11506 22372 12012
rect 22428 12002 22484 12012
rect 22540 12068 22596 12078
rect 22428 11620 22484 11630
rect 22540 11620 22596 12012
rect 22428 11618 22596 11620
rect 22428 11566 22430 11618
rect 22482 11566 22596 11618
rect 22428 11564 22596 11566
rect 22428 11554 22484 11564
rect 22316 11454 22318 11506
rect 22370 11454 22372 11506
rect 22316 11442 22372 11454
rect 22092 11396 22148 11434
rect 22092 11330 22148 11340
rect 22092 11172 22148 11182
rect 21756 10782 21758 10834
rect 21810 10782 21812 10834
rect 21756 10770 21812 10782
rect 21980 11116 22092 11172
rect 21644 9044 21700 9054
rect 21644 8258 21700 8988
rect 21644 8206 21646 8258
rect 21698 8206 21700 8258
rect 21644 8194 21700 8206
rect 21420 7362 21476 7374
rect 21420 7310 21422 7362
rect 21474 7310 21476 7362
rect 21420 6468 21476 7310
rect 21868 7362 21924 7374
rect 21868 7310 21870 7362
rect 21922 7310 21924 7362
rect 21868 7250 21924 7310
rect 21868 7198 21870 7250
rect 21922 7198 21924 7250
rect 21868 7186 21924 7198
rect 21756 7140 21812 7150
rect 21644 7084 21756 7140
rect 21532 6580 21588 6590
rect 21532 6486 21588 6524
rect 21420 6402 21476 6412
rect 21308 6188 21588 6244
rect 21532 6130 21588 6188
rect 21532 6078 21534 6130
rect 21586 6078 21588 6130
rect 21532 6066 21588 6078
rect 20748 4396 20916 4452
rect 21084 5796 21140 5806
rect 20748 4116 20804 4396
rect 20972 4340 21028 4350
rect 20748 4050 20804 4060
rect 20860 4338 21028 4340
rect 20860 4286 20974 4338
rect 21026 4286 21028 4338
rect 20860 4284 21028 4286
rect 20524 3938 20580 3948
rect 20860 2436 20916 4284
rect 20972 4274 21028 4284
rect 21084 3892 21140 5740
rect 21196 5794 21252 5806
rect 21196 5742 21198 5794
rect 21250 5742 21252 5794
rect 21196 5684 21252 5742
rect 21196 5618 21252 5628
rect 21420 5682 21476 5694
rect 21420 5630 21422 5682
rect 21474 5630 21476 5682
rect 21420 5348 21476 5630
rect 21532 5348 21588 5358
rect 21476 5346 21588 5348
rect 21476 5294 21534 5346
rect 21586 5294 21588 5346
rect 21476 5292 21588 5294
rect 21420 5254 21476 5292
rect 21532 5282 21588 5292
rect 21196 5236 21252 5246
rect 21196 4562 21252 5180
rect 21196 4510 21198 4562
rect 21250 4510 21252 4562
rect 21196 4498 21252 4510
rect 21308 4564 21364 4574
rect 21308 4450 21364 4508
rect 21308 4398 21310 4450
rect 21362 4398 21364 4450
rect 21308 4386 21364 4398
rect 21084 3554 21140 3836
rect 21084 3502 21086 3554
rect 21138 3502 21140 3554
rect 21084 3490 21140 3502
rect 21196 4228 21252 4238
rect 21196 3388 21252 4172
rect 21644 3778 21700 7084
rect 21756 7074 21812 7084
rect 21868 6804 21924 6814
rect 21868 6690 21924 6748
rect 21868 6638 21870 6690
rect 21922 6638 21924 6690
rect 21868 6580 21924 6638
rect 21868 6514 21924 6524
rect 21980 6244 22036 11116
rect 22092 11106 22148 11116
rect 22204 10610 22260 10622
rect 22204 10558 22206 10610
rect 22258 10558 22260 10610
rect 22204 8484 22260 10558
rect 22204 8418 22260 8428
rect 22316 10498 22372 10510
rect 22316 10446 22318 10498
rect 22370 10446 22372 10498
rect 22316 8372 22372 10446
rect 22540 10500 22596 10510
rect 22540 10406 22596 10444
rect 22540 9268 22596 9278
rect 22652 9268 22708 15092
rect 23436 13748 23492 13758
rect 23436 13654 23492 13692
rect 23660 13634 23716 13646
rect 23660 13582 23662 13634
rect 23714 13582 23716 13634
rect 22988 13412 23044 13422
rect 22988 12962 23044 13356
rect 23660 13074 23716 13582
rect 23660 13022 23662 13074
rect 23714 13022 23716 13074
rect 23660 13010 23716 13022
rect 23772 13522 23828 13534
rect 23772 13470 23774 13522
rect 23826 13470 23828 13522
rect 23772 13076 23828 13470
rect 25004 13412 25060 16046
rect 25004 13346 25060 13356
rect 23772 13010 23828 13020
rect 25452 13300 25508 13310
rect 22988 12910 22990 12962
rect 23042 12910 23044 12962
rect 22988 12898 23044 12910
rect 25452 12402 25508 13244
rect 25676 12964 25732 19852
rect 26012 19842 26068 19852
rect 26124 19236 26180 20526
rect 26124 19170 26180 19180
rect 26460 20018 26516 20030
rect 26460 19966 26462 20018
rect 26514 19966 26516 20018
rect 25900 19122 25956 19134
rect 25900 19070 25902 19122
rect 25954 19070 25956 19122
rect 25788 18452 25844 18462
rect 25788 18358 25844 18396
rect 25900 18340 25956 19070
rect 26236 19124 26292 19134
rect 26236 19030 26292 19068
rect 26348 19010 26404 19022
rect 26348 18958 26350 19010
rect 26402 18958 26404 19010
rect 26348 18900 26404 18958
rect 26124 18844 26404 18900
rect 26012 18564 26068 18574
rect 26124 18564 26180 18844
rect 26460 18788 26516 19966
rect 26572 19348 26628 20748
rect 26684 20132 26740 21532
rect 26908 20580 26964 20590
rect 26908 20578 27636 20580
rect 26908 20526 26910 20578
rect 26962 20526 27636 20578
rect 26908 20524 27636 20526
rect 26908 20514 26964 20524
rect 26684 20066 26740 20076
rect 27132 19908 27188 19918
rect 27132 19906 27524 19908
rect 27132 19854 27134 19906
rect 27186 19854 27524 19906
rect 27132 19852 27524 19854
rect 27132 19842 27188 19852
rect 26572 19282 26628 19292
rect 27468 19346 27524 19852
rect 27468 19294 27470 19346
rect 27522 19294 27524 19346
rect 27468 19282 27524 19294
rect 26908 19236 26964 19246
rect 26908 19142 26964 19180
rect 27580 19236 27636 20524
rect 28588 19348 28644 19358
rect 29036 19348 29092 19358
rect 28588 19346 29092 19348
rect 28588 19294 28590 19346
rect 28642 19294 29038 19346
rect 29090 19294 29092 19346
rect 28588 19292 29092 19294
rect 28588 19282 28644 19292
rect 29036 19282 29092 19292
rect 27580 19142 27636 19180
rect 26572 19012 26628 19022
rect 26572 18918 26628 18956
rect 27356 19010 27412 19022
rect 27356 18958 27358 19010
rect 27410 18958 27412 19010
rect 26068 18508 26180 18564
rect 26348 18732 26516 18788
rect 27356 18788 27412 18958
rect 28476 19010 28532 19022
rect 28476 18958 28478 19010
rect 28530 18958 28532 19010
rect 26012 18498 26068 18508
rect 26348 18452 26404 18732
rect 27356 18722 27412 18732
rect 27916 18788 27972 18798
rect 26348 18386 26404 18396
rect 25900 16884 25956 18284
rect 26460 18340 26516 18350
rect 26460 18338 26740 18340
rect 26460 18286 26462 18338
rect 26514 18286 26740 18338
rect 26460 18284 26740 18286
rect 26460 18274 26516 18284
rect 26348 17332 26404 17342
rect 26348 17106 26404 17276
rect 26348 17054 26350 17106
rect 26402 17054 26404 17106
rect 26348 17042 26404 17054
rect 26684 17106 26740 18284
rect 27916 17778 27972 18732
rect 28476 18788 28532 18958
rect 28476 18722 28532 18732
rect 27916 17726 27918 17778
rect 27970 17726 27972 17778
rect 27916 17714 27972 17726
rect 28140 18452 28196 18462
rect 27244 17666 27300 17678
rect 27244 17614 27246 17666
rect 27298 17614 27300 17666
rect 26684 17054 26686 17106
rect 26738 17054 26740 17106
rect 26684 17042 26740 17054
rect 26796 17332 26852 17342
rect 26796 17106 26852 17276
rect 26796 17054 26798 17106
rect 26850 17054 26852 17106
rect 26796 17042 26852 17054
rect 27244 17108 27300 17614
rect 27580 17108 27636 17118
rect 28140 17108 28196 18396
rect 28588 18338 28644 18350
rect 28588 18286 28590 18338
rect 28642 18286 28644 18338
rect 28588 17778 28644 18286
rect 28588 17726 28590 17778
rect 28642 17726 28644 17778
rect 28588 17714 28644 17726
rect 28700 18340 28756 18350
rect 29148 18340 29204 21532
rect 29260 20132 29316 22094
rect 29932 21476 29988 21486
rect 29820 21474 29988 21476
rect 29820 21422 29934 21474
rect 29986 21422 29988 21474
rect 29820 21420 29988 21422
rect 29820 20914 29876 21420
rect 29932 21410 29988 21420
rect 29820 20862 29822 20914
rect 29874 20862 29876 20914
rect 29820 20850 29876 20862
rect 29484 20580 29540 20590
rect 29484 20486 29540 20524
rect 29708 20578 29764 20590
rect 29708 20526 29710 20578
rect 29762 20526 29764 20578
rect 29708 20244 29764 20526
rect 29708 20178 29764 20188
rect 29932 20578 29988 20590
rect 29932 20526 29934 20578
rect 29986 20526 29988 20578
rect 29260 20066 29316 20076
rect 29596 20020 29652 20030
rect 29372 20018 29652 20020
rect 29372 19966 29598 20018
rect 29650 19966 29652 20018
rect 29372 19964 29652 19966
rect 29260 19906 29316 19918
rect 29260 19854 29262 19906
rect 29314 19854 29316 19906
rect 29260 19346 29316 19854
rect 29260 19294 29262 19346
rect 29314 19294 29316 19346
rect 29260 19282 29316 19294
rect 28756 18284 29204 18340
rect 29372 18450 29428 19964
rect 29596 19954 29652 19964
rect 29932 19236 29988 20526
rect 30492 20580 30548 20590
rect 31836 20580 31892 25452
rect 34636 25284 34692 27132
rect 34860 27076 34916 27114
rect 34748 27020 34860 27076
rect 34748 26178 34804 27020
rect 34860 27010 34916 27020
rect 35532 27076 35588 27806
rect 35980 27858 36036 28028
rect 35980 27806 35982 27858
rect 36034 27806 36036 27858
rect 35980 27794 36036 27806
rect 36092 27746 36148 27758
rect 36092 27694 36094 27746
rect 36146 27694 36148 27746
rect 35532 27010 35588 27020
rect 35868 27186 35924 27198
rect 35868 27134 35870 27186
rect 35922 27134 35924 27186
rect 34860 26850 34916 26862
rect 34860 26798 34862 26850
rect 34914 26798 34916 26850
rect 34860 26404 34916 26798
rect 34860 26338 34916 26348
rect 35532 26404 35588 26414
rect 35532 26310 35588 26348
rect 35756 26404 35812 26414
rect 35196 26292 35252 26302
rect 35196 26198 35252 26236
rect 34748 26126 34750 26178
rect 34802 26126 34804 26178
rect 34748 25508 34804 26126
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 34972 25508 35028 25518
rect 34748 25506 35028 25508
rect 34748 25454 34974 25506
rect 35026 25454 35028 25506
rect 34748 25452 35028 25454
rect 34972 25442 35028 25452
rect 35532 25506 35588 25518
rect 35532 25454 35534 25506
rect 35586 25454 35588 25506
rect 34748 25284 34804 25294
rect 34636 25228 34748 25284
rect 34748 25190 34804 25228
rect 35532 25284 35588 25454
rect 35756 25394 35812 26348
rect 35756 25342 35758 25394
rect 35810 25342 35812 25394
rect 35756 25330 35812 25342
rect 35532 25218 35588 25228
rect 32620 24948 32676 24958
rect 32396 21588 32452 21598
rect 32060 21586 32452 21588
rect 32060 21534 32398 21586
rect 32450 21534 32452 21586
rect 32060 21532 32452 21534
rect 32060 21474 32116 21532
rect 32396 21522 32452 21532
rect 32060 21422 32062 21474
rect 32114 21422 32116 21474
rect 32060 21410 32116 21422
rect 32508 21364 32564 21374
rect 30492 20578 30660 20580
rect 30492 20526 30494 20578
rect 30546 20526 30660 20578
rect 30492 20524 30660 20526
rect 30492 20514 30548 20524
rect 30156 20132 30212 20142
rect 30156 19460 30212 20076
rect 30156 19394 30212 19404
rect 30380 19906 30436 19918
rect 30380 19854 30382 19906
rect 30434 19854 30436 19906
rect 30380 19346 30436 19854
rect 30380 19294 30382 19346
rect 30434 19294 30436 19346
rect 30380 19282 30436 19294
rect 30268 19236 30324 19246
rect 29988 19234 30324 19236
rect 29988 19182 30270 19234
rect 30322 19182 30324 19234
rect 29988 19180 30324 19182
rect 29932 19142 29988 19180
rect 30268 19170 30324 19180
rect 30492 19236 30548 19246
rect 30492 19142 30548 19180
rect 29708 19124 29764 19134
rect 29708 19030 29764 19068
rect 30604 19124 30660 20524
rect 31724 20524 31892 20580
rect 32284 21362 32564 21364
rect 32284 21310 32510 21362
rect 32562 21310 32564 21362
rect 32284 21308 32564 21310
rect 31276 20132 31332 20142
rect 31276 19346 31332 20076
rect 31276 19294 31278 19346
rect 31330 19294 31332 19346
rect 31276 19236 31332 19294
rect 31276 19170 31332 19180
rect 30604 19058 30660 19068
rect 29484 19012 29540 19022
rect 29484 18918 29540 18956
rect 29820 19010 29876 19022
rect 29820 18958 29822 19010
rect 29874 18958 29876 19010
rect 29820 18564 29876 18958
rect 30716 19012 30772 19022
rect 30716 18918 30772 18956
rect 31724 18676 31780 20524
rect 31836 20356 31892 20366
rect 31836 18900 31892 20300
rect 32284 20244 32340 21308
rect 32508 21298 32564 21308
rect 32508 21026 32564 21038
rect 32508 20974 32510 21026
rect 32562 20974 32564 21026
rect 32284 20178 32340 20188
rect 32396 20578 32452 20590
rect 32396 20526 32398 20578
rect 32450 20526 32452 20578
rect 32172 19458 32228 19470
rect 32172 19406 32174 19458
rect 32226 19406 32228 19458
rect 31836 18834 31892 18844
rect 31948 19010 32004 19022
rect 31948 18958 31950 19010
rect 32002 18958 32004 19010
rect 31724 18620 31892 18676
rect 30044 18564 30100 18574
rect 29820 18562 30100 18564
rect 29820 18510 30046 18562
rect 30098 18510 30100 18562
rect 29820 18508 30100 18510
rect 30044 18498 30100 18508
rect 29372 18398 29374 18450
rect 29426 18398 29428 18450
rect 28700 17556 28756 18284
rect 28476 17444 28532 17454
rect 28476 17350 28532 17388
rect 27244 17106 28196 17108
rect 27244 17054 27582 17106
rect 27634 17054 28142 17106
rect 28194 17054 28196 17106
rect 27244 17052 28196 17054
rect 27020 16994 27076 17006
rect 27020 16942 27022 16994
rect 27074 16942 27076 16994
rect 25900 16818 25956 16828
rect 26572 16882 26628 16894
rect 26572 16830 26574 16882
rect 26626 16830 26628 16882
rect 25788 15986 25844 15998
rect 25788 15934 25790 15986
rect 25842 15934 25844 15986
rect 25788 15148 25844 15934
rect 26572 15316 26628 16830
rect 26908 15876 26964 15886
rect 26572 15260 26852 15316
rect 25788 15092 26740 15148
rect 26684 14642 26740 15092
rect 26684 14590 26686 14642
rect 26738 14590 26740 14642
rect 26684 14578 26740 14590
rect 26124 14532 26180 14542
rect 25900 14530 26180 14532
rect 25900 14478 26126 14530
rect 26178 14478 26180 14530
rect 25900 14476 26180 14478
rect 25900 13970 25956 14476
rect 26124 14466 26180 14476
rect 26796 14420 26852 15260
rect 26796 14326 26852 14364
rect 26572 14308 26628 14318
rect 26572 14214 26628 14252
rect 25900 13918 25902 13970
rect 25954 13918 25956 13970
rect 25900 13906 25956 13918
rect 26124 13858 26180 13870
rect 26124 13806 26126 13858
rect 26178 13806 26180 13858
rect 26124 13300 26180 13806
rect 26684 13860 26740 13870
rect 26684 13858 26852 13860
rect 26684 13806 26686 13858
rect 26738 13806 26852 13858
rect 26684 13804 26852 13806
rect 26684 13794 26740 13804
rect 26236 13748 26292 13758
rect 26572 13748 26628 13758
rect 26236 13746 26572 13748
rect 26236 13694 26238 13746
rect 26290 13694 26572 13746
rect 26236 13692 26572 13694
rect 26236 13682 26292 13692
rect 26572 13654 26628 13692
rect 26684 13524 26740 13534
rect 26684 13430 26740 13468
rect 26796 13300 26852 13804
rect 26124 13234 26180 13244
rect 26460 13244 26852 13300
rect 25788 13076 25844 13086
rect 26460 13076 26516 13244
rect 25788 13074 26516 13076
rect 25788 13022 25790 13074
rect 25842 13022 26516 13074
rect 25788 13020 26516 13022
rect 25788 13010 25844 13020
rect 25676 12898 25732 12908
rect 26460 12962 26516 13020
rect 26572 13076 26628 13086
rect 26572 12982 26628 13020
rect 26460 12910 26462 12962
rect 26514 12910 26516 12962
rect 26460 12898 26516 12910
rect 25452 12350 25454 12402
rect 25506 12350 25508 12402
rect 24556 12292 24612 12302
rect 24556 12066 24612 12236
rect 25452 12292 25508 12350
rect 25452 12226 25508 12236
rect 26236 12738 26292 12750
rect 26236 12686 26238 12738
rect 26290 12686 26292 12738
rect 24556 12014 24558 12066
rect 24610 12014 24612 12066
rect 24556 12002 24612 12014
rect 25228 12178 25284 12190
rect 25228 12126 25230 12178
rect 25282 12126 25284 12178
rect 24332 11844 24388 11854
rect 24108 11732 24164 11742
rect 24108 10834 24164 11676
rect 24108 10782 24110 10834
rect 24162 10782 24164 10834
rect 24108 10770 24164 10782
rect 24332 10836 24388 11788
rect 25228 11732 25284 12126
rect 25900 12180 25956 12190
rect 26236 12180 26292 12686
rect 26684 12738 26740 12750
rect 26684 12686 26686 12738
rect 26738 12686 26740 12738
rect 25900 12178 26292 12180
rect 25900 12126 25902 12178
rect 25954 12126 26292 12178
rect 25900 12124 26292 12126
rect 25900 12114 25956 12124
rect 25340 12068 25396 12078
rect 25340 11974 25396 12012
rect 25228 11666 25284 11676
rect 25676 11732 25732 11742
rect 25340 11394 25396 11406
rect 25340 11342 25342 11394
rect 25394 11342 25396 11394
rect 24892 11284 24948 11294
rect 24892 11190 24948 11228
rect 25004 11282 25060 11294
rect 25004 11230 25006 11282
rect 25058 11230 25060 11282
rect 24780 11172 24836 11182
rect 24780 11078 24836 11116
rect 25004 10836 25060 11230
rect 24332 10834 24612 10836
rect 24332 10782 24334 10834
rect 24386 10782 24612 10834
rect 24332 10780 24612 10782
rect 24332 10770 24388 10780
rect 24220 10500 24276 10510
rect 24220 10406 24276 10444
rect 22764 10388 22820 10398
rect 22764 9940 22820 10332
rect 22764 9826 22820 9884
rect 22764 9774 22766 9826
rect 22818 9774 22820 9826
rect 22764 9762 22820 9774
rect 22540 9266 22708 9268
rect 22540 9214 22542 9266
rect 22594 9214 22708 9266
rect 22540 9212 22708 9214
rect 23548 9716 23604 9726
rect 22428 8372 22484 8382
rect 22316 8370 22484 8372
rect 22316 8318 22430 8370
rect 22482 8318 22484 8370
rect 22316 8316 22484 8318
rect 22428 8306 22484 8316
rect 22540 8372 22596 9212
rect 22764 9044 22820 9054
rect 22540 8306 22596 8316
rect 22652 8988 22764 9044
rect 22204 7700 22260 7710
rect 21868 6188 22036 6244
rect 22092 7250 22148 7262
rect 22092 7198 22094 7250
rect 22146 7198 22148 7250
rect 21756 5908 21812 5946
rect 21756 5842 21812 5852
rect 21868 5684 21924 6188
rect 22092 5908 22148 7198
rect 22204 6578 22260 7644
rect 22540 7476 22596 7486
rect 22204 6526 22206 6578
rect 22258 6526 22260 6578
rect 22204 6514 22260 6526
rect 22316 7362 22372 7374
rect 22316 7310 22318 7362
rect 22370 7310 22372 7362
rect 22316 6132 22372 7310
rect 22316 6066 22372 6076
rect 22428 7250 22484 7262
rect 22428 7198 22430 7250
rect 22482 7198 22484 7250
rect 22316 5908 22372 5918
rect 22092 5906 22372 5908
rect 22092 5854 22318 5906
rect 22370 5854 22372 5906
rect 22092 5852 22372 5854
rect 21756 5628 21924 5684
rect 21980 5796 22036 5806
rect 21756 5234 21812 5628
rect 21756 5182 21758 5234
rect 21810 5182 21812 5234
rect 21756 5170 21812 5182
rect 21868 5460 21924 5470
rect 21868 5122 21924 5404
rect 21868 5070 21870 5122
rect 21922 5070 21924 5122
rect 21868 5058 21924 5070
rect 21868 4564 21924 4574
rect 21756 4452 21812 4462
rect 21756 4358 21812 4396
rect 21756 4228 21812 4238
rect 21756 4134 21812 4172
rect 21644 3726 21646 3778
rect 21698 3726 21700 3778
rect 21644 3714 21700 3726
rect 21756 4004 21812 4014
rect 20860 2370 20916 2380
rect 21084 3332 21252 3388
rect 21644 3554 21700 3566
rect 21644 3502 21646 3554
rect 21698 3502 21700 3554
rect 21644 3444 21700 3502
rect 21644 3378 21700 3388
rect 21084 800 21140 3332
rect 21308 3330 21364 3342
rect 21308 3278 21310 3330
rect 21362 3278 21364 3330
rect 21308 1652 21364 3278
rect 21308 1586 21364 1596
rect 21756 800 21812 3948
rect 21868 3780 21924 4508
rect 21980 4450 22036 5740
rect 22316 5348 22372 5852
rect 22316 5282 22372 5292
rect 22428 5234 22484 7198
rect 22540 6804 22596 7420
rect 22540 6738 22596 6748
rect 22652 6692 22708 8988
rect 22764 8978 22820 8988
rect 23548 9044 23604 9660
rect 23548 8978 23604 8988
rect 23436 8930 23492 8942
rect 23436 8878 23438 8930
rect 23490 8878 23492 8930
rect 23100 8708 23156 8718
rect 23100 7700 23156 8652
rect 23436 7700 23492 8878
rect 23884 8932 23940 8942
rect 24332 8932 24388 8942
rect 23884 8930 24276 8932
rect 23884 8878 23886 8930
rect 23938 8878 24276 8930
rect 23884 8876 24276 8878
rect 23884 8866 23940 8876
rect 23436 7644 23716 7700
rect 23100 7606 23156 7644
rect 23436 7476 23492 7486
rect 23212 7474 23492 7476
rect 23212 7422 23438 7474
rect 23490 7422 23492 7474
rect 23212 7420 23492 7422
rect 22764 7364 22820 7374
rect 22764 7362 23044 7364
rect 22764 7310 22766 7362
rect 22818 7310 23044 7362
rect 22764 7308 23044 7310
rect 22764 7298 22820 7308
rect 22652 6690 22932 6692
rect 22652 6638 22654 6690
rect 22706 6638 22932 6690
rect 22652 6636 22932 6638
rect 22652 6626 22708 6636
rect 22652 6018 22708 6030
rect 22652 5966 22654 6018
rect 22706 5966 22708 6018
rect 22652 5572 22708 5966
rect 22652 5506 22708 5516
rect 22428 5182 22430 5234
rect 22482 5182 22484 5234
rect 22428 5170 22484 5182
rect 22876 5124 22932 6636
rect 22988 6244 23044 7308
rect 23212 7250 23268 7420
rect 23436 7410 23492 7420
rect 23212 7198 23214 7250
rect 23266 7198 23268 7250
rect 23212 7186 23268 7198
rect 23436 7250 23492 7262
rect 23436 7198 23438 7250
rect 23490 7198 23492 7250
rect 23324 6804 23380 6814
rect 22988 6178 23044 6188
rect 23100 6468 23156 6478
rect 22988 5906 23044 5918
rect 22988 5854 22990 5906
rect 23042 5854 23044 5906
rect 22988 5236 23044 5854
rect 23100 5348 23156 6412
rect 23324 6018 23380 6748
rect 23436 6690 23492 7198
rect 23436 6638 23438 6690
rect 23490 6638 23492 6690
rect 23436 6626 23492 6638
rect 23324 5966 23326 6018
rect 23378 5966 23380 6018
rect 23324 5954 23380 5966
rect 23660 6020 23716 7644
rect 23772 7364 23828 7374
rect 23772 7270 23828 7308
rect 23996 6020 24052 6030
rect 23660 6018 23940 6020
rect 23660 5966 23662 6018
rect 23714 5966 23940 6018
rect 23660 5964 23940 5966
rect 23660 5954 23716 5964
rect 23212 5794 23268 5806
rect 23212 5742 23214 5794
rect 23266 5742 23268 5794
rect 23212 5460 23268 5742
rect 23660 5684 23716 5694
rect 23716 5628 23828 5684
rect 23660 5618 23716 5628
rect 23212 5404 23716 5460
rect 23100 5292 23380 5348
rect 22988 5170 23044 5180
rect 22876 5030 22932 5068
rect 22428 5012 22484 5022
rect 22316 4900 22372 4910
rect 21980 4398 21982 4450
rect 22034 4398 22036 4450
rect 21980 4386 22036 4398
rect 22204 4898 22372 4900
rect 22204 4846 22318 4898
rect 22370 4846 22372 4898
rect 22204 4844 22372 4846
rect 21980 3780 22036 3790
rect 21868 3778 22036 3780
rect 21868 3726 21982 3778
rect 22034 3726 22036 3778
rect 21868 3724 22036 3726
rect 21980 3714 22036 3724
rect 22204 2996 22260 4844
rect 22316 4834 22372 4844
rect 22428 4338 22484 4956
rect 22540 5012 22596 5022
rect 22540 5010 22820 5012
rect 22540 4958 22542 5010
rect 22594 4958 22820 5010
rect 22540 4956 22820 4958
rect 22540 4946 22596 4956
rect 22764 4564 22820 4956
rect 22876 4564 22932 4574
rect 22764 4508 22876 4564
rect 22932 4508 23044 4564
rect 22876 4470 22932 4508
rect 22652 4452 22708 4462
rect 22652 4450 22820 4452
rect 22652 4398 22654 4450
rect 22706 4398 22820 4450
rect 22652 4396 22820 4398
rect 22652 4386 22708 4396
rect 22428 4286 22430 4338
rect 22482 4286 22484 4338
rect 22428 4004 22484 4286
rect 22428 3938 22484 3948
rect 22316 3442 22372 3454
rect 22316 3390 22318 3442
rect 22370 3390 22372 3442
rect 22316 3220 22372 3390
rect 22652 3444 22708 3482
rect 22652 3378 22708 3388
rect 22316 3154 22372 3164
rect 22204 2930 22260 2940
rect 22428 2994 22484 3006
rect 22428 2942 22430 2994
rect 22482 2942 22484 2994
rect 22428 800 22484 2942
rect 22764 1428 22820 4396
rect 22988 4450 23044 4508
rect 22988 4398 22990 4450
rect 23042 4398 23044 4450
rect 22988 4386 23044 4398
rect 23100 4452 23156 4462
rect 23100 4358 23156 4396
rect 23212 4450 23268 4462
rect 23212 4398 23214 4450
rect 23266 4398 23268 4450
rect 22876 4340 22932 4350
rect 22876 3388 22932 4284
rect 22988 4116 23044 4126
rect 22988 3780 23044 4060
rect 22988 3554 23044 3724
rect 22988 3502 22990 3554
rect 23042 3502 23044 3554
rect 22988 3490 23044 3502
rect 22876 3332 23156 3388
rect 22764 1362 22820 1372
rect 23100 800 23156 3332
rect 23212 2884 23268 4398
rect 23212 2818 23268 2828
rect 23324 3220 23380 5292
rect 23548 5236 23604 5246
rect 23324 2660 23380 3164
rect 23324 2594 23380 2604
rect 23436 3666 23492 3678
rect 23436 3614 23438 3666
rect 23490 3614 23492 3666
rect 23436 2436 23492 3614
rect 23548 3388 23604 5180
rect 23660 5234 23716 5404
rect 23660 5182 23662 5234
rect 23714 5182 23716 5234
rect 23660 5170 23716 5182
rect 23772 4676 23828 5628
rect 23772 4338 23828 4620
rect 23772 4286 23774 4338
rect 23826 4286 23828 4338
rect 23772 4274 23828 4286
rect 23884 3388 23940 5964
rect 23996 5926 24052 5964
rect 23996 4452 24052 4462
rect 24220 4452 24276 8876
rect 24332 8930 24500 8932
rect 24332 8878 24334 8930
rect 24386 8878 24500 8930
rect 24332 8876 24500 8878
rect 24332 8866 24388 8876
rect 24332 7362 24388 7374
rect 24332 7310 24334 7362
rect 24386 7310 24388 7362
rect 24332 6916 24388 7310
rect 24444 7028 24500 8876
rect 24556 8370 24612 10780
rect 25004 10770 25060 10780
rect 24780 10612 24836 10622
rect 24780 10518 24836 10556
rect 25228 10612 25284 10622
rect 24668 10052 24724 10062
rect 24668 9268 24724 9996
rect 24668 9174 24724 9212
rect 25228 9266 25284 10556
rect 25340 9716 25396 11342
rect 25676 10834 25732 11676
rect 25900 11508 25956 11518
rect 25676 10782 25678 10834
rect 25730 10782 25732 10834
rect 25676 10770 25732 10782
rect 25788 10836 25844 10846
rect 25788 10742 25844 10780
rect 25900 10834 25956 11452
rect 26124 11284 26180 11294
rect 26124 11190 26180 11228
rect 25900 10782 25902 10834
rect 25954 10782 25956 10834
rect 25900 10770 25956 10782
rect 26236 10612 26292 12124
rect 26236 10518 26292 10556
rect 26348 12180 26404 12190
rect 25340 9650 25396 9660
rect 26124 9716 26180 9726
rect 25676 9492 25732 9502
rect 25564 9436 25676 9492
rect 25228 9214 25230 9266
rect 25282 9214 25284 9266
rect 25228 9202 25284 9214
rect 25452 9268 25508 9278
rect 24556 8318 24558 8370
rect 24610 8318 24612 8370
rect 24556 8306 24612 8318
rect 25004 9044 25060 9054
rect 24780 7700 24836 7710
rect 24780 7606 24836 7644
rect 24444 6962 24500 6972
rect 24332 6850 24388 6860
rect 24332 6132 24388 6142
rect 24332 6020 24388 6076
rect 24332 6018 24612 6020
rect 24332 5966 24334 6018
rect 24386 5966 24612 6018
rect 24332 5964 24612 5966
rect 24332 5954 24388 5964
rect 24332 4452 24388 4462
rect 24220 4450 24388 4452
rect 24220 4398 24334 4450
rect 24386 4398 24388 4450
rect 24220 4396 24388 4398
rect 23996 4358 24052 4396
rect 24332 4116 24388 4396
rect 24332 4050 24388 4060
rect 23548 3332 23828 3388
rect 23884 3332 24052 3388
rect 23436 2370 23492 2380
rect 23772 800 23828 3332
rect 23996 1764 24052 3332
rect 24108 3330 24164 3342
rect 24108 3278 24110 3330
rect 24162 3278 24164 3330
rect 24108 3108 24164 3278
rect 24108 3042 24164 3052
rect 23996 1708 24500 1764
rect 24444 800 24500 1708
rect 24556 980 24612 5964
rect 24668 6018 24724 6030
rect 24668 5966 24670 6018
rect 24722 5966 24724 6018
rect 24668 5348 24724 5966
rect 24668 5282 24724 5292
rect 24668 4450 24724 4462
rect 24668 4398 24670 4450
rect 24722 4398 24724 4450
rect 24668 2772 24724 4398
rect 25004 3666 25060 8988
rect 25452 9042 25508 9212
rect 25452 8990 25454 9042
rect 25506 8990 25508 9042
rect 25452 8978 25508 8990
rect 25340 8036 25396 8046
rect 25228 8034 25396 8036
rect 25228 7982 25342 8034
rect 25394 7982 25396 8034
rect 25228 7980 25396 7982
rect 25116 5684 25172 5694
rect 25116 3778 25172 5628
rect 25228 5348 25284 7980
rect 25340 7970 25396 7980
rect 25564 7588 25620 9436
rect 25676 9426 25732 9436
rect 26124 9042 26180 9660
rect 26124 8990 26126 9042
rect 26178 8990 26180 9042
rect 26124 8978 26180 8990
rect 26348 8820 26404 12124
rect 26684 11732 26740 12686
rect 26684 10276 26740 11676
rect 26908 11172 26964 15820
rect 27020 13970 27076 16942
rect 27020 13918 27022 13970
rect 27074 13918 27076 13970
rect 27020 13906 27076 13918
rect 27132 16884 27188 16894
rect 27132 12852 27188 16828
rect 27244 15876 27300 17052
rect 27580 17042 27636 17052
rect 28140 17042 28196 17052
rect 28588 16884 28644 16894
rect 28700 16884 28756 17500
rect 29372 17108 29428 18398
rect 29596 17556 29652 17566
rect 29596 17462 29652 17500
rect 29372 17042 29428 17052
rect 28476 16882 28756 16884
rect 28476 16830 28590 16882
rect 28642 16830 28756 16882
rect 28476 16828 28756 16830
rect 30156 16996 30212 17006
rect 27916 16212 27972 16222
rect 28252 16212 28308 16222
rect 27916 16210 28308 16212
rect 27916 16158 27918 16210
rect 27970 16158 28254 16210
rect 28306 16158 28308 16210
rect 27916 16156 28308 16158
rect 27916 16146 27972 16156
rect 28252 16146 28308 16156
rect 27244 15426 27300 15820
rect 27244 15374 27246 15426
rect 27298 15374 27300 15426
rect 27244 15362 27300 15374
rect 27356 15988 27412 15998
rect 27356 15148 27412 15932
rect 28364 15988 28420 15998
rect 27244 15092 27412 15148
rect 28140 15876 28196 15886
rect 27244 14308 27300 15092
rect 27244 14214 27300 14252
rect 28140 13970 28196 15820
rect 28364 15874 28420 15932
rect 28364 15822 28366 15874
rect 28418 15822 28420 15874
rect 28364 15810 28420 15822
rect 28252 14420 28308 14430
rect 28252 14326 28308 14364
rect 28140 13918 28142 13970
rect 28194 13918 28196 13970
rect 28140 13906 28196 13918
rect 27132 12786 27188 12796
rect 27244 13858 27300 13870
rect 27244 13806 27246 13858
rect 27298 13806 27300 13858
rect 27244 11844 27300 13806
rect 27916 13860 27972 13870
rect 27916 13858 28084 13860
rect 27916 13806 27918 13858
rect 27970 13806 28084 13858
rect 27916 13804 28084 13806
rect 27916 13794 27972 13804
rect 27356 13748 27412 13758
rect 27356 13654 27412 13692
rect 27804 13748 27860 13758
rect 27804 12850 27860 13692
rect 27804 12798 27806 12850
rect 27858 12798 27860 12850
rect 27804 12786 27860 12798
rect 27916 12852 27972 12862
rect 27916 12178 27972 12796
rect 27916 12126 27918 12178
rect 27970 12126 27972 12178
rect 27468 11844 27524 11854
rect 27244 11778 27300 11788
rect 27356 11788 27468 11844
rect 26796 10836 26852 10846
rect 26908 10836 26964 11116
rect 26796 10834 26964 10836
rect 26796 10782 26798 10834
rect 26850 10782 26964 10834
rect 26796 10780 26964 10782
rect 26796 10770 26852 10780
rect 26908 10612 26964 10780
rect 26908 10546 26964 10556
rect 26684 10220 26964 10276
rect 26908 9714 26964 10220
rect 26908 9662 26910 9714
rect 26962 9662 26964 9714
rect 26908 9650 26964 9662
rect 27244 9604 27300 9614
rect 27020 9602 27300 9604
rect 27020 9550 27246 9602
rect 27298 9550 27300 9602
rect 27020 9548 27300 9550
rect 26572 9156 26628 9166
rect 27020 9156 27076 9548
rect 27244 9538 27300 9548
rect 27356 9156 27412 11788
rect 27468 11778 27524 11788
rect 27916 11284 27972 12126
rect 28028 12068 28084 13804
rect 28476 13746 28532 16828
rect 28588 16818 28644 16828
rect 29260 16770 29316 16782
rect 29260 16718 29262 16770
rect 29314 16718 29316 16770
rect 29260 16210 29316 16718
rect 30156 16212 30212 16940
rect 31388 16772 31444 16782
rect 31724 16772 31780 16782
rect 31388 16770 31780 16772
rect 31388 16718 31390 16770
rect 31442 16718 31726 16770
rect 31778 16718 31780 16770
rect 31388 16716 31780 16718
rect 31388 16706 31444 16716
rect 31724 16706 31780 16716
rect 29260 16158 29262 16210
rect 29314 16158 29316 16210
rect 29260 16146 29316 16158
rect 29372 16210 30212 16212
rect 29372 16158 30158 16210
rect 30210 16158 30212 16210
rect 29372 16156 30212 16158
rect 29372 16098 29428 16156
rect 30156 16146 30212 16156
rect 29372 16046 29374 16098
rect 29426 16046 29428 16098
rect 29372 16034 29428 16046
rect 31500 16100 31556 16110
rect 29148 15874 29204 15886
rect 29148 15822 29150 15874
rect 29202 15822 29204 15874
rect 29148 14420 29204 15822
rect 29596 15876 29652 15886
rect 29596 15782 29652 15820
rect 30828 15314 30884 15326
rect 30828 15262 30830 15314
rect 30882 15262 30884 15314
rect 30828 15148 30884 15262
rect 31388 15202 31444 15214
rect 31388 15150 31390 15202
rect 31442 15150 31444 15202
rect 31388 15148 31444 15150
rect 30828 15092 31444 15148
rect 29148 14326 29204 14364
rect 30940 14420 30996 14430
rect 30940 14418 31220 14420
rect 30940 14366 30942 14418
rect 30994 14366 31220 14418
rect 30940 14364 31220 14366
rect 30940 14354 30996 14364
rect 28588 14308 28644 14318
rect 28588 14214 28644 14252
rect 29260 14306 29316 14318
rect 29260 14254 29262 14306
rect 29314 14254 29316 14306
rect 29148 13860 29204 13870
rect 29260 13860 29316 14254
rect 29372 14306 29428 14318
rect 29372 14254 29374 14306
rect 29426 14254 29428 14306
rect 29372 14196 29428 14254
rect 29372 14130 29428 14140
rect 29484 14308 29540 14318
rect 29148 13858 29316 13860
rect 29148 13806 29150 13858
rect 29202 13806 29316 13858
rect 29148 13804 29316 13806
rect 29148 13794 29204 13804
rect 28476 13694 28478 13746
rect 28530 13694 28532 13746
rect 28476 13682 28532 13694
rect 28140 12852 28196 12862
rect 29148 12852 29204 12862
rect 28140 12850 28308 12852
rect 28140 12798 28142 12850
rect 28194 12798 28308 12850
rect 28140 12796 28308 12798
rect 28140 12786 28196 12796
rect 28252 12516 28308 12796
rect 29148 12758 29204 12796
rect 29484 12850 29540 14252
rect 29596 14306 29652 14318
rect 29596 14254 29598 14306
rect 29650 14254 29652 14306
rect 29596 13524 29652 14254
rect 30156 14306 30212 14318
rect 30156 14254 30158 14306
rect 30210 14254 30212 14306
rect 30156 14196 30212 14254
rect 30156 14130 30212 14140
rect 30828 14306 30884 14318
rect 30828 14254 30830 14306
rect 30882 14254 30884 14306
rect 30828 14196 30884 14254
rect 30828 14130 30884 14140
rect 31164 13636 31220 14364
rect 31276 14308 31332 15092
rect 31388 14532 31444 14542
rect 31500 14532 31556 16044
rect 31388 14530 31556 14532
rect 31388 14478 31390 14530
rect 31442 14478 31556 14530
rect 31388 14476 31556 14478
rect 31388 14466 31444 14476
rect 31276 14252 31444 14308
rect 31276 13636 31332 13646
rect 31164 13634 31332 13636
rect 31164 13582 31278 13634
rect 31330 13582 31332 13634
rect 31164 13580 31332 13582
rect 31276 13570 31332 13580
rect 29596 13458 29652 13468
rect 29484 12798 29486 12850
rect 29538 12798 29540 12850
rect 29484 12786 29540 12798
rect 31388 12740 31444 14252
rect 31388 12674 31444 12684
rect 28252 12402 28308 12460
rect 28252 12350 28254 12402
rect 28306 12350 28308 12402
rect 28252 12338 28308 12350
rect 31500 12292 31556 12302
rect 29260 12180 29316 12190
rect 29260 12178 29428 12180
rect 29260 12126 29262 12178
rect 29314 12126 29428 12178
rect 29260 12124 29428 12126
rect 29260 12114 29316 12124
rect 28028 12012 28308 12068
rect 28252 11508 28308 12012
rect 28252 11414 28308 11452
rect 27916 11228 28420 11284
rect 28140 10724 28196 10734
rect 28140 10610 28196 10668
rect 28140 10558 28142 10610
rect 28194 10558 28196 10610
rect 28140 10546 28196 10558
rect 27804 10500 27860 10510
rect 27804 10498 27972 10500
rect 27804 10446 27806 10498
rect 27858 10446 27972 10498
rect 27804 10444 27972 10446
rect 27804 10434 27860 10444
rect 27804 9604 27860 9614
rect 25900 8764 26404 8820
rect 26460 9100 26572 9156
rect 25788 8036 25844 8046
rect 25788 7942 25844 7980
rect 25452 7532 25620 7588
rect 25676 7698 25732 7710
rect 25676 7646 25678 7698
rect 25730 7646 25732 7698
rect 25676 7588 25732 7646
rect 25900 7698 25956 8764
rect 26348 8258 26404 8270
rect 26348 8206 26350 8258
rect 26402 8206 26404 8258
rect 25900 7646 25902 7698
rect 25954 7646 25956 7698
rect 25788 7588 25844 7598
rect 25676 7532 25788 7588
rect 25340 7476 25396 7486
rect 25340 7382 25396 7420
rect 25340 7028 25396 7038
rect 25340 5572 25396 6972
rect 25452 5794 25508 7532
rect 25788 7522 25844 7532
rect 25788 7364 25844 7374
rect 25788 7270 25844 7308
rect 25564 6804 25620 6814
rect 25900 6804 25956 7646
rect 26236 8034 26292 8046
rect 26236 7982 26238 8034
rect 26290 7982 26292 8034
rect 26236 7700 26292 7982
rect 26236 7634 26292 7644
rect 25564 6802 25956 6804
rect 25564 6750 25566 6802
rect 25618 6750 25956 6802
rect 25564 6748 25956 6750
rect 26012 7588 26068 7598
rect 25564 6738 25620 6748
rect 26012 6692 26068 7532
rect 26348 7474 26404 8206
rect 26348 7422 26350 7474
rect 26402 7422 26404 7474
rect 26348 7028 26404 7422
rect 26348 6962 26404 6972
rect 26236 6804 26292 6814
rect 26236 6710 26292 6748
rect 26124 6692 26180 6702
rect 26012 6690 26180 6692
rect 26012 6638 26126 6690
rect 26178 6638 26180 6690
rect 26012 6636 26180 6638
rect 25900 6580 25956 6590
rect 25564 6018 25620 6030
rect 25564 5966 25566 6018
rect 25618 5966 25620 6018
rect 25564 5908 25620 5966
rect 25564 5842 25620 5852
rect 25452 5742 25454 5794
rect 25506 5742 25508 5794
rect 25452 5730 25508 5742
rect 25788 5684 25844 5694
rect 25340 5516 25508 5572
rect 25228 5292 25396 5348
rect 25228 5124 25284 5134
rect 25228 4338 25284 5068
rect 25228 4286 25230 4338
rect 25282 4286 25284 4338
rect 25228 4274 25284 4286
rect 25116 3726 25118 3778
rect 25170 3726 25172 3778
rect 25116 3714 25172 3726
rect 25004 3614 25006 3666
rect 25058 3614 25060 3666
rect 25004 3602 25060 3614
rect 24780 3556 24836 3566
rect 24780 3462 24836 3500
rect 25340 3556 25396 5292
rect 25340 3490 25396 3500
rect 25452 4788 25508 5516
rect 25788 5460 25844 5628
rect 25788 5394 25844 5404
rect 25788 5236 25844 5246
rect 25900 5236 25956 6524
rect 26124 6018 26180 6636
rect 26348 6692 26404 6702
rect 26460 6692 26516 9100
rect 26572 9090 26628 9100
rect 26684 9100 27076 9156
rect 27132 9100 27412 9156
rect 27692 9602 27860 9604
rect 27692 9550 27806 9602
rect 27858 9550 27860 9602
rect 27692 9548 27860 9550
rect 26572 7588 26628 7598
rect 26572 7494 26628 7532
rect 26684 7476 26740 9100
rect 26908 8932 26964 8942
rect 26908 8838 26964 8876
rect 26796 8484 26852 8494
rect 26796 8258 26852 8428
rect 26908 8372 26964 8382
rect 26908 8278 26964 8316
rect 26796 8206 26798 8258
rect 26850 8206 26852 8258
rect 26796 8194 26852 8206
rect 27020 8034 27076 8046
rect 27020 7982 27022 8034
rect 27074 7982 27076 8034
rect 27020 7700 27076 7982
rect 27020 7634 27076 7644
rect 26908 7476 26964 7486
rect 26684 7474 26964 7476
rect 26684 7422 26910 7474
rect 26962 7422 26964 7474
rect 26684 7420 26964 7422
rect 26348 6690 26516 6692
rect 26348 6638 26350 6690
rect 26402 6638 26516 6690
rect 26348 6636 26516 6638
rect 26796 7028 26852 7038
rect 26796 6690 26852 6972
rect 26908 6804 26964 7420
rect 26908 6738 26964 6748
rect 26796 6638 26798 6690
rect 26850 6638 26852 6690
rect 26348 6580 26404 6636
rect 26348 6514 26404 6524
rect 26796 6580 26852 6638
rect 27020 6580 27076 6590
rect 26796 6578 27076 6580
rect 26796 6526 27022 6578
rect 27074 6526 27076 6578
rect 26796 6524 27076 6526
rect 26460 6356 26516 6366
rect 26348 6132 26404 6142
rect 26348 6038 26404 6076
rect 26124 5966 26126 6018
rect 26178 5966 26180 6018
rect 26124 5954 26180 5966
rect 26236 5794 26292 5806
rect 26236 5742 26238 5794
rect 26290 5742 26292 5794
rect 26236 5684 26292 5742
rect 26236 5618 26292 5628
rect 25788 5234 25956 5236
rect 25788 5182 25790 5234
rect 25842 5182 25956 5234
rect 25788 5180 25956 5182
rect 26460 5234 26516 6300
rect 26796 5906 26852 6524
rect 27020 6514 27076 6524
rect 26796 5854 26798 5906
rect 26850 5854 26852 5906
rect 26796 5842 26852 5854
rect 27020 6244 27076 6254
rect 26908 5796 26964 5806
rect 26684 5684 26740 5694
rect 26572 5460 26628 5470
rect 26572 5346 26628 5404
rect 26572 5294 26574 5346
rect 26626 5294 26628 5346
rect 26572 5282 26628 5294
rect 26460 5182 26462 5234
rect 26514 5182 26516 5234
rect 25788 5170 25844 5180
rect 26460 5170 26516 5182
rect 26348 4900 26404 4910
rect 25452 3554 25508 4732
rect 26236 4898 26404 4900
rect 26236 4846 26350 4898
rect 26402 4846 26404 4898
rect 26236 4844 26404 4846
rect 25788 4340 25844 4350
rect 25452 3502 25454 3554
rect 25506 3502 25508 3554
rect 25452 3490 25508 3502
rect 25676 3668 25732 3678
rect 24668 2706 24724 2716
rect 25676 1764 25732 3612
rect 25788 3442 25844 4284
rect 26012 4228 26068 4238
rect 26012 4134 26068 4172
rect 26124 3780 26180 3790
rect 26124 3556 26180 3724
rect 26124 3462 26180 3500
rect 25788 3390 25790 3442
rect 25842 3390 25844 3442
rect 25788 3378 25844 3390
rect 26236 2884 26292 4844
rect 26348 4834 26404 4844
rect 26236 2818 26292 2828
rect 26348 4116 26404 4126
rect 26348 1764 26404 4060
rect 26460 3444 26516 3454
rect 26684 3444 26740 5628
rect 26796 5460 26852 5470
rect 26796 5348 26852 5404
rect 26908 5348 26964 5740
rect 26796 5292 26964 5348
rect 26908 5010 26964 5292
rect 26908 4958 26910 5010
rect 26962 4958 26964 5010
rect 26908 4946 26964 4958
rect 27020 4788 27076 6188
rect 27132 6132 27188 9100
rect 27580 8932 27636 8942
rect 27244 8708 27300 8718
rect 27244 7812 27300 8652
rect 27356 8372 27412 8382
rect 27356 8278 27412 8316
rect 27580 8370 27636 8876
rect 27580 8318 27582 8370
rect 27634 8318 27636 8370
rect 27580 8306 27636 8318
rect 27244 6690 27300 7756
rect 27580 8034 27636 8046
rect 27580 7982 27582 8034
rect 27634 7982 27636 8034
rect 27468 7362 27524 7374
rect 27468 7310 27470 7362
rect 27522 7310 27524 7362
rect 27468 7252 27524 7310
rect 27468 7186 27524 7196
rect 27580 7140 27636 7982
rect 27580 7074 27636 7084
rect 27244 6638 27246 6690
rect 27298 6638 27300 6690
rect 27244 6626 27300 6638
rect 27692 6468 27748 9548
rect 27804 9538 27860 9548
rect 27804 7700 27860 7710
rect 27804 7606 27860 7644
rect 27916 6916 27972 10444
rect 27916 6850 27972 6860
rect 28028 10164 28084 10174
rect 27468 6412 27748 6468
rect 27804 6804 27860 6814
rect 27468 6244 27524 6412
rect 27132 5124 27188 6076
rect 27356 6188 27524 6244
rect 27244 5796 27300 5806
rect 27244 5702 27300 5740
rect 27132 5058 27188 5068
rect 27244 5460 27300 5470
rect 27244 5122 27300 5404
rect 27244 5070 27246 5122
rect 27298 5070 27300 5122
rect 27244 5058 27300 5070
rect 26908 4732 27076 4788
rect 27132 4900 27188 4910
rect 26908 3668 26964 4732
rect 26908 3554 26964 3612
rect 26908 3502 26910 3554
rect 26962 3502 26964 3554
rect 26908 3490 26964 3502
rect 27020 4004 27076 4014
rect 26460 3442 26740 3444
rect 26460 3390 26462 3442
rect 26514 3390 26740 3442
rect 26460 3388 26740 3390
rect 26460 3378 26516 3388
rect 27020 1764 27076 3948
rect 27132 3442 27188 4844
rect 27356 4788 27412 6188
rect 27804 6132 27860 6748
rect 27916 6692 27972 6702
rect 27916 6598 27972 6636
rect 27916 6132 27972 6142
rect 27804 6130 27972 6132
rect 27804 6078 27918 6130
rect 27970 6078 27972 6130
rect 27804 6076 27972 6078
rect 27916 6066 27972 6076
rect 27132 3390 27134 3442
rect 27186 3390 27188 3442
rect 27132 3378 27188 3390
rect 27244 4732 27412 4788
rect 27468 6018 27524 6030
rect 27468 5966 27470 6018
rect 27522 5966 27524 6018
rect 27244 3108 27300 4732
rect 27468 3388 27524 5966
rect 27580 5796 27636 5806
rect 28028 5796 28084 10108
rect 28252 9602 28308 9614
rect 28252 9550 28254 9602
rect 28306 9550 28308 9602
rect 28252 8708 28308 9550
rect 28252 8642 28308 8652
rect 28140 8484 28196 8494
rect 28140 8390 28196 8428
rect 28252 8146 28308 8158
rect 28252 8094 28254 8146
rect 28306 8094 28308 8146
rect 28140 8034 28196 8046
rect 28140 7982 28142 8034
rect 28194 7982 28196 8034
rect 28140 7924 28196 7982
rect 28140 7252 28196 7868
rect 28252 7588 28308 8094
rect 28364 7698 28420 11228
rect 29372 10724 29428 12124
rect 29932 12066 29988 12078
rect 29932 12014 29934 12066
rect 29986 12014 29988 12066
rect 29932 11506 29988 12014
rect 29932 11454 29934 11506
rect 29986 11454 29988 11506
rect 29932 11442 29988 11454
rect 31500 11394 31556 12236
rect 31724 11956 31780 11966
rect 31500 11342 31502 11394
rect 31554 11342 31556 11394
rect 31500 11330 31556 11342
rect 31612 11900 31724 11956
rect 30044 11284 30100 11294
rect 30044 11190 30100 11228
rect 31388 11284 31444 11294
rect 31388 11190 31444 11228
rect 29820 11170 29876 11182
rect 29820 11118 29822 11170
rect 29874 11118 29876 11170
rect 29484 10724 29540 10734
rect 29372 10668 29484 10724
rect 28812 10500 28868 10510
rect 28812 10498 29204 10500
rect 28812 10446 28814 10498
rect 28866 10446 29204 10498
rect 28812 10444 29204 10446
rect 28812 10434 28868 10444
rect 29148 10050 29204 10444
rect 29148 9998 29150 10050
rect 29202 9998 29204 10050
rect 29148 9986 29204 9998
rect 28812 9828 28868 9838
rect 28868 9772 28980 9828
rect 28812 9762 28868 9772
rect 28700 9604 28756 9614
rect 28588 9602 28756 9604
rect 28588 9550 28702 9602
rect 28754 9550 28756 9602
rect 28588 9548 28756 9550
rect 28364 7646 28366 7698
rect 28418 7646 28420 7698
rect 28364 7634 28420 7646
rect 28476 8036 28532 8046
rect 28252 7522 28308 7532
rect 28140 7186 28196 7196
rect 28476 7028 28532 7980
rect 28588 7476 28644 9548
rect 28700 9538 28756 9548
rect 28700 8708 28756 8718
rect 28700 7476 28756 8652
rect 28812 8372 28868 8382
rect 28812 7700 28868 8316
rect 28924 8260 28980 9772
rect 29260 9602 29316 9614
rect 29260 9550 29262 9602
rect 29314 9550 29316 9602
rect 29036 9380 29092 9390
rect 29092 9324 29204 9380
rect 29036 9314 29092 9324
rect 29036 8932 29092 8942
rect 29036 8484 29092 8876
rect 29036 8418 29092 8428
rect 29036 8260 29092 8270
rect 28924 8258 29092 8260
rect 28924 8206 29038 8258
rect 29090 8206 29092 8258
rect 28924 8204 29092 8206
rect 29036 8194 29092 8204
rect 28812 7588 28868 7644
rect 29036 7924 29092 7934
rect 28812 7532 28980 7588
rect 28700 7420 28868 7476
rect 28588 7410 28644 7420
rect 28364 6972 28532 7028
rect 28588 7252 28644 7262
rect 28140 6916 28196 6926
rect 28140 6580 28196 6860
rect 28140 6514 28196 6524
rect 28252 6804 28308 6814
rect 28252 6690 28308 6748
rect 28252 6638 28254 6690
rect 28306 6638 28308 6690
rect 28252 5906 28308 6638
rect 28252 5854 28254 5906
rect 28306 5854 28308 5906
rect 28252 5842 28308 5854
rect 27580 5794 28084 5796
rect 27580 5742 27582 5794
rect 27634 5742 28084 5794
rect 27580 5740 28084 5742
rect 27580 5730 27636 5740
rect 28028 5572 28084 5582
rect 28084 5516 28196 5572
rect 28028 5506 28084 5516
rect 27804 5348 27860 5358
rect 27580 5236 27636 5246
rect 27580 5122 27636 5180
rect 27804 5234 27860 5292
rect 27804 5182 27806 5234
rect 27858 5182 27860 5234
rect 27804 5170 27860 5182
rect 27916 5236 27972 5246
rect 27916 5142 27972 5180
rect 27580 5070 27582 5122
rect 27634 5070 27636 5122
rect 27580 5058 27636 5070
rect 28028 5124 28084 5134
rect 28140 5124 28196 5516
rect 28364 5234 28420 6972
rect 28588 6916 28644 7196
rect 28476 6860 28644 6916
rect 28700 7250 28756 7262
rect 28700 7198 28702 7250
rect 28754 7198 28756 7250
rect 28476 6802 28532 6860
rect 28476 6750 28478 6802
rect 28530 6750 28532 6802
rect 28476 6738 28532 6750
rect 28588 6692 28644 6702
rect 28476 6580 28532 6590
rect 28476 5906 28532 6524
rect 28476 5854 28478 5906
rect 28530 5854 28532 5906
rect 28476 5842 28532 5854
rect 28588 5572 28644 6636
rect 28700 6468 28756 7198
rect 28700 6402 28756 6412
rect 28364 5182 28366 5234
rect 28418 5182 28420 5234
rect 28364 5170 28420 5182
rect 28476 5516 28644 5572
rect 28252 5124 28308 5134
rect 28140 5122 28308 5124
rect 28140 5070 28254 5122
rect 28306 5070 28308 5122
rect 28140 5068 28308 5070
rect 28476 5124 28532 5516
rect 28588 5348 28644 5358
rect 28588 5346 28756 5348
rect 28588 5294 28590 5346
rect 28642 5294 28756 5346
rect 28588 5292 28756 5294
rect 28588 5282 28644 5292
rect 28700 5236 28756 5292
rect 28700 5170 28756 5180
rect 28476 5068 28644 5124
rect 28028 4228 28084 5068
rect 28252 5058 28308 5068
rect 28140 4228 28196 4238
rect 28028 4226 28196 4228
rect 28028 4174 28142 4226
rect 28194 4174 28196 4226
rect 28028 4172 28196 4174
rect 28140 4162 28196 4172
rect 27692 3892 27748 3902
rect 27356 3332 27524 3388
rect 27580 3554 27636 3566
rect 27580 3502 27582 3554
rect 27634 3502 27636 3554
rect 27356 3266 27412 3276
rect 27580 3108 27636 3502
rect 27244 3052 27636 3108
rect 27580 2324 27636 3052
rect 27580 2258 27636 2268
rect 27692 1764 27748 3836
rect 28588 3892 28644 5068
rect 28812 5012 28868 7420
rect 28924 7474 28980 7532
rect 28924 7422 28926 7474
rect 28978 7422 28980 7474
rect 28924 7410 28980 7422
rect 28924 7028 28980 7038
rect 28924 6130 28980 6972
rect 29036 6356 29092 7868
rect 29148 7700 29204 9324
rect 29260 9044 29316 9550
rect 29260 8978 29316 8988
rect 29372 9044 29428 10668
rect 29484 10658 29540 10668
rect 29484 10500 29540 10510
rect 29484 10050 29540 10444
rect 29820 10164 29876 11118
rect 31276 11170 31332 11182
rect 31276 11118 31278 11170
rect 31330 11118 31332 11170
rect 31276 11060 31332 11118
rect 30940 10836 30996 10846
rect 29820 10098 29876 10108
rect 30156 10612 30212 10622
rect 29484 9998 29486 10050
rect 29538 9998 29540 10050
rect 29484 9986 29540 9998
rect 30156 9940 30212 10556
rect 30940 10498 30996 10780
rect 30940 10446 30942 10498
rect 30994 10446 30996 10498
rect 30940 10434 30996 10446
rect 31276 10610 31332 11004
rect 31500 10836 31556 10846
rect 31612 10836 31668 11900
rect 31724 11890 31780 11900
rect 31836 11508 31892 18620
rect 31948 18452 32004 18958
rect 31948 18386 32004 18396
rect 32172 18338 32228 19406
rect 32172 18286 32174 18338
rect 32226 18286 32228 18338
rect 32172 18274 32228 18286
rect 32284 19012 32340 19022
rect 32284 17780 32340 18956
rect 31948 17724 32340 17780
rect 31948 14532 32004 17724
rect 32396 17108 32452 20526
rect 32508 19906 32564 20974
rect 32508 19854 32510 19906
rect 32562 19854 32564 19906
rect 32508 19842 32564 19854
rect 32508 17108 32564 17118
rect 32172 17052 32508 17108
rect 32060 16996 32116 17006
rect 32060 16902 32116 16940
rect 32172 16100 32228 17052
rect 32508 17014 32564 17052
rect 32172 16006 32228 16044
rect 32620 15764 32676 24892
rect 35308 24834 35364 24846
rect 35308 24782 35310 24834
rect 35362 24782 35364 24834
rect 34972 24724 35028 24734
rect 35196 24724 35252 24734
rect 34972 24630 35028 24668
rect 35084 24722 35252 24724
rect 35084 24670 35198 24722
rect 35250 24670 35252 24722
rect 35084 24668 35252 24670
rect 34076 24164 34132 24174
rect 34076 24050 34132 24108
rect 35084 24052 35140 24668
rect 35196 24658 35252 24668
rect 35308 24724 35364 24782
rect 35532 24836 35588 24846
rect 35532 24742 35588 24780
rect 35308 24658 35364 24668
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 34076 23998 34078 24050
rect 34130 23998 34132 24050
rect 34076 23986 34132 23998
rect 34636 23996 35140 24052
rect 35756 24164 35812 24174
rect 34524 23940 34580 23950
rect 34524 23846 34580 23884
rect 34076 23156 34132 23166
rect 34076 23062 34132 23100
rect 33852 23044 33908 23054
rect 33628 23042 33908 23044
rect 33628 22990 33854 23042
rect 33906 22990 33908 23042
rect 33628 22988 33908 22990
rect 33404 21588 33460 21598
rect 32956 21028 33012 21038
rect 32956 21026 33236 21028
rect 32956 20974 32958 21026
rect 33010 20974 33236 21026
rect 32956 20972 33236 20974
rect 32956 20962 33012 20972
rect 33180 20914 33236 20972
rect 33180 20862 33182 20914
rect 33234 20862 33236 20914
rect 33180 20850 33236 20862
rect 32956 20580 33012 20590
rect 32956 20486 33012 20524
rect 33404 20242 33460 21532
rect 33404 20190 33406 20242
rect 33458 20190 33460 20242
rect 33404 20178 33460 20190
rect 33516 20690 33572 20702
rect 33516 20638 33518 20690
rect 33570 20638 33572 20690
rect 33516 20132 33572 20638
rect 33516 20066 33572 20076
rect 33292 19906 33348 19918
rect 33292 19854 33294 19906
rect 33346 19854 33348 19906
rect 32844 19458 32900 19470
rect 32844 19406 32846 19458
rect 32898 19406 32900 19458
rect 32844 19348 32900 19406
rect 33068 19348 33124 19358
rect 32844 19346 33124 19348
rect 32844 19294 33070 19346
rect 33122 19294 33124 19346
rect 32844 19292 33124 19294
rect 33068 19282 33124 19292
rect 32732 19012 32788 19022
rect 33292 19012 33348 19854
rect 32732 19010 33348 19012
rect 32732 18958 32734 19010
rect 32786 18958 33348 19010
rect 32732 18956 33348 18958
rect 33404 19124 33460 19134
rect 33628 19124 33684 22988
rect 33852 22978 33908 22988
rect 34636 22596 34692 23996
rect 35644 23940 35700 23950
rect 35084 23938 35700 23940
rect 35084 23886 35646 23938
rect 35698 23886 35700 23938
rect 35084 23884 35700 23886
rect 34860 23714 34916 23726
rect 34860 23662 34862 23714
rect 34914 23662 34916 23714
rect 34860 23604 34916 23662
rect 34860 23538 34916 23548
rect 34860 23380 34916 23390
rect 34524 22540 34692 22596
rect 34748 23324 34860 23380
rect 34412 22484 34468 22494
rect 34412 22390 34468 22428
rect 33964 22148 34020 22158
rect 33964 22054 34020 22092
rect 33964 20916 34020 20926
rect 33852 20860 33964 20916
rect 33852 20242 33908 20860
rect 33964 20850 34020 20860
rect 34300 20690 34356 20702
rect 34300 20638 34302 20690
rect 34354 20638 34356 20690
rect 33852 20190 33854 20242
rect 33906 20190 33908 20242
rect 33852 20178 33908 20190
rect 34076 20578 34132 20590
rect 34076 20526 34078 20578
rect 34130 20526 34132 20578
rect 33740 20020 33796 20030
rect 33740 19926 33796 19964
rect 34076 19908 34132 20526
rect 34300 20242 34356 20638
rect 34524 20578 34580 22540
rect 34748 22372 34804 23324
rect 34860 23314 34916 23324
rect 34972 23154 35028 23166
rect 34972 23102 34974 23154
rect 35026 23102 35028 23154
rect 34972 23044 35028 23102
rect 34972 22978 35028 22988
rect 34636 22316 34804 22372
rect 34860 22820 34916 22830
rect 34636 20916 34692 22316
rect 34748 22148 34804 22158
rect 34860 22148 34916 22764
rect 34748 22146 34916 22148
rect 34748 22094 34750 22146
rect 34802 22094 34916 22146
rect 34748 22092 34916 22094
rect 34972 22146 35028 22158
rect 34972 22094 34974 22146
rect 35026 22094 35028 22146
rect 34748 22082 34804 22092
rect 34972 21812 35028 22094
rect 34748 21756 35028 21812
rect 34748 21364 34804 21756
rect 35084 21700 35140 23884
rect 35644 23874 35700 23884
rect 35756 23826 35812 24108
rect 35756 23774 35758 23826
rect 35810 23774 35812 23826
rect 35756 23762 35812 23774
rect 35420 23716 35476 23726
rect 35420 23622 35476 23660
rect 35868 23492 35924 27134
rect 36092 26908 36148 27694
rect 36204 27074 36260 29036
rect 37100 28754 37156 29036
rect 37100 28702 37102 28754
rect 37154 28702 37156 28754
rect 37100 28690 37156 28702
rect 36988 28084 37044 28094
rect 36988 27990 37044 28028
rect 37436 28084 37492 67172
rect 37996 55468 38052 76300
rect 38108 76290 38164 76300
rect 38220 75684 38276 76524
rect 38668 76356 38724 76366
rect 38668 76262 38724 76300
rect 38556 75908 38612 75918
rect 38556 75794 38612 75852
rect 38556 75742 38558 75794
rect 38610 75742 38612 75794
rect 38556 75730 38612 75742
rect 39004 75796 39060 76636
rect 39228 76690 40068 76692
rect 39228 76638 39230 76690
rect 39282 76638 40068 76690
rect 39228 76636 40068 76638
rect 39228 76626 39284 76636
rect 38220 75590 38276 75628
rect 38892 75684 38948 75694
rect 38892 75122 38948 75628
rect 39004 75682 39060 75740
rect 40012 75794 40068 76636
rect 40012 75742 40014 75794
rect 40066 75742 40068 75794
rect 40012 75730 40068 75742
rect 40124 76690 40180 79200
rect 40124 76638 40126 76690
rect 40178 76638 40180 76690
rect 39004 75630 39006 75682
rect 39058 75630 39060 75682
rect 39004 75618 39060 75630
rect 39564 75684 39620 75694
rect 40124 75684 40180 76638
rect 40796 76692 40852 79200
rect 41020 76692 41076 76702
rect 40796 76636 41020 76692
rect 41020 76598 41076 76636
rect 41468 76580 41524 79200
rect 42028 76692 42084 76702
rect 42140 76692 42196 79200
rect 42812 77026 42868 79200
rect 42812 76974 42814 77026
rect 42866 76974 42868 77026
rect 42812 76962 42868 76974
rect 43484 77028 43540 79200
rect 43484 76962 43540 76972
rect 43596 77026 43652 77038
rect 43596 76974 43598 77026
rect 43650 76974 43652 77026
rect 42364 76692 42420 76702
rect 43596 76692 43652 76974
rect 42140 76690 42532 76692
rect 42140 76638 42366 76690
rect 42418 76638 42532 76690
rect 42140 76636 42532 76638
rect 42028 76598 42084 76636
rect 42364 76626 42420 76636
rect 41468 76524 41748 76580
rect 39564 75682 39956 75684
rect 39564 75630 39566 75682
rect 39618 75630 39956 75682
rect 39564 75628 39956 75630
rect 39564 75618 39620 75628
rect 38892 75070 38894 75122
rect 38946 75070 38948 75122
rect 38892 75058 38948 75070
rect 37884 55412 38052 55468
rect 39788 74788 39844 74798
rect 37884 43708 37940 55412
rect 37884 43652 38164 43708
rect 38108 28084 38164 43652
rect 39788 38668 39844 74732
rect 39900 67228 39956 75628
rect 40124 75618 40180 75628
rect 40684 76354 40740 76366
rect 40684 76302 40686 76354
rect 40738 76302 40740 76354
rect 39900 67172 40180 67228
rect 39788 38612 39956 38668
rect 39788 28532 39844 28542
rect 37436 28082 37828 28084
rect 37436 28030 37438 28082
rect 37490 28030 37828 28082
rect 37436 28028 37828 28030
rect 37436 28018 37492 28028
rect 36204 27022 36206 27074
rect 36258 27022 36260 27074
rect 36204 27010 36260 27022
rect 36428 27970 36484 27982
rect 36428 27918 36430 27970
rect 36482 27918 36484 27970
rect 36428 26962 36484 27918
rect 37772 27858 37828 28028
rect 37772 27806 37774 27858
rect 37826 27806 37828 27858
rect 37772 27794 37828 27806
rect 37548 27074 37604 27086
rect 37548 27022 37550 27074
rect 37602 27022 37604 27074
rect 36428 26910 36430 26962
rect 36482 26910 36484 26962
rect 36092 26852 36260 26908
rect 36092 26290 36148 26302
rect 36092 26238 36094 26290
rect 36146 26238 36148 26290
rect 35980 25618 36036 25630
rect 35980 25566 35982 25618
rect 36034 25566 36036 25618
rect 35980 25284 36036 25566
rect 35980 25218 36036 25228
rect 35980 24836 36036 24846
rect 35980 24722 36036 24780
rect 35980 24670 35982 24722
rect 36034 24670 36036 24722
rect 35980 24658 36036 24670
rect 35980 23940 36036 23950
rect 36092 23940 36148 26238
rect 36204 24834 36260 26852
rect 36204 24782 36206 24834
rect 36258 24782 36260 24834
rect 36204 24770 36260 24782
rect 36316 26852 36372 26862
rect 35980 23938 36148 23940
rect 35980 23886 35982 23938
rect 36034 23886 36148 23938
rect 35980 23884 36148 23886
rect 35980 23874 36036 23884
rect 36204 23826 36260 23838
rect 36204 23774 36206 23826
rect 36258 23774 36260 23826
rect 35868 23436 36036 23492
rect 35756 23156 35812 23166
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 35756 22594 35812 23100
rect 35756 22542 35758 22594
rect 35810 22542 35812 22594
rect 35756 22530 35812 22542
rect 35196 22372 35252 22382
rect 35196 22258 35252 22316
rect 35196 22206 35198 22258
rect 35250 22206 35252 22258
rect 35196 22194 35252 22206
rect 35308 22258 35364 22270
rect 35308 22206 35310 22258
rect 35362 22206 35364 22258
rect 35196 21700 35252 21710
rect 35084 21698 35252 21700
rect 35084 21646 35198 21698
rect 35250 21646 35252 21698
rect 35084 21644 35252 21646
rect 35196 21634 35252 21644
rect 34972 21588 35028 21598
rect 34972 21494 35028 21532
rect 34860 21476 34916 21486
rect 34860 21382 34916 21420
rect 35308 21364 35364 22206
rect 35868 22260 35924 22270
rect 35868 22166 35924 22204
rect 35756 22148 35812 22158
rect 35756 22054 35812 22092
rect 35980 22036 36036 23436
rect 36204 23380 36260 23774
rect 36204 23314 36260 23324
rect 36316 23826 36372 26796
rect 36428 26404 36484 26910
rect 36988 26962 37044 26974
rect 36988 26910 36990 26962
rect 37042 26910 37044 26962
rect 36428 26338 36484 26348
rect 36652 26514 36708 26526
rect 36652 26462 36654 26514
rect 36706 26462 36708 26514
rect 36652 25508 36708 26462
rect 36988 26516 37044 26910
rect 37548 26908 37604 27022
rect 38108 27074 38164 28028
rect 38668 28084 38724 28094
rect 39340 28084 39396 28094
rect 38668 28082 38948 28084
rect 38668 28030 38670 28082
rect 38722 28030 38948 28082
rect 38668 28028 38948 28030
rect 38668 28018 38724 28028
rect 38108 27022 38110 27074
rect 38162 27022 38164 27074
rect 38108 27010 38164 27022
rect 38220 27970 38276 27982
rect 38220 27918 38222 27970
rect 38274 27918 38276 27970
rect 38220 26962 38276 27918
rect 38780 27858 38836 27870
rect 38780 27806 38782 27858
rect 38834 27806 38836 27858
rect 38668 27636 38724 27646
rect 38220 26910 38222 26962
rect 38274 26910 38276 26962
rect 38220 26908 38276 26910
rect 37548 26852 38276 26908
rect 36988 26180 37044 26460
rect 37996 26402 38052 26414
rect 37996 26350 37998 26402
rect 38050 26350 38052 26402
rect 36988 26114 37044 26124
rect 37212 26292 37268 26302
rect 36652 25442 36708 25452
rect 37212 25620 37268 26236
rect 37660 26290 37716 26302
rect 37660 26238 37662 26290
rect 37714 26238 37716 26290
rect 37212 25506 37268 25564
rect 37212 25454 37214 25506
rect 37266 25454 37268 25506
rect 37212 25442 37268 25454
rect 37324 25844 37380 25854
rect 36652 25284 36708 25294
rect 36652 24276 36708 25228
rect 36876 24948 36932 24958
rect 36876 24854 36932 24892
rect 36540 24220 36708 24276
rect 37212 24276 37268 24286
rect 36540 24164 36596 24220
rect 36316 23774 36318 23826
rect 36370 23774 36372 23826
rect 36316 23268 36372 23774
rect 36316 23202 36372 23212
rect 36428 24108 36596 24164
rect 36428 23266 36484 24108
rect 36652 24052 36708 24062
rect 36428 23214 36430 23266
rect 36482 23214 36484 23266
rect 36428 23202 36484 23214
rect 36540 23714 36596 23726
rect 36540 23662 36542 23714
rect 36594 23662 36596 23714
rect 36540 23154 36596 23662
rect 36540 23102 36542 23154
rect 36594 23102 36596 23154
rect 36540 23090 36596 23102
rect 36316 23044 36372 23054
rect 36316 22484 36372 22988
rect 35868 21980 36036 22036
rect 36204 22258 36260 22270
rect 36204 22206 36206 22258
rect 36258 22206 36260 22258
rect 35420 21588 35476 21598
rect 35420 21494 35476 21532
rect 35644 21586 35700 21598
rect 35644 21534 35646 21586
rect 35698 21534 35700 21586
rect 35308 21308 35588 21364
rect 34748 21298 34804 21308
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 35532 21028 35588 21308
rect 35308 20972 35588 21028
rect 35084 20916 35140 20926
rect 34636 20860 35028 20916
rect 34636 20692 34692 20702
rect 34636 20598 34692 20636
rect 34860 20692 34916 20702
rect 34860 20598 34916 20636
rect 34524 20526 34526 20578
rect 34578 20526 34580 20578
rect 34524 20514 34580 20526
rect 34300 20190 34302 20242
rect 34354 20190 34356 20242
rect 34300 20178 34356 20190
rect 34636 20356 34692 20366
rect 34188 19908 34244 19918
rect 34076 19906 34244 19908
rect 34076 19854 34190 19906
rect 34242 19854 34244 19906
rect 34076 19852 34244 19854
rect 34188 19796 34244 19852
rect 34188 19730 34244 19740
rect 34076 19684 34132 19694
rect 33964 19628 34076 19684
rect 33964 19458 34020 19628
rect 34076 19618 34132 19628
rect 33964 19406 33966 19458
rect 34018 19406 34020 19458
rect 33964 19394 34020 19406
rect 34636 19234 34692 20300
rect 34972 20132 35028 20860
rect 35084 20802 35140 20860
rect 35308 20914 35364 20972
rect 35308 20862 35310 20914
rect 35362 20862 35364 20914
rect 35308 20850 35364 20862
rect 35084 20750 35086 20802
rect 35138 20750 35140 20802
rect 35084 20738 35140 20750
rect 35196 20804 35252 20814
rect 35084 20132 35140 20142
rect 34972 20130 35140 20132
rect 34972 20078 35086 20130
rect 35138 20078 35140 20130
rect 34972 20076 35140 20078
rect 35084 20066 35140 20076
rect 34860 20018 34916 20030
rect 34860 19966 34862 20018
rect 34914 19966 34916 20018
rect 34860 19684 34916 19966
rect 35196 20018 35252 20748
rect 35532 20804 35588 20814
rect 35532 20710 35588 20748
rect 35644 20802 35700 21534
rect 35644 20750 35646 20802
rect 35698 20750 35700 20802
rect 35644 20692 35700 20750
rect 35532 20132 35588 20142
rect 35644 20132 35700 20636
rect 35532 20130 35700 20132
rect 35532 20078 35534 20130
rect 35586 20078 35700 20130
rect 35532 20076 35700 20078
rect 35756 20580 35812 20590
rect 35532 20066 35588 20076
rect 35196 19966 35198 20018
rect 35250 19966 35252 20018
rect 35196 19954 35252 19966
rect 34860 19618 34916 19628
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 35644 19460 35700 19470
rect 35420 19404 35644 19460
rect 35420 19346 35476 19404
rect 35644 19394 35700 19404
rect 35420 19294 35422 19346
rect 35474 19294 35476 19346
rect 35420 19282 35476 19294
rect 34636 19182 34638 19234
rect 34690 19182 34692 19234
rect 34636 19170 34692 19182
rect 34972 19236 35028 19246
rect 33628 19068 33796 19124
rect 32732 18676 32788 18956
rect 33404 18788 33460 19068
rect 33404 18722 33460 18732
rect 32732 18610 32788 18620
rect 33628 18452 33684 18462
rect 32956 17668 33012 17678
rect 32956 17332 33012 17612
rect 33628 17666 33684 18396
rect 33628 17614 33630 17666
rect 33682 17614 33684 17666
rect 33628 17602 33684 17614
rect 32956 17266 33012 17276
rect 33740 16996 33796 19068
rect 33852 19122 33908 19134
rect 33852 19070 33854 19122
rect 33906 19070 33908 19122
rect 33852 19012 33908 19070
rect 33852 18946 33908 18956
rect 34300 19124 34356 19134
rect 33852 17556 33908 17566
rect 33852 17106 33908 17500
rect 33852 17054 33854 17106
rect 33906 17054 33908 17106
rect 33852 17042 33908 17054
rect 34300 17106 34356 19068
rect 34972 19122 35028 19180
rect 35644 19236 35700 19246
rect 34972 19070 34974 19122
rect 35026 19070 35028 19122
rect 34972 19058 35028 19070
rect 35308 19124 35364 19134
rect 35308 19030 35364 19068
rect 35196 18340 35252 18350
rect 35084 18284 35196 18340
rect 34300 17054 34302 17106
rect 34354 17054 34356 17106
rect 34300 17042 34356 17054
rect 34524 17108 34580 17118
rect 35084 17108 35140 18284
rect 35196 18274 35252 18284
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 35420 17780 35476 17790
rect 35308 17556 35364 17566
rect 35308 17462 35364 17500
rect 35420 17332 35476 17724
rect 35644 17780 35700 19180
rect 35644 17666 35700 17724
rect 35644 17614 35646 17666
rect 35698 17614 35700 17666
rect 35644 17602 35700 17614
rect 35532 17444 35588 17454
rect 35756 17444 35812 20524
rect 35868 20130 35924 21980
rect 35980 21698 36036 21710
rect 35980 21646 35982 21698
rect 36034 21646 36036 21698
rect 35980 21588 36036 21646
rect 35980 20804 36036 21532
rect 35980 20738 36036 20748
rect 36092 20692 36148 20702
rect 36092 20598 36148 20636
rect 35868 20078 35870 20130
rect 35922 20078 35924 20130
rect 35868 20066 35924 20078
rect 36204 19460 36260 22206
rect 36316 22258 36372 22428
rect 36316 22206 36318 22258
rect 36370 22206 36372 22258
rect 36316 22194 36372 22206
rect 36540 22146 36596 22158
rect 36540 22094 36542 22146
rect 36594 22094 36596 22146
rect 36316 21588 36372 21598
rect 36540 21588 36596 22094
rect 36316 21586 36484 21588
rect 36316 21534 36318 21586
rect 36370 21534 36484 21586
rect 36316 21532 36484 21534
rect 36316 21522 36372 21532
rect 36316 21364 36372 21374
rect 36428 21364 36484 21532
rect 36540 21522 36596 21532
rect 36428 21308 36596 21364
rect 36316 20018 36372 21308
rect 36428 20916 36484 20926
rect 36428 20802 36484 20860
rect 36428 20750 36430 20802
rect 36482 20750 36484 20802
rect 36428 20738 36484 20750
rect 36540 20356 36596 21308
rect 36540 20290 36596 20300
rect 36316 19966 36318 20018
rect 36370 19966 36372 20018
rect 36316 19954 36372 19966
rect 35980 19404 36260 19460
rect 36652 19460 36708 23996
rect 37212 23940 37268 24220
rect 37100 23826 37156 23838
rect 37100 23774 37102 23826
rect 37154 23774 37156 23826
rect 36988 23492 37044 23502
rect 36764 23268 36820 23278
rect 36764 21700 36820 23212
rect 36988 22708 37044 23436
rect 36988 22642 37044 22652
rect 36876 22260 36932 22270
rect 36876 21924 36932 22204
rect 36876 21868 37044 21924
rect 36876 21700 36932 21710
rect 36764 21698 36932 21700
rect 36764 21646 36878 21698
rect 36930 21646 36932 21698
rect 36764 21644 36932 21646
rect 36876 21634 36932 21644
rect 35532 17442 35812 17444
rect 35532 17390 35534 17442
rect 35586 17390 35812 17442
rect 35532 17388 35812 17390
rect 35868 19124 35924 19134
rect 35868 17666 35924 19068
rect 35868 17614 35870 17666
rect 35922 17614 35924 17666
rect 35532 17378 35588 17388
rect 35420 17266 35476 17276
rect 35196 17108 35252 17118
rect 34580 17106 35252 17108
rect 34580 17054 35198 17106
rect 35250 17054 35252 17106
rect 34580 17052 35252 17054
rect 33628 16940 33796 16996
rect 33516 16884 33572 16894
rect 33516 16212 33572 16828
rect 33628 16548 33684 16940
rect 33740 16772 33796 16782
rect 33740 16770 33908 16772
rect 33740 16718 33742 16770
rect 33794 16718 33908 16770
rect 33740 16716 33908 16718
rect 33740 16706 33796 16716
rect 33628 16492 33796 16548
rect 33516 16146 33572 16156
rect 32844 15988 32900 15998
rect 32844 15986 33124 15988
rect 32844 15934 32846 15986
rect 32898 15934 33124 15986
rect 32844 15932 33124 15934
rect 32844 15922 32900 15932
rect 32620 15708 32900 15764
rect 32844 15540 32900 15708
rect 33068 15652 33124 15932
rect 33068 15596 33572 15652
rect 32844 15484 33348 15540
rect 32956 15314 33012 15326
rect 32956 15262 32958 15314
rect 33010 15262 33012 15314
rect 32508 15204 32564 15242
rect 32956 15148 33012 15262
rect 32508 15138 32564 15148
rect 31948 14466 32004 14476
rect 32620 15092 33012 15148
rect 32060 14420 32116 14430
rect 32060 14326 32116 14364
rect 32508 13188 32564 13198
rect 32620 13188 32676 15092
rect 32508 13186 32676 13188
rect 32508 13134 32510 13186
rect 32562 13134 32676 13186
rect 32508 13132 32676 13134
rect 33068 13746 33124 13758
rect 33068 13694 33070 13746
rect 33122 13694 33124 13746
rect 33068 13186 33124 13694
rect 33068 13134 33070 13186
rect 33122 13134 33124 13186
rect 32508 13122 32564 13132
rect 33068 13122 33124 13134
rect 32620 12964 32676 12974
rect 33180 12964 33236 12974
rect 32620 12962 33180 12964
rect 32620 12910 32622 12962
rect 32674 12910 33180 12962
rect 32620 12908 33180 12910
rect 32620 12898 32676 12908
rect 33180 12870 33236 12908
rect 32508 12740 32564 12750
rect 32508 12738 32788 12740
rect 32508 12686 32510 12738
rect 32562 12686 32788 12738
rect 32508 12684 32788 12686
rect 32508 12674 32564 12684
rect 32060 12292 32116 12302
rect 32060 12066 32116 12236
rect 32060 12014 32062 12066
rect 32114 12014 32116 12066
rect 32060 12002 32116 12014
rect 31836 11442 31892 11452
rect 31556 10780 31668 10836
rect 31948 11394 32004 11406
rect 31948 11342 31950 11394
rect 32002 11342 32004 11394
rect 31948 11284 32004 11342
rect 32396 11396 32452 11406
rect 32396 11302 32452 11340
rect 31500 10742 31556 10780
rect 31276 10558 31278 10610
rect 31330 10558 31332 10610
rect 30156 9874 30212 9884
rect 30268 10050 30324 10062
rect 30268 9998 30270 10050
rect 30322 9998 30324 10050
rect 30044 9604 30100 9614
rect 29932 9602 30100 9604
rect 29932 9550 30046 9602
rect 30098 9550 30100 9602
rect 29932 9548 30100 9550
rect 29372 9042 29764 9044
rect 29372 8990 29374 9042
rect 29426 8990 29764 9042
rect 29372 8988 29764 8990
rect 29372 8978 29428 8988
rect 29484 8820 29540 8830
rect 29260 8260 29316 8270
rect 29260 8146 29316 8204
rect 29260 8094 29262 8146
rect 29314 8094 29316 8146
rect 29260 8082 29316 8094
rect 29372 8146 29428 8158
rect 29372 8094 29374 8146
rect 29426 8094 29428 8146
rect 29260 7700 29316 7710
rect 29148 7698 29316 7700
rect 29148 7646 29262 7698
rect 29314 7646 29316 7698
rect 29148 7644 29316 7646
rect 29260 7634 29316 7644
rect 29260 7476 29316 7486
rect 29148 7420 29260 7476
rect 29148 6468 29204 7420
rect 29260 7410 29316 7420
rect 29372 6916 29428 8094
rect 29484 7700 29540 8764
rect 29484 7634 29540 7644
rect 29260 6860 29428 6916
rect 29596 7250 29652 7262
rect 29596 7198 29598 7250
rect 29650 7198 29652 7250
rect 29596 6916 29652 7198
rect 29260 6804 29316 6860
rect 29260 6738 29316 6748
rect 29372 6692 29428 6702
rect 29596 6692 29652 6860
rect 29372 6690 29652 6692
rect 29372 6638 29374 6690
rect 29426 6638 29652 6690
rect 29372 6636 29652 6638
rect 29372 6626 29428 6636
rect 29596 6468 29652 6478
rect 29148 6466 29652 6468
rect 29148 6414 29598 6466
rect 29650 6414 29652 6466
rect 29148 6412 29652 6414
rect 29596 6402 29652 6412
rect 29036 6290 29092 6300
rect 28924 6078 28926 6130
rect 28978 6078 28980 6130
rect 28924 5236 28980 6078
rect 29036 6020 29092 6030
rect 29092 5964 29204 6020
rect 29036 5954 29092 5964
rect 28924 5170 28980 5180
rect 29148 5124 29204 5964
rect 29260 5908 29316 5918
rect 29260 5460 29316 5852
rect 29708 5906 29764 8988
rect 29820 8260 29876 8270
rect 29820 7474 29876 8204
rect 29820 7422 29822 7474
rect 29874 7422 29876 7474
rect 29820 7410 29876 7422
rect 29932 6804 29988 9548
rect 30044 9538 30100 9548
rect 30156 8930 30212 8942
rect 30156 8878 30158 8930
rect 30210 8878 30212 8930
rect 30156 8370 30212 8878
rect 30268 8482 30324 9998
rect 31276 9828 31332 10558
rect 31948 10610 32004 11228
rect 32620 11284 32676 11294
rect 32620 11190 32676 11228
rect 32172 11170 32228 11182
rect 32172 11118 32174 11170
rect 32226 11118 32228 11170
rect 32172 11060 32228 11118
rect 32284 11172 32340 11182
rect 32508 11172 32564 11182
rect 32284 11170 32452 11172
rect 32284 11118 32286 11170
rect 32338 11118 32452 11170
rect 32284 11116 32452 11118
rect 32284 11106 32340 11116
rect 32172 10994 32228 11004
rect 31948 10558 31950 10610
rect 32002 10558 32004 10610
rect 31388 10500 31444 10510
rect 31388 10406 31444 10444
rect 31388 10050 31444 10062
rect 31388 9998 31390 10050
rect 31442 9998 31444 10050
rect 31388 9940 31444 9998
rect 31836 10052 31892 10062
rect 31724 9940 31780 9950
rect 31388 9938 31780 9940
rect 31388 9886 31726 9938
rect 31778 9886 31780 9938
rect 31388 9884 31780 9886
rect 31724 9874 31780 9884
rect 31276 9772 31444 9828
rect 30492 9602 30548 9614
rect 30492 9550 30494 9602
rect 30546 9550 30548 9602
rect 30268 8430 30270 8482
rect 30322 8430 30324 8482
rect 30268 8418 30324 8430
rect 30380 8484 30436 8494
rect 30156 8318 30158 8370
rect 30210 8318 30212 8370
rect 30156 8306 30212 8318
rect 30044 8034 30100 8046
rect 30044 7982 30046 8034
rect 30098 7982 30100 8034
rect 30044 7924 30100 7982
rect 30044 7858 30100 7868
rect 30380 7812 30436 8428
rect 30268 7756 30436 7812
rect 30044 7700 30100 7710
rect 30044 7606 30100 7644
rect 30268 7698 30324 7756
rect 30268 7646 30270 7698
rect 30322 7646 30324 7698
rect 30268 7028 30324 7646
rect 30380 7588 30436 7598
rect 30380 7494 30436 7532
rect 30156 6972 30324 7028
rect 30492 7476 30548 9550
rect 30940 9602 30996 9614
rect 30940 9550 30942 9602
rect 30994 9550 30996 9602
rect 30828 8034 30884 8046
rect 30828 7982 30830 8034
rect 30882 7982 30884 8034
rect 30716 7476 30772 7486
rect 30492 7474 30772 7476
rect 30492 7422 30718 7474
rect 30770 7422 30772 7474
rect 30492 7420 30772 7422
rect 29708 5854 29710 5906
rect 29762 5854 29764 5906
rect 29708 5842 29764 5854
rect 29820 6748 29988 6804
rect 30044 6916 30100 6926
rect 29820 5460 29876 6748
rect 30044 6690 30100 6860
rect 30044 6638 30046 6690
rect 30098 6638 30100 6690
rect 30044 6468 30100 6638
rect 30156 6580 30212 6972
rect 30156 6514 30212 6524
rect 30268 6804 30324 6814
rect 30268 6578 30324 6748
rect 30268 6526 30270 6578
rect 30322 6526 30324 6578
rect 30268 6514 30324 6526
rect 30044 6402 30100 6412
rect 30492 6356 30548 7420
rect 30716 7410 30772 7420
rect 30604 7140 30660 7150
rect 30604 6690 30660 7084
rect 30828 6916 30884 7982
rect 30940 7364 30996 9550
rect 31276 9602 31332 9614
rect 31276 9550 31278 9602
rect 31330 9550 31332 9602
rect 31276 9380 31332 9550
rect 31388 9604 31444 9772
rect 31836 9826 31892 9996
rect 31836 9774 31838 9826
rect 31890 9774 31892 9826
rect 31724 9716 31780 9726
rect 31612 9604 31668 9614
rect 31388 9602 31668 9604
rect 31388 9550 31614 9602
rect 31666 9550 31668 9602
rect 31388 9548 31668 9550
rect 31276 8260 31332 9324
rect 31276 8194 31332 8204
rect 31500 8146 31556 9548
rect 31612 9538 31668 9548
rect 31500 8094 31502 8146
rect 31554 8094 31556 8146
rect 31500 8082 31556 8094
rect 31276 8034 31332 8046
rect 31276 7982 31278 8034
rect 31330 7982 31332 8034
rect 31052 7588 31108 7598
rect 31052 7586 31220 7588
rect 31052 7534 31054 7586
rect 31106 7534 31220 7586
rect 31052 7532 31220 7534
rect 31052 7522 31108 7532
rect 30940 7298 30996 7308
rect 30828 6850 30884 6860
rect 31164 6804 31220 7532
rect 31276 7476 31332 7982
rect 31724 7698 31780 9660
rect 31836 9380 31892 9774
rect 31948 9828 32004 10558
rect 32396 10050 32452 11116
rect 32508 10834 32564 11116
rect 32508 10782 32510 10834
rect 32562 10782 32564 10834
rect 32508 10770 32564 10782
rect 32396 9998 32398 10050
rect 32450 9998 32452 10050
rect 32396 9986 32452 9998
rect 32284 9828 32340 9838
rect 31948 9826 32340 9828
rect 31948 9774 32286 9826
rect 32338 9774 32340 9826
rect 31948 9772 32340 9774
rect 32284 9716 32340 9772
rect 32284 9650 32340 9660
rect 31836 9324 32340 9380
rect 32284 8930 32340 9324
rect 32284 8878 32286 8930
rect 32338 8878 32340 8930
rect 32284 8866 32340 8878
rect 32396 9268 32452 9278
rect 32284 8372 32340 8382
rect 32396 8372 32452 9212
rect 32732 8932 32788 12684
rect 33068 12738 33124 12750
rect 33068 12686 33070 12738
rect 33122 12686 33124 12738
rect 33068 12180 33124 12686
rect 33068 12114 33124 12124
rect 33292 11620 33348 15484
rect 33516 15538 33572 15596
rect 33516 15486 33518 15538
rect 33570 15486 33572 15538
rect 33516 15474 33572 15486
rect 33404 15428 33460 15438
rect 33404 15334 33460 15372
rect 33628 15314 33684 15326
rect 33628 15262 33630 15314
rect 33682 15262 33684 15314
rect 33404 14420 33460 14430
rect 33460 14364 33572 14420
rect 33404 14354 33460 14364
rect 33404 13972 33460 13982
rect 33404 13878 33460 13916
rect 33516 13970 33572 14364
rect 33516 13918 33518 13970
rect 33570 13918 33572 13970
rect 33516 13906 33572 13918
rect 33628 13970 33684 15262
rect 33628 13918 33630 13970
rect 33682 13918 33684 13970
rect 33628 13860 33684 13918
rect 33628 13794 33684 13804
rect 33740 13076 33796 16492
rect 33852 15204 33908 16716
rect 34188 16770 34244 16782
rect 34188 16718 34190 16770
rect 34242 16718 34244 16770
rect 34076 15652 34132 15662
rect 34188 15652 34244 16718
rect 34132 15596 34244 15652
rect 34076 15538 34132 15596
rect 34076 15486 34078 15538
rect 34130 15486 34132 15538
rect 34076 15474 34132 15486
rect 34524 15538 34580 17052
rect 35196 17042 35252 17052
rect 34636 16882 34692 16894
rect 34636 16830 34638 16882
rect 34690 16830 34692 16882
rect 34636 16772 34692 16830
rect 34748 16884 34804 16894
rect 34748 16790 34804 16828
rect 35644 16882 35700 16894
rect 35644 16830 35646 16882
rect 35698 16830 35700 16882
rect 34636 16706 34692 16716
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 34972 16212 35028 16222
rect 34972 16210 35364 16212
rect 34972 16158 34974 16210
rect 35026 16158 35364 16210
rect 34972 16156 35364 16158
rect 34972 16146 35028 16156
rect 35308 16098 35364 16156
rect 35308 16046 35310 16098
rect 35362 16046 35364 16098
rect 35308 16034 35364 16046
rect 34524 15486 34526 15538
rect 34578 15486 34580 15538
rect 34524 15474 34580 15486
rect 34636 15988 34692 15998
rect 33852 15138 33908 15148
rect 34188 14644 34244 14654
rect 34524 14644 34580 14654
rect 34188 14642 34580 14644
rect 34188 14590 34190 14642
rect 34242 14590 34526 14642
rect 34578 14590 34580 14642
rect 34188 14588 34580 14590
rect 34188 14578 34244 14588
rect 34524 14578 34580 14588
rect 34076 14532 34132 14542
rect 33964 14476 34076 14532
rect 33964 13186 34020 14476
rect 34076 14466 34132 14476
rect 34412 14308 34468 14318
rect 34188 13972 34244 13982
rect 34188 13878 34244 13916
rect 34412 13970 34468 14252
rect 34636 14084 34692 15932
rect 35420 15874 35476 15886
rect 35420 15822 35422 15874
rect 35474 15822 35476 15874
rect 34972 15764 35028 15774
rect 34636 14018 34692 14028
rect 34860 15092 34916 15102
rect 34860 14642 34916 15036
rect 34860 14590 34862 14642
rect 34914 14590 34916 14642
rect 34412 13918 34414 13970
rect 34466 13918 34468 13970
rect 34412 13748 34468 13918
rect 34860 13972 34916 14590
rect 34860 13906 34916 13916
rect 34748 13860 34804 13870
rect 34748 13766 34804 13804
rect 34412 13682 34468 13692
rect 33964 13134 33966 13186
rect 34018 13134 34020 13186
rect 33964 13122 34020 13134
rect 33292 11554 33348 11564
rect 33628 13020 33796 13076
rect 33180 11396 33236 11406
rect 33180 11394 33348 11396
rect 33180 11342 33182 11394
rect 33234 11342 33348 11394
rect 33180 11340 33348 11342
rect 33180 11330 33236 11340
rect 33180 10948 33236 10958
rect 32844 10052 32900 10062
rect 33068 10052 33124 10062
rect 32844 10050 33124 10052
rect 32844 9998 32846 10050
rect 32898 9998 33070 10050
rect 33122 9998 33124 10050
rect 32844 9996 33124 9998
rect 32844 9986 32900 9996
rect 33068 9986 33124 9996
rect 33180 9938 33236 10892
rect 33292 10724 33348 11340
rect 33628 11060 33684 13020
rect 33852 12964 33908 12974
rect 33740 12908 33852 12964
rect 33740 12402 33796 12908
rect 33852 12870 33908 12908
rect 34412 12964 34468 12974
rect 34412 12870 34468 12908
rect 34748 12964 34804 12974
rect 34748 12870 34804 12908
rect 33964 12740 34020 12750
rect 33740 12350 33742 12402
rect 33794 12350 33796 12402
rect 33740 12338 33796 12350
rect 33852 12738 34020 12740
rect 33852 12686 33966 12738
rect 34018 12686 34020 12738
rect 33852 12684 34020 12686
rect 33852 11844 33908 12684
rect 33964 12674 34020 12684
rect 34524 12738 34580 12750
rect 34524 12686 34526 12738
rect 34578 12686 34580 12738
rect 33964 12516 34020 12526
rect 33964 12178 34020 12460
rect 33964 12126 33966 12178
rect 34018 12126 34020 12178
rect 33964 12068 34020 12126
rect 33964 12002 34020 12012
rect 33852 11778 33908 11788
rect 33852 11282 33908 11294
rect 33852 11230 33854 11282
rect 33906 11230 33908 11282
rect 33740 11060 33796 11070
rect 33628 11004 33740 11060
rect 33740 10994 33796 11004
rect 33852 10948 33908 11230
rect 33852 10882 33908 10892
rect 33348 10668 34020 10724
rect 33292 10630 33348 10668
rect 33180 9886 33182 9938
rect 33234 9886 33236 9938
rect 33180 9874 33236 9886
rect 33740 9716 33796 9726
rect 33740 9622 33796 9660
rect 32844 9602 32900 9614
rect 32844 9550 32846 9602
rect 32898 9550 32900 9602
rect 32844 9268 32900 9550
rect 33292 9604 33348 9614
rect 33292 9510 33348 9548
rect 32844 9202 32900 9212
rect 32732 8866 32788 8876
rect 33292 9042 33348 9054
rect 33292 8990 33294 9042
rect 33346 8990 33348 9042
rect 32284 8370 32676 8372
rect 32284 8318 32286 8370
rect 32338 8318 32676 8370
rect 32284 8316 32676 8318
rect 32284 8306 32340 8316
rect 32620 8258 32676 8316
rect 32620 8206 32622 8258
rect 32674 8206 32676 8258
rect 32620 8194 32676 8206
rect 32844 8148 32900 8158
rect 31836 8036 31892 8046
rect 31836 8034 32004 8036
rect 31836 7982 31838 8034
rect 31890 7982 32004 8034
rect 31836 7980 32004 7982
rect 31836 7970 31892 7980
rect 31724 7646 31726 7698
rect 31778 7646 31780 7698
rect 31724 7634 31780 7646
rect 31836 7812 31892 7822
rect 31276 7420 31780 7476
rect 31500 7250 31556 7262
rect 31500 7198 31502 7250
rect 31554 7198 31556 7250
rect 31500 7028 31556 7198
rect 31500 6962 31556 6972
rect 31052 6748 31220 6804
rect 31500 6804 31556 6814
rect 30604 6638 30606 6690
rect 30658 6638 30660 6690
rect 30604 6626 30660 6638
rect 30828 6692 30884 6702
rect 30828 6598 30884 6636
rect 30268 6300 30548 6356
rect 29260 5394 29316 5404
rect 29372 5404 29876 5460
rect 29932 6132 29988 6142
rect 29260 5124 29316 5134
rect 29148 5122 29316 5124
rect 29148 5070 29262 5122
rect 29314 5070 29316 5122
rect 29148 5068 29316 5070
rect 29260 5058 29316 5068
rect 28812 4946 28868 4956
rect 28812 4452 28868 4462
rect 28812 4358 28868 4396
rect 28476 3556 28532 3566
rect 27804 3330 27860 3342
rect 27804 3278 27806 3330
rect 27858 3278 27860 3330
rect 27804 2996 27860 3278
rect 27804 2930 27860 2940
rect 25676 1708 25844 1764
rect 26348 1708 26516 1764
rect 27020 1708 27188 1764
rect 27692 1708 27860 1764
rect 24556 924 25172 980
rect 25116 800 25172 924
rect 25788 800 25844 1708
rect 26460 800 26516 1708
rect 27132 800 27188 1708
rect 27804 800 27860 1708
rect 28476 800 28532 3500
rect 28588 3554 28644 3836
rect 28588 3502 28590 3554
rect 28642 3502 28644 3554
rect 28588 3490 28644 3502
rect 28700 4338 28756 4350
rect 28700 4286 28702 4338
rect 28754 4286 28756 4338
rect 28700 3444 28756 4286
rect 29372 3554 29428 5404
rect 29596 5236 29652 5246
rect 29932 5236 29988 6076
rect 29596 5142 29652 5180
rect 29708 5180 29988 5236
rect 30044 5908 30100 5918
rect 29484 5124 29540 5134
rect 29484 5030 29540 5068
rect 29372 3502 29374 3554
rect 29426 3502 29428 3554
rect 29372 3388 29428 3502
rect 28700 3378 28756 3388
rect 28924 3330 28980 3342
rect 28924 3278 28926 3330
rect 28978 3278 28980 3330
rect 28924 3108 28980 3278
rect 28924 3042 28980 3052
rect 29260 3332 29428 3388
rect 29596 3444 29652 3454
rect 29708 3444 29764 5180
rect 29932 5012 29988 5022
rect 29596 3442 29764 3444
rect 29596 3390 29598 3442
rect 29650 3390 29764 3442
rect 29596 3388 29764 3390
rect 29820 4676 29876 4686
rect 29596 3378 29652 3388
rect 29148 2660 29204 2670
rect 29148 800 29204 2604
rect 29260 1876 29316 3332
rect 29260 1810 29316 1820
rect 29820 800 29876 4620
rect 29932 4116 29988 4956
rect 30044 4452 30100 5852
rect 30268 5796 30324 6300
rect 30604 6244 30660 6254
rect 30380 6188 30604 6244
rect 30380 6018 30436 6188
rect 30604 6178 30660 6188
rect 30380 5966 30382 6018
rect 30434 5966 30436 6018
rect 30380 5954 30436 5966
rect 30828 5908 30884 5918
rect 30268 5740 30436 5796
rect 30268 5012 30324 5022
rect 30268 4918 30324 4956
rect 30268 4676 30324 4686
rect 30044 4386 30100 4396
rect 30156 4620 30268 4676
rect 29932 4050 29988 4060
rect 30044 3556 30100 3566
rect 30156 3556 30212 4620
rect 30268 4610 30324 4620
rect 30044 3554 30212 3556
rect 30044 3502 30046 3554
rect 30098 3502 30212 3554
rect 30044 3500 30212 3502
rect 30268 4228 30324 4238
rect 30044 3490 30100 3500
rect 30268 3442 30324 4172
rect 30268 3390 30270 3442
rect 30322 3390 30324 3442
rect 30268 3378 30324 3390
rect 30380 3388 30436 5740
rect 30828 5234 30884 5852
rect 30940 5796 30996 5806
rect 30940 5346 30996 5740
rect 30940 5294 30942 5346
rect 30994 5294 30996 5346
rect 30940 5282 30996 5294
rect 30828 5182 30830 5234
rect 30882 5182 30884 5234
rect 30828 5170 30884 5182
rect 30604 5124 30660 5134
rect 30604 5030 30660 5068
rect 30716 4788 30772 4798
rect 30604 3442 30660 3454
rect 30604 3390 30606 3442
rect 30658 3390 30660 3442
rect 30380 3332 30548 3388
rect 30492 800 30548 3332
rect 30604 3220 30660 3390
rect 30716 3388 30772 4732
rect 31052 4452 31108 6748
rect 31500 6710 31556 6748
rect 31164 6580 31220 6618
rect 31164 6514 31220 6524
rect 31612 6466 31668 6478
rect 31612 6414 31614 6466
rect 31666 6414 31668 6466
rect 31164 6356 31220 6366
rect 31220 6300 31556 6356
rect 31164 6290 31220 6300
rect 31388 5236 31444 5246
rect 31388 5122 31444 5180
rect 31388 5070 31390 5122
rect 31442 5070 31444 5122
rect 31388 5058 31444 5070
rect 31388 4452 31444 4462
rect 31052 4450 31444 4452
rect 31052 4398 31390 4450
rect 31442 4398 31444 4450
rect 31052 4396 31444 4398
rect 31388 4386 31444 4396
rect 30828 4340 30884 4350
rect 30828 4246 30884 4284
rect 31388 3556 31444 3566
rect 31500 3556 31556 6300
rect 31612 5348 31668 6414
rect 31612 5282 31668 5292
rect 31724 5236 31780 7420
rect 31836 7362 31892 7756
rect 31948 7476 32004 7980
rect 32508 7586 32564 7598
rect 32508 7534 32510 7586
rect 32562 7534 32564 7586
rect 32172 7476 32228 7486
rect 31948 7474 32228 7476
rect 31948 7422 32174 7474
rect 32226 7422 32228 7474
rect 31948 7420 32228 7422
rect 31836 7310 31838 7362
rect 31890 7310 31892 7362
rect 31836 7298 31892 7310
rect 32172 6916 32228 7420
rect 32172 6850 32228 6860
rect 31836 6804 31892 6814
rect 31836 6710 31892 6748
rect 32508 6692 32564 7534
rect 32732 6804 32788 6814
rect 32732 6710 32788 6748
rect 32620 6692 32676 6702
rect 32508 6636 32620 6692
rect 32620 6598 32676 6636
rect 32844 6690 32900 8092
rect 32956 8034 33012 8046
rect 32956 7982 32958 8034
rect 33010 7982 33012 8034
rect 32956 7588 33012 7982
rect 33292 8036 33348 8990
rect 33964 9044 34020 10668
rect 34076 9602 34132 9614
rect 34076 9550 34078 9602
rect 34130 9550 34132 9602
rect 34076 9268 34132 9550
rect 34076 9202 34132 9212
rect 34524 9156 34580 12686
rect 34972 10164 35028 15708
rect 35420 15428 35476 15822
rect 35644 15764 35700 16830
rect 35868 16884 35924 17614
rect 35980 17106 36036 19404
rect 36652 19394 36708 19404
rect 36428 19236 36484 19246
rect 36428 19142 36484 19180
rect 36316 19122 36372 19134
rect 36316 19070 36318 19122
rect 36370 19070 36372 19122
rect 36316 18900 36372 19070
rect 35980 17054 35982 17106
rect 36034 17054 36036 17106
rect 35980 17042 36036 17054
rect 36092 17780 36148 17790
rect 36092 16994 36148 17724
rect 36316 17778 36372 18844
rect 36316 17726 36318 17778
rect 36370 17726 36372 17778
rect 36316 17714 36372 17726
rect 36540 18228 36596 18238
rect 36092 16942 36094 16994
rect 36146 16942 36148 16994
rect 36092 16930 36148 16942
rect 35868 16828 36036 16884
rect 35980 16772 36036 16828
rect 36204 16882 36260 16894
rect 36204 16830 36206 16882
rect 36258 16830 36260 16882
rect 36204 16772 36260 16830
rect 35980 16716 36260 16772
rect 36540 16772 36596 18172
rect 36988 17780 37044 21868
rect 37100 20580 37156 23774
rect 37212 23826 37268 23884
rect 37212 23774 37214 23826
rect 37266 23774 37268 23826
rect 37212 23762 37268 23774
rect 37324 23380 37380 25788
rect 37660 25732 37716 26238
rect 37660 25666 37716 25676
rect 37772 25508 37828 25518
rect 37772 25414 37828 25452
rect 37772 25284 37828 25294
rect 37548 25228 37772 25284
rect 37212 23324 37380 23380
rect 37436 23714 37492 23726
rect 37436 23662 37438 23714
rect 37490 23662 37492 23714
rect 37212 22148 37268 23324
rect 37324 23156 37380 23166
rect 37324 23062 37380 23100
rect 37212 22082 37268 22092
rect 37324 22932 37380 22942
rect 37324 22482 37380 22876
rect 37324 22430 37326 22482
rect 37378 22430 37380 22482
rect 37212 21924 37268 21934
rect 37212 20914 37268 21868
rect 37324 21364 37380 22430
rect 37436 22372 37492 23662
rect 37548 23266 37604 25228
rect 37772 25218 37828 25228
rect 37996 24834 38052 26350
rect 38220 26404 38276 26852
rect 38220 26338 38276 26348
rect 38556 27186 38612 27198
rect 38556 27134 38558 27186
rect 38610 27134 38612 27186
rect 38332 25508 38388 25518
rect 38332 25414 38388 25452
rect 38220 25284 38276 25294
rect 38220 25190 38276 25228
rect 37996 24782 37998 24834
rect 38050 24782 38052 24834
rect 37884 24722 37940 24734
rect 37884 24670 37886 24722
rect 37938 24670 37940 24722
rect 37884 24612 37940 24670
rect 37884 24546 37940 24556
rect 37772 24500 37828 24510
rect 37660 24052 37716 24062
rect 37660 23938 37716 23996
rect 37660 23886 37662 23938
rect 37714 23886 37716 23938
rect 37660 23874 37716 23886
rect 37772 23826 37828 24444
rect 37996 24052 38052 24782
rect 37772 23774 37774 23826
rect 37826 23774 37828 23826
rect 37772 23716 37828 23774
rect 37772 23650 37828 23660
rect 37884 23996 38052 24052
rect 37548 23214 37550 23266
rect 37602 23214 37604 23266
rect 37548 23202 37604 23214
rect 37884 22932 37940 23996
rect 38444 23940 38500 23950
rect 37996 23938 38500 23940
rect 37996 23886 38446 23938
rect 38498 23886 38500 23938
rect 37996 23884 38500 23886
rect 37996 23826 38052 23884
rect 38444 23874 38500 23884
rect 37996 23774 37998 23826
rect 38050 23774 38052 23826
rect 37996 23762 38052 23774
rect 38556 23826 38612 27134
rect 38668 25506 38724 27580
rect 38668 25454 38670 25506
rect 38722 25454 38724 25506
rect 38668 25284 38724 25454
rect 38780 27074 38836 27806
rect 38780 27022 38782 27074
rect 38834 27022 38836 27074
rect 38780 26292 38836 27022
rect 38780 25508 38836 26236
rect 38780 25442 38836 25452
rect 38668 25218 38724 25228
rect 38556 23774 38558 23826
rect 38610 23774 38612 23826
rect 38556 23762 38612 23774
rect 38892 23548 38948 28028
rect 39340 27990 39396 28028
rect 39452 27244 39732 27300
rect 39452 26908 39508 27244
rect 39676 27186 39732 27244
rect 39676 27134 39678 27186
rect 39730 27134 39732 27186
rect 39676 27122 39732 27134
rect 39788 27074 39844 28476
rect 39788 27022 39790 27074
rect 39842 27022 39844 27074
rect 39788 27010 39844 27022
rect 39452 26852 39620 26908
rect 39116 26404 39172 26414
rect 39116 25394 39172 26348
rect 39116 25342 39118 25394
rect 39170 25342 39172 25394
rect 39116 25330 39172 25342
rect 38444 23492 38948 23548
rect 39340 24834 39396 24846
rect 39340 24782 39342 24834
rect 39394 24782 39396 24834
rect 37884 22866 37940 22876
rect 38220 23378 38276 23390
rect 38220 23326 38222 23378
rect 38274 23326 38276 23378
rect 37436 22306 37492 22316
rect 37548 22708 37604 22718
rect 37548 21924 37604 22652
rect 37548 21858 37604 21868
rect 37772 22146 37828 22158
rect 37772 22094 37774 22146
rect 37826 22094 37828 22146
rect 37660 21812 37716 21822
rect 37660 21586 37716 21756
rect 37660 21534 37662 21586
rect 37714 21534 37716 21586
rect 37660 21522 37716 21534
rect 37324 21308 37716 21364
rect 37436 20916 37492 20926
rect 37212 20862 37214 20914
rect 37266 20862 37268 20914
rect 37212 20850 37268 20862
rect 37324 20860 37436 20916
rect 37100 20514 37156 20524
rect 37100 19684 37156 19694
rect 37100 19348 37156 19628
rect 37100 19282 37156 19292
rect 37324 19234 37380 20860
rect 37436 20850 37492 20860
rect 37436 20578 37492 20590
rect 37436 20526 37438 20578
rect 37490 20526 37492 20578
rect 37436 20356 37492 20526
rect 37436 20290 37492 20300
rect 37324 19182 37326 19234
rect 37378 19182 37380 19234
rect 37324 19170 37380 19182
rect 37548 20242 37604 20254
rect 37548 20190 37550 20242
rect 37602 20190 37604 20242
rect 37100 19124 37156 19134
rect 37100 19030 37156 19068
rect 37100 17780 37156 17790
rect 36988 17778 37156 17780
rect 36988 17726 37102 17778
rect 37154 17726 37156 17778
rect 36988 17724 37156 17726
rect 37100 17714 37156 17724
rect 37212 17780 37268 17790
rect 37548 17780 37604 20190
rect 37660 20018 37716 21308
rect 37772 20804 37828 22094
rect 38108 22036 38164 22046
rect 37772 20738 37828 20748
rect 37996 21980 38108 22036
rect 37772 20580 37828 20590
rect 37772 20578 37940 20580
rect 37772 20526 37774 20578
rect 37826 20526 37940 20578
rect 37772 20524 37940 20526
rect 37772 20514 37828 20524
rect 37660 19966 37662 20018
rect 37714 19966 37716 20018
rect 37660 19954 37716 19966
rect 37884 20020 37940 20524
rect 37996 20468 38052 21980
rect 38108 21970 38164 21980
rect 38108 20916 38164 20926
rect 38108 20802 38164 20860
rect 38108 20750 38110 20802
rect 38162 20750 38164 20802
rect 38108 20738 38164 20750
rect 37996 20412 38164 20468
rect 37772 19460 37828 19470
rect 37212 17666 37268 17724
rect 37212 17614 37214 17666
rect 37266 17614 37268 17666
rect 37212 17602 37268 17614
rect 37436 17724 37604 17780
rect 37660 19124 37716 19134
rect 36988 17554 37044 17566
rect 36988 17502 36990 17554
rect 37042 17502 37044 17554
rect 36988 16884 37044 17502
rect 37100 17332 37156 17342
rect 37436 17332 37492 17724
rect 37548 17556 37604 17566
rect 37660 17556 37716 19068
rect 37548 17554 37716 17556
rect 37548 17502 37550 17554
rect 37602 17502 37716 17554
rect 37548 17500 37716 17502
rect 37548 17490 37604 17500
rect 37100 17106 37156 17276
rect 37324 17276 37492 17332
rect 37100 17054 37102 17106
rect 37154 17054 37156 17106
rect 37100 16996 37156 17054
rect 37100 16930 37156 16940
rect 37212 17220 37268 17230
rect 36988 16818 37044 16828
rect 36092 16324 36148 16334
rect 36092 16210 36148 16268
rect 36092 16158 36094 16210
rect 36146 16158 36148 16210
rect 36092 16146 36148 16158
rect 36540 16210 36596 16716
rect 36540 16158 36542 16210
rect 36594 16158 36596 16210
rect 36540 16146 36596 16158
rect 36988 16324 37044 16334
rect 36988 16210 37044 16268
rect 37100 16324 37156 16334
rect 37212 16324 37268 17164
rect 37100 16322 37268 16324
rect 37100 16270 37102 16322
rect 37154 16270 37268 16322
rect 37100 16268 37268 16270
rect 37100 16258 37156 16268
rect 36988 16158 36990 16210
rect 37042 16158 37044 16210
rect 36988 16146 37044 16158
rect 35644 15698 35700 15708
rect 35420 15362 35476 15372
rect 35196 15314 35252 15326
rect 35196 15262 35198 15314
rect 35250 15262 35252 15314
rect 35196 15148 35252 15262
rect 35084 15092 35252 15148
rect 35980 15202 36036 15214
rect 35980 15150 35982 15202
rect 36034 15150 36036 15202
rect 35084 13746 35140 15092
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35980 14642 36036 15150
rect 37324 15148 37380 17276
rect 37548 17108 37604 17118
rect 37772 17108 37828 19404
rect 37884 19348 37940 19964
rect 37996 20018 38052 20030
rect 37996 19966 37998 20018
rect 38050 19966 38052 20018
rect 37996 19684 38052 19966
rect 37996 19618 38052 19628
rect 37884 19282 37940 19292
rect 38108 19346 38164 20412
rect 38108 19294 38110 19346
rect 38162 19294 38164 19346
rect 38108 19282 38164 19294
rect 37996 19236 38052 19246
rect 37996 19142 38052 19180
rect 38220 18900 38276 23326
rect 38332 22372 38388 22382
rect 38332 22278 38388 22316
rect 38444 22258 38500 23492
rect 38444 22206 38446 22258
rect 38498 22206 38500 22258
rect 38444 22194 38500 22206
rect 38668 23268 38724 23278
rect 38556 21588 38612 21598
rect 38668 21588 38724 23212
rect 39228 23154 39284 23166
rect 39228 23102 39230 23154
rect 39282 23102 39284 23154
rect 39228 22932 39284 23102
rect 39228 22866 39284 22876
rect 39228 21810 39284 21822
rect 39228 21758 39230 21810
rect 39282 21758 39284 21810
rect 39116 21588 39172 21598
rect 38556 21586 38836 21588
rect 38556 21534 38558 21586
rect 38610 21534 38836 21586
rect 38556 21532 38836 21534
rect 38556 21522 38612 21532
rect 38780 21026 38836 21532
rect 39116 21494 39172 21532
rect 39228 21252 39284 21758
rect 39228 21186 39284 21196
rect 38780 20974 38782 21026
rect 38834 20974 38836 21026
rect 38780 20962 38836 20974
rect 38892 20916 38948 20926
rect 38444 20578 38500 20590
rect 38444 20526 38446 20578
rect 38498 20526 38500 20578
rect 38332 19348 38388 19358
rect 38332 19234 38388 19292
rect 38332 19182 38334 19234
rect 38386 19182 38388 19234
rect 38332 19012 38388 19182
rect 38444 19234 38500 20526
rect 38892 20580 38948 20860
rect 38892 20514 38948 20524
rect 38444 19182 38446 19234
rect 38498 19182 38500 19234
rect 38444 19124 38500 19182
rect 38780 20356 38836 20366
rect 38668 19124 38724 19134
rect 38444 19068 38668 19124
rect 38332 18956 38500 19012
rect 38220 18844 38388 18900
rect 38220 18340 38276 18350
rect 38220 18246 38276 18284
rect 37548 17106 37828 17108
rect 37548 17054 37550 17106
rect 37602 17054 37828 17106
rect 37548 17052 37828 17054
rect 37996 17666 38052 17678
rect 37996 17614 37998 17666
rect 38050 17614 38052 17666
rect 37996 17106 38052 17614
rect 38220 17444 38276 17454
rect 37996 17054 37998 17106
rect 38050 17054 38052 17106
rect 37548 17042 37604 17052
rect 37996 17042 38052 17054
rect 38108 17442 38276 17444
rect 38108 17390 38222 17442
rect 38274 17390 38276 17442
rect 38108 17388 38276 17390
rect 37436 16882 37492 16894
rect 37436 16830 37438 16882
rect 37490 16830 37492 16882
rect 37436 16772 37492 16830
rect 37772 16884 37828 16894
rect 37772 16772 37828 16828
rect 37884 16772 37940 16782
rect 37772 16770 37940 16772
rect 37772 16718 37886 16770
rect 37938 16718 37940 16770
rect 37772 16716 37940 16718
rect 37436 16706 37492 16716
rect 37884 16706 37940 16716
rect 38108 16660 38164 17388
rect 38220 17378 38276 17388
rect 38332 17220 38388 18844
rect 38444 17666 38500 18956
rect 38444 17614 38446 17666
rect 38498 17614 38500 17666
rect 38444 17602 38500 17614
rect 38556 18452 38612 18462
rect 38108 16594 38164 16604
rect 38220 17164 38388 17220
rect 37996 16324 38052 16334
rect 37996 16230 38052 16268
rect 37548 15988 37604 15998
rect 37884 15988 37940 15998
rect 37548 15986 37828 15988
rect 37548 15934 37550 15986
rect 37602 15934 37828 15986
rect 37548 15932 37828 15934
rect 37548 15922 37604 15932
rect 35980 14590 35982 14642
rect 36034 14590 36036 14642
rect 35980 14578 36036 14590
rect 37100 15092 37380 15148
rect 37436 15874 37492 15886
rect 37436 15822 37438 15874
rect 37490 15822 37492 15874
rect 35420 14532 35476 14542
rect 35420 14438 35476 14476
rect 35868 14532 35924 14542
rect 35868 14438 35924 14476
rect 35084 13694 35086 13746
rect 35138 13694 35140 13746
rect 35084 13188 35140 13694
rect 36092 14306 36148 14318
rect 36092 14254 36094 14306
rect 36146 14254 36148 14306
rect 36092 13860 36148 14254
rect 35868 13634 35924 13646
rect 35868 13582 35870 13634
rect 35922 13582 35924 13634
rect 35756 13524 35812 13534
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35084 13122 35140 13132
rect 35420 12964 35476 12974
rect 35420 12870 35476 12908
rect 35756 12962 35812 13468
rect 35868 13074 35924 13582
rect 35868 13022 35870 13074
rect 35922 13022 35924 13074
rect 35868 13010 35924 13022
rect 35756 12910 35758 12962
rect 35810 12910 35812 12962
rect 35756 12898 35812 12910
rect 35980 12964 36036 12974
rect 36092 12964 36148 13804
rect 35980 12962 36148 12964
rect 35980 12910 35982 12962
rect 36034 12910 36148 12962
rect 35980 12908 36148 12910
rect 36204 12964 36260 12974
rect 35980 12898 36036 12908
rect 36204 12402 36260 12908
rect 36204 12350 36206 12402
rect 36258 12350 36260 12402
rect 36204 12338 36260 12350
rect 36428 12292 36484 12302
rect 36316 12290 36484 12292
rect 36316 12238 36430 12290
rect 36482 12238 36484 12290
rect 36316 12236 36484 12238
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35980 11508 36036 11518
rect 36316 11508 36372 12236
rect 36428 12226 36484 12236
rect 36988 12292 37044 12302
rect 36988 12198 37044 12236
rect 36540 12180 36596 12190
rect 36876 12180 36932 12190
rect 36540 12178 36876 12180
rect 36540 12126 36542 12178
rect 36594 12126 36876 12178
rect 36540 12124 36876 12126
rect 37100 12180 37156 15092
rect 37436 14532 37492 15822
rect 37772 15204 37828 15932
rect 37884 15894 37940 15932
rect 38108 15204 38164 15214
rect 37772 15202 38164 15204
rect 37772 15150 38110 15202
rect 38162 15150 38164 15202
rect 37772 15148 38164 15150
rect 38108 15138 38164 15148
rect 38220 14532 38276 17164
rect 38444 16324 38500 16334
rect 38556 16324 38612 18396
rect 38668 17666 38724 19068
rect 38668 17614 38670 17666
rect 38722 17614 38724 17666
rect 38668 17602 38724 17614
rect 38668 16884 38724 16894
rect 38668 16790 38724 16828
rect 38444 16322 38612 16324
rect 38444 16270 38446 16322
rect 38498 16270 38612 16322
rect 38444 16268 38612 16270
rect 38444 16258 38500 16268
rect 38780 16100 38836 20300
rect 39340 20356 39396 24782
rect 39452 20804 39508 20814
rect 39452 20710 39508 20748
rect 39340 20290 39396 20300
rect 39452 20020 39508 20030
rect 39340 20018 39508 20020
rect 39340 19966 39454 20018
rect 39506 19966 39508 20018
rect 39340 19964 39508 19966
rect 39228 19572 39284 19582
rect 39228 19348 39284 19516
rect 39116 19236 39172 19246
rect 39116 19142 39172 19180
rect 38892 19122 38948 19134
rect 38892 19070 38894 19122
rect 38946 19070 38948 19122
rect 38892 17220 38948 19070
rect 39116 19012 39172 19022
rect 39116 18918 39172 18956
rect 39116 18564 39172 18574
rect 38892 17154 38948 17164
rect 39004 18508 39116 18564
rect 39004 17106 39060 18508
rect 39116 18498 39172 18508
rect 39228 18450 39284 19292
rect 39340 19234 39396 19964
rect 39452 19954 39508 19964
rect 39340 19182 39342 19234
rect 39394 19182 39396 19234
rect 39340 19124 39396 19182
rect 39564 19236 39620 26852
rect 39676 26290 39732 26302
rect 39676 26238 39678 26290
rect 39730 26238 39732 26290
rect 39676 25730 39732 26238
rect 39676 25678 39678 25730
rect 39730 25678 39732 25730
rect 39676 25666 39732 25678
rect 39788 26178 39844 26190
rect 39788 26126 39790 26178
rect 39842 26126 39844 26178
rect 39676 25284 39732 25294
rect 39676 25190 39732 25228
rect 39676 24722 39732 24734
rect 39676 24670 39678 24722
rect 39730 24670 39732 24722
rect 39676 24612 39732 24670
rect 39676 24546 39732 24556
rect 39676 23268 39732 23278
rect 39676 23174 39732 23212
rect 39788 21700 39844 26126
rect 39900 21924 39956 38612
rect 40012 26964 40068 27002
rect 40012 26898 40068 26908
rect 40012 26292 40068 26302
rect 40012 26198 40068 26236
rect 40124 25730 40180 67172
rect 40684 28532 40740 76302
rect 41468 75794 41524 76524
rect 41468 75742 41470 75794
rect 41522 75742 41524 75794
rect 41468 75730 41524 75742
rect 41580 76354 41636 76366
rect 41580 76302 41582 76354
rect 41634 76302 41636 76354
rect 40908 75684 40964 75694
rect 40908 75590 40964 75628
rect 41580 67228 41636 76302
rect 41692 75682 41748 76524
rect 42476 75794 42532 76636
rect 43372 76690 43652 76692
rect 43372 76638 43598 76690
rect 43650 76638 43652 76690
rect 43372 76636 43652 76638
rect 42476 75742 42478 75794
rect 42530 75742 42532 75794
rect 42476 75730 42532 75742
rect 42812 76354 42868 76366
rect 42812 76302 42814 76354
rect 42866 76302 42868 76354
rect 41692 75630 41694 75682
rect 41746 75630 41748 75682
rect 41692 75618 41748 75630
rect 42028 75458 42084 75470
rect 42028 75406 42030 75458
rect 42082 75406 42084 75458
rect 42028 67228 42084 75406
rect 41580 67172 41748 67228
rect 42028 67172 42196 67228
rect 41244 38948 41300 38958
rect 41244 38854 41300 38892
rect 41468 38946 41524 38958
rect 41468 38894 41470 38946
rect 41522 38894 41524 38946
rect 41132 38724 41188 38734
rect 41468 38724 41524 38894
rect 41580 38836 41636 38846
rect 41580 38742 41636 38780
rect 41132 38722 41468 38724
rect 41132 38670 41134 38722
rect 41186 38670 41468 38722
rect 41132 38668 41468 38670
rect 41132 38658 41188 38668
rect 41468 38658 41524 38668
rect 40684 28466 40740 28476
rect 41020 28084 41076 28094
rect 40572 28082 41076 28084
rect 40572 28030 41022 28082
rect 41074 28030 41076 28082
rect 40572 28028 41076 28030
rect 40124 25678 40126 25730
rect 40178 25678 40180 25730
rect 40124 25618 40180 25678
rect 40124 25566 40126 25618
rect 40178 25566 40180 25618
rect 40124 25554 40180 25566
rect 40236 27972 40292 27982
rect 40124 24724 40180 24734
rect 40236 24724 40292 27916
rect 40348 27860 40404 27870
rect 40348 27766 40404 27804
rect 40460 25620 40516 25630
rect 40460 25506 40516 25564
rect 40460 25454 40462 25506
rect 40514 25454 40516 25506
rect 40460 25442 40516 25454
rect 40124 24722 40292 24724
rect 40124 24670 40126 24722
rect 40178 24670 40292 24722
rect 40124 24668 40292 24670
rect 40348 24836 40404 24846
rect 40124 24388 40180 24668
rect 40124 24322 40180 24332
rect 40348 24164 40404 24780
rect 40236 24108 40404 24164
rect 40236 24052 40292 24108
rect 40124 23996 40292 24052
rect 40012 23044 40068 23054
rect 40012 22146 40068 22988
rect 40012 22094 40014 22146
rect 40066 22094 40068 22146
rect 40012 22082 40068 22094
rect 39900 21868 40068 21924
rect 39900 21700 39956 21710
rect 39788 21698 39956 21700
rect 39788 21646 39902 21698
rect 39954 21646 39956 21698
rect 39788 21644 39956 21646
rect 39900 21634 39956 21644
rect 40012 21252 40068 21868
rect 39788 21196 40068 21252
rect 39676 20020 39732 20030
rect 39676 19926 39732 19964
rect 39564 19170 39620 19180
rect 39340 19058 39396 19068
rect 39788 19012 39844 21196
rect 40124 20802 40180 23996
rect 40348 23940 40404 23950
rect 40348 23846 40404 23884
rect 40236 23828 40292 23838
rect 40236 23714 40292 23772
rect 40236 23662 40238 23714
rect 40290 23662 40292 23714
rect 40236 23650 40292 23662
rect 40460 23826 40516 23838
rect 40460 23774 40462 23826
rect 40514 23774 40516 23826
rect 40460 23268 40516 23774
rect 40348 22708 40404 22718
rect 40348 22370 40404 22652
rect 40348 22318 40350 22370
rect 40402 22318 40404 22370
rect 40348 22306 40404 22318
rect 40460 22258 40516 23212
rect 40460 22206 40462 22258
rect 40514 22206 40516 22258
rect 40460 22194 40516 22206
rect 40124 20750 40126 20802
rect 40178 20750 40180 20802
rect 40124 20738 40180 20750
rect 39900 20580 39956 20590
rect 39900 20486 39956 20524
rect 39900 20244 39956 20254
rect 39900 20242 40180 20244
rect 39900 20190 39902 20242
rect 39954 20190 40180 20242
rect 39900 20188 40180 20190
rect 39900 20178 39956 20188
rect 40012 20018 40068 20030
rect 40012 19966 40014 20018
rect 40066 19966 40068 20018
rect 40012 19460 40068 19966
rect 40012 19394 40068 19404
rect 39452 18956 39844 19012
rect 39900 19122 39956 19134
rect 39900 19070 39902 19122
rect 39954 19070 39956 19122
rect 39228 18398 39230 18450
rect 39282 18398 39284 18450
rect 39228 18386 39284 18398
rect 39340 18452 39396 18462
rect 39340 18358 39396 18396
rect 39452 18228 39508 18956
rect 39900 18564 39956 19070
rect 40012 19010 40068 19022
rect 40012 18958 40014 19010
rect 40066 18958 40068 19010
rect 40012 18900 40068 18958
rect 40012 18834 40068 18844
rect 39900 18498 39956 18508
rect 39676 18452 39732 18462
rect 39452 18162 39508 18172
rect 39564 18338 39620 18350
rect 39564 18286 39566 18338
rect 39618 18286 39620 18338
rect 39116 18116 39172 18126
rect 39116 17780 39172 18060
rect 39116 17686 39172 17724
rect 39340 17668 39396 17678
rect 39340 17574 39396 17612
rect 39564 17444 39620 18286
rect 39564 17378 39620 17388
rect 39676 17442 39732 18396
rect 39676 17390 39678 17442
rect 39730 17390 39732 17442
rect 39676 17378 39732 17390
rect 39788 18450 39844 18462
rect 39788 18398 39790 18450
rect 39842 18398 39844 18450
rect 39788 17666 39844 18398
rect 39788 17614 39790 17666
rect 39842 17614 39844 17666
rect 39788 17332 39844 17614
rect 40012 18450 40068 18462
rect 40012 18398 40014 18450
rect 40066 18398 40068 18450
rect 40012 17668 40068 18398
rect 40124 18004 40180 20188
rect 40572 20132 40628 28028
rect 41020 28018 41076 28028
rect 41692 28084 41748 67172
rect 42028 39060 42084 39098
rect 42028 38994 42084 39004
rect 41692 28018 41748 28028
rect 41804 38836 41860 38846
rect 42028 38836 42084 38846
rect 41860 38834 42084 38836
rect 41860 38782 42030 38834
rect 42082 38782 42084 38834
rect 41860 38780 42084 38782
rect 41356 27972 41412 27982
rect 41020 27858 41076 27870
rect 41020 27806 41022 27858
rect 41074 27806 41076 27858
rect 40684 27074 40740 27086
rect 40684 27022 40686 27074
rect 40738 27022 40740 27074
rect 40684 26908 40740 27022
rect 41020 27074 41076 27806
rect 41020 27022 41022 27074
rect 41074 27022 41076 27074
rect 41020 26908 41076 27022
rect 40684 26852 41076 26908
rect 41356 26908 41412 27916
rect 41580 27970 41636 27982
rect 41580 27918 41582 27970
rect 41634 27918 41636 27970
rect 41468 27860 41524 27870
rect 41468 27766 41524 27804
rect 41580 27300 41636 27918
rect 41580 27244 41748 27300
rect 41692 26964 41748 27244
rect 40908 26290 40964 26852
rect 40908 26238 40910 26290
rect 40962 26238 40964 26290
rect 40908 25618 40964 26238
rect 40908 25566 40910 25618
rect 40962 25566 40964 25618
rect 40908 25554 40964 25566
rect 41132 26850 41188 26862
rect 41356 26852 41636 26908
rect 41132 26798 41134 26850
rect 41186 26798 41188 26850
rect 41020 25508 41076 25518
rect 40908 24948 40964 24958
rect 41020 24948 41076 25452
rect 40908 24946 41076 24948
rect 40908 24894 40910 24946
rect 40962 24894 41076 24946
rect 40908 24892 41076 24894
rect 40908 24882 40964 24892
rect 41020 23154 41076 23166
rect 41020 23102 41022 23154
rect 41074 23102 41076 23154
rect 41020 21474 41076 23102
rect 41020 21422 41022 21474
rect 41074 21422 41076 21474
rect 41020 21028 41076 21422
rect 40796 20972 41076 21028
rect 40684 20578 40740 20590
rect 40684 20526 40686 20578
rect 40738 20526 40740 20578
rect 40684 20468 40740 20526
rect 40684 20402 40740 20412
rect 40572 20066 40628 20076
rect 40236 20020 40292 20030
rect 40796 20020 40852 20972
rect 41132 20690 41188 26798
rect 41356 26516 41412 26526
rect 41356 25508 41412 26460
rect 41356 25414 41412 25452
rect 41468 26178 41524 26190
rect 41468 26126 41470 26178
rect 41522 26126 41524 26178
rect 41244 24836 41300 24846
rect 41244 24742 41300 24780
rect 41356 21588 41412 21598
rect 41356 20916 41412 21532
rect 41356 20850 41412 20860
rect 41132 20638 41134 20690
rect 41186 20638 41188 20690
rect 41132 20626 41188 20638
rect 41244 20802 41300 20814
rect 41244 20750 41246 20802
rect 41298 20750 41300 20802
rect 40908 20132 40964 20142
rect 40908 20038 40964 20076
rect 40236 19234 40292 19964
rect 40684 19964 40852 20020
rect 41132 20020 41188 20030
rect 40236 19182 40238 19234
rect 40290 19182 40292 19234
rect 40236 19170 40292 19182
rect 40572 19684 40628 19694
rect 40460 19124 40516 19162
rect 40460 19058 40516 19068
rect 40572 19122 40628 19628
rect 40572 19070 40574 19122
rect 40626 19070 40628 19122
rect 40572 19058 40628 19070
rect 40124 17938 40180 17948
rect 40460 18900 40516 18910
rect 40460 17780 40516 18844
rect 40572 18340 40628 18350
rect 40684 18340 40740 19964
rect 41132 19926 41188 19964
rect 41132 19684 41188 19694
rect 40796 19460 40852 19470
rect 40796 19234 40852 19404
rect 40796 19182 40798 19234
rect 40850 19182 40852 19234
rect 40796 19170 40852 19182
rect 41020 19236 41076 19246
rect 41020 19142 41076 19180
rect 40628 18284 40740 18340
rect 40572 18274 40628 18284
rect 40460 17724 40628 17780
rect 40012 17574 40068 17612
rect 40348 17668 40404 17678
rect 40348 17554 40404 17612
rect 40348 17502 40350 17554
rect 40402 17502 40404 17554
rect 40348 17490 40404 17502
rect 39788 17276 40068 17332
rect 39004 17054 39006 17106
rect 39058 17054 39060 17106
rect 39004 17042 39060 17054
rect 39228 17052 39620 17108
rect 38892 16996 38948 17006
rect 38892 16884 38948 16940
rect 38892 16882 39172 16884
rect 38892 16830 38894 16882
rect 38946 16830 39172 16882
rect 38892 16828 39172 16830
rect 38892 16818 38948 16828
rect 38892 16100 38948 16110
rect 38780 16098 38948 16100
rect 38780 16046 38894 16098
rect 38946 16046 38948 16098
rect 38780 16044 38948 16046
rect 38892 16034 38948 16044
rect 38332 15986 38388 15998
rect 38332 15934 38334 15986
rect 38386 15934 38388 15986
rect 38332 15540 38388 15934
rect 39116 15988 39172 16828
rect 39228 16882 39284 17052
rect 39452 16884 39508 16894
rect 39228 16830 39230 16882
rect 39282 16830 39284 16882
rect 39228 16818 39284 16830
rect 39340 16882 39508 16884
rect 39340 16830 39454 16882
rect 39506 16830 39508 16882
rect 39340 16828 39508 16830
rect 39228 15988 39284 15998
rect 39116 15986 39284 15988
rect 39116 15934 39230 15986
rect 39282 15934 39284 15986
rect 39116 15932 39284 15934
rect 39228 15922 39284 15932
rect 39340 15764 39396 16828
rect 39452 16818 39508 16828
rect 39564 15988 39620 17052
rect 39788 17106 39844 17118
rect 39788 17054 39790 17106
rect 39842 17054 39844 17106
rect 39788 16772 39844 17054
rect 39900 16996 39956 17006
rect 40012 16996 40068 17276
rect 39956 16940 40068 16996
rect 39900 16902 39956 16940
rect 40124 16884 40180 16894
rect 40124 16790 40180 16828
rect 39788 16706 39844 16716
rect 39676 16212 39732 16222
rect 39676 16118 39732 16156
rect 40460 16212 40516 16222
rect 40572 16212 40628 17724
rect 40684 17668 40740 17678
rect 40684 17574 40740 17612
rect 41020 17668 41076 17678
rect 40460 16210 40628 16212
rect 40460 16158 40462 16210
rect 40514 16158 40628 16210
rect 40460 16156 40628 16158
rect 40908 16212 40964 16222
rect 41020 16212 41076 17612
rect 41132 17106 41188 19628
rect 41244 19460 41300 20750
rect 41244 19394 41300 19404
rect 41356 19124 41412 19134
rect 41356 18674 41412 19068
rect 41356 18622 41358 18674
rect 41410 18622 41412 18674
rect 41356 18610 41412 18622
rect 41244 18452 41300 18462
rect 41244 18358 41300 18396
rect 41132 17054 41134 17106
rect 41186 17054 41188 17106
rect 41132 17042 41188 17054
rect 41244 18228 41300 18238
rect 41244 16548 41300 18172
rect 41356 18226 41412 18238
rect 41356 18174 41358 18226
rect 41410 18174 41412 18226
rect 41356 17666 41412 18174
rect 41356 17614 41358 17666
rect 41410 17614 41412 17666
rect 41356 17602 41412 17614
rect 41468 17554 41524 26126
rect 41580 20692 41636 26852
rect 41692 26292 41748 26908
rect 41692 26226 41748 26236
rect 41692 24612 41748 24622
rect 41692 24518 41748 24556
rect 41804 24050 41860 38780
rect 42028 38770 42084 38780
rect 41916 28084 41972 28094
rect 41916 26290 41972 28028
rect 42140 27188 42196 67172
rect 42812 55468 42868 76302
rect 43372 75794 43428 76636
rect 43596 76626 43652 76636
rect 43932 77028 43988 77038
rect 43372 75742 43374 75794
rect 43426 75742 43428 75794
rect 43372 75730 43428 75742
rect 43932 75794 43988 76972
rect 44156 76692 44212 79200
rect 44156 76626 44212 76636
rect 44492 77028 44548 77038
rect 44492 76690 44548 76972
rect 44828 76804 44884 79200
rect 45500 77026 45556 79200
rect 45500 76974 45502 77026
rect 45554 76974 45556 77026
rect 45500 76962 45556 76974
rect 44492 76638 44494 76690
rect 44546 76638 44548 76690
rect 44492 76626 44548 76638
rect 44604 76748 45220 76804
rect 44604 76468 44660 76748
rect 44380 76412 44660 76468
rect 43932 75742 43934 75794
rect 43986 75742 43988 75794
rect 43932 75730 43988 75742
rect 44156 76354 44212 76366
rect 44156 76302 44158 76354
rect 44210 76302 44212 76354
rect 42140 27074 42196 27132
rect 42140 27022 42142 27074
rect 42194 27022 42196 27074
rect 42140 27010 42196 27022
rect 42364 55412 42868 55468
rect 43820 75684 43876 75694
rect 41916 26238 41918 26290
rect 41970 26238 41972 26290
rect 41916 26226 41972 26238
rect 42028 26962 42084 26974
rect 42028 26910 42030 26962
rect 42082 26910 42084 26962
rect 42028 26402 42084 26910
rect 42364 26908 42420 55412
rect 43596 41860 43652 41870
rect 43148 40628 43204 40638
rect 42588 40404 42644 40414
rect 42588 38946 42644 40348
rect 42588 38894 42590 38946
rect 42642 38894 42644 38946
rect 42588 38882 42644 38894
rect 43036 38948 43092 38958
rect 43036 38854 43092 38892
rect 42924 38836 42980 38846
rect 42924 38742 42980 38780
rect 42588 28532 42644 28542
rect 42476 28084 42532 28094
rect 42476 27990 42532 28028
rect 42028 26350 42030 26402
rect 42082 26350 42084 26402
rect 42028 26292 42084 26350
rect 42028 26226 42084 26236
rect 42252 26852 42420 26908
rect 42476 27636 42532 27646
rect 41916 25732 41972 25742
rect 41916 25618 41972 25676
rect 41916 25566 41918 25618
rect 41970 25566 41972 25618
rect 41916 25554 41972 25566
rect 42028 25620 42084 25630
rect 42028 24946 42084 25564
rect 42252 25284 42308 26852
rect 42364 26516 42420 26526
rect 42364 26422 42420 26460
rect 42252 25218 42308 25228
rect 42476 24948 42532 27580
rect 42588 27186 42644 28476
rect 42588 27134 42590 27186
rect 42642 27134 42644 27186
rect 42588 27122 42644 27134
rect 43036 27188 43092 27198
rect 43036 27094 43092 27132
rect 42924 26292 42980 26302
rect 42924 26198 42980 26236
rect 43036 25732 43092 25742
rect 42812 25506 42868 25518
rect 42812 25454 42814 25506
rect 42866 25454 42868 25506
rect 42700 25394 42756 25406
rect 42700 25342 42702 25394
rect 42754 25342 42756 25394
rect 42700 25060 42756 25342
rect 42812 25284 42868 25454
rect 42812 25218 42868 25228
rect 43036 25060 43092 25676
rect 42700 25004 43092 25060
rect 42028 24894 42030 24946
rect 42082 24894 42084 24946
rect 42028 24882 42084 24894
rect 42140 24892 42532 24948
rect 41804 23998 41806 24050
rect 41858 23998 41860 24050
rect 41692 23268 41748 23278
rect 41804 23268 41860 23998
rect 41692 23266 41860 23268
rect 41692 23214 41694 23266
rect 41746 23214 41860 23266
rect 41692 23212 41860 23214
rect 41692 23202 41748 23212
rect 42140 22482 42196 24892
rect 43036 24834 43092 25004
rect 43036 24782 43038 24834
rect 43090 24782 43092 24834
rect 43036 24770 43092 24782
rect 42364 24724 42420 24734
rect 42140 22430 42142 22482
rect 42194 22430 42196 22482
rect 42140 22418 42196 22430
rect 42252 24722 42644 24724
rect 42252 24670 42366 24722
rect 42418 24670 42644 24722
rect 42252 24668 42644 24670
rect 42140 21364 42196 21374
rect 42140 21270 42196 21308
rect 42252 20692 42308 24668
rect 42364 24658 42420 24668
rect 42588 24162 42644 24668
rect 42588 24110 42590 24162
rect 42642 24110 42644 24162
rect 42588 24098 42644 24110
rect 42700 24388 42756 24398
rect 42364 23716 42420 23726
rect 42700 23716 42756 24332
rect 42812 23716 42868 23726
rect 42364 23714 42644 23716
rect 42364 23662 42366 23714
rect 42418 23662 42644 23714
rect 42364 23660 42644 23662
rect 42364 23650 42420 23660
rect 42588 23548 42644 23660
rect 42476 23492 42644 23548
rect 42700 23714 42868 23716
rect 42700 23662 42814 23714
rect 42866 23662 42868 23714
rect 42700 23660 42868 23662
rect 42476 22372 42532 23492
rect 42476 22278 42532 22316
rect 42364 22258 42420 22270
rect 42364 22206 42366 22258
rect 42418 22206 42420 22258
rect 42364 21140 42420 22206
rect 42476 21588 42532 21598
rect 42476 21494 42532 21532
rect 42364 21074 42420 21084
rect 41580 20636 41972 20692
rect 42252 20636 42420 20692
rect 41580 19460 41636 19470
rect 41580 18900 41636 19404
rect 41580 18834 41636 18844
rect 41692 19234 41748 19246
rect 41692 19182 41694 19234
rect 41746 19182 41748 19234
rect 41468 17502 41470 17554
rect 41522 17502 41524 17554
rect 41468 17490 41524 17502
rect 41356 17444 41412 17454
rect 41356 16994 41412 17388
rect 41692 17106 41748 19182
rect 41804 19012 41860 19022
rect 41804 18562 41860 18956
rect 41804 18510 41806 18562
rect 41858 18510 41860 18562
rect 41804 18498 41860 18510
rect 41916 18674 41972 20636
rect 42140 20580 42196 20590
rect 42140 20578 42308 20580
rect 42140 20526 42142 20578
rect 42194 20526 42308 20578
rect 42140 20524 42308 20526
rect 42140 20514 42196 20524
rect 41916 18622 41918 18674
rect 41970 18622 41972 18674
rect 41916 18452 41972 18622
rect 41916 18386 41972 18396
rect 42140 19124 42196 19134
rect 41916 18228 41972 18238
rect 41916 18134 41972 18172
rect 41692 17054 41694 17106
rect 41746 17054 41748 17106
rect 41692 17042 41748 17054
rect 42140 17106 42196 19068
rect 42140 17054 42142 17106
rect 42194 17054 42196 17106
rect 42140 17042 42196 17054
rect 41356 16942 41358 16994
rect 41410 16942 41412 16994
rect 41356 16930 41412 16942
rect 41468 16994 41524 17006
rect 41468 16942 41470 16994
rect 41522 16942 41524 16994
rect 41468 16884 41524 16942
rect 41468 16818 41524 16828
rect 41916 16884 41972 16894
rect 40908 16210 41076 16212
rect 40908 16158 40910 16210
rect 40962 16158 41076 16210
rect 40908 16156 41076 16158
rect 41132 16492 41300 16548
rect 40460 16146 40516 16156
rect 40908 16146 40964 16156
rect 39564 15932 39844 15988
rect 39004 15708 39396 15764
rect 38556 15540 38612 15550
rect 38332 15538 38612 15540
rect 38332 15486 38558 15538
rect 38610 15486 38612 15538
rect 38332 15484 38612 15486
rect 38556 14868 38612 15484
rect 38892 15540 38948 15550
rect 38892 15426 38948 15484
rect 39004 15538 39060 15708
rect 39004 15486 39006 15538
rect 39058 15486 39060 15538
rect 39004 15474 39060 15486
rect 39452 15540 39508 15550
rect 39452 15446 39508 15484
rect 38892 15374 38894 15426
rect 38946 15374 38948 15426
rect 38892 15362 38948 15374
rect 39676 15314 39732 15326
rect 39676 15262 39678 15314
rect 39730 15262 39732 15314
rect 38556 14802 38612 14812
rect 39228 15204 39284 15214
rect 38220 14476 38612 14532
rect 37436 14466 37492 14476
rect 37212 14420 37268 14430
rect 37212 12402 37268 14364
rect 38444 14308 38500 14318
rect 37660 13972 37716 13982
rect 37436 13188 37492 13198
rect 37492 13132 37604 13188
rect 37436 13122 37492 13132
rect 37212 12350 37214 12402
rect 37266 12350 37268 12402
rect 37212 12338 37268 12350
rect 37324 12850 37380 12862
rect 37324 12798 37326 12850
rect 37378 12798 37380 12850
rect 37324 12180 37380 12798
rect 37100 12124 37268 12180
rect 36540 12114 36596 12124
rect 36876 12086 36932 12124
rect 35980 11506 36372 11508
rect 35980 11454 35982 11506
rect 36034 11454 36372 11506
rect 35980 11452 36372 11454
rect 36988 12068 37044 12078
rect 35980 11396 36036 11452
rect 35980 11330 36036 11340
rect 36988 11394 37044 12012
rect 37212 11732 37268 12124
rect 37212 11666 37268 11676
rect 36988 11342 36990 11394
rect 37042 11342 37044 11394
rect 36428 11172 36484 11182
rect 36428 11078 36484 11116
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 34972 10108 35140 10164
rect 35196 10154 35460 10164
rect 35084 10052 35140 10108
rect 35196 10052 35252 10062
rect 35084 10050 35252 10052
rect 35084 9998 35198 10050
rect 35250 9998 35252 10050
rect 35084 9996 35252 9998
rect 35196 9986 35252 9996
rect 34860 9940 34916 9950
rect 34916 9884 35140 9940
rect 34860 9846 34916 9884
rect 35084 9826 35140 9884
rect 35084 9774 35086 9826
rect 35138 9774 35140 9826
rect 35084 9762 35140 9774
rect 36876 9828 36932 9838
rect 34524 9090 34580 9100
rect 33964 9042 34468 9044
rect 33964 8990 33966 9042
rect 34018 8990 34468 9042
rect 33964 8988 34468 8990
rect 33964 8978 34020 8988
rect 33516 8932 33572 8942
rect 33516 8838 33572 8876
rect 33628 8820 33684 8830
rect 34300 8820 34356 8830
rect 33628 8818 34244 8820
rect 33628 8766 33630 8818
rect 33682 8766 34244 8818
rect 33628 8764 34244 8766
rect 33628 8754 33684 8764
rect 34188 8370 34244 8764
rect 34188 8318 34190 8370
rect 34242 8318 34244 8370
rect 34188 8306 34244 8318
rect 34300 8258 34356 8764
rect 34300 8206 34302 8258
rect 34354 8206 34356 8258
rect 34300 8194 34356 8206
rect 33292 7970 33348 7980
rect 33516 8034 33572 8046
rect 33516 7982 33518 8034
rect 33570 7982 33572 8034
rect 32956 7532 33460 7588
rect 33404 7474 33460 7532
rect 33404 7422 33406 7474
rect 33458 7422 33460 7474
rect 32844 6638 32846 6690
rect 32898 6638 32900 6690
rect 32396 6466 32452 6478
rect 32844 6468 32900 6638
rect 32396 6414 32398 6466
rect 32450 6414 32452 6466
rect 32172 5908 32228 5918
rect 31724 5170 31780 5180
rect 31836 5348 31892 5358
rect 31836 5234 31892 5292
rect 31836 5182 31838 5234
rect 31890 5182 31892 5234
rect 31836 5170 31892 5182
rect 31388 3554 31556 3556
rect 31388 3502 31390 3554
rect 31442 3502 31556 3554
rect 31388 3500 31556 3502
rect 31388 3490 31444 3500
rect 30716 3332 30884 3388
rect 30604 2212 30660 3164
rect 30604 2146 30660 2156
rect 30828 980 30884 3332
rect 30940 3332 30996 3342
rect 30940 3238 30996 3276
rect 31500 1764 31556 3500
rect 31836 3780 31892 3790
rect 31500 1698 31556 1708
rect 31612 3330 31668 3342
rect 31612 3278 31614 3330
rect 31666 3278 31668 3330
rect 31612 1540 31668 3278
rect 31612 1474 31668 1484
rect 30828 924 31220 980
rect 31164 800 31220 924
rect 31836 800 31892 3724
rect 32172 3556 32228 5852
rect 32284 5124 32340 5134
rect 32284 5030 32340 5068
rect 32396 4788 32452 6414
rect 32508 6412 32900 6468
rect 33068 7364 33124 7374
rect 33292 7364 33348 7374
rect 33068 7140 33124 7308
rect 32508 5794 32564 6412
rect 32508 5742 32510 5794
rect 32562 5742 32564 5794
rect 32508 5730 32564 5742
rect 32620 5684 32676 5694
rect 32620 5122 32676 5628
rect 33068 5460 33124 7084
rect 33180 7362 33348 7364
rect 33180 7310 33294 7362
rect 33346 7310 33348 7362
rect 33180 7308 33348 7310
rect 33180 5572 33236 7308
rect 33292 7298 33348 7308
rect 33292 6804 33348 6814
rect 33404 6804 33460 7422
rect 33348 6748 33460 6804
rect 33292 6690 33348 6748
rect 33292 6638 33294 6690
rect 33346 6638 33348 6690
rect 33292 6626 33348 6638
rect 33516 5908 33572 7982
rect 34076 8036 34132 8046
rect 34076 8034 34244 8036
rect 34076 7982 34078 8034
rect 34130 7982 34244 8034
rect 34076 7980 34244 7982
rect 34076 7970 34132 7980
rect 33964 7700 34020 7710
rect 33964 7606 34020 7644
rect 33852 7588 33908 7598
rect 34188 7588 34244 7980
rect 33852 7494 33908 7532
rect 34076 7532 34244 7588
rect 33740 7476 33796 7486
rect 33628 7420 33740 7476
rect 33628 6690 33684 7420
rect 33740 7410 33796 7420
rect 34076 7474 34132 7532
rect 34076 7422 34078 7474
rect 34130 7422 34132 7474
rect 34076 7028 34132 7422
rect 34412 7476 34468 8988
rect 34748 8932 34804 8942
rect 34748 8838 34804 8876
rect 36876 8930 36932 9772
rect 36988 9826 37044 11342
rect 37324 11284 37380 12124
rect 37436 12738 37492 12750
rect 37436 12686 37438 12738
rect 37490 12686 37492 12738
rect 37436 11956 37492 12686
rect 37548 12178 37604 13132
rect 37660 12962 37716 13916
rect 37884 13748 37940 13758
rect 38332 13748 38388 13758
rect 37884 13300 37940 13692
rect 37996 13746 38388 13748
rect 37996 13694 38334 13746
rect 38386 13694 38388 13746
rect 37996 13692 38388 13694
rect 37996 13634 38052 13692
rect 38332 13682 38388 13692
rect 37996 13582 37998 13634
rect 38050 13582 38052 13634
rect 37996 13570 38052 13582
rect 38444 13524 38500 14252
rect 38444 13430 38500 13468
rect 37884 13244 38500 13300
rect 37660 12910 37662 12962
rect 37714 12910 37716 12962
rect 37660 12898 37716 12910
rect 38444 12962 38500 13244
rect 38444 12910 38446 12962
rect 38498 12910 38500 12962
rect 38444 12898 38500 12910
rect 37548 12126 37550 12178
rect 37602 12126 37604 12178
rect 37548 12114 37604 12126
rect 37996 12516 38052 12526
rect 37436 11890 37492 11900
rect 37996 11618 38052 12460
rect 37996 11566 37998 11618
rect 38050 11566 38052 11618
rect 37996 11554 38052 11566
rect 38220 12066 38276 12078
rect 38220 12014 38222 12066
rect 38274 12014 38276 12066
rect 38220 11396 38276 12014
rect 38220 11330 38276 11340
rect 37884 11284 37940 11294
rect 37324 11282 37940 11284
rect 37324 11230 37326 11282
rect 37378 11230 37886 11282
rect 37938 11230 37940 11282
rect 37324 11228 37940 11230
rect 37324 11218 37380 11228
rect 37884 11218 37940 11228
rect 37996 11170 38052 11182
rect 37996 11118 37998 11170
rect 38050 11118 38052 11170
rect 37996 10052 38052 11118
rect 38556 11060 38612 14476
rect 39228 14530 39284 15148
rect 39228 14478 39230 14530
rect 39282 14478 39284 14530
rect 39004 13748 39060 13758
rect 39004 13654 39060 13692
rect 39228 13188 39284 14478
rect 39340 14084 39396 14094
rect 39340 13970 39396 14028
rect 39340 13918 39342 13970
rect 39394 13918 39396 13970
rect 39340 13906 39396 13918
rect 39676 13972 39732 15262
rect 39676 13906 39732 13916
rect 39228 12962 39284 13132
rect 39228 12910 39230 12962
rect 39282 12910 39284 12962
rect 38780 12740 38836 12750
rect 38780 12738 39172 12740
rect 38780 12686 38782 12738
rect 38834 12686 39172 12738
rect 38780 12684 39172 12686
rect 38780 12674 38836 12684
rect 39116 11620 39172 12684
rect 39228 12068 39284 12910
rect 39564 13746 39620 13758
rect 39564 13694 39566 13746
rect 39618 13694 39620 13746
rect 39564 12516 39620 13694
rect 39788 13524 39844 15932
rect 40124 15876 40180 15886
rect 40124 15538 40180 15820
rect 40124 15486 40126 15538
rect 40178 15486 40180 15538
rect 40124 15474 40180 15486
rect 40348 15314 40404 15326
rect 40348 15262 40350 15314
rect 40402 15262 40404 15314
rect 40236 15202 40292 15214
rect 40236 15150 40238 15202
rect 40290 15150 40292 15202
rect 40236 15148 40292 15150
rect 40012 15092 40292 15148
rect 40012 14642 40068 15092
rect 40012 14590 40014 14642
rect 40066 14590 40068 14642
rect 40012 14578 40068 14590
rect 40236 13972 40292 13982
rect 40348 13972 40404 15262
rect 40292 13916 40404 13972
rect 40236 13878 40292 13916
rect 40012 13860 40068 13870
rect 40012 13766 40068 13804
rect 39788 13458 39844 13468
rect 40124 13634 40180 13646
rect 40124 13582 40126 13634
rect 40178 13582 40180 13634
rect 40124 13188 40180 13582
rect 39900 13132 40180 13188
rect 40796 13524 40852 13534
rect 39900 13074 39956 13132
rect 39900 13022 39902 13074
rect 39954 13022 39956 13074
rect 39900 13010 39956 13022
rect 39564 12450 39620 12460
rect 40684 12180 40740 12190
rect 39228 12002 39284 12012
rect 40348 12124 40684 12180
rect 40348 12066 40404 12124
rect 40684 12114 40740 12124
rect 40348 12014 40350 12066
rect 40402 12014 40404 12066
rect 40348 12002 40404 12014
rect 40796 11956 40852 13468
rect 40908 12516 40964 12526
rect 40908 12180 40964 12460
rect 40908 12124 41076 12180
rect 41020 12066 41076 12124
rect 41020 12014 41022 12066
rect 41074 12014 41076 12066
rect 41020 12002 41076 12014
rect 40908 11956 40964 11966
rect 40796 11954 40964 11956
rect 40796 11902 40910 11954
rect 40962 11902 40964 11954
rect 40796 11900 40964 11902
rect 40908 11890 40964 11900
rect 41132 11844 41188 16492
rect 41468 16212 41524 16222
rect 41468 16118 41524 16156
rect 41916 16210 41972 16828
rect 41916 16158 41918 16210
rect 41970 16158 41972 16210
rect 41916 16146 41972 16158
rect 41020 11788 41188 11844
rect 41244 16100 41300 16110
rect 42252 16100 42308 20524
rect 42364 18674 42420 20636
rect 42700 20020 42756 23660
rect 42812 23650 42868 23660
rect 43148 23716 43204 40572
rect 43596 40404 43652 41804
rect 43260 39396 43316 39406
rect 43260 38946 43316 39340
rect 43596 39058 43652 40348
rect 43596 39006 43598 39058
rect 43650 39006 43652 39058
rect 43596 38994 43652 39006
rect 43260 38894 43262 38946
rect 43314 38894 43316 38946
rect 43260 38882 43316 38894
rect 43820 27412 43876 75628
rect 44156 67228 44212 76302
rect 44380 75794 44436 76412
rect 45052 76356 45108 76366
rect 44380 75742 44382 75794
rect 44434 75742 44436 75794
rect 44380 75730 44436 75742
rect 44940 76354 45108 76356
rect 44940 76302 45054 76354
rect 45106 76302 45108 76354
rect 44940 76300 45108 76302
rect 44940 67228 44996 76300
rect 45052 76290 45108 76300
rect 45164 75682 45220 76748
rect 45388 76692 45444 76702
rect 45388 76598 45444 76636
rect 45836 76692 45892 76702
rect 45836 75796 45892 76636
rect 46172 76692 46228 79200
rect 46172 76626 46228 76636
rect 46284 77026 46340 77038
rect 46284 76974 46286 77026
rect 46338 76974 46340 77026
rect 46284 76692 46340 76974
rect 46284 76690 46564 76692
rect 46284 76638 46286 76690
rect 46338 76638 46564 76690
rect 46284 76636 46564 76638
rect 46284 76626 46340 76636
rect 45948 76356 46004 76366
rect 45948 76354 46228 76356
rect 45948 76302 45950 76354
rect 46002 76302 46228 76354
rect 45948 76300 46228 76302
rect 45948 76290 46004 76300
rect 46060 75796 46116 75806
rect 45836 75794 46116 75796
rect 45836 75742 46062 75794
rect 46114 75742 46116 75794
rect 45836 75740 46116 75742
rect 46060 75730 46116 75740
rect 45164 75630 45166 75682
rect 45218 75630 45220 75682
rect 45164 75618 45220 75630
rect 45612 75682 45668 75694
rect 45612 75630 45614 75682
rect 45666 75630 45668 75682
rect 45612 67228 45668 75630
rect 46172 67228 46228 76300
rect 46508 75794 46564 76636
rect 46844 76580 46900 79200
rect 47516 77026 47572 79200
rect 47516 76974 47518 77026
rect 47570 76974 47572 77026
rect 47516 76962 47572 76974
rect 47404 76692 47460 76702
rect 47404 76598 47460 76636
rect 47852 76692 47908 76702
rect 48188 76692 48244 79200
rect 47908 76636 48132 76692
rect 47852 76626 47908 76636
rect 46844 76524 47124 76580
rect 46844 76354 46900 76366
rect 46844 76302 46846 76354
rect 46898 76302 46900 76354
rect 46844 75908 46900 76302
rect 46844 75842 46900 75852
rect 46508 75742 46510 75794
rect 46562 75742 46564 75794
rect 46508 75730 46564 75742
rect 47068 75684 47124 76524
rect 47852 76356 47908 76366
rect 47852 76262 47908 76300
rect 48076 75794 48132 76636
rect 48188 76626 48244 76636
rect 48300 77026 48356 77038
rect 48300 76974 48302 77026
rect 48354 76974 48356 77026
rect 48300 76692 48356 76974
rect 48860 77026 48916 79200
rect 48860 76974 48862 77026
rect 48914 76974 48916 77026
rect 48860 76962 48916 76974
rect 49196 76692 49252 76702
rect 48300 76690 48580 76692
rect 48300 76638 48302 76690
rect 48354 76638 48580 76690
rect 48300 76636 48580 76638
rect 48300 76626 48356 76636
rect 48076 75742 48078 75794
rect 48130 75742 48132 75794
rect 48076 75730 48132 75742
rect 48412 75908 48468 75918
rect 46844 75682 47124 75684
rect 46844 75630 47070 75682
rect 47122 75630 47124 75682
rect 46844 75628 47124 75630
rect 46844 75122 46900 75628
rect 47068 75618 47124 75628
rect 47628 75682 47684 75694
rect 47628 75630 47630 75682
rect 47682 75630 47684 75682
rect 46844 75070 46846 75122
rect 46898 75070 46900 75122
rect 46844 75058 46900 75070
rect 44156 67172 44324 67228
rect 44940 67172 45108 67228
rect 45612 67172 46004 67228
rect 46172 67172 46788 67228
rect 44268 43708 44324 67172
rect 43820 27346 43876 27356
rect 43932 43652 44324 43708
rect 43484 26402 43540 26414
rect 43484 26350 43486 26402
rect 43538 26350 43540 26402
rect 43484 25732 43540 26350
rect 43484 25666 43540 25676
rect 43708 25620 43764 25630
rect 43372 25508 43428 25518
rect 43372 25414 43428 25452
rect 43708 25506 43764 25564
rect 43708 25454 43710 25506
rect 43762 25454 43764 25506
rect 43708 25442 43764 25454
rect 43260 25284 43316 25294
rect 43260 25282 43540 25284
rect 43260 25230 43262 25282
rect 43314 25230 43540 25282
rect 43260 25228 43540 25230
rect 43260 25218 43316 25228
rect 43372 24162 43428 24174
rect 43372 24110 43374 24162
rect 43426 24110 43428 24162
rect 43260 23716 43316 23726
rect 43148 23714 43316 23716
rect 43148 23662 43262 23714
rect 43314 23662 43316 23714
rect 43148 23660 43316 23662
rect 43036 22146 43092 22158
rect 43036 22094 43038 22146
rect 43090 22094 43092 22146
rect 43036 21588 43092 22094
rect 43036 21522 43092 21532
rect 42812 21476 42868 21486
rect 42812 20242 42868 21420
rect 42812 20190 42814 20242
rect 42866 20190 42868 20242
rect 42812 20178 42868 20190
rect 42924 21364 42980 21374
rect 42924 20690 42980 21308
rect 43148 21140 43204 23660
rect 43260 23650 43316 23660
rect 43372 22370 43428 24110
rect 43372 22318 43374 22370
rect 43426 22318 43428 22370
rect 43372 22306 43428 22318
rect 43260 21700 43316 21710
rect 43260 21606 43316 21644
rect 43260 21140 43316 21150
rect 43148 21084 43260 21140
rect 43260 21074 43316 21084
rect 42924 20638 42926 20690
rect 42978 20638 42980 20690
rect 42924 20130 42980 20638
rect 43148 20802 43204 20814
rect 43148 20750 43150 20802
rect 43202 20750 43204 20802
rect 43148 20468 43204 20750
rect 43148 20402 43204 20412
rect 42924 20078 42926 20130
rect 42978 20078 42980 20130
rect 42700 19964 42868 20020
rect 42364 18622 42366 18674
rect 42418 18622 42420 18674
rect 42364 16548 42420 18622
rect 42588 18452 42644 18462
rect 42588 17106 42644 18396
rect 42588 17054 42590 17106
rect 42642 17054 42644 17106
rect 42588 17042 42644 17054
rect 42700 18450 42756 18462
rect 42700 18398 42702 18450
rect 42754 18398 42756 18450
rect 42364 16482 42420 16492
rect 42700 16996 42756 18398
rect 42812 16996 42868 19964
rect 42924 19122 42980 20078
rect 43484 20132 43540 25228
rect 43596 24724 43652 24734
rect 43932 24724 43988 43652
rect 44044 38836 44100 38846
rect 44044 38742 44100 38780
rect 44828 36372 44884 36382
rect 44828 36278 44884 36316
rect 44268 36260 44324 36270
rect 44268 35924 44324 36204
rect 44940 36260 44996 36270
rect 44940 36166 44996 36204
rect 44268 35922 44660 35924
rect 44268 35870 44270 35922
rect 44322 35870 44660 35922
rect 44268 35868 44660 35870
rect 44268 35858 44324 35868
rect 44604 35810 44660 35868
rect 44604 35758 44606 35810
rect 44658 35758 44660 35810
rect 44604 35746 44660 35758
rect 44716 35700 44772 35710
rect 44716 35606 44772 35644
rect 45052 35140 45108 67172
rect 45948 38668 46004 67172
rect 45724 38612 46004 38668
rect 46508 38948 46564 38958
rect 45388 36372 45444 36382
rect 45388 36278 45444 36316
rect 45388 35700 45444 35710
rect 45388 35606 45444 35644
rect 45612 35588 45668 35598
rect 45612 35494 45668 35532
rect 44716 35084 45108 35140
rect 44380 34692 44436 34702
rect 44380 34598 44436 34636
rect 44156 34244 44212 34254
rect 44380 34244 44436 34254
rect 44212 34242 44436 34244
rect 44212 34190 44382 34242
rect 44434 34190 44436 34242
rect 44212 34188 44436 34190
rect 44156 34150 44212 34188
rect 44380 34178 44436 34188
rect 44492 33906 44548 33918
rect 44492 33854 44494 33906
rect 44546 33854 44548 33906
rect 44492 33348 44548 33854
rect 44492 33282 44548 33292
rect 44380 31668 44436 31678
rect 44380 31574 44436 31612
rect 44156 31108 44212 31118
rect 44380 31108 44436 31118
rect 44212 31106 44436 31108
rect 44212 31054 44382 31106
rect 44434 31054 44436 31106
rect 44212 31052 44436 31054
rect 44156 31014 44212 31052
rect 44380 31042 44436 31052
rect 44492 30770 44548 30782
rect 44492 30718 44494 30770
rect 44546 30718 44548 30770
rect 44492 30212 44548 30718
rect 44716 30324 44772 35084
rect 44940 34916 44996 34926
rect 45388 34916 45444 34926
rect 44940 34914 45444 34916
rect 44940 34862 44942 34914
rect 44994 34862 45390 34914
rect 45442 34862 45444 34914
rect 44940 34860 45444 34862
rect 44940 34850 44996 34860
rect 45388 34850 45444 34860
rect 45612 34916 45668 34926
rect 45612 34822 45668 34860
rect 44828 34802 44884 34814
rect 44828 34750 44830 34802
rect 44882 34750 44884 34802
rect 44828 34692 44884 34750
rect 44828 34626 44884 34636
rect 45724 34356 45780 38612
rect 45612 34300 45780 34356
rect 45836 35812 45892 35822
rect 45836 34914 45892 35756
rect 45836 34862 45838 34914
rect 45890 34862 45892 34914
rect 45388 33348 45444 33358
rect 45388 33254 45444 33292
rect 45500 32788 45556 32798
rect 45388 32732 45500 32788
rect 45612 32788 45668 34300
rect 45724 34132 45780 34142
rect 45724 33122 45780 34076
rect 45836 33348 45892 34862
rect 45836 33254 45892 33292
rect 45948 35700 46004 35710
rect 46396 35700 46452 35710
rect 45948 35698 46452 35700
rect 45948 35646 45950 35698
rect 46002 35646 46398 35698
rect 46450 35646 46452 35698
rect 45948 35644 46452 35646
rect 45948 34914 46004 35644
rect 46396 35634 46452 35644
rect 45948 34862 45950 34914
rect 46002 34862 46004 34914
rect 45948 33236 46004 34862
rect 46396 33348 46452 33358
rect 46060 33236 46116 33246
rect 45948 33234 46116 33236
rect 45948 33182 46062 33234
rect 46114 33182 46116 33234
rect 45948 33180 46116 33182
rect 45724 33070 45726 33122
rect 45778 33070 45780 33122
rect 45724 33058 45780 33070
rect 45612 32732 46004 32788
rect 45388 32674 45444 32732
rect 45500 32722 45556 32732
rect 45388 32622 45390 32674
rect 45442 32622 45444 32674
rect 45388 32610 45444 32622
rect 45836 32562 45892 32574
rect 45836 32510 45838 32562
rect 45890 32510 45892 32562
rect 45052 32450 45108 32462
rect 45052 32398 45054 32450
rect 45106 32398 45108 32450
rect 45052 31892 45108 32398
rect 45276 31892 45332 31902
rect 45052 31836 45276 31892
rect 45276 31798 45332 31836
rect 44940 31780 44996 31790
rect 44940 31686 44996 31724
rect 45724 31780 45780 31790
rect 45724 31686 45780 31724
rect 44828 31668 44884 31678
rect 44828 31574 44884 31612
rect 45388 31668 45444 31678
rect 45388 31666 45668 31668
rect 45388 31614 45390 31666
rect 45442 31614 45668 31666
rect 45388 31612 45668 31614
rect 45388 31602 45444 31612
rect 45612 31556 45668 31612
rect 45612 31500 45780 31556
rect 45500 31108 45556 31118
rect 45500 31014 45556 31052
rect 45276 30996 45332 31006
rect 45276 30902 45332 30940
rect 45612 30996 45668 31006
rect 45500 30772 45556 30782
rect 44716 30268 45108 30324
rect 44492 30146 44548 30156
rect 44940 30100 44996 30110
rect 44940 29650 44996 30044
rect 44940 29598 44942 29650
rect 44994 29598 44996 29650
rect 44940 29586 44996 29598
rect 44604 29540 44660 29550
rect 44828 29540 44884 29550
rect 44660 29538 44884 29540
rect 44660 29486 44830 29538
rect 44882 29486 44884 29538
rect 44660 29484 44884 29486
rect 44604 29446 44660 29484
rect 44828 29474 44884 29484
rect 44716 28532 44772 28542
rect 44716 28084 44772 28476
rect 45052 28532 45108 30268
rect 45052 28466 45108 28476
rect 44716 28082 45108 28084
rect 44716 28030 44718 28082
rect 44770 28030 45108 28082
rect 44716 28028 45108 28030
rect 44716 28018 44772 28028
rect 45052 27970 45108 28028
rect 45052 27918 45054 27970
rect 45106 27918 45108 27970
rect 45052 27906 45108 27918
rect 45164 27634 45220 27646
rect 45164 27582 45166 27634
rect 45218 27582 45220 27634
rect 44828 27300 44884 27310
rect 44044 27188 44100 27198
rect 44044 26290 44100 27132
rect 44828 27186 44884 27244
rect 45164 27298 45220 27582
rect 45164 27246 45166 27298
rect 45218 27246 45220 27298
rect 45164 27234 45220 27246
rect 45388 27300 45444 27310
rect 44828 27134 44830 27186
rect 44882 27134 44884 27186
rect 44828 27122 44884 27134
rect 45388 27186 45444 27244
rect 45388 27134 45390 27186
rect 45442 27134 45444 27186
rect 45388 27122 45444 27134
rect 44940 26964 44996 27002
rect 45500 26908 45556 30716
rect 44940 26898 44996 26908
rect 45388 26852 45556 26908
rect 45612 30772 45668 30940
rect 45724 30994 45780 31500
rect 45724 30942 45726 30994
rect 45778 30942 45780 30994
rect 45724 30930 45780 30942
rect 45836 30772 45892 32510
rect 45948 32004 46004 32732
rect 46060 32786 46116 33180
rect 46396 33234 46452 33292
rect 46396 33182 46398 33234
rect 46450 33182 46452 33234
rect 46396 33170 46452 33182
rect 46060 32734 46062 32786
rect 46114 32734 46116 32786
rect 46060 32722 46116 32734
rect 46508 32788 46564 38892
rect 46620 35812 46676 35822
rect 46620 35718 46676 35756
rect 46732 35308 46788 67172
rect 47628 43708 47684 75630
rect 47628 43652 48020 43708
rect 46956 36260 47012 36270
rect 46956 35810 47012 36204
rect 46956 35758 46958 35810
rect 47010 35758 47012 35810
rect 46956 35746 47012 35758
rect 46844 35588 46900 35598
rect 46844 35494 46900 35532
rect 46508 32562 46564 32732
rect 46508 32510 46510 32562
rect 46562 32510 46564 32562
rect 45948 31948 46116 32004
rect 45948 31780 46004 31790
rect 45948 31686 46004 31724
rect 45948 30884 46004 30894
rect 45948 30790 46004 30828
rect 45612 30716 45892 30772
rect 44492 26514 44548 26526
rect 44492 26462 44494 26514
rect 44546 26462 44548 26514
rect 44380 26292 44436 26302
rect 44044 26238 44046 26290
rect 44098 26238 44100 26290
rect 44044 26226 44100 26238
rect 44268 26290 44436 26292
rect 44268 26238 44382 26290
rect 44434 26238 44436 26290
rect 44268 26236 44436 26238
rect 44268 25618 44324 26236
rect 44380 26226 44436 26236
rect 44268 25566 44270 25618
rect 44322 25566 44324 25618
rect 44268 25508 44324 25566
rect 43596 24722 43988 24724
rect 43596 24670 43598 24722
rect 43650 24670 43988 24722
rect 43596 24668 43988 24670
rect 44044 24946 44100 24958
rect 44044 24894 44046 24946
rect 44098 24894 44100 24946
rect 43596 24052 43652 24668
rect 43596 23986 43652 23996
rect 44044 23940 44100 24894
rect 44156 24724 44212 24734
rect 44268 24724 44324 25452
rect 44156 24722 44324 24724
rect 44156 24670 44158 24722
rect 44210 24670 44324 24722
rect 44156 24668 44324 24670
rect 44156 24658 44212 24668
rect 44044 23884 44436 23940
rect 44268 23714 44324 23726
rect 44268 23662 44270 23714
rect 44322 23662 44324 23714
rect 43708 23380 43764 23390
rect 43708 22820 43764 23324
rect 44268 23380 44324 23662
rect 44268 23314 44324 23324
rect 44268 23156 44324 23166
rect 43820 23154 44324 23156
rect 43820 23102 44270 23154
rect 44322 23102 44324 23154
rect 43820 23100 44324 23102
rect 43820 23042 43876 23100
rect 43820 22990 43822 23042
rect 43874 22990 43876 23042
rect 43820 22978 43876 22990
rect 43820 22820 43876 22830
rect 43708 22764 43820 22820
rect 43708 22260 43764 22270
rect 43708 22166 43764 22204
rect 43820 22258 43876 22764
rect 44268 22484 44324 23100
rect 44380 22596 44436 23884
rect 44492 22708 44548 26462
rect 45052 26292 45108 26302
rect 45052 26198 45108 26236
rect 44940 26178 44996 26190
rect 44940 26126 44942 26178
rect 44994 26126 44996 26178
rect 44940 26068 44996 26126
rect 44940 26002 44996 26012
rect 45276 25618 45332 25630
rect 45276 25566 45278 25618
rect 45330 25566 45332 25618
rect 44940 25508 44996 25546
rect 44940 25442 44996 25452
rect 44604 25284 44660 25294
rect 44604 24946 44660 25228
rect 44604 24894 44606 24946
rect 44658 24894 44660 24946
rect 44604 24882 44660 24894
rect 44828 24836 44884 24846
rect 44716 24780 44828 24836
rect 44604 24612 44660 24622
rect 44604 23156 44660 24556
rect 44716 23268 44772 24780
rect 44828 24770 44884 24780
rect 45164 24836 45220 24846
rect 45164 24742 45220 24780
rect 44940 24052 44996 24062
rect 44940 23958 44996 23996
rect 44828 23940 44884 23950
rect 44828 23548 44884 23884
rect 45164 23940 45220 23950
rect 45052 23716 45108 23726
rect 45052 23548 45108 23660
rect 44828 23492 45108 23548
rect 44716 23212 44884 23268
rect 44604 23100 44772 23156
rect 44716 23042 44772 23100
rect 44716 22990 44718 23042
rect 44770 22990 44772 23042
rect 44716 22978 44772 22990
rect 44828 23044 44884 23212
rect 45052 23266 45108 23492
rect 45164 23378 45220 23884
rect 45164 23326 45166 23378
rect 45218 23326 45220 23378
rect 45164 23314 45220 23326
rect 45052 23214 45054 23266
rect 45106 23214 45108 23266
rect 45052 23202 45108 23214
rect 44828 22988 45220 23044
rect 44492 22652 44884 22708
rect 44380 22540 44660 22596
rect 44268 22428 44436 22484
rect 43820 22206 43822 22258
rect 43874 22206 43876 22258
rect 43820 22194 43876 22206
rect 44044 22146 44100 22158
rect 44044 22094 44046 22146
rect 44098 22094 44100 22146
rect 43484 20066 43540 20076
rect 43932 22036 43988 22046
rect 43036 20018 43092 20030
rect 43036 19966 43038 20018
rect 43090 19966 43092 20018
rect 43036 19348 43092 19966
rect 43036 19282 43092 19292
rect 42924 19070 42926 19122
rect 42978 19070 42980 19122
rect 42924 17666 42980 19070
rect 43372 19234 43428 19246
rect 43372 19182 43374 19234
rect 43426 19182 43428 19234
rect 43036 19012 43092 19022
rect 43036 19010 43316 19012
rect 43036 18958 43038 19010
rect 43090 18958 43316 19010
rect 43036 18956 43316 18958
rect 43036 18946 43092 18956
rect 43036 18338 43092 18350
rect 43036 18286 43038 18338
rect 43090 18286 43092 18338
rect 43036 17780 43092 18286
rect 43148 18340 43204 18350
rect 43148 18246 43204 18284
rect 43036 17714 43092 17724
rect 42924 17614 42926 17666
rect 42978 17614 42980 17666
rect 42924 17602 42980 17614
rect 43148 17668 43204 17678
rect 43148 17574 43204 17612
rect 43036 17444 43092 17454
rect 43036 17442 43204 17444
rect 43036 17390 43038 17442
rect 43090 17390 43204 17442
rect 43036 17388 43204 17390
rect 43036 17378 43092 17388
rect 42924 16996 42980 17006
rect 42812 16994 42980 16996
rect 42812 16942 42926 16994
rect 42978 16942 42980 16994
rect 42812 16940 42980 16942
rect 42588 16436 42644 16446
rect 42252 16044 42420 16100
rect 39116 11564 39844 11620
rect 38780 11396 38836 11406
rect 38556 10994 38612 11004
rect 38668 11394 38836 11396
rect 38668 11342 38782 11394
rect 38834 11342 38836 11394
rect 38668 11340 38836 11342
rect 38668 11172 38724 11340
rect 38780 11330 38836 11340
rect 39676 11396 39732 11406
rect 38668 10836 38724 11116
rect 38332 10780 38724 10836
rect 39564 10948 39620 10958
rect 39564 10834 39620 10892
rect 39564 10782 39566 10834
rect 39618 10782 39620 10834
rect 38332 10610 38388 10780
rect 39564 10770 39620 10782
rect 39676 10834 39732 11340
rect 39676 10782 39678 10834
rect 39730 10782 39732 10834
rect 39676 10770 39732 10782
rect 39788 10834 39844 11564
rect 39788 10782 39790 10834
rect 39842 10782 39844 10834
rect 38780 10722 38836 10734
rect 38780 10670 38782 10722
rect 38834 10670 38836 10722
rect 38332 10558 38334 10610
rect 38386 10558 38388 10610
rect 38332 10546 38388 10558
rect 38668 10610 38724 10622
rect 38668 10558 38670 10610
rect 38722 10558 38724 10610
rect 37996 9986 38052 9996
rect 36988 9774 36990 9826
rect 37042 9774 37044 9826
rect 36988 9762 37044 9774
rect 37548 9940 37604 9950
rect 37324 9716 37380 9726
rect 37324 9622 37380 9660
rect 37548 9044 37604 9884
rect 37660 9828 37716 9838
rect 38220 9828 38276 9838
rect 38668 9828 38724 10558
rect 38780 10052 38836 10670
rect 39004 10722 39060 10734
rect 39004 10670 39006 10722
rect 39058 10670 39060 10722
rect 39004 10612 39060 10670
rect 39116 10612 39172 10622
rect 39004 10610 39172 10612
rect 39004 10558 39118 10610
rect 39170 10558 39172 10610
rect 39004 10556 39172 10558
rect 39116 10546 39172 10556
rect 38780 9986 38836 9996
rect 38780 9828 38836 9838
rect 37660 9826 38836 9828
rect 37660 9774 37662 9826
rect 37714 9774 38222 9826
rect 38274 9774 38782 9826
rect 38834 9774 38836 9826
rect 37660 9772 38836 9774
rect 37660 9716 37716 9772
rect 38220 9762 38276 9772
rect 38780 9762 38836 9772
rect 39788 9828 39844 10782
rect 40348 11396 40404 11406
rect 40348 10948 40404 11340
rect 40348 10834 40404 10892
rect 40348 10782 40350 10834
rect 40402 10782 40404 10834
rect 40348 10770 40404 10782
rect 37660 9650 37716 9660
rect 39004 9716 39060 9726
rect 36876 8878 36878 8930
rect 36930 8878 36932 8930
rect 36876 8820 36932 8878
rect 36876 8754 36932 8764
rect 37436 9042 37604 9044
rect 37436 8990 37550 9042
rect 37602 8990 37604 9042
rect 37436 8988 37604 8990
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 34412 7382 34468 7420
rect 34636 8258 34692 8270
rect 34636 8206 34638 8258
rect 34690 8206 34692 8258
rect 34076 6972 34244 7028
rect 33628 6638 33630 6690
rect 33682 6638 33684 6690
rect 33628 6626 33684 6638
rect 34188 6692 34244 6972
rect 34188 6130 34244 6636
rect 34412 6916 34468 6926
rect 34188 6078 34190 6130
rect 34242 6078 34244 6130
rect 34188 6066 34244 6078
rect 34300 6578 34356 6590
rect 34300 6526 34302 6578
rect 34354 6526 34356 6578
rect 34300 6020 34356 6526
rect 34412 6130 34468 6860
rect 34412 6078 34414 6130
rect 34466 6078 34468 6130
rect 34412 6066 34468 6078
rect 34636 6804 34692 8206
rect 35308 8258 35364 8270
rect 35308 8206 35310 8258
rect 35362 8206 35364 8258
rect 34972 8146 35028 8158
rect 34972 8094 34974 8146
rect 35026 8094 35028 8146
rect 34972 7700 35028 8094
rect 34972 7634 35028 7644
rect 35084 8034 35140 8046
rect 35084 7982 35086 8034
rect 35138 7982 35140 8034
rect 35084 7588 35140 7982
rect 35308 7812 35364 8206
rect 37324 8260 37380 8270
rect 35308 7746 35364 7756
rect 35868 8034 35924 8046
rect 35868 7982 35870 8034
rect 35922 7982 35924 8034
rect 35196 7588 35252 7598
rect 35084 7586 35252 7588
rect 35084 7534 35198 7586
rect 35250 7534 35252 7586
rect 35084 7532 35252 7534
rect 35196 7522 35252 7532
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 34636 6130 34692 6748
rect 34636 6078 34638 6130
rect 34690 6078 34692 6130
rect 34636 6066 34692 6078
rect 35644 6132 35700 6142
rect 34300 5954 34356 5964
rect 35644 6018 35700 6076
rect 35644 5966 35646 6018
rect 35698 5966 35700 6018
rect 35644 5954 35700 5966
rect 33852 5908 33908 5946
rect 35084 5908 35140 5918
rect 33516 5842 33572 5852
rect 33628 5852 33852 5908
rect 33292 5796 33348 5806
rect 33292 5794 33460 5796
rect 33292 5742 33294 5794
rect 33346 5742 33460 5794
rect 33292 5740 33460 5742
rect 33292 5730 33348 5740
rect 33292 5572 33348 5582
rect 33180 5516 33292 5572
rect 33292 5506 33348 5516
rect 33068 5404 33236 5460
rect 32620 5070 32622 5122
rect 32674 5070 32676 5122
rect 32620 5058 32676 5070
rect 33180 5124 33236 5404
rect 32396 4732 33124 4788
rect 32396 4564 32452 4574
rect 32396 4470 32452 4508
rect 32732 4452 32788 4462
rect 32508 3668 32564 3678
rect 32396 3556 32452 3566
rect 32172 3500 32396 3556
rect 32396 3462 32452 3500
rect 32508 800 32564 3612
rect 32732 3442 32788 4396
rect 32956 4340 33012 4350
rect 32956 4246 33012 4284
rect 32732 3390 32734 3442
rect 32786 3390 32788 3442
rect 32732 3378 32788 3390
rect 33068 3554 33124 4732
rect 33180 4562 33236 5068
rect 33292 5010 33348 5022
rect 33292 4958 33294 5010
rect 33346 4958 33348 5010
rect 33292 4900 33348 4958
rect 33292 4834 33348 4844
rect 33404 4676 33460 5740
rect 33404 4610 33460 4620
rect 33516 5682 33572 5694
rect 33516 5630 33518 5682
rect 33570 5630 33572 5682
rect 33516 5124 33572 5630
rect 33180 4510 33182 4562
rect 33234 4510 33236 4562
rect 33180 4498 33236 4510
rect 33292 4450 33348 4462
rect 33292 4398 33294 4450
rect 33346 4398 33348 4450
rect 33180 4340 33236 4350
rect 33292 4340 33348 4398
rect 33236 4284 33348 4340
rect 33404 4340 33460 4350
rect 33180 4274 33236 4284
rect 33068 3502 33070 3554
rect 33122 3502 33124 3554
rect 33068 2884 33124 3502
rect 33068 2818 33124 2828
rect 33180 4116 33236 4126
rect 33180 800 33236 4060
rect 33404 3442 33460 4284
rect 33404 3390 33406 3442
rect 33458 3390 33460 3442
rect 33404 3378 33460 3390
rect 33516 2772 33572 5068
rect 33516 2706 33572 2716
rect 33628 1428 33684 5852
rect 33852 5842 33908 5852
rect 34972 5906 35140 5908
rect 34972 5854 35086 5906
rect 35138 5854 35140 5906
rect 34972 5852 35140 5854
rect 34300 5796 34356 5806
rect 34300 5702 34356 5740
rect 33852 5684 33908 5694
rect 33852 5590 33908 5628
rect 33740 5572 33796 5582
rect 33740 3668 33796 5516
rect 33740 3554 33796 3612
rect 33740 3502 33742 3554
rect 33794 3502 33796 3554
rect 33740 3490 33796 3502
rect 33852 5236 33908 5246
rect 33628 1362 33684 1372
rect 33852 800 33908 5180
rect 34076 5236 34132 5246
rect 33964 4898 34020 4910
rect 33964 4846 33966 4898
rect 34018 4846 34020 4898
rect 33964 4338 34020 4846
rect 33964 4286 33966 4338
rect 34018 4286 34020 4338
rect 33964 4274 34020 4286
rect 34076 3442 34132 5180
rect 34524 4676 34580 4686
rect 34188 4564 34244 4574
rect 34188 4450 34244 4508
rect 34188 4398 34190 4450
rect 34242 4398 34244 4450
rect 34188 4386 34244 4398
rect 34524 3556 34580 4620
rect 34972 4228 35028 5852
rect 35084 5842 35140 5852
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 35308 5012 35364 5022
rect 35308 4918 35364 4956
rect 34972 4162 35028 4172
rect 35084 4226 35140 4238
rect 35084 4174 35086 4226
rect 35138 4174 35140 4226
rect 34524 3462 34580 3500
rect 34748 4116 34804 4126
rect 34076 3390 34078 3442
rect 34130 3390 34132 3442
rect 34076 3378 34132 3390
rect 34748 3442 34804 4060
rect 34748 3390 34750 3442
rect 34802 3390 34804 3442
rect 34748 3378 34804 3390
rect 34860 3892 34916 3902
rect 34860 3388 34916 3836
rect 34972 3780 35028 3790
rect 35084 3780 35140 4174
rect 35532 4228 35588 4238
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 35084 3724 35252 3780
rect 34972 3556 35028 3724
rect 35084 3556 35140 3566
rect 34972 3554 35140 3556
rect 34972 3502 35086 3554
rect 35138 3502 35140 3554
rect 34972 3500 35140 3502
rect 35084 3490 35140 3500
rect 35196 3388 35252 3724
rect 34860 3332 35028 3388
rect 34524 2324 34580 2334
rect 34524 800 34580 2268
rect 34972 980 35028 3332
rect 35084 3332 35252 3388
rect 35420 3444 35476 3454
rect 35532 3444 35588 4172
rect 35868 3780 35924 7982
rect 37100 8036 37156 8046
rect 37100 7942 37156 7980
rect 37324 7588 37380 8204
rect 36428 7476 36484 7486
rect 36428 6916 36484 7420
rect 37324 7362 37380 7532
rect 37324 7310 37326 7362
rect 37378 7310 37380 7362
rect 37324 7298 37380 7310
rect 36428 6802 36484 6860
rect 36428 6750 36430 6802
rect 36482 6750 36484 6802
rect 36428 6738 36484 6750
rect 36540 6692 36596 6702
rect 36092 6130 36148 6142
rect 36092 6078 36094 6130
rect 36146 6078 36148 6130
rect 36092 4564 36148 6078
rect 36540 5348 36596 6636
rect 37324 6692 37380 6702
rect 37436 6692 37492 8988
rect 37548 8978 37604 8988
rect 37772 9602 37828 9614
rect 37772 9550 37774 9602
rect 37826 9550 37828 9602
rect 37660 8034 37716 8046
rect 37660 7982 37662 8034
rect 37714 7982 37716 8034
rect 37660 7924 37716 7982
rect 37660 7858 37716 7868
rect 37772 7476 37828 9550
rect 37996 9604 38052 9614
rect 37996 9510 38052 9548
rect 38332 9602 38388 9614
rect 38332 9550 38334 9602
rect 38386 9550 38388 9602
rect 38220 8930 38276 8942
rect 38220 8878 38222 8930
rect 38274 8878 38276 8930
rect 38108 8258 38164 8270
rect 38108 8206 38110 8258
rect 38162 8206 38164 8258
rect 37772 7410 37828 7420
rect 37884 8034 37940 8046
rect 37884 7982 37886 8034
rect 37938 7982 37940 8034
rect 37884 6804 37940 7982
rect 38108 7698 38164 8206
rect 38220 8036 38276 8878
rect 38332 8260 38388 9550
rect 38556 9602 38612 9614
rect 38556 9550 38558 9602
rect 38610 9550 38612 9602
rect 38556 9492 38612 9550
rect 38556 9426 38612 9436
rect 38892 9602 38948 9614
rect 38892 9550 38894 9602
rect 38946 9550 38948 9602
rect 38332 8194 38388 8204
rect 38668 9156 38724 9166
rect 38668 8258 38724 9100
rect 38668 8206 38670 8258
rect 38722 8206 38724 8258
rect 38668 8194 38724 8206
rect 38892 8260 38948 9550
rect 38892 8194 38948 8204
rect 38780 8036 38836 8046
rect 38220 8034 38836 8036
rect 38220 7982 38782 8034
rect 38834 7982 38836 8034
rect 38220 7980 38836 7982
rect 38780 7970 38836 7980
rect 38892 8036 38948 8046
rect 39004 8036 39060 9660
rect 39452 9716 39508 9726
rect 39452 9622 39508 9660
rect 39116 9602 39172 9614
rect 39116 9550 39118 9602
rect 39170 9550 39172 9602
rect 39116 8146 39172 9550
rect 39788 9156 39844 9772
rect 40796 9716 40852 9726
rect 40348 9714 40852 9716
rect 40348 9662 40798 9714
rect 40850 9662 40852 9714
rect 40348 9660 40852 9662
rect 40012 9604 40068 9614
rect 39788 9090 39844 9100
rect 39900 9602 40068 9604
rect 39900 9550 40014 9602
rect 40066 9550 40068 9602
rect 39900 9548 40068 9550
rect 39900 8484 39956 9548
rect 40012 9538 40068 9548
rect 40348 8930 40404 9660
rect 40796 9650 40852 9660
rect 40908 9716 40964 9726
rect 40908 9602 40964 9660
rect 40908 9550 40910 9602
rect 40962 9550 40964 9602
rect 40908 9538 40964 9550
rect 40348 8878 40350 8930
rect 40402 8878 40404 8930
rect 40348 8866 40404 8878
rect 41020 8930 41076 11788
rect 41244 10388 41300 16044
rect 42140 15986 42196 15998
rect 42140 15934 42142 15986
rect 42194 15934 42196 15986
rect 41692 15314 41748 15326
rect 41692 15262 41694 15314
rect 41746 15262 41748 15314
rect 41692 15204 41748 15262
rect 41692 15138 41748 15148
rect 42028 15204 42084 15214
rect 41468 14084 41524 14094
rect 41468 12516 41524 14028
rect 41580 13970 41636 13982
rect 41580 13918 41582 13970
rect 41634 13918 41636 13970
rect 41580 13860 41636 13918
rect 41580 13794 41636 13804
rect 42028 13746 42084 15148
rect 42140 14642 42196 15934
rect 42252 15876 42308 15886
rect 42252 15782 42308 15820
rect 42140 14590 42142 14642
rect 42194 14590 42196 14642
rect 42140 14578 42196 14590
rect 42028 13694 42030 13746
rect 42082 13694 42084 13746
rect 42028 13682 42084 13694
rect 42364 13748 42420 16044
rect 42588 15876 42644 16380
rect 42588 15810 42644 15820
rect 42700 15652 42756 16940
rect 42924 16212 42980 16940
rect 42924 16146 42980 16156
rect 43036 16100 43092 16110
rect 43036 16006 43092 16044
rect 43148 15876 43204 17388
rect 42700 15586 42756 15596
rect 43036 15820 43204 15876
rect 43260 15876 43316 18956
rect 43372 18116 43428 19182
rect 43932 18564 43988 21980
rect 44044 21588 44100 22094
rect 44268 21700 44324 21710
rect 44268 21606 44324 21644
rect 44044 21522 44100 21532
rect 44156 21586 44212 21598
rect 44156 21534 44158 21586
rect 44210 21534 44212 21586
rect 44156 20244 44212 21534
rect 44156 20178 44212 20188
rect 44044 18564 44100 18574
rect 43372 18050 43428 18060
rect 43708 18562 44100 18564
rect 43708 18510 44046 18562
rect 44098 18510 44100 18562
rect 43708 18508 44100 18510
rect 43372 16660 43428 16670
rect 43372 16098 43428 16604
rect 43708 16660 43764 18508
rect 44044 18498 44100 18508
rect 44268 18450 44324 18462
rect 44268 18398 44270 18450
rect 44322 18398 44324 18450
rect 44044 18228 44100 18238
rect 44044 18226 44212 18228
rect 44044 18174 44046 18226
rect 44098 18174 44212 18226
rect 44044 18172 44212 18174
rect 44044 18162 44100 18172
rect 43932 18004 43988 18014
rect 43708 16594 43764 16604
rect 43820 17780 43876 17790
rect 43820 17220 43876 17724
rect 43596 16324 43652 16334
rect 43372 16046 43374 16098
rect 43426 16046 43428 16098
rect 43372 16034 43428 16046
rect 43484 16212 43540 16222
rect 43484 15986 43540 16156
rect 43596 16100 43652 16268
rect 43708 16100 43764 16110
rect 43596 16098 43764 16100
rect 43596 16046 43710 16098
rect 43762 16046 43764 16098
rect 43596 16044 43764 16046
rect 43708 16034 43764 16044
rect 43484 15934 43486 15986
rect 43538 15934 43540 15986
rect 43484 15922 43540 15934
rect 43260 15820 43428 15876
rect 42476 15202 42532 15214
rect 42476 15150 42478 15202
rect 42530 15150 42532 15202
rect 42476 15148 42532 15150
rect 43036 15148 43092 15820
rect 43260 15652 43316 15662
rect 42476 15092 42644 15148
rect 43036 15092 43204 15148
rect 42588 14642 42644 15092
rect 42588 14590 42590 14642
rect 42642 14590 42644 14642
rect 42588 14578 42644 14590
rect 42700 14756 42756 14766
rect 42700 14530 42756 14700
rect 42700 14478 42702 14530
rect 42754 14478 42756 14530
rect 42700 14466 42756 14478
rect 42924 14420 42980 14430
rect 42924 14326 42980 14364
rect 42476 14306 42532 14318
rect 42476 14254 42478 14306
rect 42530 14254 42532 14306
rect 42476 13972 42532 14254
rect 42532 13916 43092 13972
rect 42476 13878 42532 13916
rect 42700 13748 42756 13758
rect 42364 13692 42644 13748
rect 41692 13636 41748 13646
rect 41692 13634 41972 13636
rect 41692 13582 41694 13634
rect 41746 13582 41972 13634
rect 41692 13580 41972 13582
rect 41692 13570 41748 13580
rect 41916 13076 41972 13580
rect 42028 13076 42084 13086
rect 41916 13074 42084 13076
rect 41916 13022 42030 13074
rect 42082 13022 42084 13074
rect 41916 13020 42084 13022
rect 42028 13010 42084 13020
rect 42364 12964 42420 12974
rect 42364 12870 42420 12908
rect 42028 12852 42084 12862
rect 41468 12460 41748 12516
rect 41692 12402 41748 12460
rect 41692 12350 41694 12402
rect 41746 12350 41748 12402
rect 41580 12180 41636 12190
rect 41580 12086 41636 12124
rect 41468 12068 41524 12078
rect 41468 11282 41524 12012
rect 41692 11396 41748 12350
rect 41692 11330 41748 11340
rect 41468 11230 41470 11282
rect 41522 11230 41524 11282
rect 41468 10612 41524 11230
rect 41468 10610 41636 10612
rect 41468 10558 41470 10610
rect 41522 10558 41636 10610
rect 41468 10556 41636 10558
rect 41468 10546 41524 10556
rect 41020 8878 41022 8930
rect 41074 8878 41076 8930
rect 41020 8866 41076 8878
rect 41132 10332 41300 10388
rect 39788 8428 39956 8484
rect 39116 8094 39118 8146
rect 39170 8094 39172 8146
rect 39116 8082 39172 8094
rect 39564 8258 39620 8270
rect 39564 8206 39566 8258
rect 39618 8206 39620 8258
rect 38892 8034 39060 8036
rect 38892 7982 38894 8034
rect 38946 7982 39060 8034
rect 38892 7980 39060 7982
rect 38892 7970 38948 7980
rect 38108 7646 38110 7698
rect 38162 7646 38164 7698
rect 38108 7634 38164 7646
rect 38892 7812 38948 7822
rect 38668 7588 38724 7598
rect 38668 7494 38724 7532
rect 38444 7250 38500 7262
rect 38444 7198 38446 7250
rect 38498 7198 38500 7250
rect 37996 6804 38052 6814
rect 37884 6802 38052 6804
rect 37884 6750 37998 6802
rect 38050 6750 38052 6802
rect 37884 6748 38052 6750
rect 37996 6738 38052 6748
rect 38444 6804 38500 7198
rect 38444 6738 38500 6748
rect 37324 6690 37492 6692
rect 37324 6638 37326 6690
rect 37378 6638 37492 6690
rect 37324 6636 37492 6638
rect 37324 6626 37380 6636
rect 37660 6018 37716 6030
rect 37660 5966 37662 6018
rect 37714 5966 37716 6018
rect 37100 5908 37156 5918
rect 37548 5908 37604 5918
rect 37100 5906 37268 5908
rect 37100 5854 37102 5906
rect 37154 5854 37268 5906
rect 37100 5852 37268 5854
rect 37100 5842 37156 5852
rect 36428 5124 36484 5134
rect 36540 5124 36596 5292
rect 36428 5122 36596 5124
rect 36428 5070 36430 5122
rect 36482 5070 36596 5122
rect 36428 5068 36596 5070
rect 36764 5684 36820 5694
rect 36428 5058 36484 5068
rect 35980 4340 36036 4350
rect 36092 4340 36148 4508
rect 35980 4338 36148 4340
rect 35980 4286 35982 4338
rect 36034 4286 36148 4338
rect 35980 4284 36148 4286
rect 36428 4788 36484 4798
rect 35980 4274 36036 4284
rect 35868 3714 35924 3724
rect 36316 3892 36372 3902
rect 36428 3892 36484 4732
rect 36652 4452 36708 4462
rect 36652 4358 36708 4396
rect 36540 4340 36596 4350
rect 36540 4246 36596 4284
rect 36428 3836 36596 3892
rect 35420 3442 35588 3444
rect 35420 3390 35422 3442
rect 35474 3390 35588 3442
rect 35420 3388 35588 3390
rect 36316 3388 36372 3836
rect 35420 3378 35476 3388
rect 35980 3332 36372 3388
rect 35084 3220 35140 3332
rect 35084 3154 35140 3164
rect 35980 2436 36036 3332
rect 35980 2370 36036 2380
rect 35868 1876 35924 1886
rect 34972 924 35252 980
rect 35196 800 35252 924
rect 35868 800 35924 1820
rect 36540 800 36596 3836
rect 36764 3442 36820 5628
rect 37100 5124 37156 5134
rect 36876 5122 37156 5124
rect 36876 5070 37102 5122
rect 37154 5070 37156 5122
rect 36876 5068 37156 5070
rect 36876 3892 36932 5068
rect 37100 5058 37156 5068
rect 36876 3554 36932 3836
rect 36876 3502 36878 3554
rect 36930 3502 36932 3554
rect 36876 3490 36932 3502
rect 36764 3390 36766 3442
rect 36818 3390 36820 3442
rect 36764 3378 36820 3390
rect 37212 3388 37268 5852
rect 37324 5124 37380 5134
rect 37324 5030 37380 5068
rect 37548 5122 37604 5852
rect 37548 5070 37550 5122
rect 37602 5070 37604 5122
rect 37548 5058 37604 5070
rect 37660 4676 37716 5966
rect 38108 5796 38164 5806
rect 37884 5124 37940 5134
rect 36988 3332 37268 3388
rect 37436 4620 37716 4676
rect 37772 5068 37884 5124
rect 36988 2996 37044 3332
rect 37436 3108 37492 4620
rect 37660 3556 37716 3566
rect 37772 3556 37828 5068
rect 37884 5058 37940 5068
rect 37660 3554 37828 3556
rect 37660 3502 37662 3554
rect 37714 3502 37828 3554
rect 37660 3500 37828 3502
rect 37660 3490 37716 3500
rect 37548 3442 37604 3454
rect 37548 3390 37550 3442
rect 37602 3390 37604 3442
rect 37548 3388 37604 3390
rect 38108 3388 38164 5740
rect 38332 5348 38388 5358
rect 38332 5010 38388 5292
rect 38332 4958 38334 5010
rect 38386 4958 38388 5010
rect 38332 4946 38388 4958
rect 38892 5010 38948 7756
rect 38892 4958 38894 5010
rect 38946 4958 38948 5010
rect 38892 4676 38948 4958
rect 39116 7700 39172 7710
rect 39116 5010 39172 7644
rect 39228 7586 39284 7598
rect 39228 7534 39230 7586
rect 39282 7534 39284 7586
rect 39228 7028 39284 7534
rect 39228 6962 39284 6972
rect 39564 6692 39620 8206
rect 39788 8260 39844 8428
rect 39788 8194 39844 8204
rect 39900 8260 39956 8270
rect 39900 8258 40292 8260
rect 39900 8206 39902 8258
rect 39954 8206 40292 8258
rect 39900 8204 40292 8206
rect 39900 8194 39956 8204
rect 39676 8036 39732 8046
rect 39676 8034 39844 8036
rect 39676 7982 39678 8034
rect 39730 7982 39844 8034
rect 39676 7980 39844 7982
rect 39676 7970 39732 7980
rect 39676 7700 39732 7710
rect 39676 7606 39732 7644
rect 39564 6626 39620 6636
rect 39788 6244 39844 7980
rect 39788 6178 39844 6188
rect 40012 7474 40068 7486
rect 40012 7422 40014 7474
rect 40066 7422 40068 7474
rect 39564 6020 39620 6030
rect 39564 6018 39732 6020
rect 39564 5966 39566 6018
rect 39618 5966 39732 6018
rect 39564 5964 39732 5966
rect 39564 5954 39620 5964
rect 39340 5908 39396 5918
rect 39340 5906 39508 5908
rect 39340 5854 39342 5906
rect 39394 5854 39508 5906
rect 39340 5852 39508 5854
rect 39340 5842 39396 5852
rect 39452 5348 39508 5852
rect 39452 5124 39508 5292
rect 39564 5124 39620 5134
rect 39452 5122 39620 5124
rect 39452 5070 39566 5122
rect 39618 5070 39620 5122
rect 39452 5068 39620 5070
rect 39564 5058 39620 5068
rect 39676 5124 39732 5964
rect 40012 6018 40068 7422
rect 40124 7028 40180 7038
rect 40124 6802 40180 6972
rect 40124 6750 40126 6802
rect 40178 6750 40180 6802
rect 40124 6738 40180 6750
rect 40236 6692 40292 8204
rect 40796 8258 40852 8270
rect 40796 8206 40798 8258
rect 40850 8206 40852 8258
rect 40796 7700 40852 8206
rect 40908 8148 40964 8158
rect 40908 8054 40964 8092
rect 41020 8146 41076 8158
rect 41020 8094 41022 8146
rect 41074 8094 41076 8146
rect 41020 7812 41076 8094
rect 41020 7746 41076 7756
rect 40908 7700 40964 7710
rect 40796 7644 40908 7700
rect 40908 7586 40964 7644
rect 40908 7534 40910 7586
rect 40962 7534 40964 7586
rect 40908 7522 40964 7534
rect 40460 6692 40516 6702
rect 40236 6636 40404 6692
rect 40348 6244 40404 6636
rect 40460 6690 40964 6692
rect 40460 6638 40462 6690
rect 40514 6638 40964 6690
rect 40460 6636 40964 6638
rect 40460 6626 40516 6636
rect 40684 6468 40740 6478
rect 40684 6374 40740 6412
rect 40348 6188 40740 6244
rect 40012 5966 40014 6018
rect 40066 5966 40068 6018
rect 40012 5796 40068 5966
rect 40012 5730 40068 5740
rect 40236 6130 40292 6142
rect 40236 6078 40238 6130
rect 40290 6078 40292 6130
rect 39676 5058 39732 5068
rect 40012 5124 40068 5134
rect 40012 5030 40068 5068
rect 39116 4958 39118 5010
rect 39170 4958 39172 5010
rect 39116 4946 39172 4958
rect 39788 5010 39844 5022
rect 39788 4958 39790 5010
rect 39842 4958 39844 5010
rect 39788 4900 39844 4958
rect 39788 4834 39844 4844
rect 40124 5010 40180 5022
rect 40124 4958 40126 5010
rect 40178 4958 40180 5010
rect 40124 4676 40180 4958
rect 40236 5012 40292 6078
rect 40460 5124 40516 5134
rect 40460 5030 40516 5068
rect 40236 4946 40292 4956
rect 40572 5010 40628 5022
rect 40572 4958 40574 5010
rect 40626 4958 40628 5010
rect 38892 4620 40180 4676
rect 38668 4338 38724 4350
rect 38668 4286 38670 4338
rect 38722 4286 38724 4338
rect 37548 3332 38164 3388
rect 38556 3444 38612 3454
rect 37436 3042 37492 3052
rect 36988 2930 37044 2940
rect 37212 2212 37268 2222
rect 37212 800 37268 2156
rect 37884 1764 37940 1774
rect 37884 800 37940 1708
rect 38556 800 38612 3388
rect 38668 3332 38724 4286
rect 38668 3266 38724 3276
rect 38892 1652 38948 4620
rect 40236 4562 40292 4574
rect 40236 4510 40238 4562
rect 40290 4510 40292 4562
rect 39116 4450 39172 4462
rect 39116 4398 39118 4450
rect 39170 4398 39172 4450
rect 39116 3388 39172 4398
rect 39340 4004 39396 4014
rect 39340 3666 39396 3948
rect 39340 3614 39342 3666
rect 39394 3614 39396 3666
rect 39340 3602 39396 3614
rect 39900 3668 39956 3678
rect 38892 1586 38948 1596
rect 39004 3332 39172 3388
rect 39004 1540 39060 3332
rect 39004 1474 39060 1484
rect 39228 2884 39284 2894
rect 39228 800 39284 2828
rect 39900 800 39956 3612
rect 40236 3668 40292 4510
rect 40572 4116 40628 4958
rect 40684 4116 40740 6188
rect 40908 4452 40964 6636
rect 41132 6130 41188 10332
rect 41580 9940 41636 10556
rect 41468 9042 41524 9054
rect 41468 8990 41470 9042
rect 41522 8990 41524 9042
rect 41468 8596 41524 8990
rect 41580 9044 41636 9884
rect 41804 9940 41860 9950
rect 41804 9846 41860 9884
rect 41804 9044 41860 9054
rect 41580 9042 41860 9044
rect 41580 8990 41806 9042
rect 41858 8990 41860 9042
rect 41580 8988 41860 8990
rect 41804 8978 41860 8988
rect 41468 8540 41748 8596
rect 41692 8482 41748 8540
rect 41692 8430 41694 8482
rect 41746 8430 41748 8482
rect 41692 8418 41748 8430
rect 41356 8258 41412 8270
rect 41356 8206 41358 8258
rect 41410 8206 41412 8258
rect 41244 7812 41300 7822
rect 41244 7474 41300 7756
rect 41244 7422 41246 7474
rect 41298 7422 41300 7474
rect 41244 7410 41300 7422
rect 41356 7476 41412 8206
rect 42028 7698 42084 12796
rect 42364 12404 42420 12414
rect 42364 12310 42420 12348
rect 42140 10500 42196 10510
rect 42140 10498 42532 10500
rect 42140 10446 42142 10498
rect 42194 10446 42532 10498
rect 42140 10444 42532 10446
rect 42140 10434 42196 10444
rect 42364 10276 42420 10286
rect 42364 9940 42420 10220
rect 42364 9826 42420 9884
rect 42476 9938 42532 10444
rect 42588 10052 42644 13692
rect 42700 12852 42756 13692
rect 42812 13634 42868 13646
rect 42812 13582 42814 13634
rect 42866 13582 42868 13634
rect 42812 13076 42868 13582
rect 42924 13076 42980 13086
rect 42812 13074 42980 13076
rect 42812 13022 42926 13074
rect 42978 13022 42980 13074
rect 42812 13020 42980 13022
rect 42924 13010 42980 13020
rect 43036 12962 43092 13916
rect 43036 12910 43038 12962
rect 43090 12910 43092 12962
rect 43036 12898 43092 12910
rect 42812 12852 42868 12862
rect 42700 12850 42868 12852
rect 42700 12798 42814 12850
rect 42866 12798 42868 12850
rect 42700 12796 42868 12798
rect 42812 12786 42868 12796
rect 43148 12852 43204 15092
rect 43148 12786 43204 12796
rect 42588 9986 42644 9996
rect 42476 9886 42478 9938
rect 42530 9886 42532 9938
rect 42476 9874 42532 9886
rect 42364 9774 42366 9826
rect 42418 9774 42420 9826
rect 42364 9762 42420 9774
rect 42588 9828 42644 9838
rect 42924 9828 42980 9838
rect 42644 9826 42980 9828
rect 42644 9774 42926 9826
rect 42978 9774 42980 9826
rect 42644 9772 42980 9774
rect 42588 9734 42644 9772
rect 42924 9762 42980 9772
rect 42140 9604 42196 9614
rect 42140 9510 42196 9548
rect 43036 9602 43092 9614
rect 43036 9550 43038 9602
rect 43090 9550 43092 9602
rect 43036 9380 43092 9550
rect 43148 9604 43204 9614
rect 43148 9510 43204 9548
rect 42588 9324 43092 9380
rect 42588 9154 42644 9324
rect 42588 9102 42590 9154
rect 42642 9102 42644 9154
rect 42588 9090 42644 9102
rect 42476 8258 42532 8270
rect 42476 8206 42478 8258
rect 42530 8206 42532 8258
rect 42364 8148 42420 8158
rect 42364 8054 42420 8092
rect 42476 7812 42532 8206
rect 43036 8260 43092 8270
rect 43036 8166 43092 8204
rect 42924 8036 42980 8046
rect 43260 8036 43316 15596
rect 43372 10052 43428 15820
rect 43372 9986 43428 9996
rect 43372 9602 43428 9614
rect 43372 9550 43374 9602
rect 43426 9550 43428 9602
rect 43372 9492 43428 9550
rect 43372 9426 43428 9436
rect 42924 8034 43316 8036
rect 42924 7982 42926 8034
rect 42978 7982 43316 8034
rect 42924 7980 43316 7982
rect 43596 8148 43652 8158
rect 43708 8148 43764 8158
rect 43652 8146 43764 8148
rect 43652 8094 43710 8146
rect 43762 8094 43764 8146
rect 43652 8092 43764 8094
rect 42924 7970 42980 7980
rect 42476 7746 42532 7756
rect 42028 7646 42030 7698
rect 42082 7646 42084 7698
rect 42028 7634 42084 7646
rect 41356 7410 41412 7420
rect 41468 7588 41524 7598
rect 41132 6078 41134 6130
rect 41186 6078 41188 6130
rect 41132 6066 41188 6078
rect 41468 4452 41524 7532
rect 43036 7586 43092 7598
rect 43036 7534 43038 7586
rect 43090 7534 43092 7586
rect 41916 7476 41972 7486
rect 41580 7474 41972 7476
rect 41580 7422 41918 7474
rect 41970 7422 41972 7474
rect 41580 7420 41972 7422
rect 41580 7362 41636 7420
rect 41916 7410 41972 7420
rect 43036 7476 43092 7534
rect 41580 7310 41582 7362
rect 41634 7310 41636 7362
rect 41580 6578 41636 7310
rect 43036 6804 43092 7420
rect 43036 6738 43092 6748
rect 41580 6526 41582 6578
rect 41634 6526 41636 6578
rect 41580 6514 41636 6526
rect 43596 6578 43652 8092
rect 43708 8082 43764 8092
rect 43596 6526 43598 6578
rect 43650 6526 43652 6578
rect 43596 6514 43652 6526
rect 43820 6132 43876 17164
rect 43932 16098 43988 17948
rect 44044 17892 44100 17902
rect 44044 16322 44100 17836
rect 44044 16270 44046 16322
rect 44098 16270 44100 16322
rect 44044 16258 44100 16270
rect 43932 16046 43934 16098
rect 43986 16046 43988 16098
rect 43932 16034 43988 16046
rect 44044 15876 44100 15886
rect 44044 15782 44100 15820
rect 43932 14754 43988 14766
rect 43932 14702 43934 14754
rect 43986 14702 43988 14754
rect 43932 14642 43988 14702
rect 43932 14590 43934 14642
rect 43986 14590 43988 14642
rect 43932 14578 43988 14590
rect 43932 9604 43988 9614
rect 43932 8932 43988 9548
rect 43932 8866 43988 8876
rect 44156 8372 44212 18172
rect 44268 17106 44324 18398
rect 44380 17556 44436 22428
rect 44492 20132 44548 20142
rect 44492 20038 44548 20076
rect 44604 17668 44660 22540
rect 44716 20018 44772 20030
rect 44716 19966 44718 20018
rect 44770 19966 44772 20018
rect 44716 18228 44772 19966
rect 44828 19234 44884 22652
rect 45164 22370 45220 22988
rect 45164 22318 45166 22370
rect 45218 22318 45220 22370
rect 45164 22306 45220 22318
rect 45276 21812 45332 25566
rect 45388 24612 45444 26852
rect 45500 26178 45556 26190
rect 45500 26126 45502 26178
rect 45554 26126 45556 26178
rect 45500 26068 45556 26126
rect 45500 26002 45556 26012
rect 45500 25732 45556 25742
rect 45500 25394 45556 25676
rect 45500 25342 45502 25394
rect 45554 25342 45556 25394
rect 45500 25330 45556 25342
rect 45612 25508 45668 30716
rect 46060 30660 46116 31948
rect 46284 31778 46340 31790
rect 46284 31726 46286 31778
rect 46338 31726 46340 31778
rect 45948 30604 46116 30660
rect 46172 31666 46228 31678
rect 46172 31614 46174 31666
rect 46226 31614 46228 31666
rect 46172 31106 46228 31614
rect 46172 31054 46174 31106
rect 46226 31054 46228 31106
rect 45724 30212 45780 30222
rect 45724 30118 45780 30156
rect 45948 29988 46004 30604
rect 45500 24948 45556 24958
rect 45612 24948 45668 25452
rect 45500 24946 45668 24948
rect 45500 24894 45502 24946
rect 45554 24894 45668 24946
rect 45500 24892 45668 24894
rect 45724 29932 46004 29988
rect 46060 30436 46116 30446
rect 46060 29986 46116 30380
rect 46172 30212 46228 31054
rect 46172 30118 46228 30156
rect 46284 31108 46340 31726
rect 46284 30994 46340 31052
rect 46284 30942 46286 30994
rect 46338 30942 46340 30994
rect 46284 30324 46340 30942
rect 46508 30772 46564 32510
rect 46508 30706 46564 30716
rect 46620 35252 46788 35308
rect 46284 30210 46340 30268
rect 46620 30212 46676 35252
rect 46732 33122 46788 33134
rect 46732 33070 46734 33122
rect 46786 33070 46788 33122
rect 46732 32674 46788 33070
rect 46732 32622 46734 32674
rect 46786 32622 46788 32674
rect 46732 30996 46788 32622
rect 47068 31106 47124 31118
rect 47068 31054 47070 31106
rect 47122 31054 47124 31106
rect 46844 30996 46900 31006
rect 46732 30994 46900 30996
rect 46732 30942 46846 30994
rect 46898 30942 46900 30994
rect 46732 30940 46900 30942
rect 46284 30158 46286 30210
rect 46338 30158 46340 30210
rect 46284 30146 46340 30158
rect 46396 30156 46676 30212
rect 46732 30324 46788 30334
rect 46732 30210 46788 30268
rect 46732 30158 46734 30210
rect 46786 30158 46788 30210
rect 46060 29934 46062 29986
rect 46114 29934 46116 29986
rect 45500 24882 45556 24892
rect 45388 24546 45444 24556
rect 45724 24164 45780 29932
rect 46060 29922 46116 29934
rect 45836 28532 45892 28542
rect 45836 27188 45892 28476
rect 46396 27412 46452 30156
rect 46732 30146 46788 30158
rect 46844 29876 46900 30940
rect 46956 30212 47012 30222
rect 47068 30212 47124 31054
rect 47012 30156 47124 30212
rect 47180 30212 47236 30222
rect 46956 30118 47012 30156
rect 47180 30118 47236 30156
rect 47292 30100 47348 30110
rect 47292 30006 47348 30044
rect 46732 29820 46900 29876
rect 46396 27356 46564 27412
rect 46284 27300 46340 27310
rect 46284 27298 46452 27300
rect 46284 27246 46286 27298
rect 46338 27246 46452 27298
rect 46284 27244 46452 27246
rect 46284 27234 46340 27244
rect 45836 27094 45892 27132
rect 46396 27074 46452 27244
rect 46396 27022 46398 27074
rect 46450 27022 46452 27074
rect 46396 27010 46452 27022
rect 46060 26516 46116 26526
rect 45948 26292 46004 26302
rect 46060 26292 46116 26460
rect 46172 26404 46228 26414
rect 46172 26310 46228 26348
rect 45948 26290 46116 26292
rect 45948 26238 45950 26290
rect 46002 26238 46116 26290
rect 45948 26236 46116 26238
rect 46396 26292 46452 26302
rect 45836 25620 45892 25630
rect 45836 25506 45892 25564
rect 45836 25454 45838 25506
rect 45890 25454 45892 25506
rect 45836 25442 45892 25454
rect 45612 24108 45780 24164
rect 45836 25284 45892 25294
rect 45388 23716 45444 23726
rect 45388 23622 45444 23660
rect 45500 22146 45556 22158
rect 45500 22094 45502 22146
rect 45554 22094 45556 22146
rect 45388 21812 45444 21822
rect 45276 21756 45388 21812
rect 45388 21746 45444 21756
rect 45500 21364 45556 22094
rect 45612 22148 45668 24108
rect 45724 23940 45780 23950
rect 45724 23846 45780 23884
rect 45836 23268 45892 25228
rect 45948 24722 46004 26236
rect 46396 26198 46452 26236
rect 46508 25620 46564 27356
rect 46620 27300 46676 27310
rect 46620 27186 46676 27244
rect 46620 27134 46622 27186
rect 46674 27134 46676 27186
rect 46620 27122 46676 27134
rect 46732 26516 46788 29820
rect 47292 27074 47348 27086
rect 47292 27022 47294 27074
rect 47346 27022 47348 27074
rect 46732 26450 46788 26460
rect 46844 26962 46900 26974
rect 46844 26910 46846 26962
rect 46898 26910 46900 26962
rect 46844 26404 46900 26910
rect 47068 26962 47124 26974
rect 47068 26910 47070 26962
rect 47122 26910 47124 26962
rect 47068 26908 47124 26910
rect 46844 26310 46900 26348
rect 46956 26852 47124 26908
rect 47292 26964 47348 27022
rect 47516 27076 47572 27086
rect 47516 26982 47572 27020
rect 47852 27074 47908 27086
rect 47852 27022 47854 27074
rect 47906 27022 47908 27074
rect 47292 26898 47348 26908
rect 47740 26962 47796 26974
rect 47740 26910 47742 26962
rect 47794 26910 47796 26962
rect 46620 26292 46676 26302
rect 46620 26198 46676 26236
rect 46956 26290 47012 26852
rect 47740 26404 47796 26910
rect 47740 26310 47796 26348
rect 47292 26292 47348 26302
rect 46956 26238 46958 26290
rect 47010 26238 47012 26290
rect 46956 26180 47012 26238
rect 46060 25508 46116 25518
rect 46284 25508 46340 25518
rect 46116 25506 46340 25508
rect 46116 25454 46286 25506
rect 46338 25454 46340 25506
rect 46116 25452 46340 25454
rect 46060 25442 46116 25452
rect 45948 24670 45950 24722
rect 46002 24670 46004 24722
rect 45948 24658 46004 24670
rect 46172 24834 46228 24846
rect 46172 24782 46174 24834
rect 46226 24782 46228 24834
rect 46060 23940 46116 23950
rect 46172 23940 46228 24782
rect 46284 24052 46340 25452
rect 46508 24948 46564 25564
rect 46844 26124 46956 26180
rect 46620 25396 46676 25406
rect 46844 25396 46900 26124
rect 46956 26086 47012 26124
rect 47180 26290 47348 26292
rect 47180 26238 47294 26290
rect 47346 26238 47348 26290
rect 47180 26236 47348 26238
rect 47068 25732 47124 25742
rect 47180 25732 47236 26236
rect 47292 26226 47348 26236
rect 47852 26290 47908 27022
rect 47852 26238 47854 26290
rect 47906 26238 47908 26290
rect 47516 26178 47572 26190
rect 47516 26126 47518 26178
rect 47570 26126 47572 26178
rect 47516 26068 47572 26126
rect 47852 26180 47908 26238
rect 47852 26114 47908 26124
rect 47516 26002 47572 26012
rect 47068 25730 47236 25732
rect 47068 25678 47070 25730
rect 47122 25678 47236 25730
rect 47068 25676 47236 25678
rect 47068 25666 47124 25676
rect 46620 25394 46900 25396
rect 46620 25342 46622 25394
rect 46674 25342 46900 25394
rect 46620 25340 46900 25342
rect 46956 25396 47012 25406
rect 46620 25330 46676 25340
rect 46956 25302 47012 25340
rect 47516 25396 47572 25406
rect 47516 25302 47572 25340
rect 46620 24948 46676 24958
rect 46508 24946 46676 24948
rect 46508 24894 46622 24946
rect 46674 24894 46676 24946
rect 46508 24892 46676 24894
rect 46620 24882 46676 24892
rect 47068 24612 47124 24622
rect 46956 24610 47124 24612
rect 46956 24558 47070 24610
rect 47122 24558 47124 24610
rect 46956 24556 47124 24558
rect 46284 23996 46788 24052
rect 45948 23938 46228 23940
rect 45948 23886 46062 23938
rect 46114 23886 46228 23938
rect 45948 23884 46228 23886
rect 46732 23938 46788 23996
rect 46732 23886 46734 23938
rect 46786 23886 46788 23938
rect 45948 23492 46004 23884
rect 46060 23874 46116 23884
rect 46732 23874 46788 23886
rect 46396 23826 46452 23838
rect 46396 23774 46398 23826
rect 46450 23774 46452 23826
rect 46060 23716 46116 23726
rect 46060 23622 46116 23660
rect 46396 23604 46452 23774
rect 46396 23538 46452 23548
rect 45948 23436 46116 23492
rect 45836 23202 45892 23212
rect 45948 23154 46004 23166
rect 45948 23102 45950 23154
rect 46002 23102 46004 23154
rect 45948 22372 46004 23102
rect 46060 23156 46116 23436
rect 46284 23380 46340 23390
rect 46844 23380 46900 23390
rect 46284 23378 46788 23380
rect 46284 23326 46286 23378
rect 46338 23326 46788 23378
rect 46284 23324 46788 23326
rect 46284 23314 46340 23324
rect 46732 23266 46788 23324
rect 46844 23286 46900 23324
rect 46732 23214 46734 23266
rect 46786 23214 46788 23266
rect 46732 23202 46788 23214
rect 46172 23156 46228 23166
rect 46060 23154 46228 23156
rect 46060 23102 46174 23154
rect 46226 23102 46228 23154
rect 46060 23100 46228 23102
rect 45948 22278 46004 22316
rect 46172 22370 46228 23100
rect 46284 23156 46340 23166
rect 46284 22482 46340 23100
rect 46508 23154 46564 23166
rect 46508 23102 46510 23154
rect 46562 23102 46564 23154
rect 46508 22596 46564 23102
rect 46844 22932 46900 22942
rect 46844 22838 46900 22876
rect 46732 22596 46788 22606
rect 46508 22594 46788 22596
rect 46508 22542 46734 22594
rect 46786 22542 46788 22594
rect 46508 22540 46788 22542
rect 46732 22530 46788 22540
rect 46956 22596 47012 24556
rect 47068 24546 47124 24556
rect 47964 24388 48020 43652
rect 47964 24322 48020 24332
rect 48076 29204 48132 29214
rect 48076 24052 48132 29148
rect 47516 24050 48132 24052
rect 47516 23998 48078 24050
rect 48130 23998 48132 24050
rect 47516 23996 48132 23998
rect 47292 23940 47348 23950
rect 46284 22430 46286 22482
rect 46338 22430 46340 22482
rect 46284 22418 46340 22430
rect 46172 22318 46174 22370
rect 46226 22318 46228 22370
rect 45612 22092 45892 22148
rect 45724 21810 45780 21822
rect 45724 21758 45726 21810
rect 45778 21758 45780 21810
rect 45612 21588 45668 21598
rect 45612 21494 45668 21532
rect 45052 20802 45108 20814
rect 45052 20750 45054 20802
rect 45106 20750 45108 20802
rect 45052 20244 45108 20750
rect 45500 20802 45556 21308
rect 45500 20750 45502 20802
rect 45554 20750 45556 20802
rect 45500 20738 45556 20750
rect 45052 20178 45108 20188
rect 44828 19182 44830 19234
rect 44882 19182 44884 19234
rect 44828 19170 44884 19182
rect 45388 19234 45444 19246
rect 45388 19182 45390 19234
rect 45442 19182 45444 19234
rect 44716 18162 44772 18172
rect 45052 18788 45108 18798
rect 44940 17780 44996 17790
rect 44828 17668 44884 17678
rect 44604 17666 44884 17668
rect 44604 17614 44830 17666
rect 44882 17614 44884 17666
rect 44604 17612 44884 17614
rect 44828 17602 44884 17612
rect 44380 17500 44660 17556
rect 44268 17054 44270 17106
rect 44322 17054 44324 17106
rect 44268 17042 44324 17054
rect 44604 16882 44660 17500
rect 44604 16830 44606 16882
rect 44658 16830 44660 16882
rect 44604 16818 44660 16830
rect 44940 17220 44996 17724
rect 44268 16212 44324 16222
rect 44268 14754 44324 16156
rect 44940 16210 44996 17164
rect 44940 16158 44942 16210
rect 44994 16158 44996 16210
rect 44940 16146 44996 16158
rect 45052 17668 45108 18732
rect 45388 17892 45444 19182
rect 45612 18452 45668 18462
rect 45612 18358 45668 18396
rect 45500 18340 45556 18350
rect 45500 18246 45556 18284
rect 45388 17826 45444 17836
rect 45052 15988 45108 17612
rect 45388 17666 45444 17678
rect 45388 17614 45390 17666
rect 45442 17614 45444 17666
rect 45388 16324 45444 17614
rect 45612 16996 45668 17006
rect 45612 16902 45668 16940
rect 45724 16772 45780 21758
rect 45836 20804 45892 22092
rect 46172 21700 46228 22318
rect 46396 22258 46452 22270
rect 46396 22206 46398 22258
rect 46450 22206 46452 22258
rect 46396 22148 46452 22206
rect 46844 22260 46900 22270
rect 46956 22260 47012 22540
rect 47068 23714 47124 23726
rect 47068 23662 47070 23714
rect 47122 23662 47124 23714
rect 47068 23604 47124 23662
rect 47068 22372 47124 23548
rect 47292 23380 47348 23884
rect 47404 23826 47460 23838
rect 47404 23774 47406 23826
rect 47458 23774 47460 23826
rect 47404 23716 47460 23774
rect 47516 23826 47572 23996
rect 48076 23986 48132 23996
rect 47516 23774 47518 23826
rect 47570 23774 47572 23826
rect 47516 23762 47572 23774
rect 47404 23650 47460 23660
rect 47740 23714 47796 23726
rect 47740 23662 47742 23714
rect 47794 23662 47796 23714
rect 47740 23492 47796 23662
rect 47740 23436 48356 23492
rect 47404 23380 47460 23390
rect 47292 23378 47460 23380
rect 47292 23326 47406 23378
rect 47458 23326 47460 23378
rect 47292 23324 47460 23326
rect 47404 23314 47460 23324
rect 47964 23268 48020 23278
rect 47964 23174 48020 23212
rect 47292 23156 47348 23166
rect 47852 23156 47908 23166
rect 47292 23062 47348 23100
rect 47628 23154 47908 23156
rect 47628 23102 47854 23154
rect 47906 23102 47908 23154
rect 47628 23100 47908 23102
rect 47404 22932 47460 22942
rect 47292 22930 47460 22932
rect 47292 22878 47406 22930
rect 47458 22878 47460 22930
rect 47292 22876 47460 22878
rect 47068 22306 47124 22316
rect 47180 22370 47236 22382
rect 47180 22318 47182 22370
rect 47234 22318 47236 22370
rect 46844 22258 47012 22260
rect 46844 22206 46846 22258
rect 46898 22206 47012 22258
rect 46844 22204 47012 22206
rect 46844 22194 46900 22204
rect 47180 22148 47236 22318
rect 46396 22082 46452 22092
rect 47012 22092 47236 22148
rect 47012 22036 47068 22092
rect 46956 21980 47068 22036
rect 46172 21634 46228 21644
rect 46396 21812 46452 21822
rect 46396 21698 46452 21756
rect 46396 21646 46398 21698
rect 46450 21646 46452 21698
rect 46396 21634 46452 21646
rect 46284 21588 46340 21598
rect 46172 21140 46228 21150
rect 45948 20804 46004 20814
rect 45836 20802 46004 20804
rect 45836 20750 45950 20802
rect 46002 20750 46004 20802
rect 45836 20748 46004 20750
rect 45948 19572 46004 20748
rect 45948 19506 46004 19516
rect 45612 16716 45780 16772
rect 45388 16258 45444 16268
rect 45500 16548 45556 16558
rect 45500 16098 45556 16492
rect 45500 16046 45502 16098
rect 45554 16046 45556 16098
rect 45500 16034 45556 16046
rect 44268 14702 44270 14754
rect 44322 14702 44324 14754
rect 44268 14690 44324 14702
rect 44380 15932 45108 15988
rect 44380 14642 44436 15932
rect 45500 15314 45556 15326
rect 45500 15262 45502 15314
rect 45554 15262 45556 15314
rect 44604 15202 44660 15214
rect 44604 15150 44606 15202
rect 44658 15150 44660 15202
rect 44604 15148 44660 15150
rect 44604 15092 45108 15148
rect 44380 14590 44382 14642
rect 44434 14590 44436 14642
rect 44380 14578 44436 14590
rect 45052 14530 45108 15092
rect 45164 14756 45220 14766
rect 45164 14662 45220 14700
rect 45052 14478 45054 14530
rect 45106 14478 45108 14530
rect 45052 14466 45108 14478
rect 45500 14308 45556 15262
rect 45500 14242 45556 14252
rect 45276 13748 45332 13758
rect 44940 13746 45332 13748
rect 44940 13694 45278 13746
rect 45330 13694 45332 13746
rect 44940 13692 45332 13694
rect 44940 13634 44996 13692
rect 45276 13682 45332 13692
rect 45388 13748 45444 13758
rect 45388 13654 45444 13692
rect 44940 13582 44942 13634
rect 44994 13582 44996 13634
rect 44940 13570 44996 13582
rect 45276 13524 45332 13534
rect 44828 11284 44884 11294
rect 44268 11282 44884 11284
rect 44268 11230 44830 11282
rect 44882 11230 44884 11282
rect 44268 11228 44884 11230
rect 44268 10498 44324 11228
rect 44828 11218 44884 11228
rect 45164 11282 45220 11294
rect 45164 11230 45166 11282
rect 45218 11230 45220 11282
rect 44268 10446 44270 10498
rect 44322 10446 44324 10498
rect 44268 10434 44324 10446
rect 45164 11172 45220 11230
rect 45164 10276 45220 11116
rect 45164 10210 45220 10220
rect 45276 10052 45332 13468
rect 45612 11844 45668 16716
rect 46060 16548 46116 16558
rect 45836 16324 45892 16334
rect 45724 15874 45780 15886
rect 45724 15822 45726 15874
rect 45778 15822 45780 15874
rect 45724 15764 45780 15822
rect 45724 15698 45780 15708
rect 45836 15876 45892 16268
rect 46060 16098 46116 16492
rect 46060 16046 46062 16098
rect 46114 16046 46116 16098
rect 46060 16034 46116 16046
rect 45836 15148 45892 15820
rect 45724 15092 45892 15148
rect 45724 14642 45780 15092
rect 45724 14590 45726 14642
rect 45778 14590 45780 14642
rect 45724 14578 45780 14590
rect 45612 11778 45668 11788
rect 45164 9996 45332 10052
rect 44716 8932 44772 8942
rect 45052 8932 45108 8942
rect 44716 8930 45108 8932
rect 44716 8878 44718 8930
rect 44770 8878 45054 8930
rect 45106 8878 45108 8930
rect 44716 8876 45108 8878
rect 44716 8866 44772 8876
rect 45052 8866 45108 8876
rect 45164 8708 45220 9996
rect 45836 9828 45892 9838
rect 45276 8932 45332 8942
rect 45276 8838 45332 8876
rect 45164 8652 45332 8708
rect 43932 8316 44212 8372
rect 43932 8036 43988 8316
rect 44716 8260 44772 8270
rect 44716 8166 44772 8204
rect 43932 7474 43988 7980
rect 44044 8146 44100 8158
rect 44044 8094 44046 8146
rect 44098 8094 44100 8146
rect 44044 7588 44100 8094
rect 44044 7522 44100 7532
rect 44380 8148 44436 8158
rect 43932 7422 43934 7474
rect 43986 7422 43988 7474
rect 43932 7410 43988 7422
rect 44380 7140 44436 8092
rect 45052 8148 45108 8158
rect 45052 8054 45108 8092
rect 44940 8034 44996 8046
rect 44940 7982 44942 8034
rect 44994 7982 44996 8034
rect 44940 7700 44996 7982
rect 44940 7634 44996 7644
rect 44492 7588 44548 7598
rect 44492 7494 44548 7532
rect 44268 7084 44436 7140
rect 44268 7028 44324 7084
rect 44268 6690 44324 6972
rect 44268 6638 44270 6690
rect 44322 6638 44324 6690
rect 44268 6626 44324 6638
rect 44380 6244 44436 6254
rect 44044 6132 44100 6142
rect 43820 6130 44100 6132
rect 43820 6078 44046 6130
rect 44098 6078 44100 6130
rect 43820 6076 44100 6078
rect 44044 6066 44100 6076
rect 42252 6020 42308 6030
rect 43148 6020 43204 6030
rect 42252 5926 42308 5964
rect 43036 6018 43204 6020
rect 43036 5966 43150 6018
rect 43202 5966 43204 6018
rect 43036 5964 43204 5966
rect 41804 5908 41860 5918
rect 42476 5908 42532 5918
rect 41804 5814 41860 5852
rect 42364 5852 42476 5908
rect 41580 5682 41636 5694
rect 41580 5630 41582 5682
rect 41634 5630 41636 5682
rect 41580 4900 41636 5630
rect 42028 5682 42084 5694
rect 42028 5630 42030 5682
rect 42082 5630 42084 5682
rect 41580 4834 41636 4844
rect 41804 5124 41860 5134
rect 42028 5124 42084 5630
rect 41860 5068 42084 5124
rect 42140 5236 42196 5246
rect 41580 4452 41636 4462
rect 40908 4450 41412 4452
rect 40908 4398 40910 4450
rect 40962 4398 41412 4450
rect 40908 4396 41412 4398
rect 40908 4386 40964 4396
rect 41244 4226 41300 4238
rect 41244 4174 41246 4226
rect 41298 4174 41300 4226
rect 40796 4116 40852 4126
rect 40684 4060 40796 4116
rect 40572 4050 40628 4060
rect 40796 4050 40852 4060
rect 41244 4116 41300 4174
rect 41244 4050 41300 4060
rect 40236 3602 40292 3612
rect 41132 3892 41188 3902
rect 40572 3556 40628 3566
rect 40572 800 40628 3500
rect 41132 3388 41188 3836
rect 41356 3554 41412 4396
rect 41356 3502 41358 3554
rect 41410 3502 41412 3554
rect 41356 3490 41412 3502
rect 41468 4450 41636 4452
rect 41468 4398 41582 4450
rect 41634 4398 41636 4450
rect 41468 4396 41636 4398
rect 41468 3442 41524 4396
rect 41580 4386 41636 4396
rect 41804 3666 41860 5068
rect 42140 4562 42196 5180
rect 42140 4510 42142 4562
rect 42194 4510 42196 4562
rect 42140 4498 42196 4510
rect 41804 3614 41806 3666
rect 41858 3614 41860 3666
rect 41804 3602 41860 3614
rect 41916 3892 41972 3902
rect 41468 3390 41470 3442
rect 41522 3390 41524 3442
rect 41132 3332 41300 3388
rect 41468 3378 41524 3390
rect 41244 800 41300 3332
rect 41916 800 41972 3836
rect 42252 3556 42308 3566
rect 42252 3442 42308 3500
rect 42252 3390 42254 3442
rect 42306 3390 42308 3442
rect 42252 3378 42308 3390
rect 42364 3388 42420 5852
rect 42476 5842 42532 5852
rect 42700 5122 42756 5134
rect 42700 5070 42702 5122
rect 42754 5070 42756 5122
rect 42476 5012 42532 5022
rect 42476 4900 42532 4956
rect 42476 4844 42644 4900
rect 42588 4450 42644 4844
rect 42588 4398 42590 4450
rect 42642 4398 42644 4450
rect 42588 4386 42644 4398
rect 42700 4340 42756 5070
rect 42700 4274 42756 4284
rect 42812 4898 42868 4910
rect 42812 4846 42814 4898
rect 42866 4846 42868 4898
rect 42588 3780 42644 3790
rect 42364 3332 42532 3388
rect 42476 3220 42532 3332
rect 42476 3154 42532 3164
rect 42588 800 42644 3724
rect 42812 3556 42868 4846
rect 43036 4004 43092 5964
rect 43148 5954 43204 5964
rect 44268 5908 44324 5918
rect 43260 5236 43316 5246
rect 43148 5010 43204 5022
rect 43148 4958 43150 5010
rect 43202 4958 43204 5010
rect 43148 4228 43204 4958
rect 43148 4162 43204 4172
rect 43036 3938 43092 3948
rect 43036 3556 43092 3566
rect 42812 3554 43092 3556
rect 42812 3502 43038 3554
rect 43090 3502 43092 3554
rect 42812 3500 43092 3502
rect 43036 3444 43092 3500
rect 43036 3378 43092 3388
rect 43260 800 43316 5180
rect 43708 4564 43764 4574
rect 43708 3554 43764 4508
rect 44156 4340 44212 4350
rect 44268 4340 44324 5852
rect 44156 4338 44324 4340
rect 44156 4286 44158 4338
rect 44210 4286 44324 4338
rect 44156 4284 44324 4286
rect 44156 4274 44212 4284
rect 43708 3502 43710 3554
rect 43762 3502 43764 3554
rect 43708 3490 43764 3502
rect 43932 4004 43988 4014
rect 43932 800 43988 3948
rect 44380 3442 44436 6188
rect 45164 6020 45220 6030
rect 45164 5926 45220 5964
rect 44828 5908 44884 5918
rect 44828 5122 44884 5852
rect 44828 5070 44830 5122
rect 44882 5070 44884 5122
rect 44828 5058 44884 5070
rect 45164 5572 45220 5582
rect 44380 3390 44382 3442
rect 44434 3390 44436 3442
rect 44380 3378 44436 3390
rect 44604 3668 44660 3678
rect 44604 800 44660 3612
rect 45164 3332 45220 5516
rect 45276 4226 45332 8652
rect 45500 8034 45556 8046
rect 45500 7982 45502 8034
rect 45554 7982 45556 8034
rect 45500 5236 45556 7982
rect 45724 6804 45780 6814
rect 45500 5170 45556 5180
rect 45612 6020 45668 6030
rect 45388 5010 45444 5022
rect 45388 4958 45390 5010
rect 45442 4958 45444 5010
rect 45388 4900 45444 4958
rect 45388 4834 45444 4844
rect 45612 4564 45668 5964
rect 45612 4450 45668 4508
rect 45612 4398 45614 4450
rect 45666 4398 45668 4450
rect 45612 4386 45668 4398
rect 45276 4174 45278 4226
rect 45330 4174 45332 4226
rect 45276 4162 45332 4174
rect 45724 3666 45780 6748
rect 45836 4898 45892 9772
rect 46172 8260 46228 21084
rect 46284 20018 46340 21532
rect 46956 20804 47012 21980
rect 47180 21698 47236 21710
rect 47180 21646 47182 21698
rect 47234 21646 47236 21698
rect 47180 21588 47236 21646
rect 47180 21522 47236 21532
rect 47068 20804 47124 20814
rect 46956 20748 47068 20804
rect 47068 20710 47124 20748
rect 46396 20690 46452 20702
rect 46396 20638 46398 20690
rect 46450 20638 46452 20690
rect 46396 20244 46452 20638
rect 46396 20178 46452 20188
rect 46844 20578 46900 20590
rect 46844 20526 46846 20578
rect 46898 20526 46900 20578
rect 46284 19966 46286 20018
rect 46338 19966 46340 20018
rect 46284 19236 46340 19966
rect 46732 20018 46788 20030
rect 46732 19966 46734 20018
rect 46786 19966 46788 20018
rect 46732 19348 46788 19966
rect 46284 19170 46340 19180
rect 46620 19236 46676 19274
rect 46620 19170 46676 19180
rect 46620 19012 46676 19022
rect 46620 18918 46676 18956
rect 46620 18676 46676 18686
rect 46732 18676 46788 19292
rect 46676 18620 46788 18676
rect 46620 18610 46676 18620
rect 46284 18564 46340 18574
rect 46284 15988 46340 18508
rect 46284 15922 46340 15932
rect 46732 17780 46788 17790
rect 46732 16882 46788 17724
rect 46732 16830 46734 16882
rect 46786 16830 46788 16882
rect 46396 15876 46452 15886
rect 46396 15782 46452 15820
rect 46396 15652 46452 15662
rect 46396 15314 46452 15596
rect 46396 15262 46398 15314
rect 46450 15262 46452 15314
rect 46396 15250 46452 15262
rect 46508 15538 46564 15550
rect 46508 15486 46510 15538
rect 46562 15486 46564 15538
rect 46508 11284 46564 15486
rect 46732 13636 46788 16830
rect 46844 14418 46900 20526
rect 47068 19796 47124 19806
rect 47124 19740 47236 19796
rect 47068 19730 47124 19740
rect 46956 19236 47012 19246
rect 47012 19180 47124 19236
rect 46956 19170 47012 19180
rect 46956 17668 47012 17678
rect 46956 17574 47012 17612
rect 47068 17554 47124 19180
rect 47180 19234 47236 19740
rect 47180 19182 47182 19234
rect 47234 19182 47236 19234
rect 47180 18900 47236 19182
rect 47180 18834 47236 18844
rect 47068 17502 47070 17554
rect 47122 17502 47124 17554
rect 47068 17490 47124 17502
rect 47180 18226 47236 18238
rect 47180 18174 47182 18226
rect 47234 18174 47236 18226
rect 47068 16884 47124 16894
rect 47068 14644 47124 16828
rect 47180 16772 47236 18174
rect 47180 16706 47236 16716
rect 47292 16548 47348 22876
rect 47404 22866 47460 22876
rect 47628 22932 47684 23100
rect 47852 23090 47908 23100
rect 47628 22866 47684 22876
rect 47964 22930 48020 22942
rect 47964 22878 47966 22930
rect 48018 22878 48020 22930
rect 47964 22708 48020 22878
rect 47964 22642 48020 22652
rect 47628 22596 47684 22606
rect 47628 21924 47684 22540
rect 47516 21868 47684 21924
rect 47740 22428 48132 22484
rect 47740 22146 47796 22428
rect 48076 22370 48132 22428
rect 48076 22318 48078 22370
rect 48130 22318 48132 22370
rect 48076 22306 48132 22318
rect 47740 22094 47742 22146
rect 47794 22094 47796 22146
rect 47404 21700 47460 21710
rect 47404 21606 47460 21644
rect 47404 20244 47460 20254
rect 47404 20130 47460 20188
rect 47404 20078 47406 20130
rect 47458 20078 47460 20130
rect 47404 20066 47460 20078
rect 47404 19908 47460 19918
rect 47404 16994 47460 19852
rect 47404 16942 47406 16994
rect 47458 16942 47460 16994
rect 47404 16930 47460 16942
rect 47180 16492 47348 16548
rect 47180 15314 47236 16492
rect 47292 16098 47348 16110
rect 47292 16046 47294 16098
rect 47346 16046 47348 16098
rect 47292 15428 47348 16046
rect 47292 15362 47348 15372
rect 47180 15262 47182 15314
rect 47234 15262 47236 15314
rect 47180 15250 47236 15262
rect 47068 14578 47124 14588
rect 47516 14530 47572 21868
rect 47628 21700 47684 21710
rect 47628 21606 47684 21644
rect 47628 20804 47684 20842
rect 47628 20738 47684 20748
rect 47628 20578 47684 20590
rect 47628 20526 47630 20578
rect 47682 20526 47684 20578
rect 47628 15428 47684 20526
rect 47740 19012 47796 22094
rect 48076 22148 48132 22158
rect 48076 21810 48132 22092
rect 48076 21758 48078 21810
rect 48130 21758 48132 21810
rect 48076 21746 48132 21758
rect 48188 21812 48244 21822
rect 48188 21698 48244 21756
rect 48188 21646 48190 21698
rect 48242 21646 48244 21698
rect 48188 21634 48244 21646
rect 47852 21588 47908 21598
rect 47852 21586 48020 21588
rect 47852 21534 47854 21586
rect 47906 21534 48020 21586
rect 47852 21532 48020 21534
rect 47852 21522 47908 21532
rect 47852 20804 47908 20814
rect 47852 19908 47908 20748
rect 47964 20244 48020 21532
rect 48188 21028 48244 21038
rect 48188 20580 48244 20972
rect 48076 20244 48132 20254
rect 47964 20242 48132 20244
rect 47964 20190 48078 20242
rect 48130 20190 48132 20242
rect 47964 20188 48132 20190
rect 48076 20178 48132 20188
rect 48188 20130 48244 20524
rect 48188 20078 48190 20130
rect 48242 20078 48244 20130
rect 48188 20066 48244 20078
rect 48076 20020 48132 20030
rect 48076 19908 48132 19964
rect 47852 19852 48244 19908
rect 47740 18956 48020 19012
rect 47852 18450 47908 18462
rect 47852 18398 47854 18450
rect 47906 18398 47908 18450
rect 47740 18004 47796 18014
rect 47740 17778 47796 17948
rect 47740 17726 47742 17778
rect 47794 17726 47796 17778
rect 47740 17714 47796 17726
rect 47740 16772 47796 16782
rect 47740 15986 47796 16716
rect 47740 15934 47742 15986
rect 47794 15934 47796 15986
rect 47740 15652 47796 15934
rect 47852 15764 47908 18398
rect 47964 16660 48020 18956
rect 48076 17106 48132 17118
rect 48076 17054 48078 17106
rect 48130 17054 48132 17106
rect 48076 16884 48132 17054
rect 48076 16818 48132 16828
rect 48188 16882 48244 19852
rect 48300 18788 48356 23436
rect 48412 21028 48468 75852
rect 48524 75794 48580 76636
rect 48524 75742 48526 75794
rect 48578 75742 48580 75794
rect 48524 75730 48580 75742
rect 48860 76354 48916 76366
rect 48860 76302 48862 76354
rect 48914 76302 48916 76354
rect 48860 38668 48916 76302
rect 49084 75796 49140 75806
rect 49196 75796 49252 76636
rect 49084 75794 49252 75796
rect 49084 75742 49086 75794
rect 49138 75742 49252 75794
rect 49084 75740 49252 75742
rect 49532 75796 49588 79200
rect 50092 77026 50148 77038
rect 50092 76974 50094 77026
rect 50146 76974 50148 77026
rect 50092 76690 50148 76974
rect 50092 76638 50094 76690
rect 50146 76638 50148 76690
rect 49756 76356 49812 76366
rect 49756 76354 49924 76356
rect 49756 76302 49758 76354
rect 49810 76302 49924 76354
rect 49756 76300 49924 76302
rect 49756 76290 49812 76300
rect 49532 75794 49812 75796
rect 49532 75742 49534 75794
rect 49586 75742 49812 75794
rect 49532 75740 49812 75742
rect 49084 75730 49140 75740
rect 49532 75730 49588 75740
rect 49756 75682 49812 75740
rect 49756 75630 49758 75682
rect 49810 75630 49812 75682
rect 49756 75618 49812 75630
rect 49868 55468 49924 76300
rect 50092 75796 50148 76638
rect 50204 76692 50260 79200
rect 50876 77138 50932 79200
rect 50876 77086 50878 77138
rect 50930 77086 50932 77138
rect 50876 77074 50932 77086
rect 51548 77026 51604 79200
rect 51548 76974 51550 77026
rect 51602 76974 51604 77026
rect 51548 76962 51604 76974
rect 51772 77138 51828 77150
rect 51772 77086 51774 77138
rect 51826 77086 51828 77138
rect 50556 76860 50820 76870
rect 50612 76804 50660 76860
rect 50716 76804 50764 76860
rect 50556 76794 50820 76804
rect 50204 76626 50260 76636
rect 51212 76692 51268 76702
rect 50540 76354 50596 76366
rect 50540 76302 50542 76354
rect 50594 76302 50596 76354
rect 50092 75730 50148 75740
rect 50204 75794 50260 75806
rect 50204 75742 50206 75794
rect 50258 75742 50260 75794
rect 48748 38612 48916 38668
rect 49756 55412 49924 55468
rect 48748 35308 48804 38612
rect 48636 35252 48804 35308
rect 48636 26740 48692 35252
rect 49756 29428 49812 55412
rect 50204 43708 50260 75742
rect 50540 75684 50596 76302
rect 50764 75796 50820 75806
rect 50764 75702 50820 75740
rect 51212 75794 51268 76636
rect 51212 75742 51214 75794
rect 51266 75742 51268 75794
rect 51212 75730 51268 75742
rect 51660 76354 51716 76366
rect 51660 76302 51662 76354
rect 51714 76302 51716 76354
rect 50540 75618 50596 75628
rect 50556 75292 50820 75302
rect 50612 75236 50660 75292
rect 50716 75236 50764 75292
rect 50556 75226 50820 75236
rect 50556 73724 50820 73734
rect 50612 73668 50660 73724
rect 50716 73668 50764 73724
rect 50556 73658 50820 73668
rect 50556 72156 50820 72166
rect 50612 72100 50660 72156
rect 50716 72100 50764 72156
rect 50556 72090 50820 72100
rect 50556 70588 50820 70598
rect 50612 70532 50660 70588
rect 50716 70532 50764 70588
rect 50556 70522 50820 70532
rect 50556 69020 50820 69030
rect 50612 68964 50660 69020
rect 50716 68964 50764 69020
rect 50556 68954 50820 68964
rect 50556 67452 50820 67462
rect 50612 67396 50660 67452
rect 50716 67396 50764 67452
rect 50556 67386 50820 67396
rect 50556 65884 50820 65894
rect 50612 65828 50660 65884
rect 50716 65828 50764 65884
rect 50556 65818 50820 65828
rect 50556 64316 50820 64326
rect 50612 64260 50660 64316
rect 50716 64260 50764 64316
rect 50556 64250 50820 64260
rect 50556 62748 50820 62758
rect 50612 62692 50660 62748
rect 50716 62692 50764 62748
rect 50556 62682 50820 62692
rect 50556 61180 50820 61190
rect 50612 61124 50660 61180
rect 50716 61124 50764 61180
rect 50556 61114 50820 61124
rect 50556 59612 50820 59622
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50556 59546 50820 59556
rect 50556 58044 50820 58054
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50556 57978 50820 57988
rect 50556 56476 50820 56486
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50556 56410 50820 56420
rect 51660 55468 51716 76302
rect 51772 75794 51828 77086
rect 52108 77138 52164 77150
rect 52108 77086 52110 77138
rect 52162 77086 52164 77138
rect 52108 76690 52164 77086
rect 52108 76638 52110 76690
rect 52162 76638 52164 76690
rect 52108 76626 52164 76638
rect 51772 75742 51774 75794
rect 51826 75742 51828 75794
rect 51772 75730 51828 75742
rect 52220 75796 52276 79200
rect 52892 76692 52948 79200
rect 52892 76626 52948 76636
rect 53004 77026 53060 77038
rect 53004 76974 53006 77026
rect 53058 76974 53060 77026
rect 53004 76690 53060 76974
rect 53004 76638 53006 76690
rect 53058 76638 53060 76690
rect 52668 76356 52724 76366
rect 52668 76354 52948 76356
rect 52668 76302 52670 76354
rect 52722 76302 52948 76354
rect 52668 76300 52948 76302
rect 52668 76290 52724 76300
rect 52220 75794 52724 75796
rect 52220 75742 52222 75794
rect 52274 75742 52724 75794
rect 52220 75740 52724 75742
rect 52220 75730 52276 75740
rect 52668 75682 52724 75740
rect 52668 75630 52670 75682
rect 52722 75630 52724 75682
rect 52668 75618 52724 75630
rect 52780 75124 52836 75134
rect 52780 75030 52836 75068
rect 52892 73892 52948 76300
rect 53004 75124 53060 76638
rect 53564 76580 53620 79200
rect 53900 76692 53956 76702
rect 53900 76598 53956 76636
rect 54236 76580 54292 79200
rect 53564 76524 53844 76580
rect 54236 76524 54740 76580
rect 53452 76356 53508 76366
rect 53004 75058 53060 75068
rect 53116 76354 53508 76356
rect 53116 76302 53454 76354
rect 53506 76302 53508 76354
rect 53116 76300 53508 76302
rect 52892 73826 52948 73836
rect 53116 68292 53172 76300
rect 53452 76290 53508 76300
rect 53228 75684 53284 75694
rect 53788 75684 53844 76524
rect 54348 76354 54404 76366
rect 54348 76302 54350 76354
rect 54402 76302 54404 76354
rect 54236 75796 54292 75806
rect 53228 75682 53508 75684
rect 53228 75630 53230 75682
rect 53282 75630 53508 75682
rect 53228 75628 53508 75630
rect 53228 75618 53284 75628
rect 51100 55412 51716 55468
rect 52668 68236 53172 68292
rect 53340 73892 53396 73902
rect 50556 54908 50820 54918
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50556 54842 50820 54852
rect 50556 53340 50820 53350
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50556 53274 50820 53284
rect 50556 51772 50820 51782
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50556 51706 50820 51716
rect 50556 50204 50820 50214
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50556 50138 50820 50148
rect 50556 48636 50820 48646
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50556 48570 50820 48580
rect 50556 47068 50820 47078
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50556 47002 50820 47012
rect 50556 45500 50820 45510
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50556 45434 50820 45444
rect 50556 43932 50820 43942
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50556 43866 50820 43876
rect 50204 43652 50372 43708
rect 49756 29362 49812 29372
rect 50092 30548 50148 30558
rect 49196 28644 49252 28654
rect 48972 27300 49028 27310
rect 48972 27074 49028 27244
rect 48972 27022 48974 27074
rect 49026 27022 49028 27074
rect 48972 27010 49028 27022
rect 49084 27188 49140 27198
rect 49084 26962 49140 27132
rect 49084 26910 49086 26962
rect 49138 26910 49140 26962
rect 49084 26898 49140 26910
rect 49196 26740 49252 28588
rect 49644 27300 49700 27310
rect 49420 27298 49700 27300
rect 49420 27246 49646 27298
rect 49698 27246 49700 27298
rect 49420 27244 49700 27246
rect 48636 26684 49028 26740
rect 48860 26516 48916 26554
rect 48860 26450 48916 26460
rect 48748 26292 48804 26302
rect 48748 26198 48804 26236
rect 48860 26068 48916 26078
rect 48748 26066 48916 26068
rect 48748 26014 48862 26066
rect 48914 26014 48916 26066
rect 48748 26012 48916 26014
rect 48524 23940 48580 23950
rect 48524 23846 48580 23884
rect 48636 22372 48692 22382
rect 48636 22278 48692 22316
rect 48412 20802 48468 20972
rect 48412 20750 48414 20802
rect 48466 20750 48468 20802
rect 48412 20738 48468 20750
rect 48524 20690 48580 20702
rect 48524 20638 48526 20690
rect 48578 20638 48580 20690
rect 48524 20132 48580 20638
rect 48748 20356 48804 26012
rect 48860 26002 48916 26012
rect 48972 25844 49028 26684
rect 48860 25788 49028 25844
rect 49084 26684 49252 26740
rect 49308 26850 49364 26862
rect 49308 26798 49310 26850
rect 49362 26798 49364 26850
rect 48860 22596 48916 25788
rect 48972 24388 49028 24398
rect 48972 23716 49028 24332
rect 48972 23622 49028 23660
rect 48972 23380 49028 23390
rect 49084 23380 49140 26684
rect 49308 26516 49364 26798
rect 49420 26628 49476 27244
rect 49644 27234 49700 27244
rect 49532 27076 49588 27086
rect 49532 26982 49588 27020
rect 49644 26964 49700 27002
rect 49644 26898 49700 26908
rect 49420 26572 49588 26628
rect 49028 23324 49140 23380
rect 49196 26460 49364 26516
rect 48972 23286 49028 23324
rect 48860 21140 48916 22540
rect 48860 21074 48916 21084
rect 48972 22372 49028 22382
rect 48972 21586 49028 22316
rect 48972 21534 48974 21586
rect 49026 21534 49028 21586
rect 48972 20804 49028 21534
rect 48972 20738 49028 20748
rect 49084 22146 49140 22158
rect 49084 22094 49086 22146
rect 49138 22094 49140 22146
rect 48524 19908 48580 20076
rect 48524 19842 48580 19852
rect 48636 20300 48804 20356
rect 48972 20578 49028 20590
rect 48972 20526 48974 20578
rect 49026 20526 49028 20578
rect 48972 20356 49028 20526
rect 48524 19348 48580 19358
rect 48524 19254 48580 19292
rect 48300 18722 48356 18732
rect 48524 18900 48580 18910
rect 48524 17778 48580 18844
rect 48636 18340 48692 20300
rect 48972 20290 49028 20300
rect 48748 20020 48804 20030
rect 48748 19926 48804 19964
rect 49084 19684 49140 22094
rect 49196 22148 49252 26460
rect 49420 26404 49476 26414
rect 49420 26310 49476 26348
rect 49308 26290 49364 26302
rect 49308 26238 49310 26290
rect 49362 26238 49364 26290
rect 49308 26068 49364 26238
rect 49308 26002 49364 26012
rect 49532 25172 49588 26572
rect 50092 26516 50148 30492
rect 50204 27188 50260 27198
rect 50204 27094 50260 27132
rect 50092 26422 50148 26460
rect 49644 26292 49700 26302
rect 49644 26198 49700 26236
rect 49980 26292 50036 26302
rect 49756 26180 49812 26190
rect 49532 25116 49700 25172
rect 49532 23714 49588 23726
rect 49532 23662 49534 23714
rect 49586 23662 49588 23714
rect 49420 23268 49476 23278
rect 49420 22932 49476 23212
rect 49420 22866 49476 22876
rect 49420 22372 49476 22382
rect 49532 22372 49588 23662
rect 49644 22820 49700 25116
rect 49756 23380 49812 26124
rect 49756 23314 49812 23324
rect 49756 23042 49812 23054
rect 49756 22990 49758 23042
rect 49810 22990 49812 23042
rect 49756 22932 49812 22990
rect 49868 22932 49924 22942
rect 49756 22930 49924 22932
rect 49756 22878 49870 22930
rect 49922 22878 49924 22930
rect 49756 22876 49924 22878
rect 49868 22866 49924 22876
rect 49644 22764 49812 22820
rect 49476 22316 49588 22372
rect 49420 22306 49476 22316
rect 49196 22092 49700 22148
rect 49532 21588 49588 21598
rect 49532 21494 49588 21532
rect 49196 21474 49252 21486
rect 49196 21422 49198 21474
rect 49250 21422 49252 21474
rect 49196 19796 49252 21422
rect 49532 21140 49588 21150
rect 49532 20802 49588 21084
rect 49532 20750 49534 20802
rect 49586 20750 49588 20802
rect 49532 20738 49588 20750
rect 49420 20132 49476 20142
rect 49420 20038 49476 20076
rect 49308 20020 49364 20030
rect 49308 19926 49364 19964
rect 49532 19906 49588 19918
rect 49532 19854 49534 19906
rect 49586 19854 49588 19906
rect 49196 19740 49476 19796
rect 49084 19628 49252 19684
rect 48972 19236 49028 19246
rect 48860 19180 48972 19236
rect 48860 18562 48916 19180
rect 48972 19170 49028 19180
rect 48860 18510 48862 18562
rect 48914 18510 48916 18562
rect 48860 18498 48916 18510
rect 48972 18788 49028 18798
rect 48748 18340 48804 18350
rect 48636 18284 48748 18340
rect 48748 18274 48804 18284
rect 48524 17726 48526 17778
rect 48578 17726 48580 17778
rect 48524 17714 48580 17726
rect 48188 16830 48190 16882
rect 48242 16830 48244 16882
rect 48188 16818 48244 16830
rect 48748 16884 48804 16894
rect 48748 16660 48804 16828
rect 47964 16604 48132 16660
rect 48748 16604 48916 16660
rect 47852 15698 47908 15708
rect 47964 15874 48020 15886
rect 47964 15822 47966 15874
rect 48018 15822 48020 15874
rect 47740 15586 47796 15596
rect 47740 15428 47796 15438
rect 47628 15426 47796 15428
rect 47628 15374 47742 15426
rect 47794 15374 47796 15426
rect 47628 15372 47796 15374
rect 47740 15362 47796 15372
rect 47516 14478 47518 14530
rect 47570 14478 47572 14530
rect 47516 14466 47572 14478
rect 46844 14366 46846 14418
rect 46898 14366 46900 14418
rect 46844 14354 46900 14366
rect 46956 13636 47012 13646
rect 46732 13634 47012 13636
rect 46732 13582 46958 13634
rect 47010 13582 47012 13634
rect 46732 13580 47012 13582
rect 46956 13524 47012 13580
rect 46956 13458 47012 13468
rect 46508 11218 46564 11228
rect 45948 8036 46004 8046
rect 45948 7942 46004 7980
rect 46172 7362 46228 8204
rect 47292 10948 47348 10958
rect 46732 7812 46788 7822
rect 46172 7310 46174 7362
rect 46226 7310 46228 7362
rect 46172 7298 46228 7310
rect 46508 7474 46564 7486
rect 46508 7422 46510 7474
rect 46562 7422 46564 7474
rect 46508 7364 46564 7422
rect 46508 7298 46564 7308
rect 46620 6690 46676 6702
rect 46620 6638 46622 6690
rect 46674 6638 46676 6690
rect 46060 6578 46116 6590
rect 46060 6526 46062 6578
rect 46114 6526 46116 6578
rect 46060 6132 46116 6526
rect 46060 6066 46116 6076
rect 46396 5906 46452 5918
rect 46396 5854 46398 5906
rect 46450 5854 46452 5906
rect 45836 4846 45838 4898
rect 45890 4846 45892 4898
rect 45836 4834 45892 4846
rect 45948 5348 46004 5358
rect 45724 3614 45726 3666
rect 45778 3614 45780 3666
rect 45724 3602 45780 3614
rect 45276 3556 45332 3566
rect 45276 3462 45332 3500
rect 45388 3444 45444 3482
rect 45388 3378 45444 3388
rect 45164 3276 45332 3332
rect 45276 800 45332 3276
rect 45948 800 46004 5292
rect 46396 5124 46452 5854
rect 46284 5068 46396 5124
rect 46284 4338 46340 5068
rect 46396 5058 46452 5068
rect 46620 4900 46676 6638
rect 46732 6130 46788 7756
rect 47068 7364 47124 7374
rect 47068 7270 47124 7308
rect 47068 6692 47124 6702
rect 47068 6690 47236 6692
rect 47068 6638 47070 6690
rect 47122 6638 47236 6690
rect 47068 6636 47236 6638
rect 47068 6626 47124 6636
rect 46732 6078 46734 6130
rect 46786 6078 46788 6130
rect 46732 6066 46788 6078
rect 47068 6466 47124 6478
rect 47068 6414 47070 6466
rect 47122 6414 47124 6466
rect 47068 5908 47124 6414
rect 46956 5906 47124 5908
rect 46956 5854 47070 5906
rect 47122 5854 47124 5906
rect 46956 5852 47124 5854
rect 46844 5124 46900 5134
rect 46844 5030 46900 5068
rect 46620 4834 46676 4844
rect 46620 4564 46676 4574
rect 46620 4450 46676 4508
rect 46620 4398 46622 4450
rect 46674 4398 46676 4450
rect 46620 4386 46676 4398
rect 46956 4450 47012 5852
rect 47068 5842 47124 5852
rect 47180 4564 47236 6636
rect 47292 6468 47348 10892
rect 47964 9604 48020 15822
rect 48076 15876 48132 16604
rect 48076 15810 48132 15820
rect 48188 15652 48244 15662
rect 48188 14530 48244 15596
rect 48860 15426 48916 16604
rect 48972 16098 49028 18732
rect 49084 18340 49140 18350
rect 49084 16882 49140 18284
rect 49196 17554 49252 19628
rect 49308 19236 49364 19246
rect 49308 19122 49364 19180
rect 49308 19070 49310 19122
rect 49362 19070 49364 19122
rect 49308 19058 49364 19070
rect 49196 17502 49198 17554
rect 49250 17502 49252 17554
rect 49196 17490 49252 17502
rect 49308 17444 49364 17454
rect 49308 17220 49364 17388
rect 49084 16830 49086 16882
rect 49138 16830 49140 16882
rect 49084 16818 49140 16830
rect 49196 17164 49364 17220
rect 48972 16046 48974 16098
rect 49026 16046 49028 16098
rect 48972 16034 49028 16046
rect 48860 15374 48862 15426
rect 48914 15374 48916 15426
rect 48860 15362 48916 15374
rect 48972 15316 49028 15326
rect 48972 15222 49028 15260
rect 49196 15148 49252 17164
rect 49308 16996 49364 17006
rect 49420 16996 49476 19740
rect 49308 16994 49476 16996
rect 49308 16942 49310 16994
rect 49362 16942 49476 16994
rect 49308 16940 49476 16942
rect 49308 16930 49364 16940
rect 49532 15986 49588 19854
rect 49644 17666 49700 22092
rect 49756 19234 49812 22764
rect 49868 22258 49924 22270
rect 49868 22206 49870 22258
rect 49922 22206 49924 22258
rect 49868 21700 49924 22206
rect 49980 21812 50036 26236
rect 50316 23380 50372 43652
rect 50556 42364 50820 42374
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50556 42298 50820 42308
rect 50556 40796 50820 40806
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50556 40730 50820 40740
rect 50556 39228 50820 39238
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50556 39162 50820 39172
rect 50556 37660 50820 37670
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50556 37594 50820 37604
rect 50556 36092 50820 36102
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50556 36026 50820 36036
rect 50556 34524 50820 34534
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50556 34458 50820 34468
rect 50556 32956 50820 32966
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50556 32890 50820 32900
rect 50556 31388 50820 31398
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50556 31322 50820 31332
rect 50540 30772 50596 30782
rect 50428 30716 50540 30772
rect 50428 26516 50484 30716
rect 50540 30706 50596 30716
rect 50876 30212 50932 30222
rect 50876 30118 50932 30156
rect 50556 29820 50820 29830
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50556 29754 50820 29764
rect 50556 28252 50820 28262
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50556 28186 50820 28196
rect 50876 27412 50932 27422
rect 50932 27356 51044 27412
rect 50876 27346 50932 27356
rect 50652 26964 50708 26974
rect 50652 26870 50708 26908
rect 50556 26684 50820 26694
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50556 26618 50820 26628
rect 50540 26516 50596 26526
rect 50484 26514 50596 26516
rect 50484 26462 50542 26514
rect 50594 26462 50596 26514
rect 50484 26460 50596 26462
rect 50428 26422 50484 26460
rect 50540 26450 50596 26460
rect 50556 25116 50820 25126
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50556 25050 50820 25060
rect 50556 23548 50820 23558
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50556 23482 50820 23492
rect 50988 23492 51044 27356
rect 50988 23426 51044 23436
rect 50092 23378 50372 23380
rect 50092 23326 50318 23378
rect 50370 23326 50372 23378
rect 50092 23324 50372 23326
rect 50092 22370 50148 23324
rect 50316 23314 50372 23324
rect 50764 23380 50820 23390
rect 50764 23286 50820 23324
rect 50092 22318 50094 22370
rect 50146 22318 50148 22370
rect 50092 22306 50148 22318
rect 50204 22930 50260 22942
rect 50204 22878 50206 22930
rect 50258 22878 50260 22930
rect 50204 21812 50260 22878
rect 50876 22370 50932 22382
rect 50876 22318 50878 22370
rect 50930 22318 50932 22370
rect 50556 21980 50820 21990
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50556 21914 50820 21924
rect 49980 21756 50148 21812
rect 49868 21698 50036 21700
rect 49868 21646 49870 21698
rect 49922 21646 50036 21698
rect 49868 21644 50036 21646
rect 49868 21634 49924 21644
rect 49980 20692 50036 21644
rect 49980 20598 50036 20636
rect 49756 19182 49758 19234
rect 49810 19182 49812 19234
rect 49756 19170 49812 19182
rect 49980 19012 50036 19022
rect 49644 17614 49646 17666
rect 49698 17614 49700 17666
rect 49644 17602 49700 17614
rect 49756 19010 50036 19012
rect 49756 18958 49982 19010
rect 50034 18958 50036 19010
rect 49756 18956 50036 18958
rect 49532 15934 49534 15986
rect 49586 15934 49588 15986
rect 49532 15922 49588 15934
rect 48188 14478 48190 14530
rect 48242 14478 48244 14530
rect 48188 14466 48244 14478
rect 48300 15092 48356 15102
rect 48300 13970 48356 15036
rect 48972 15092 49252 15148
rect 48748 14532 48804 14542
rect 48748 14438 48804 14476
rect 48300 13918 48302 13970
rect 48354 13918 48356 13970
rect 48300 13906 48356 13918
rect 48412 14306 48468 14318
rect 48412 14254 48414 14306
rect 48466 14254 48468 14306
rect 47964 9538 48020 9548
rect 48412 9156 48468 14254
rect 48972 13970 49028 15092
rect 48972 13918 48974 13970
rect 49026 13918 49028 13970
rect 48972 13906 49028 13918
rect 49420 14868 49476 14878
rect 49420 14196 49476 14812
rect 49420 13970 49476 14140
rect 49420 13918 49422 13970
rect 49474 13918 49476 13970
rect 49420 13906 49476 13918
rect 48412 9090 48468 9100
rect 48860 11844 48916 11854
rect 47292 6402 47348 6412
rect 47628 7362 47684 7374
rect 47628 7310 47630 7362
rect 47682 7310 47684 7362
rect 47516 5908 47572 5918
rect 47180 4498 47236 4508
rect 47292 5794 47348 5806
rect 47292 5742 47294 5794
rect 47346 5742 47348 5794
rect 46956 4398 46958 4450
rect 47010 4398 47012 4450
rect 46956 4386 47012 4398
rect 46284 4286 46286 4338
rect 46338 4286 46340 4338
rect 46284 4274 46340 4286
rect 47292 4340 47348 5742
rect 47404 5010 47460 5022
rect 47404 4958 47406 5010
rect 47458 4958 47460 5010
rect 47404 4676 47460 4958
rect 47404 4610 47460 4620
rect 47292 4338 47460 4340
rect 47292 4286 47294 4338
rect 47346 4286 47460 4338
rect 47292 4284 47460 4286
rect 47292 4274 47348 4284
rect 46620 4228 46676 4238
rect 46620 800 46676 4172
rect 47404 3666 47460 4284
rect 47404 3614 47406 3666
rect 47458 3614 47460 3666
rect 47404 3602 47460 3614
rect 47516 3388 47572 5852
rect 47628 5906 47684 7310
rect 48636 6578 48692 6590
rect 48636 6526 48638 6578
rect 48690 6526 48692 6578
rect 47964 6132 48020 6142
rect 47964 6038 48020 6076
rect 48636 6132 48692 6526
rect 48636 6066 48692 6076
rect 47628 5854 47630 5906
rect 47682 5854 47684 5906
rect 47628 5572 47684 5854
rect 47628 5506 47684 5516
rect 48748 6018 48804 6030
rect 48748 5966 48750 6018
rect 48802 5966 48804 6018
rect 48076 5460 48132 5470
rect 47964 5236 48020 5246
rect 47964 3554 48020 5180
rect 47964 3502 47966 3554
rect 48018 3502 48020 3554
rect 47964 3490 48020 3502
rect 47292 3332 47572 3388
rect 48076 3332 48132 5404
rect 48748 5236 48804 5966
rect 48860 6020 48916 11788
rect 49532 8036 49588 8046
rect 48860 5954 48916 5964
rect 49084 6466 49140 6478
rect 49084 6414 49086 6466
rect 49138 6414 49140 6466
rect 48748 5170 48804 5180
rect 49084 5906 49140 6414
rect 49084 5854 49086 5906
rect 49138 5854 49140 5906
rect 48188 5124 48244 5134
rect 48188 3554 48244 5068
rect 48972 5124 49028 5134
rect 48972 5010 49028 5068
rect 48972 4958 48974 5010
rect 49026 4958 49028 5010
rect 48972 4946 49028 4958
rect 49084 4788 49140 5854
rect 49196 5348 49252 5358
rect 49196 5122 49252 5292
rect 49196 5070 49198 5122
rect 49250 5070 49252 5122
rect 49196 5058 49252 5070
rect 48972 4732 49140 4788
rect 48748 4564 48804 4574
rect 48748 4470 48804 4508
rect 48188 3502 48190 3554
rect 48242 3502 48244 3554
rect 48188 3490 48244 3502
rect 48524 4340 48580 4350
rect 48524 3442 48580 4284
rect 48972 4228 49028 4732
rect 48972 4162 49028 4172
rect 49084 4340 49140 4350
rect 48860 4116 48916 4126
rect 48748 3892 48804 3902
rect 48748 3554 48804 3836
rect 48748 3502 48750 3554
rect 48802 3502 48804 3554
rect 48748 3490 48804 3502
rect 48524 3390 48526 3442
rect 48578 3390 48580 3442
rect 48524 3378 48580 3390
rect 48860 3444 48916 4060
rect 48972 4004 49028 4014
rect 49084 4004 49140 4284
rect 49532 4338 49588 7980
rect 49756 8036 49812 18956
rect 49980 18946 50036 18956
rect 49868 18674 49924 18686
rect 49868 18622 49870 18674
rect 49922 18622 49924 18674
rect 49868 13412 49924 18622
rect 49980 18452 50036 18462
rect 50092 18452 50148 21756
rect 50204 21746 50260 21756
rect 50876 21700 50932 22318
rect 50764 21644 50932 21700
rect 50204 21586 50260 21598
rect 50204 21534 50206 21586
rect 50258 21534 50260 21586
rect 50204 21364 50260 21534
rect 50204 21298 50260 21308
rect 50652 21474 50708 21486
rect 50652 21422 50654 21474
rect 50706 21422 50708 21474
rect 50316 20804 50372 20814
rect 50316 20710 50372 20748
rect 50652 20692 50708 21422
rect 50764 21364 50820 21644
rect 50764 21298 50820 21308
rect 51100 21140 51156 55412
rect 51660 38836 51716 38846
rect 51324 38724 51380 38734
rect 51212 30100 51268 30110
rect 51212 30006 51268 30044
rect 51324 26908 51380 38668
rect 51436 31780 51492 31790
rect 51436 31686 51492 31724
rect 51548 31668 51604 31678
rect 51548 31574 51604 31612
rect 51436 30994 51492 31006
rect 51436 30942 51438 30994
rect 51490 30942 51492 30994
rect 51436 30884 51492 30942
rect 51436 30818 51492 30828
rect 50652 20626 50708 20636
rect 50876 21084 51156 21140
rect 51212 26852 51380 26908
rect 51436 29986 51492 29998
rect 51436 29934 51438 29986
rect 51490 29934 51492 29986
rect 50428 20578 50484 20590
rect 50428 20526 50430 20578
rect 50482 20526 50484 20578
rect 50316 19906 50372 19918
rect 50316 19854 50318 19906
rect 50370 19854 50372 19906
rect 50204 19572 50260 19582
rect 50316 19572 50372 19854
rect 50260 19516 50372 19572
rect 50204 19506 50260 19516
rect 50428 19236 50484 20526
rect 50556 20412 50820 20422
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50556 20346 50820 20356
rect 50876 20018 50932 21084
rect 50988 20692 51044 20702
rect 50988 20598 51044 20636
rect 51100 20132 51156 20142
rect 51100 20038 51156 20076
rect 50876 19966 50878 20018
rect 50930 19966 50932 20018
rect 50876 19908 50932 19966
rect 50876 19842 50932 19852
rect 50428 19170 50484 19180
rect 50988 19234 51044 19246
rect 50988 19182 50990 19234
rect 51042 19182 51044 19234
rect 50556 18844 50820 18854
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50556 18778 50820 18788
rect 50988 18564 51044 19182
rect 50988 18498 51044 18508
rect 51100 19122 51156 19134
rect 51100 19070 51102 19122
rect 51154 19070 51156 19122
rect 51100 18562 51156 19070
rect 51100 18510 51102 18562
rect 51154 18510 51156 18562
rect 49980 18450 50148 18452
rect 49980 18398 49982 18450
rect 50034 18398 50148 18450
rect 49980 18396 50148 18398
rect 50876 18450 50932 18462
rect 50876 18398 50878 18450
rect 50930 18398 50932 18450
rect 49980 18386 50036 18396
rect 50876 17444 50932 18398
rect 50876 17378 50932 17388
rect 51100 17554 51156 18510
rect 51100 17502 51102 17554
rect 51154 17502 51156 17554
rect 50556 17276 50820 17286
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50556 17210 50820 17220
rect 49868 13346 49924 13356
rect 49980 17106 50036 17118
rect 49980 17054 49982 17106
rect 50034 17054 50036 17106
rect 49756 7970 49812 7980
rect 49980 7588 50036 17054
rect 50988 17108 51044 17118
rect 50988 16882 51044 17052
rect 50988 16830 50990 16882
rect 51042 16830 51044 16882
rect 50428 16098 50484 16110
rect 50428 16046 50430 16098
rect 50482 16046 50484 16098
rect 50316 15764 50372 15774
rect 50428 15764 50484 16046
rect 50372 15708 50484 15764
rect 50316 15698 50372 15708
rect 50092 14644 50148 14654
rect 50092 14550 50148 14588
rect 50316 14644 50372 14654
rect 50316 14084 50372 14588
rect 50428 14532 50484 15708
rect 50556 15708 50820 15718
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50556 15642 50820 15652
rect 50988 15540 51044 16830
rect 51100 16994 51156 17502
rect 51100 16942 51102 16994
rect 51154 16942 51156 16994
rect 51100 16322 51156 16942
rect 51100 16270 51102 16322
rect 51154 16270 51156 16322
rect 51100 16258 51156 16270
rect 50764 15484 51044 15540
rect 50652 15428 50708 15438
rect 50652 15334 50708 15372
rect 50764 15148 50820 15484
rect 50652 15092 50820 15148
rect 50876 15314 50932 15326
rect 50876 15262 50878 15314
rect 50930 15262 50932 15314
rect 50876 15092 50932 15262
rect 50652 14642 50708 15092
rect 50876 15026 50932 15036
rect 50652 14590 50654 14642
rect 50706 14590 50708 14642
rect 50652 14578 50708 14590
rect 51212 14532 51268 26852
rect 51436 22708 51492 29934
rect 51436 22642 51492 22652
rect 51548 23492 51604 23502
rect 51324 22370 51380 22382
rect 51324 22318 51326 22370
rect 51378 22318 51380 22370
rect 51324 21698 51380 22318
rect 51324 21646 51326 21698
rect 51378 21646 51380 21698
rect 51324 20132 51380 21646
rect 51548 21812 51604 23436
rect 51436 20804 51492 20814
rect 51548 20804 51604 21756
rect 51436 20802 51604 20804
rect 51436 20750 51438 20802
rect 51490 20750 51604 20802
rect 51436 20748 51604 20750
rect 51436 20738 51492 20748
rect 51548 20244 51604 20254
rect 51324 20066 51380 20076
rect 51436 20242 51604 20244
rect 51436 20190 51550 20242
rect 51602 20190 51604 20242
rect 51436 20188 51604 20190
rect 51324 17666 51380 17678
rect 51324 17614 51326 17666
rect 51378 17614 51380 17666
rect 51324 14868 51380 17614
rect 51436 16100 51492 20188
rect 51548 20178 51604 20188
rect 51660 19796 51716 38780
rect 52332 34580 52388 34590
rect 51772 31556 51828 31566
rect 51772 31554 51940 31556
rect 51772 31502 51774 31554
rect 51826 31502 51940 31554
rect 51772 31500 51940 31502
rect 51772 31490 51828 31500
rect 51772 31106 51828 31118
rect 51772 31054 51774 31106
rect 51826 31054 51828 31106
rect 51772 30324 51828 31054
rect 51772 30258 51828 30268
rect 51772 22596 51828 22606
rect 51772 22482 51828 22540
rect 51772 22430 51774 22482
rect 51826 22430 51828 22482
rect 51772 22418 51828 22430
rect 51884 21924 51940 31500
rect 51996 30882 52052 30894
rect 51996 30830 51998 30882
rect 52050 30830 52052 30882
rect 51996 30324 52052 30830
rect 52332 30324 52388 34524
rect 52556 32004 52612 32014
rect 52556 31106 52612 31948
rect 52556 31054 52558 31106
rect 52610 31054 52612 31106
rect 52556 31042 52612 31054
rect 52444 30994 52500 31006
rect 52444 30942 52446 30994
rect 52498 30942 52500 30994
rect 52444 30436 52500 30942
rect 52444 30370 52500 30380
rect 51996 30268 52164 30324
rect 51996 30100 52052 30110
rect 51996 30006 52052 30044
rect 51772 21868 51940 21924
rect 51772 20692 51828 21868
rect 51884 21588 51940 21598
rect 51884 21494 51940 21532
rect 51996 21474 52052 21486
rect 51996 21422 51998 21474
rect 52050 21422 52052 21474
rect 51884 21028 51940 21038
rect 51884 20914 51940 20972
rect 51884 20862 51886 20914
rect 51938 20862 51940 20914
rect 51884 20850 51940 20862
rect 51772 20636 51940 20692
rect 51436 16034 51492 16044
rect 51548 19740 51716 19796
rect 51772 20020 51828 20030
rect 51436 15876 51492 15886
rect 51436 15782 51492 15820
rect 51324 14802 51380 14812
rect 50428 14466 50484 14476
rect 51100 14476 51268 14532
rect 51324 14532 51380 14542
rect 50556 14140 50820 14150
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50556 14074 50820 14084
rect 51100 14084 51156 14476
rect 51324 14438 51380 14476
rect 51100 14028 51268 14084
rect 50316 14018 50372 14028
rect 50556 12572 50820 12582
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50556 12506 50820 12516
rect 50556 11004 50820 11014
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50556 10938 50820 10948
rect 50556 9436 50820 9446
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50556 9370 50820 9380
rect 50988 8484 51044 8494
rect 50556 7868 50820 7878
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50556 7802 50820 7812
rect 49980 7522 50036 7532
rect 49980 6692 50036 6702
rect 49644 6468 49700 6478
rect 49644 6466 49812 6468
rect 49644 6414 49646 6466
rect 49698 6414 49812 6466
rect 49644 6412 49812 6414
rect 49644 6402 49700 6412
rect 49644 6132 49700 6142
rect 49644 6038 49700 6076
rect 49756 5908 49812 6412
rect 49980 6132 50036 6636
rect 50988 6690 51044 8428
rect 51212 8428 51268 14028
rect 51324 13748 51380 13758
rect 51324 13654 51380 13692
rect 51548 8428 51604 19740
rect 51772 19236 51828 19964
rect 51772 19170 51828 19180
rect 51772 17554 51828 17566
rect 51772 17502 51774 17554
rect 51826 17502 51828 17554
rect 51772 17444 51828 17502
rect 51772 17378 51828 17388
rect 51884 16884 51940 20636
rect 51996 19796 52052 21422
rect 52108 21140 52164 30268
rect 52332 30258 52388 30268
rect 52668 26908 52724 68236
rect 53340 55468 53396 73836
rect 53228 55412 53396 55468
rect 52780 36036 52836 36046
rect 52780 31778 52836 35980
rect 53004 34132 53060 34142
rect 53004 34038 53060 34076
rect 53116 33906 53172 33918
rect 53116 33854 53118 33906
rect 53170 33854 53172 33906
rect 52780 31726 52782 31778
rect 52834 31726 52836 31778
rect 52780 31668 52836 31726
rect 52780 31602 52836 31612
rect 53004 33796 53060 33806
rect 52892 30884 52948 30894
rect 52892 30790 52948 30828
rect 52892 30324 52948 30334
rect 52892 30230 52948 30268
rect 52668 26852 52948 26908
rect 52780 23492 52836 23502
rect 52556 22708 52612 22718
rect 52444 21586 52500 21598
rect 52444 21534 52446 21586
rect 52498 21534 52500 21586
rect 52108 21084 52276 21140
rect 52108 20020 52164 20030
rect 52108 19926 52164 19964
rect 52108 19796 52164 19806
rect 51996 19740 52108 19796
rect 52108 19730 52164 19740
rect 51884 16818 51940 16828
rect 51996 19236 52052 19246
rect 51996 16210 52052 19180
rect 51996 16158 51998 16210
rect 52050 16158 52052 16210
rect 51996 16146 52052 16158
rect 51996 15316 52052 15326
rect 51660 15204 51716 15242
rect 51660 15138 51716 15148
rect 51996 14306 52052 15260
rect 52220 15204 52276 21084
rect 52332 20242 52388 20254
rect 52332 20190 52334 20242
rect 52386 20190 52388 20242
rect 52332 15426 52388 20190
rect 52444 20020 52500 21534
rect 52444 19954 52500 19964
rect 52444 19796 52500 19806
rect 52556 19796 52612 22652
rect 52780 22484 52836 23436
rect 52668 22482 52836 22484
rect 52668 22430 52782 22482
rect 52834 22430 52836 22482
rect 52668 22428 52836 22430
rect 52668 21588 52724 22428
rect 52780 22418 52836 22428
rect 52668 21522 52724 21532
rect 52780 21586 52836 21598
rect 52780 21534 52782 21586
rect 52834 21534 52836 21586
rect 52780 21364 52836 21534
rect 52780 21298 52836 21308
rect 52780 20580 52836 20590
rect 52780 20486 52836 20524
rect 52892 20020 52948 26852
rect 52892 19926 52948 19964
rect 52556 19740 52948 19796
rect 52444 16994 52500 19740
rect 52668 19236 52724 19246
rect 52668 19142 52724 19180
rect 52556 18338 52612 18350
rect 52556 18286 52558 18338
rect 52610 18286 52612 18338
rect 52556 18228 52612 18286
rect 52556 18162 52612 18172
rect 52444 16942 52446 16994
rect 52498 16942 52500 16994
rect 52444 16930 52500 16942
rect 52780 17444 52836 17454
rect 52668 16884 52724 16894
rect 52668 16790 52724 16828
rect 52668 16100 52724 16110
rect 52668 16006 52724 16044
rect 52332 15374 52334 15426
rect 52386 15374 52388 15426
rect 52332 15362 52388 15374
rect 52556 15316 52612 15326
rect 52444 15314 52612 15316
rect 52444 15262 52558 15314
rect 52610 15262 52612 15314
rect 52444 15260 52612 15262
rect 52444 15204 52500 15260
rect 52556 15250 52612 15260
rect 52220 15148 52500 15204
rect 52668 14532 52724 14542
rect 52668 14438 52724 14476
rect 52780 14420 52836 17388
rect 52892 16098 52948 19740
rect 53004 18450 53060 33740
rect 53004 18398 53006 18450
rect 53058 18398 53060 18450
rect 53004 18386 53060 18398
rect 53116 17668 53172 33854
rect 53228 21364 53284 55412
rect 53340 34244 53396 34254
rect 53340 34150 53396 34188
rect 53452 33572 53508 75628
rect 53564 75682 53844 75684
rect 53564 75630 53790 75682
rect 53842 75630 53844 75682
rect 53564 75628 53844 75630
rect 53564 75122 53620 75628
rect 53788 75618 53844 75628
rect 53900 75794 54292 75796
rect 53900 75742 54238 75794
rect 54290 75742 54292 75794
rect 53900 75740 54292 75742
rect 53564 75070 53566 75122
rect 53618 75070 53620 75122
rect 53564 75058 53620 75070
rect 53788 40852 53844 40862
rect 53788 38724 53844 40796
rect 53788 38658 53844 38668
rect 53788 36148 53844 36158
rect 53564 34916 53620 34954
rect 53564 34850 53620 34860
rect 53564 34690 53620 34702
rect 53564 34638 53566 34690
rect 53618 34638 53620 34690
rect 53564 33796 53620 34638
rect 53788 34244 53844 36092
rect 53788 34178 53844 34188
rect 53564 33730 53620 33740
rect 53452 33516 53844 33572
rect 53676 32788 53732 32798
rect 53676 32004 53732 32732
rect 53676 31218 53732 31948
rect 53676 31166 53678 31218
rect 53730 31166 53732 31218
rect 53676 31154 53732 31166
rect 53340 30884 53396 30894
rect 53396 30828 53508 30884
rect 53340 30818 53396 30828
rect 53452 26908 53508 30828
rect 53452 26852 53732 26908
rect 53340 21588 53396 21598
rect 53340 21494 53396 21532
rect 53228 21308 53396 21364
rect 53228 20132 53284 20142
rect 53228 20038 53284 20076
rect 53340 19234 53396 21308
rect 53564 20802 53620 20814
rect 53564 20750 53566 20802
rect 53618 20750 53620 20802
rect 53564 20356 53620 20750
rect 53340 19182 53342 19234
rect 53394 19182 53396 19234
rect 53228 18564 53284 18574
rect 53228 18470 53284 18508
rect 53340 18340 53396 19182
rect 53452 20132 53508 20142
rect 53452 19122 53508 20076
rect 53564 20018 53620 20300
rect 53564 19966 53566 20018
rect 53618 19966 53620 20018
rect 53564 19954 53620 19966
rect 53676 19796 53732 26852
rect 53788 23492 53844 33516
rect 53788 23426 53844 23436
rect 53788 21812 53844 21822
rect 53788 21718 53844 21756
rect 53900 20804 53956 75740
rect 54236 75730 54292 75740
rect 54348 55468 54404 76302
rect 54684 75684 54740 76524
rect 54908 76468 54964 79200
rect 55580 77812 55636 79200
rect 55580 77756 55860 77812
rect 55132 76692 55188 76702
rect 55132 76598 55188 76636
rect 54908 76412 55636 76468
rect 55132 75796 55188 75806
rect 54460 75682 54740 75684
rect 54460 75630 54686 75682
rect 54738 75630 54740 75682
rect 54460 75628 54740 75630
rect 54460 75122 54516 75628
rect 54684 75618 54740 75628
rect 54908 75794 55188 75796
rect 54908 75742 55134 75794
rect 55186 75742 55188 75794
rect 54908 75740 55188 75742
rect 54460 75070 54462 75122
rect 54514 75070 54516 75122
rect 54460 75058 54516 75070
rect 54124 55412 54404 55468
rect 54012 35474 54068 35486
rect 54012 35422 54014 35474
rect 54066 35422 54068 35474
rect 54012 34802 54068 35422
rect 54012 34750 54014 34802
rect 54066 34750 54068 34802
rect 54012 34738 54068 34750
rect 54012 34244 54068 34254
rect 54012 33458 54068 34188
rect 54012 33406 54014 33458
rect 54066 33406 54068 33458
rect 54012 33394 54068 33406
rect 54124 31948 54180 55412
rect 54908 43708 54964 75740
rect 55132 75730 55188 75740
rect 55580 75684 55636 76412
rect 55356 75682 55636 75684
rect 55356 75630 55582 75682
rect 55634 75630 55636 75682
rect 55356 75628 55636 75630
rect 55356 75122 55412 75628
rect 55580 75618 55636 75628
rect 55692 76356 55748 76366
rect 55804 76356 55860 77756
rect 56252 77364 56308 79200
rect 56252 77308 56756 77364
rect 55916 76356 55972 76366
rect 55804 76354 55972 76356
rect 55804 76302 55918 76354
rect 55970 76302 55972 76354
rect 55804 76300 55972 76302
rect 55356 75070 55358 75122
rect 55410 75070 55412 75122
rect 55356 75058 55412 75070
rect 55692 43708 55748 76300
rect 55916 76290 55972 76300
rect 56700 75906 56756 77308
rect 56924 76692 56980 79200
rect 56924 76626 56980 76636
rect 56700 75854 56702 75906
rect 56754 75854 56756 75906
rect 56700 75842 56756 75854
rect 57484 76468 57540 76478
rect 56028 75796 56084 75806
rect 54796 43652 54964 43708
rect 55468 43652 55748 43708
rect 55804 75794 56084 75796
rect 55804 75742 56030 75794
rect 56082 75742 56084 75794
rect 55804 75740 56084 75742
rect 54348 39060 54404 39070
rect 54348 35922 54404 39004
rect 54796 37828 54852 43652
rect 54908 41860 54964 41870
rect 55132 41860 55188 41870
rect 54964 41858 55188 41860
rect 54964 41806 55134 41858
rect 55186 41806 55188 41858
rect 54964 41804 55188 41806
rect 54908 41766 54964 41804
rect 55020 40962 55076 40974
rect 55020 40910 55022 40962
rect 55074 40910 55076 40962
rect 55020 40852 55076 40910
rect 55020 40786 55076 40796
rect 55132 40740 55188 41804
rect 55356 41746 55412 41758
rect 55356 41694 55358 41746
rect 55410 41694 55412 41746
rect 55356 41412 55412 41694
rect 55356 41346 55412 41356
rect 55356 41186 55412 41198
rect 55356 41134 55358 41186
rect 55410 41134 55412 41186
rect 55356 40852 55412 41134
rect 55356 40786 55412 40796
rect 55132 40674 55188 40684
rect 55468 37828 55524 43652
rect 55580 42756 55636 42766
rect 55580 42754 55748 42756
rect 55580 42702 55582 42754
rect 55634 42702 55748 42754
rect 55580 42700 55748 42702
rect 55580 42690 55636 42700
rect 55692 42194 55748 42700
rect 55692 42142 55694 42194
rect 55746 42142 55748 42194
rect 55692 42130 55748 42142
rect 55580 41412 55636 41422
rect 55580 41318 55636 41356
rect 54796 37772 54964 37828
rect 55468 37772 55748 37828
rect 54348 35870 54350 35922
rect 54402 35870 54404 35922
rect 54348 35474 54404 35870
rect 54348 35422 54350 35474
rect 54402 35422 54404 35474
rect 54348 35410 54404 35422
rect 54460 35588 54516 35598
rect 54236 35364 54292 35374
rect 54236 34130 54292 35308
rect 54460 34914 54516 35532
rect 54460 34862 54462 34914
rect 54514 34862 54516 34914
rect 54460 34850 54516 34862
rect 54796 34916 54852 34926
rect 54796 34802 54852 34860
rect 54796 34750 54798 34802
rect 54850 34750 54852 34802
rect 54796 34738 54852 34750
rect 54572 34356 54628 34366
rect 54572 34242 54628 34300
rect 54572 34190 54574 34242
rect 54626 34190 54628 34242
rect 54572 34178 54628 34190
rect 54236 34078 54238 34130
rect 54290 34078 54292 34130
rect 54236 34066 54292 34078
rect 54572 34018 54628 34030
rect 54572 33966 54574 34018
rect 54626 33966 54628 34018
rect 54124 31892 54292 31948
rect 54124 20914 54180 20926
rect 54124 20862 54126 20914
rect 54178 20862 54180 20914
rect 54012 20804 54068 20814
rect 53900 20748 54012 20804
rect 54012 20710 54068 20748
rect 53452 19070 53454 19122
rect 53506 19070 53508 19122
rect 53452 19058 53508 19070
rect 53564 19740 53732 19796
rect 54012 19906 54068 19918
rect 54012 19854 54014 19906
rect 54066 19854 54068 19906
rect 53340 18274 53396 18284
rect 53228 17668 53284 17678
rect 53116 17666 53284 17668
rect 53116 17614 53230 17666
rect 53282 17614 53284 17666
rect 53116 17612 53284 17614
rect 53228 17602 53284 17612
rect 53452 17668 53508 17678
rect 53452 17554 53508 17612
rect 53452 17502 53454 17554
rect 53506 17502 53508 17554
rect 53452 17490 53508 17502
rect 52892 16046 52894 16098
rect 52946 16046 52948 16098
rect 52892 16034 52948 16046
rect 53452 17332 53508 17342
rect 53452 14754 53508 17276
rect 53452 14702 53454 14754
rect 53506 14702 53508 14754
rect 53452 14690 53508 14702
rect 52780 14354 52836 14364
rect 51996 14254 51998 14306
rect 52050 14254 52052 14306
rect 51996 13858 52052 14254
rect 51996 13806 51998 13858
rect 52050 13806 52052 13858
rect 51996 13794 52052 13806
rect 52220 13970 52276 13982
rect 52220 13918 52222 13970
rect 52274 13918 52276 13970
rect 51884 9604 51940 9614
rect 51212 8372 51380 8428
rect 50988 6638 50990 6690
rect 51042 6638 51044 6690
rect 50988 6626 51044 6638
rect 50540 6580 50596 6590
rect 50540 6486 50596 6524
rect 51324 6580 51380 8372
rect 51436 8372 51604 8428
rect 51772 9268 51828 9278
rect 51884 9268 51940 9548
rect 51828 9212 51940 9268
rect 51436 6692 51492 8372
rect 51436 6598 51492 6636
rect 51324 6514 51380 6524
rect 50556 6300 50820 6310
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50556 6234 50820 6244
rect 49980 6066 50036 6076
rect 50764 6132 50820 6142
rect 50764 6038 50820 6076
rect 49868 5908 49924 5918
rect 49756 5852 49868 5908
rect 49868 5814 49924 5852
rect 50092 5796 50148 5806
rect 49756 5348 49812 5358
rect 49756 5234 49812 5292
rect 49756 5182 49758 5234
rect 49810 5182 49812 5234
rect 49756 5170 49812 5182
rect 50092 5234 50148 5740
rect 51212 5794 51268 5806
rect 51212 5742 51214 5794
rect 51266 5742 51268 5794
rect 50092 5182 50094 5234
rect 50146 5182 50148 5234
rect 50092 5170 50148 5182
rect 50540 5348 50596 5358
rect 50540 5122 50596 5292
rect 51212 5348 51268 5742
rect 51212 5282 51268 5292
rect 51660 5794 51716 5806
rect 51660 5742 51662 5794
rect 51714 5742 51716 5794
rect 50540 5070 50542 5122
rect 50594 5070 50596 5122
rect 50540 5058 50596 5070
rect 51100 5122 51156 5134
rect 51100 5070 51102 5122
rect 51154 5070 51156 5122
rect 49532 4286 49534 4338
rect 49586 4286 49588 4338
rect 49028 3948 49140 4004
rect 49308 4116 49364 4126
rect 48972 3938 49028 3948
rect 49196 3444 49252 3454
rect 48860 3442 49252 3444
rect 48860 3390 49198 3442
rect 49250 3390 49252 3442
rect 48860 3388 49252 3390
rect 49196 3378 49252 3388
rect 47292 800 47348 3332
rect 47964 3276 48132 3332
rect 47964 800 48020 3276
rect 49308 800 49364 4060
rect 49420 3780 49476 3790
rect 49420 3554 49476 3724
rect 49420 3502 49422 3554
rect 49474 3502 49476 3554
rect 49420 3490 49476 3502
rect 49532 3556 49588 4286
rect 49532 3490 49588 3500
rect 49868 4900 49924 4910
rect 49868 3442 49924 4844
rect 50556 4732 50820 4742
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50556 4666 50820 4676
rect 50540 4116 50596 4126
rect 50540 4022 50596 4060
rect 50092 4004 50148 4014
rect 50092 3668 50148 3948
rect 51100 3892 51156 5070
rect 51100 3826 51156 3836
rect 51548 5122 51604 5134
rect 51548 5070 51550 5122
rect 51602 5070 51604 5122
rect 51548 3780 51604 5070
rect 51548 3714 51604 3724
rect 50092 3554 50148 3612
rect 50652 3668 50708 3678
rect 50652 3574 50708 3612
rect 51324 3668 51380 3678
rect 50092 3502 50094 3554
rect 50146 3502 50148 3554
rect 50092 3490 50148 3502
rect 50876 3556 50932 3566
rect 49868 3390 49870 3442
rect 49922 3390 49924 3442
rect 49868 3378 49924 3390
rect 49980 3444 50036 3454
rect 49980 800 50036 3388
rect 50556 3164 50820 3174
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50556 3098 50820 3108
rect 50876 2996 50932 3500
rect 51212 3444 51268 3454
rect 51212 3350 51268 3388
rect 50652 2940 50932 2996
rect 50652 800 50708 2940
rect 51324 800 51380 3612
rect 51660 3444 51716 5742
rect 51772 3666 51828 9212
rect 51772 3614 51774 3666
rect 51826 3614 51828 3666
rect 51772 3602 51828 3614
rect 51884 8484 51940 8494
rect 51884 6466 51940 8428
rect 51884 6414 51886 6466
rect 51938 6414 51940 6466
rect 51660 3378 51716 3388
rect 51884 3444 51940 6414
rect 52108 4898 52164 4910
rect 52108 4846 52110 4898
rect 52162 4846 52164 4898
rect 51884 3378 51940 3388
rect 51996 3780 52052 3790
rect 51996 800 52052 3724
rect 52108 3556 52164 4846
rect 52220 4228 52276 13918
rect 53564 13746 53620 19740
rect 53676 19346 53732 19358
rect 53676 19294 53678 19346
rect 53730 19294 53732 19346
rect 53676 16772 53732 19294
rect 54012 17668 54068 19854
rect 54124 18564 54180 20862
rect 54236 20132 54292 31892
rect 54236 20018 54292 20076
rect 54348 21698 54404 21710
rect 54348 21646 54350 21698
rect 54402 21646 54404 21698
rect 54348 21588 54404 21646
rect 54348 20692 54404 21532
rect 54348 20130 54404 20636
rect 54348 20078 54350 20130
rect 54402 20078 54404 20130
rect 54348 20066 54404 20078
rect 54236 19966 54238 20018
rect 54290 19966 54292 20018
rect 54236 19954 54292 19966
rect 54572 19234 54628 33966
rect 54908 26908 54964 37772
rect 55580 35028 55636 35038
rect 55580 34934 55636 34972
rect 55020 34690 55076 34702
rect 55020 34638 55022 34690
rect 55074 34638 55076 34690
rect 55020 31948 55076 34638
rect 55468 34356 55524 34366
rect 55468 34262 55524 34300
rect 55020 31892 55300 31948
rect 54908 26852 55188 26908
rect 54908 21812 54964 21822
rect 54908 21586 54964 21756
rect 54908 21534 54910 21586
rect 54962 21534 54964 21586
rect 54908 21522 54964 21534
rect 54572 19182 54574 19234
rect 54626 19182 54628 19234
rect 54572 19170 54628 19182
rect 54796 20972 55076 21028
rect 54796 19122 54852 20972
rect 55020 20914 55076 20972
rect 55020 20862 55022 20914
rect 55074 20862 55076 20914
rect 55020 20850 55076 20862
rect 55132 20916 55188 26852
rect 55132 20802 55188 20860
rect 55132 20750 55134 20802
rect 55186 20750 55188 20802
rect 55132 20738 55188 20750
rect 55020 20692 55076 20702
rect 55020 20598 55076 20636
rect 55020 20020 55076 20030
rect 54796 19070 54798 19122
rect 54850 19070 54852 19122
rect 54796 19058 54852 19070
rect 54908 20018 55076 20020
rect 54908 19966 55022 20018
rect 55074 19966 55076 20018
rect 54908 19964 55076 19966
rect 54908 18900 54964 19964
rect 55020 19954 55076 19964
rect 54124 18498 54180 18508
rect 54684 18844 54964 18900
rect 54012 17602 54068 17612
rect 54124 17442 54180 17454
rect 54124 17390 54126 17442
rect 54178 17390 54180 17442
rect 53676 16716 53956 16772
rect 53788 15874 53844 15886
rect 53788 15822 53790 15874
rect 53842 15822 53844 15874
rect 53564 13694 53566 13746
rect 53618 13694 53620 13746
rect 53564 13682 53620 13694
rect 53676 15204 53732 15214
rect 52556 10836 52612 10846
rect 52332 6132 52388 6142
rect 52388 6076 52500 6132
rect 52332 6066 52388 6076
rect 52220 4162 52276 4172
rect 52332 3556 52388 3566
rect 52108 3500 52332 3556
rect 52332 3462 52388 3500
rect 52108 3332 52164 3342
rect 52444 3332 52500 6076
rect 52556 5796 52612 10780
rect 53676 9380 53732 15148
rect 53676 9314 53732 9324
rect 53452 7364 53508 7374
rect 52556 5794 52724 5796
rect 52556 5742 52558 5794
rect 52610 5742 52724 5794
rect 52556 5740 52724 5742
rect 52556 5730 52612 5740
rect 52556 4340 52612 4350
rect 52668 4340 52724 5740
rect 53228 4898 53284 4910
rect 53228 4846 53230 4898
rect 53282 4846 53284 4898
rect 52892 4340 52948 4350
rect 52668 4338 52948 4340
rect 52668 4286 52894 4338
rect 52946 4286 52948 4338
rect 52668 4284 52948 4286
rect 52556 4246 52612 4284
rect 52892 4274 52948 4284
rect 52108 3330 52500 3332
rect 52108 3278 52110 3330
rect 52162 3278 52500 3330
rect 52108 3276 52500 3278
rect 52668 4116 52724 4126
rect 52108 3266 52164 3276
rect 52668 800 52724 4060
rect 53228 3780 53284 4846
rect 53228 3714 53284 3724
rect 53004 3668 53060 3678
rect 53004 3554 53060 3612
rect 53004 3502 53006 3554
rect 53058 3502 53060 3554
rect 53004 3490 53060 3502
rect 53340 3668 53396 3678
rect 52780 3444 52836 3454
rect 52780 3350 52836 3388
rect 53340 800 53396 3612
rect 53452 3442 53508 7308
rect 53564 5122 53620 5134
rect 53564 5070 53566 5122
rect 53618 5070 53620 5122
rect 53564 4004 53620 5070
rect 53788 4564 53844 15822
rect 53900 13858 53956 16716
rect 53900 13806 53902 13858
rect 53954 13806 53956 13858
rect 53900 13794 53956 13806
rect 53900 11620 53956 11630
rect 53900 6132 53956 11564
rect 54124 8428 54180 17390
rect 54348 16882 54404 16894
rect 54348 16830 54350 16882
rect 54402 16830 54404 16882
rect 54348 16100 54404 16830
rect 54572 16882 54628 16894
rect 54572 16830 54574 16882
rect 54626 16830 54628 16882
rect 54572 16436 54628 16830
rect 54572 16370 54628 16380
rect 54460 16100 54516 16110
rect 54348 16098 54516 16100
rect 54348 16046 54462 16098
rect 54514 16046 54516 16098
rect 54348 16044 54516 16046
rect 54236 15316 54292 15326
rect 54348 15316 54404 16044
rect 54460 16034 54516 16044
rect 54684 15876 54740 18844
rect 54796 18676 54852 18686
rect 54796 18674 55076 18676
rect 54796 18622 54798 18674
rect 54850 18622 55076 18674
rect 54796 18620 55076 18622
rect 54796 18610 54852 18620
rect 54908 18452 54964 18462
rect 54796 18396 54908 18452
rect 54796 17332 54852 18396
rect 54908 18358 54964 18396
rect 54796 17276 54964 17332
rect 54684 15810 54740 15820
rect 54796 16098 54852 16110
rect 54796 16046 54798 16098
rect 54850 16046 54852 16098
rect 54292 15260 54404 15316
rect 54460 15314 54516 15326
rect 54460 15262 54462 15314
rect 54514 15262 54516 15314
rect 54236 15222 54292 15260
rect 54460 14756 54516 15262
rect 54460 14690 54516 14700
rect 54796 13860 54852 16046
rect 54796 13794 54852 13804
rect 54908 11172 54964 17276
rect 55020 15148 55076 18620
rect 55132 18564 55188 18574
rect 55132 17554 55188 18508
rect 55244 17668 55300 31892
rect 55356 21810 55412 21822
rect 55356 21758 55358 21810
rect 55410 21758 55412 21810
rect 55356 19572 55412 21758
rect 55468 21586 55524 21598
rect 55468 21534 55470 21586
rect 55522 21534 55524 21586
rect 55468 20356 55524 21534
rect 55692 21028 55748 37772
rect 55804 21812 55860 75740
rect 56028 75730 56084 75740
rect 57484 75122 57540 76412
rect 57484 75070 57486 75122
rect 57538 75070 57540 75122
rect 56924 73220 56980 73230
rect 56028 45332 56084 45342
rect 56028 42866 56084 45276
rect 56588 43540 56644 43550
rect 56028 42814 56030 42866
rect 56082 42814 56084 42866
rect 56028 42802 56084 42814
rect 56140 43538 56644 43540
rect 56140 43486 56590 43538
rect 56642 43486 56644 43538
rect 56140 43484 56644 43486
rect 56140 42196 56196 43484
rect 56588 43474 56644 43484
rect 56700 42530 56756 42542
rect 56700 42478 56702 42530
rect 56754 42478 56756 42530
rect 55916 42140 56196 42196
rect 56588 42196 56644 42206
rect 56700 42196 56756 42478
rect 56588 42194 56756 42196
rect 56588 42142 56590 42194
rect 56642 42142 56756 42194
rect 56588 42140 56756 42142
rect 55916 41410 55972 42140
rect 56588 42130 56644 42140
rect 56924 41972 56980 73164
rect 57484 55468 57540 75070
rect 57596 74788 57652 79200
rect 58268 76692 58324 79200
rect 58156 76636 58324 76692
rect 58716 76804 58772 76814
rect 58156 75572 58212 76636
rect 58268 76468 58324 76478
rect 58268 76466 58548 76468
rect 58268 76414 58270 76466
rect 58322 76414 58548 76466
rect 58268 76412 58548 76414
rect 58268 76402 58324 76412
rect 58156 75506 58212 75516
rect 58044 74788 58100 74798
rect 57596 74786 58100 74788
rect 57596 74734 58046 74786
rect 58098 74734 58100 74786
rect 57596 74732 58100 74734
rect 58044 74722 58100 74732
rect 57260 55412 57540 55468
rect 58492 74226 58548 76412
rect 58492 74174 58494 74226
rect 58546 74174 58548 74226
rect 57036 43428 57092 43438
rect 57036 43334 57092 43372
rect 57260 42866 57316 55412
rect 58492 45332 58548 74174
rect 58492 45266 58548 45276
rect 57260 42814 57262 42866
rect 57314 42814 57316 42866
rect 57260 42802 57316 42814
rect 58156 42868 58212 42878
rect 58156 42774 58212 42812
rect 57596 42530 57652 42542
rect 57596 42478 57598 42530
rect 57650 42478 57652 42530
rect 57484 42196 57540 42206
rect 57596 42196 57652 42478
rect 57484 42194 57652 42196
rect 57484 42142 57486 42194
rect 57538 42142 57652 42194
rect 57484 42140 57652 42142
rect 57484 42130 57540 42140
rect 56924 41916 57092 41972
rect 55916 41358 55918 41410
rect 55970 41358 55972 41410
rect 55916 41346 55972 41358
rect 56364 41748 56420 41758
rect 56364 41298 56420 41692
rect 56924 41746 56980 41758
rect 56924 41694 56926 41746
rect 56978 41694 56980 41746
rect 56924 41412 56980 41694
rect 56924 41346 56980 41356
rect 56364 41246 56366 41298
rect 56418 41246 56420 41298
rect 56364 38836 56420 41246
rect 56364 38770 56420 38780
rect 57036 37604 57092 41916
rect 57148 41858 57204 41870
rect 57148 41806 57150 41858
rect 57202 41806 57204 41858
rect 57148 41748 57204 41806
rect 58044 41860 58100 41870
rect 58044 41858 58324 41860
rect 58044 41806 58046 41858
rect 58098 41806 58324 41858
rect 58044 41804 58324 41806
rect 58044 41794 58100 41804
rect 57148 41682 57204 41692
rect 57820 41746 57876 41758
rect 57820 41694 57822 41746
rect 57874 41694 57876 41746
rect 57820 41412 57876 41694
rect 57876 41356 58212 41412
rect 57820 41346 57876 41356
rect 58156 41074 58212 41356
rect 58156 41022 58158 41074
rect 58210 41022 58212 41074
rect 58156 41010 58212 41022
rect 57148 40964 57204 40974
rect 57148 40628 57204 40908
rect 58268 40964 58324 41804
rect 58492 41188 58548 41198
rect 58492 41094 58548 41132
rect 58268 40898 58324 40908
rect 57148 40562 57204 40572
rect 58716 37716 58772 76748
rect 58828 76468 58884 76478
rect 58828 76374 58884 76412
rect 58940 75460 58996 79200
rect 59612 76468 59668 79200
rect 59836 76692 59892 76702
rect 59836 76598 59892 76636
rect 59612 76402 59668 76412
rect 58940 75394 58996 75404
rect 59052 75682 59108 75694
rect 59052 75630 59054 75682
rect 59106 75630 59108 75682
rect 59052 73892 59108 75630
rect 59388 75572 59444 75582
rect 59164 75516 59388 75572
rect 59164 74226 59220 75516
rect 59388 75478 59444 75516
rect 60284 75572 60340 79200
rect 60956 77026 61012 79200
rect 60956 76974 60958 77026
rect 61010 76974 61012 77026
rect 60956 76962 61012 76974
rect 61628 77028 61684 79200
rect 61628 76962 61684 76972
rect 61852 77026 61908 77038
rect 61852 76974 61854 77026
rect 61906 76974 61908 77026
rect 61740 76580 61796 76590
rect 61628 76578 61796 76580
rect 61628 76526 61742 76578
rect 61794 76526 61796 76578
rect 61628 76524 61796 76526
rect 60284 75506 60340 75516
rect 61180 75572 61236 75582
rect 61180 75478 61236 75516
rect 59724 75460 59780 75470
rect 60508 75460 60564 75470
rect 59724 75458 59892 75460
rect 59724 75406 59726 75458
rect 59778 75406 59892 75458
rect 59724 75404 59892 75406
rect 59724 75394 59780 75404
rect 59164 74174 59166 74226
rect 59218 74174 59220 74226
rect 59164 74162 59220 74174
rect 59500 73892 59556 73902
rect 59052 73890 59780 73892
rect 59052 73838 59502 73890
rect 59554 73838 59780 73890
rect 59052 73836 59780 73838
rect 59500 73826 59556 73836
rect 59612 70588 59668 70598
rect 59612 68068 59668 70532
rect 59052 68012 59668 68068
rect 59052 43708 59108 68012
rect 59724 62188 59780 73836
rect 59836 70644 59892 75404
rect 60508 75366 60564 75404
rect 60844 75460 60900 75470
rect 61292 75460 61348 75470
rect 60844 75458 61012 75460
rect 60844 75406 60846 75458
rect 60898 75406 61012 75458
rect 60844 75404 61012 75406
rect 60844 75394 60900 75404
rect 60396 74900 60452 74910
rect 60844 74900 60900 74910
rect 60396 74898 60900 74900
rect 60396 74846 60398 74898
rect 60450 74846 60846 74898
rect 60898 74846 60900 74898
rect 60396 74844 60900 74846
rect 60396 73948 60452 74844
rect 60844 74834 60900 74844
rect 60956 74788 61012 75404
rect 61292 75122 61348 75404
rect 61292 75070 61294 75122
rect 61346 75070 61348 75122
rect 61292 75058 61348 75070
rect 61516 75458 61572 75470
rect 61516 75406 61518 75458
rect 61570 75406 61572 75458
rect 60956 74732 61236 74788
rect 60844 74676 60900 74686
rect 59836 70578 59892 70588
rect 59948 73892 60452 73948
rect 60732 74620 60844 74676
rect 59500 62132 59780 62188
rect 59052 43652 59220 43708
rect 59164 41972 59220 43652
rect 59500 43428 59556 62132
rect 59500 43362 59556 43372
rect 59948 42868 60004 73892
rect 60396 55076 60452 55086
rect 60396 43708 60452 55020
rect 59948 42802 60004 42812
rect 60284 43652 60452 43708
rect 58940 41300 58996 41310
rect 58940 41298 59108 41300
rect 58940 41246 58942 41298
rect 58994 41246 59108 41298
rect 58940 41244 59108 41246
rect 58940 41234 58996 41244
rect 58716 37650 58772 37660
rect 57036 37538 57092 37548
rect 57036 36596 57092 36606
rect 57036 34356 57092 36540
rect 59052 36484 59108 41244
rect 59164 41074 59220 41916
rect 60172 41858 60228 41870
rect 60172 41806 60174 41858
rect 60226 41806 60228 41858
rect 59388 41188 59444 41198
rect 59388 41094 59444 41132
rect 59948 41188 60004 41198
rect 60172 41188 60228 41806
rect 59948 41186 60116 41188
rect 59948 41134 59950 41186
rect 60002 41134 60116 41186
rect 59948 41132 60116 41134
rect 59948 41122 60004 41132
rect 59164 41022 59166 41074
rect 59218 41022 59220 41074
rect 59164 41010 59220 41022
rect 59948 40626 60004 40638
rect 59948 40574 59950 40626
rect 60002 40574 60004 40626
rect 57036 34290 57092 34300
rect 58604 36428 59108 36484
rect 59612 40180 59668 40190
rect 58604 26180 58660 36428
rect 58604 26114 58660 26124
rect 56812 23828 56868 23838
rect 55916 21812 55972 21822
rect 55860 21810 55972 21812
rect 55860 21758 55918 21810
rect 55970 21758 55972 21810
rect 55860 21756 55972 21758
rect 55804 21718 55860 21756
rect 55916 21746 55972 21756
rect 55692 20972 55972 21028
rect 55804 20802 55860 20814
rect 55804 20750 55806 20802
rect 55858 20750 55860 20802
rect 55804 20356 55860 20750
rect 55524 20300 55860 20356
rect 55468 19906 55524 20300
rect 55468 19854 55470 19906
rect 55522 19854 55524 19906
rect 55468 19842 55524 19854
rect 55356 19506 55412 19516
rect 55916 18228 55972 20972
rect 56476 20804 56532 20814
rect 56476 20710 56532 20748
rect 56812 20692 56868 23772
rect 56924 20916 56980 20926
rect 56924 20822 56980 20860
rect 56812 20636 56980 20692
rect 56700 20020 56756 20030
rect 56700 19926 56756 19964
rect 56028 19908 56084 19918
rect 56028 19814 56084 19852
rect 56588 19572 56644 19582
rect 56140 19234 56196 19246
rect 56140 19182 56142 19234
rect 56194 19182 56196 19234
rect 56140 18564 56196 19182
rect 56364 19010 56420 19022
rect 56364 18958 56366 19010
rect 56418 18958 56420 19010
rect 56364 18900 56420 18958
rect 56364 18834 56420 18844
rect 56140 18498 56196 18508
rect 55916 18162 55972 18172
rect 55244 17602 55300 17612
rect 55468 17666 55524 17678
rect 55468 17614 55470 17666
rect 55522 17614 55524 17666
rect 55132 17502 55134 17554
rect 55186 17502 55188 17554
rect 55132 17332 55188 17502
rect 55132 17266 55188 17276
rect 55468 16884 55524 17614
rect 56588 17666 56644 19516
rect 56700 18452 56756 18462
rect 56700 18358 56756 18396
rect 56588 17614 56590 17666
rect 56642 17614 56644 17666
rect 56588 17602 56644 17614
rect 56812 17668 56868 17678
rect 56700 16884 56756 16894
rect 55468 16882 56756 16884
rect 55468 16830 56702 16882
rect 56754 16830 56756 16882
rect 55468 16828 56756 16830
rect 55356 16770 55412 16782
rect 55356 16718 55358 16770
rect 55410 16718 55412 16770
rect 55244 15204 55300 15242
rect 55020 15092 55188 15148
rect 55244 15138 55300 15148
rect 54908 11106 54964 11116
rect 55020 11508 55076 11518
rect 54124 8372 54404 8428
rect 53900 6130 54292 6132
rect 53900 6078 53902 6130
rect 53954 6078 54292 6130
rect 53900 6076 54292 6078
rect 53900 6066 53956 6076
rect 53788 4498 53844 4508
rect 54012 5236 54068 5246
rect 53900 4116 53956 4126
rect 53900 4022 53956 4060
rect 53564 3938 53620 3948
rect 53676 3780 53732 3790
rect 53676 3554 53732 3724
rect 53676 3502 53678 3554
rect 53730 3502 53732 3554
rect 53676 3490 53732 3502
rect 53452 3390 53454 3442
rect 53506 3390 53508 3442
rect 53452 3378 53508 3390
rect 54012 800 54068 5180
rect 54236 5122 54292 6076
rect 54348 5796 54404 8372
rect 54348 5730 54404 5740
rect 54236 5070 54238 5122
rect 54290 5070 54292 5122
rect 54236 5058 54292 5070
rect 55020 5012 55076 11452
rect 55132 8428 55188 15092
rect 55132 8372 55300 8428
rect 55244 7812 55300 8372
rect 55244 7746 55300 7756
rect 55356 5908 55412 16718
rect 55468 14644 55524 16828
rect 56700 16818 56756 16828
rect 56812 16660 56868 17612
rect 56476 16604 56868 16660
rect 56476 16210 56532 16604
rect 56476 16158 56478 16210
rect 56530 16158 56532 16210
rect 56476 16146 56532 16158
rect 55468 14578 55524 14588
rect 56588 11732 56644 11742
rect 56028 6468 56084 6478
rect 56028 6130 56084 6412
rect 56028 6078 56030 6130
rect 56082 6078 56084 6130
rect 56028 6066 56084 6078
rect 55356 5842 55412 5852
rect 55244 5236 55300 5246
rect 55244 5142 55300 5180
rect 56140 5236 56196 5246
rect 54236 3556 54292 3566
rect 54236 3462 54292 3500
rect 55020 3554 55076 4956
rect 55916 5012 55972 5022
rect 55916 4562 55972 4956
rect 55916 4510 55918 4562
rect 55970 4510 55972 4562
rect 55916 4498 55972 4510
rect 56028 3668 56084 3678
rect 56028 3574 56084 3612
rect 55020 3502 55022 3554
rect 55074 3502 55076 3554
rect 55020 3490 55076 3502
rect 55356 3556 55412 3566
rect 54684 3444 54740 3454
rect 54684 800 54740 3388
rect 55356 800 55412 3500
rect 56140 2212 56196 5180
rect 56588 4340 56644 11676
rect 56924 8428 56980 20636
rect 57260 20468 57316 20478
rect 57148 19906 57204 19918
rect 57148 19854 57150 19906
rect 57202 19854 57204 19906
rect 57036 19236 57092 19246
rect 57148 19236 57204 19854
rect 57260 19684 57316 20412
rect 57596 20132 57652 20142
rect 57596 20038 57652 20076
rect 57260 19618 57316 19628
rect 57036 19234 57204 19236
rect 57036 19182 57038 19234
rect 57090 19182 57204 19234
rect 57036 19180 57204 19182
rect 57036 9716 57092 19180
rect 58828 18452 58884 18462
rect 57148 18340 57204 18350
rect 57148 18246 57204 18284
rect 57036 9650 57092 9660
rect 57148 17668 57204 17678
rect 57148 17106 57204 17612
rect 58716 17668 58772 17678
rect 58716 17574 58772 17612
rect 58828 17554 58884 18396
rect 58828 17502 58830 17554
rect 58882 17502 58884 17554
rect 58828 17490 58884 17502
rect 57148 17054 57150 17106
rect 57202 17054 57204 17106
rect 57148 8932 57204 17054
rect 57148 8866 57204 8876
rect 57708 17442 57764 17454
rect 57708 17390 57710 17442
rect 57762 17390 57764 17442
rect 56812 8372 56980 8428
rect 56812 6466 56868 8372
rect 57708 7700 57764 17390
rect 57708 7634 57764 7644
rect 58156 13412 58212 13422
rect 56812 6414 56814 6466
rect 56866 6414 56868 6466
rect 56588 4246 56644 4284
rect 56700 5684 56756 5694
rect 56028 2156 56196 2212
rect 56028 800 56084 2156
rect 56700 800 56756 5628
rect 56812 5124 56868 6414
rect 56924 6468 56980 6478
rect 56924 5906 56980 6412
rect 58156 6244 58212 13356
rect 59500 12852 59556 12862
rect 59500 6692 59556 12796
rect 59612 9604 59668 40124
rect 59948 31948 60004 40574
rect 60060 40404 60116 41132
rect 60172 41122 60228 41132
rect 60060 40310 60116 40348
rect 59948 31892 60228 31948
rect 60172 24052 60228 31892
rect 60284 28756 60340 43652
rect 60620 41970 60676 41982
rect 60620 41918 60622 41970
rect 60674 41918 60676 41970
rect 60620 41860 60676 41918
rect 60620 41794 60676 41804
rect 60620 41298 60676 41310
rect 60620 41246 60622 41298
rect 60674 41246 60676 41298
rect 60508 41188 60564 41198
rect 60508 40402 60564 41132
rect 60508 40350 60510 40402
rect 60562 40350 60564 40402
rect 60508 40338 60564 40350
rect 60620 36372 60676 41246
rect 60732 40516 60788 74620
rect 60844 74610 60900 74620
rect 61180 74564 61236 74732
rect 60956 74508 61236 74564
rect 60956 41074 61012 74508
rect 61516 73948 61572 75406
rect 61628 74676 61684 76524
rect 61740 76514 61796 76524
rect 61852 75684 61908 76974
rect 62300 77026 62356 79200
rect 62972 77140 63028 79200
rect 62972 77074 63028 77084
rect 62300 76974 62302 77026
rect 62354 76974 62356 77026
rect 62300 76962 62356 76974
rect 62636 77028 62692 77038
rect 62636 76578 62692 76972
rect 63308 77026 63364 77038
rect 63308 76974 63310 77026
rect 63362 76974 63364 77026
rect 63308 76692 63364 76974
rect 63644 77028 63700 79200
rect 63644 76962 63700 76972
rect 63980 77140 64036 77150
rect 63308 76690 63588 76692
rect 63308 76638 63310 76690
rect 63362 76638 63588 76690
rect 63308 76636 63588 76638
rect 63308 76626 63364 76636
rect 62636 76526 62638 76578
rect 62690 76526 62692 76578
rect 62076 76468 62132 76478
rect 62132 76412 62468 76468
rect 62076 76374 62132 76412
rect 62412 75684 62468 76412
rect 62636 75906 62692 76526
rect 62636 75854 62638 75906
rect 62690 75854 62692 75906
rect 62636 75842 62692 75854
rect 62972 76578 63028 76590
rect 62972 76526 62974 76578
rect 63026 76526 63028 76578
rect 62636 75684 62692 75694
rect 61852 75682 62132 75684
rect 61852 75630 61854 75682
rect 61906 75630 62132 75682
rect 61852 75628 62132 75630
rect 62412 75682 62692 75684
rect 62412 75630 62638 75682
rect 62690 75630 62692 75682
rect 62412 75628 62692 75630
rect 61852 75618 61908 75628
rect 61740 75572 61796 75582
rect 61740 75122 61796 75516
rect 62076 75236 62132 75628
rect 62636 75618 62692 75628
rect 62188 75460 62244 75470
rect 62188 75458 62580 75460
rect 62188 75406 62190 75458
rect 62242 75406 62580 75458
rect 62188 75404 62580 75406
rect 62188 75394 62244 75404
rect 62076 75180 62244 75236
rect 61740 75070 61742 75122
rect 61794 75070 61796 75122
rect 61740 75058 61796 75070
rect 62188 75122 62244 75180
rect 62188 75070 62190 75122
rect 62242 75070 62244 75122
rect 62188 75058 62244 75070
rect 61628 74610 61684 74620
rect 61516 73892 61684 73948
rect 61628 43708 61684 73892
rect 62524 67228 62580 75404
rect 62972 67228 63028 76526
rect 63084 75906 63140 75918
rect 63084 75854 63086 75906
rect 63138 75854 63140 75906
rect 63084 75794 63140 75854
rect 63084 75742 63086 75794
rect 63138 75742 63140 75794
rect 63084 75730 63140 75742
rect 63532 75794 63588 76636
rect 63980 76690 64036 77084
rect 64316 77026 64372 79200
rect 64316 76974 64318 77026
rect 64370 76974 64372 77026
rect 64316 76962 64372 76974
rect 64652 77028 64708 77038
rect 63980 76638 63982 76690
rect 64034 76638 64036 76690
rect 63532 75742 63534 75794
rect 63586 75742 63588 75794
rect 63532 75730 63588 75742
rect 63644 76578 63700 76590
rect 63644 76526 63646 76578
rect 63698 76526 63700 76578
rect 62524 67172 62916 67228
rect 62972 67172 63140 67228
rect 62860 50428 62916 67172
rect 63084 50428 63140 67172
rect 63644 55468 63700 76526
rect 63980 75794 64036 76638
rect 64652 76690 64708 76972
rect 64988 76804 65044 79200
rect 65324 77026 65380 77038
rect 65324 76974 65326 77026
rect 65378 76974 65380 77026
rect 64988 76748 65156 76804
rect 64652 76638 64654 76690
rect 64706 76638 64708 76690
rect 64316 76580 64372 76590
rect 64316 76578 64484 76580
rect 64316 76526 64318 76578
rect 64370 76526 64484 76578
rect 64316 76524 64484 76526
rect 64316 76514 64372 76524
rect 63980 75742 63982 75794
rect 64034 75742 64036 75794
rect 63980 75730 64036 75742
rect 64316 76244 64372 76254
rect 62300 50372 62916 50428
rect 62972 50372 63140 50428
rect 63532 55412 63700 55468
rect 63756 75012 63812 75022
rect 61628 43652 62020 43708
rect 61068 41972 61124 41982
rect 61068 41878 61124 41916
rect 61628 41972 61684 41982
rect 61628 41878 61684 41916
rect 61964 41412 62020 43652
rect 62300 42868 62356 50372
rect 62300 42866 62916 42868
rect 62300 42814 62302 42866
rect 62354 42814 62916 42866
rect 62300 42812 62916 42814
rect 62300 42802 62356 42812
rect 62524 41970 62580 41982
rect 62524 41918 62526 41970
rect 62578 41918 62580 41970
rect 62076 41860 62132 41870
rect 62524 41860 62580 41918
rect 62860 41970 62916 42812
rect 62860 41918 62862 41970
rect 62914 41918 62916 41970
rect 62860 41906 62916 41918
rect 62076 41858 62580 41860
rect 62076 41806 62078 41858
rect 62130 41806 62580 41858
rect 62076 41804 62580 41806
rect 62076 41794 62132 41804
rect 60956 41022 60958 41074
rect 61010 41022 61012 41074
rect 60956 40740 61012 41022
rect 61516 41356 62020 41412
rect 60956 40684 61460 40740
rect 60732 40514 61348 40516
rect 60732 40462 60734 40514
rect 60786 40462 61348 40514
rect 60732 40460 61348 40462
rect 60732 40450 60788 40460
rect 61292 39730 61348 40460
rect 61292 39678 61294 39730
rect 61346 39678 61348 39730
rect 61292 39666 61348 39678
rect 61404 39732 61460 40684
rect 61516 40626 61572 41356
rect 61516 40574 61518 40626
rect 61570 40574 61572 40626
rect 61516 40562 61572 40574
rect 61628 41188 61684 41198
rect 61628 40404 61684 41132
rect 61964 41074 62020 41356
rect 61964 41022 61966 41074
rect 62018 41022 62020 41074
rect 61964 41010 62020 41022
rect 62412 41298 62468 41310
rect 62412 41246 62414 41298
rect 62466 41246 62468 41298
rect 61740 40404 61796 40414
rect 61684 40402 61796 40404
rect 61684 40350 61742 40402
rect 61794 40350 61796 40402
rect 61684 40348 61796 40350
rect 61628 40310 61684 40348
rect 61740 40338 61796 40348
rect 62300 40402 62356 40414
rect 62300 40350 62302 40402
rect 62354 40350 62356 40402
rect 62300 40292 62356 40350
rect 62188 40236 62300 40292
rect 61852 39732 61908 39742
rect 61404 39730 61908 39732
rect 61404 39678 61854 39730
rect 61906 39678 61908 39730
rect 61404 39676 61908 39678
rect 61852 39666 61908 39676
rect 62188 39058 62244 40236
rect 62300 40226 62356 40236
rect 62412 39844 62468 41246
rect 62524 41186 62580 41804
rect 62524 41134 62526 41186
rect 62578 41134 62580 41186
rect 62524 41076 62580 41134
rect 62524 41010 62580 41020
rect 62748 41858 62804 41870
rect 62748 41806 62750 41858
rect 62802 41806 62804 41858
rect 62748 40628 62804 41806
rect 62860 41188 62916 41226
rect 62860 41122 62916 41132
rect 62524 40572 62804 40628
rect 62860 40964 62916 40974
rect 62524 40180 62580 40572
rect 62860 40516 62916 40908
rect 62636 40460 62916 40516
rect 62972 40516 63028 50372
rect 63196 41972 63252 41982
rect 63196 41970 63364 41972
rect 63196 41918 63198 41970
rect 63250 41918 63364 41970
rect 63196 41916 63364 41918
rect 63196 41906 63252 41916
rect 63308 41188 63364 41916
rect 63532 41300 63588 55412
rect 63756 43540 63812 74956
rect 64316 67284 64372 76188
rect 64428 71652 64484 76524
rect 64540 75796 64596 75806
rect 64652 75796 64708 76638
rect 64988 76580 65044 76590
rect 64540 75794 64708 75796
rect 64540 75742 64542 75794
rect 64594 75742 64708 75794
rect 64540 75740 64708 75742
rect 64876 76578 65044 76580
rect 64876 76526 64990 76578
rect 65042 76526 65044 76578
rect 64876 76524 65044 76526
rect 64540 75730 64596 75740
rect 64876 71876 64932 76524
rect 64988 76514 65044 76524
rect 64988 75796 65044 75806
rect 65100 75796 65156 76748
rect 65324 76690 65380 76974
rect 65660 77026 65716 79200
rect 66332 77138 66388 79200
rect 66332 77086 66334 77138
rect 66386 77086 66388 77138
rect 66332 77074 66388 77086
rect 65660 76974 65662 77026
rect 65714 76974 65716 77026
rect 65660 76962 65716 76974
rect 66444 77026 66500 77038
rect 66444 76974 66446 77026
rect 66498 76974 66500 77026
rect 65324 76638 65326 76690
rect 65378 76638 65380 76690
rect 65324 75796 65380 76638
rect 66444 76690 66500 76974
rect 67004 77028 67060 79200
rect 67004 76962 67060 76972
rect 67116 77138 67172 77150
rect 67116 77086 67118 77138
rect 67170 77086 67172 77138
rect 67116 76692 67172 77086
rect 66444 76638 66446 76690
rect 66498 76638 66500 76690
rect 64988 75794 65268 75796
rect 64988 75742 64990 75794
rect 65042 75742 65268 75794
rect 64988 75740 65268 75742
rect 64988 75730 65044 75740
rect 65212 75682 65268 75740
rect 65324 75730 65380 75740
rect 65660 76578 65716 76590
rect 65660 76526 65662 76578
rect 65714 76526 65716 76578
rect 65212 75630 65214 75682
rect 65266 75630 65268 75682
rect 65212 75618 65268 75630
rect 65548 75460 65604 75470
rect 65548 75366 65604 75404
rect 64876 71820 65492 71876
rect 64428 71596 65156 71652
rect 64316 67228 64708 67284
rect 64652 67172 64820 67228
rect 63756 43474 63812 43484
rect 64540 55972 64596 55982
rect 64428 41972 64484 41982
rect 64428 41412 64484 41916
rect 64428 41346 64484 41356
rect 63308 40852 63364 41132
rect 63420 41186 63476 41198
rect 63420 41134 63422 41186
rect 63474 41134 63476 41186
rect 63420 41076 63476 41134
rect 63420 41010 63476 41020
rect 63532 41074 63588 41244
rect 64316 41188 64372 41226
rect 64372 41132 64484 41188
rect 64316 41122 64372 41132
rect 63532 41022 63534 41074
rect 63586 41022 63588 41074
rect 63532 41010 63588 41022
rect 64316 40962 64372 40974
rect 64316 40910 64318 40962
rect 64370 40910 64372 40962
rect 63308 40796 63588 40852
rect 62972 40514 63140 40516
rect 62972 40462 62974 40514
rect 63026 40462 63140 40514
rect 62972 40460 63140 40462
rect 62636 40402 62692 40460
rect 62972 40450 63028 40460
rect 62636 40350 62638 40402
rect 62690 40350 62692 40402
rect 62636 40338 62692 40350
rect 62748 40290 62804 40302
rect 62748 40238 62750 40290
rect 62802 40238 62804 40290
rect 62524 40124 62692 40180
rect 62412 39778 62468 39788
rect 62188 39006 62190 39058
rect 62242 39006 62244 39058
rect 62188 38994 62244 39006
rect 61852 38948 61908 38958
rect 61852 38854 61908 38892
rect 62524 38836 62580 38846
rect 62524 38742 62580 38780
rect 60620 36306 60676 36316
rect 61740 36260 61796 36270
rect 60284 28690 60340 28700
rect 60396 31108 60452 31118
rect 60396 27076 60452 31052
rect 60396 27010 60452 27020
rect 60172 23986 60228 23996
rect 61628 21252 61684 21262
rect 60172 10052 60228 10062
rect 59612 9538 59668 9548
rect 60060 9940 60116 9950
rect 60060 6692 60116 9884
rect 60172 7362 60228 9996
rect 60172 7310 60174 7362
rect 60226 7310 60228 7362
rect 60172 7028 60228 7310
rect 60172 6972 60676 7028
rect 60508 6692 60564 6702
rect 59500 6690 59892 6692
rect 59500 6638 59502 6690
rect 59554 6638 59892 6690
rect 59500 6636 59892 6638
rect 59500 6626 59556 6636
rect 58156 6178 58212 6188
rect 56924 5854 56926 5906
rect 56978 5854 56980 5906
rect 56924 5842 56980 5854
rect 59836 5906 59892 6636
rect 60060 6690 60564 6692
rect 60060 6638 60062 6690
rect 60114 6638 60510 6690
rect 60562 6638 60564 6690
rect 60060 6636 60564 6638
rect 60060 6626 60116 6636
rect 60508 6626 60564 6636
rect 59836 5854 59838 5906
rect 59890 5854 59892 5906
rect 59836 5842 59892 5854
rect 60060 6468 60116 6478
rect 57932 5684 57988 5694
rect 57932 5590 57988 5628
rect 59388 5684 59444 5694
rect 58156 5236 58212 5246
rect 58156 5142 58212 5180
rect 57148 5124 57204 5134
rect 56812 5122 57204 5124
rect 56812 5070 57150 5122
rect 57202 5070 57204 5122
rect 56812 5068 57204 5070
rect 57148 5058 57204 5068
rect 58716 4900 58772 4910
rect 58044 4340 58100 4350
rect 57372 4116 57428 4126
rect 57372 800 57428 4060
rect 57596 4114 57652 4126
rect 57596 4062 57598 4114
rect 57650 4062 57652 4114
rect 57596 3444 57652 4062
rect 58044 3666 58100 4284
rect 58044 3614 58046 3666
rect 58098 3614 58100 3666
rect 58044 3602 58100 3614
rect 57596 3378 57652 3388
rect 58044 3444 58100 3454
rect 58044 800 58100 3388
rect 58716 800 58772 4844
rect 59052 3668 59108 3678
rect 59052 3574 59108 3612
rect 59388 800 59444 5628
rect 59724 4116 59780 4126
rect 59724 4022 59780 4060
rect 60060 800 60116 6412
rect 60620 5122 60676 6972
rect 61516 6468 61572 6478
rect 61516 6374 61572 6412
rect 60844 5684 60900 5694
rect 60844 5590 60900 5628
rect 60620 5070 60622 5122
rect 60674 5070 60676 5122
rect 60620 5058 60676 5070
rect 60732 5236 60788 5246
rect 60732 800 60788 5180
rect 61516 4900 61572 4910
rect 61516 4806 61572 4844
rect 61628 4452 61684 21196
rect 61740 17780 61796 36204
rect 62076 33236 62132 33246
rect 62076 30100 62132 33180
rect 62076 30034 62132 30044
rect 62636 24052 62692 40124
rect 62748 35308 62804 40238
rect 62860 39844 62916 39854
rect 62860 38668 62916 39788
rect 63084 39732 63140 40460
rect 63532 40514 63588 40796
rect 63532 40462 63534 40514
rect 63586 40462 63588 40514
rect 63196 40404 63252 40414
rect 63196 40310 63252 40348
rect 63532 40404 63588 40462
rect 64204 40628 64260 40638
rect 63532 40338 63588 40348
rect 63756 40402 63812 40414
rect 63756 40350 63758 40402
rect 63810 40350 63812 40402
rect 63756 40292 63812 40350
rect 63420 39732 63476 39742
rect 63084 39730 63476 39732
rect 63084 39678 63422 39730
rect 63474 39678 63476 39730
rect 63084 39676 63476 39678
rect 63420 39666 63476 39676
rect 63756 39060 63812 40236
rect 63868 39060 63924 39070
rect 63756 39004 63868 39060
rect 63868 38994 63924 39004
rect 62860 38612 63252 38668
rect 62748 35252 63140 35308
rect 63084 24946 63140 35252
rect 63196 25172 63252 38612
rect 64204 26516 64260 40572
rect 64316 38668 64372 40910
rect 64428 40402 64484 41132
rect 64428 40350 64430 40402
rect 64482 40350 64484 40402
rect 64428 40338 64484 40350
rect 64316 38612 64484 38668
rect 64204 26450 64260 26460
rect 64428 25508 64484 38612
rect 64540 28420 64596 55916
rect 64652 40628 64708 40638
rect 64652 40534 64708 40572
rect 64652 39394 64708 39406
rect 64652 39342 64654 39394
rect 64706 39342 64708 39394
rect 64652 39060 64708 39342
rect 64652 38994 64708 39004
rect 64764 38052 64820 67172
rect 65100 41972 65156 71596
rect 64988 41858 65044 41870
rect 64988 41806 64990 41858
rect 65042 41806 65044 41858
rect 64988 41524 65044 41806
rect 64988 41458 65044 41468
rect 64988 41300 65044 41310
rect 64988 41206 65044 41244
rect 65100 40514 65156 41916
rect 65436 41972 65492 71820
rect 65660 67228 65716 76526
rect 65916 76076 66180 76086
rect 65972 76020 66020 76076
rect 66076 76020 66124 76076
rect 65916 76010 66180 76020
rect 65996 75796 66052 75806
rect 65996 75702 66052 75740
rect 66444 75794 66500 76638
rect 67004 76690 67172 76692
rect 67004 76638 67118 76690
rect 67170 76638 67172 76690
rect 67004 76636 67172 76638
rect 66444 75742 66446 75794
rect 66498 75742 66500 75794
rect 66444 75730 66500 75742
rect 66780 76578 66836 76590
rect 66780 76526 66782 76578
rect 66834 76526 66836 76578
rect 66108 75460 66164 75470
rect 66164 75404 66388 75460
rect 66108 75394 66164 75404
rect 65916 74508 66180 74518
rect 65972 74452 66020 74508
rect 66076 74452 66124 74508
rect 65916 74442 66180 74452
rect 65916 72940 66180 72950
rect 65972 72884 66020 72940
rect 66076 72884 66124 72940
rect 65916 72874 66180 72884
rect 65916 71372 66180 71382
rect 65972 71316 66020 71372
rect 66076 71316 66124 71372
rect 65916 71306 66180 71316
rect 65916 69804 66180 69814
rect 65972 69748 66020 69804
rect 66076 69748 66124 69804
rect 65916 69738 66180 69748
rect 65916 68236 66180 68246
rect 65972 68180 66020 68236
rect 66076 68180 66124 68236
rect 65916 68170 66180 68180
rect 65660 67172 65828 67228
rect 65772 42196 65828 67172
rect 65916 66668 66180 66678
rect 65972 66612 66020 66668
rect 66076 66612 66124 66668
rect 65916 66602 66180 66612
rect 65916 65100 66180 65110
rect 65972 65044 66020 65100
rect 66076 65044 66124 65100
rect 65916 65034 66180 65044
rect 65916 63532 66180 63542
rect 65972 63476 66020 63532
rect 66076 63476 66124 63532
rect 65916 63466 66180 63476
rect 65916 61964 66180 61974
rect 65972 61908 66020 61964
rect 66076 61908 66124 61964
rect 65916 61898 66180 61908
rect 65916 60396 66180 60406
rect 65972 60340 66020 60396
rect 66076 60340 66124 60396
rect 65916 60330 66180 60340
rect 65916 58828 66180 58838
rect 65972 58772 66020 58828
rect 66076 58772 66124 58828
rect 65916 58762 66180 58772
rect 65916 57260 66180 57270
rect 65972 57204 66020 57260
rect 66076 57204 66124 57260
rect 65916 57194 66180 57204
rect 65916 55692 66180 55702
rect 65972 55636 66020 55692
rect 66076 55636 66124 55692
rect 65916 55626 66180 55636
rect 65916 54124 66180 54134
rect 65972 54068 66020 54124
rect 66076 54068 66124 54124
rect 65916 54058 66180 54068
rect 65916 52556 66180 52566
rect 65972 52500 66020 52556
rect 66076 52500 66124 52556
rect 65916 52490 66180 52500
rect 65916 50988 66180 50998
rect 65972 50932 66020 50988
rect 66076 50932 66124 50988
rect 65916 50922 66180 50932
rect 65916 49420 66180 49430
rect 65972 49364 66020 49420
rect 66076 49364 66124 49420
rect 65916 49354 66180 49364
rect 65916 47852 66180 47862
rect 65972 47796 66020 47852
rect 66076 47796 66124 47852
rect 65916 47786 66180 47796
rect 65916 46284 66180 46294
rect 65972 46228 66020 46284
rect 66076 46228 66124 46284
rect 65916 46218 66180 46228
rect 65916 44716 66180 44726
rect 65972 44660 66020 44716
rect 66076 44660 66124 44716
rect 65916 44650 66180 44660
rect 65916 43148 66180 43158
rect 65972 43092 66020 43148
rect 66076 43092 66124 43148
rect 65916 43082 66180 43092
rect 65772 42130 65828 42140
rect 65884 41972 65940 41982
rect 65436 41970 65828 41972
rect 65436 41918 65438 41970
rect 65490 41918 65828 41970
rect 65436 41916 65828 41918
rect 65436 41906 65492 41916
rect 65100 40462 65102 40514
rect 65154 40462 65156 40514
rect 65100 40450 65156 40462
rect 65660 41524 65716 41534
rect 65660 41186 65716 41468
rect 65660 41134 65662 41186
rect 65714 41134 65716 41186
rect 65548 40404 65604 40414
rect 65660 40404 65716 41134
rect 65772 41074 65828 41916
rect 65884 41878 65940 41916
rect 65916 41580 66180 41590
rect 65972 41524 66020 41580
rect 66076 41524 66124 41580
rect 65916 41514 66180 41524
rect 65772 41022 65774 41074
rect 65826 41022 65828 41074
rect 65772 41010 65828 41022
rect 66332 40628 66388 75404
rect 66780 67228 66836 76526
rect 67004 75794 67060 76636
rect 67116 76626 67172 76636
rect 67452 77138 67508 77150
rect 67452 77086 67454 77138
rect 67506 77086 67508 77138
rect 67452 76578 67508 77086
rect 67676 77026 67732 79200
rect 67676 76974 67678 77026
rect 67730 76974 67732 77026
rect 67676 76962 67732 76974
rect 67788 77028 67844 77038
rect 67788 76692 67844 76972
rect 67452 76526 67454 76578
rect 67506 76526 67508 76578
rect 67452 76514 67508 76526
rect 67564 76690 67844 76692
rect 67564 76638 67790 76690
rect 67842 76638 67844 76690
rect 67564 76636 67844 76638
rect 67004 75742 67006 75794
rect 67058 75742 67060 75794
rect 67004 75730 67060 75742
rect 67564 75794 67620 76636
rect 67788 76626 67844 76636
rect 68348 76692 68404 79200
rect 69020 77250 69076 79200
rect 69020 77198 69022 77250
rect 69074 77198 69076 77250
rect 69020 77186 69076 77198
rect 68684 77138 68740 77150
rect 68684 77086 68686 77138
rect 68738 77086 68740 77138
rect 68348 76626 68404 76636
rect 68460 77026 68516 77038
rect 68460 76974 68462 77026
rect 68514 76974 68516 77026
rect 68460 76690 68516 76974
rect 68460 76638 68462 76690
rect 68514 76638 68516 76690
rect 68012 76580 68068 76590
rect 68012 76020 68068 76524
rect 67564 75742 67566 75794
rect 67618 75742 67620 75794
rect 67564 75730 67620 75742
rect 67676 75964 68068 76020
rect 68124 76578 68180 76590
rect 68124 76526 68126 76578
rect 68178 76526 68180 76578
rect 66780 67172 67060 67228
rect 67004 50428 67060 67172
rect 67004 50372 67172 50428
rect 66780 41186 66836 41198
rect 66780 41134 66782 41186
rect 66834 41134 66836 41186
rect 66332 40514 66388 40572
rect 66332 40462 66334 40514
rect 66386 40462 66388 40514
rect 66332 40450 66388 40462
rect 66556 40962 66612 40974
rect 66556 40910 66558 40962
rect 66610 40910 66612 40962
rect 65884 40404 65940 40414
rect 65548 40402 65940 40404
rect 65548 40350 65550 40402
rect 65602 40350 65886 40402
rect 65938 40350 65940 40402
rect 65548 40348 65940 40350
rect 65212 39620 65268 39630
rect 65212 39526 65268 39564
rect 65548 39618 65604 40348
rect 65884 40338 65940 40348
rect 65916 40012 66180 40022
rect 65972 39956 66020 40012
rect 66076 39956 66124 40012
rect 65916 39946 66180 39956
rect 65548 39566 65550 39618
rect 65602 39566 65604 39618
rect 65548 39554 65604 39566
rect 65772 39732 65828 39742
rect 65772 39508 65828 39676
rect 65772 39414 65828 39452
rect 66332 39620 66388 39630
rect 65884 39172 65940 39182
rect 65324 39060 65380 39070
rect 65324 38966 65380 39004
rect 65884 38834 65940 39116
rect 65884 38782 65886 38834
rect 65938 38782 65940 38834
rect 65884 38770 65940 38782
rect 66332 38834 66388 39564
rect 66332 38782 66334 38834
rect 66386 38782 66388 38834
rect 66332 38770 66388 38782
rect 66444 39394 66500 39406
rect 66444 39342 66446 39394
rect 66498 39342 66500 39394
rect 65916 38444 66180 38454
rect 65972 38388 66020 38444
rect 66076 38388 66124 38444
rect 65916 38378 66180 38388
rect 64764 37986 64820 37996
rect 65916 36876 66180 36886
rect 65972 36820 66020 36876
rect 66076 36820 66124 36876
rect 65916 36810 66180 36820
rect 65916 35308 66180 35318
rect 65972 35252 66020 35308
rect 66076 35252 66124 35308
rect 65916 35242 66180 35252
rect 64540 28354 64596 28364
rect 64652 33908 64708 33918
rect 64428 25442 64484 25452
rect 63196 25106 63252 25116
rect 63084 24894 63086 24946
rect 63138 24894 63140 24946
rect 63084 24882 63140 24894
rect 63308 25060 63364 25070
rect 63308 24946 63364 25004
rect 63308 24894 63310 24946
rect 63362 24894 63364 24946
rect 63308 24882 63364 24894
rect 64652 25060 64708 33852
rect 65916 33740 66180 33750
rect 65972 33684 66020 33740
rect 66076 33684 66124 33740
rect 65916 33674 66180 33684
rect 65916 32172 66180 32182
rect 65972 32116 66020 32172
rect 66076 32116 66124 32172
rect 65916 32106 66180 32116
rect 64652 24946 64708 25004
rect 64652 24894 64654 24946
rect 64706 24894 64708 24946
rect 64652 24882 64708 24894
rect 64764 31780 64820 31790
rect 63532 24724 63588 24734
rect 63532 24722 63812 24724
rect 63532 24670 63534 24722
rect 63586 24670 63812 24722
rect 63532 24668 63812 24670
rect 63532 24658 63588 24668
rect 63420 24612 63476 24622
rect 63420 24518 63476 24556
rect 63532 24276 63588 24286
rect 62860 24052 62916 24062
rect 63420 24052 63476 24062
rect 62636 24050 63028 24052
rect 62636 23998 62862 24050
rect 62914 23998 63028 24050
rect 62636 23996 63028 23998
rect 62860 23986 62916 23996
rect 62972 23938 63028 23996
rect 62972 23886 62974 23938
rect 63026 23886 63028 23938
rect 62972 23874 63028 23886
rect 63420 23938 63476 23996
rect 63532 24050 63588 24220
rect 63532 23998 63534 24050
rect 63586 23998 63588 24050
rect 63532 23986 63588 23998
rect 63420 23886 63422 23938
rect 63474 23886 63476 23938
rect 63420 23874 63476 23886
rect 63644 23714 63700 23726
rect 63644 23662 63646 23714
rect 63698 23662 63700 23714
rect 61740 17714 61796 17724
rect 61852 23156 61908 23166
rect 61628 4338 61684 4396
rect 61628 4286 61630 4338
rect 61682 4286 61684 4338
rect 61628 4274 61684 4286
rect 61404 3892 61460 3902
rect 61292 3836 61404 3892
rect 61292 1540 61348 3836
rect 61404 3826 61460 3836
rect 61852 3668 61908 23100
rect 63644 21812 63700 23662
rect 63756 23044 63812 24668
rect 64092 24052 64148 24062
rect 64092 23958 64148 23996
rect 63756 22978 63812 22988
rect 63644 21746 63700 21756
rect 62636 21476 62692 21486
rect 62188 8036 62244 8046
rect 62188 6356 62244 7980
rect 62188 6290 62244 6300
rect 62524 4452 62580 4462
rect 62524 4358 62580 4396
rect 62636 4114 62692 21420
rect 63532 20244 63588 20254
rect 63420 6690 63476 6702
rect 63420 6638 63422 6690
rect 63474 6638 63476 6690
rect 62636 4062 62638 4114
rect 62690 4062 62692 4114
rect 61404 3666 61908 3668
rect 61404 3614 61854 3666
rect 61906 3614 61908 3666
rect 61404 3612 61908 3614
rect 61404 3554 61460 3612
rect 61852 3602 61908 3612
rect 62076 3780 62132 3790
rect 61404 3502 61406 3554
rect 61458 3502 61460 3554
rect 61404 3490 61460 3502
rect 61292 1484 61460 1540
rect 61404 800 61460 1484
rect 62076 800 62132 3724
rect 62636 3554 62692 4062
rect 62636 3502 62638 3554
rect 62690 3502 62692 3554
rect 62636 3490 62692 3502
rect 62748 6468 62804 6478
rect 62748 800 62804 6412
rect 63196 6020 63252 6030
rect 63420 6020 63476 6638
rect 63252 5964 63476 6020
rect 63196 5926 63252 5964
rect 63532 5124 63588 20188
rect 64652 19012 64708 19022
rect 64540 18004 64596 18014
rect 63868 9156 63924 9166
rect 63868 6132 63924 9100
rect 64428 6468 64484 6478
rect 64428 6374 64484 6412
rect 63868 6130 64484 6132
rect 63868 6078 63870 6130
rect 63922 6078 64484 6130
rect 63868 6076 64484 6078
rect 63868 6066 63924 6076
rect 64428 5906 64484 6076
rect 64428 5854 64430 5906
rect 64482 5854 64484 5906
rect 64428 5842 64484 5854
rect 64428 5236 64484 5246
rect 64428 5142 64484 5180
rect 63756 5124 63812 5134
rect 63196 5122 63588 5124
rect 63196 5070 63534 5122
rect 63586 5070 63588 5122
rect 63196 5068 63588 5070
rect 63196 4562 63252 5068
rect 63532 5058 63588 5068
rect 63644 5068 63756 5124
rect 63196 4510 63198 4562
rect 63250 4510 63252 4562
rect 63196 4498 63252 4510
rect 63532 4226 63588 4238
rect 63532 4174 63534 4226
rect 63586 4174 63588 4226
rect 63532 4114 63588 4174
rect 63532 4062 63534 4114
rect 63586 4062 63588 4114
rect 63532 4050 63588 4062
rect 63644 980 63700 5068
rect 63756 5058 63812 5068
rect 64540 4340 64596 17948
rect 64652 5236 64708 18956
rect 64764 9828 64820 31724
rect 65916 30604 66180 30614
rect 65972 30548 66020 30604
rect 66076 30548 66124 30604
rect 65916 30538 66180 30548
rect 65916 29036 66180 29046
rect 65972 28980 66020 29036
rect 66076 28980 66124 29036
rect 65916 28970 66180 28980
rect 65916 27468 66180 27478
rect 65972 27412 66020 27468
rect 66076 27412 66124 27468
rect 65916 27402 66180 27412
rect 65916 25900 66180 25910
rect 65972 25844 66020 25900
rect 66076 25844 66124 25900
rect 65916 25834 66180 25844
rect 65916 24332 66180 24342
rect 65972 24276 66020 24332
rect 66076 24276 66124 24332
rect 65916 24266 66180 24276
rect 65916 22764 66180 22774
rect 65972 22708 66020 22764
rect 66076 22708 66124 22764
rect 65916 22698 66180 22708
rect 66444 21700 66500 39342
rect 66444 21634 66500 21644
rect 65916 21196 66180 21206
rect 65972 21140 66020 21196
rect 66076 21140 66124 21196
rect 65916 21130 66180 21140
rect 66556 20916 66612 40910
rect 66780 40402 66836 41134
rect 66892 40628 66948 40638
rect 66892 40626 67060 40628
rect 66892 40574 66894 40626
rect 66946 40574 67060 40626
rect 66892 40572 67060 40574
rect 66892 40562 66948 40572
rect 66780 40350 66782 40402
rect 66834 40350 66836 40402
rect 66668 39620 66724 39630
rect 66780 39620 66836 40350
rect 66724 39564 66836 39620
rect 66668 39526 66724 39564
rect 66668 38722 66724 38734
rect 66668 38670 66670 38722
rect 66722 38670 66724 38722
rect 66668 28980 66724 38670
rect 67004 32900 67060 40572
rect 67116 39956 67172 50372
rect 67452 40628 67508 40638
rect 67452 40534 67508 40572
rect 67564 40404 67620 40414
rect 67116 39900 67284 39956
rect 67116 39732 67172 39742
rect 67116 39638 67172 39676
rect 67228 39508 67284 39900
rect 67116 39452 67284 39508
rect 67116 38948 67172 39452
rect 67116 38854 67172 38892
rect 67564 39394 67620 40348
rect 67676 39508 67732 75964
rect 67900 41412 67956 41422
rect 67900 41076 67956 41356
rect 67900 40626 67956 41020
rect 67900 40574 67902 40626
rect 67954 40574 67956 40626
rect 67900 40562 67956 40574
rect 67676 39442 67732 39452
rect 67564 39342 67566 39394
rect 67618 39342 67620 39394
rect 67340 38834 67396 38846
rect 67340 38782 67342 38834
rect 67394 38782 67396 38834
rect 67340 38724 67396 38782
rect 67228 38612 67396 38668
rect 67228 38162 67284 38612
rect 67228 38110 67230 38162
rect 67282 38110 67284 38162
rect 67228 38098 67284 38110
rect 67564 36260 67620 39342
rect 68012 39060 68068 39070
rect 68012 38946 68068 39004
rect 68012 38894 68014 38946
rect 68066 38894 68068 38946
rect 68012 38882 68068 38894
rect 67900 38722 67956 38734
rect 67900 38670 67902 38722
rect 67954 38670 67956 38722
rect 67788 37828 67844 37838
rect 67788 37734 67844 37772
rect 67564 36194 67620 36204
rect 67004 32834 67060 32844
rect 66668 28914 66724 28924
rect 67900 26908 67956 38670
rect 68124 37828 68180 76526
rect 68460 75794 68516 76638
rect 68460 75742 68462 75794
rect 68514 75742 68516 75794
rect 68460 75730 68516 75742
rect 68236 40404 68292 40414
rect 68236 40310 68292 40348
rect 68572 40402 68628 40414
rect 68572 40350 68574 40402
rect 68626 40350 68628 40402
rect 68460 39844 68516 39854
rect 68348 39620 68404 39630
rect 68236 39618 68404 39620
rect 68236 39566 68350 39618
rect 68402 39566 68404 39618
rect 68236 39564 68404 39566
rect 68236 38834 68292 39564
rect 68348 39554 68404 39564
rect 68460 39508 68516 39788
rect 68460 39414 68516 39452
rect 68236 38782 68238 38834
rect 68290 38782 68292 38834
rect 68236 38724 68292 38782
rect 68572 39172 68628 40350
rect 68572 38834 68628 39116
rect 68684 39060 68740 77086
rect 69132 76692 69188 76702
rect 68796 76580 68852 76590
rect 68796 76486 68852 76524
rect 69020 75796 69076 75806
rect 69132 75796 69188 76636
rect 69468 76580 69524 76590
rect 69020 75794 69188 75796
rect 69020 75742 69022 75794
rect 69074 75742 69188 75794
rect 69020 75740 69188 75742
rect 69244 76578 69524 76580
rect 69244 76526 69470 76578
rect 69522 76526 69524 76578
rect 69244 76524 69524 76526
rect 69020 75730 69076 75740
rect 68684 38994 68740 39004
rect 68908 58212 68964 58222
rect 68572 38782 68574 38834
rect 68626 38782 68628 38834
rect 68572 38770 68628 38782
rect 68236 38612 68404 38668
rect 68348 38050 68404 38612
rect 68348 37998 68350 38050
rect 68402 37998 68404 38050
rect 68348 37986 68404 37998
rect 68460 37938 68516 37950
rect 68460 37886 68462 37938
rect 68514 37886 68516 37938
rect 68460 37828 68516 37886
rect 68124 37772 68516 37828
rect 68684 37828 68740 37838
rect 68124 37490 68180 37772
rect 68124 37438 68126 37490
rect 68178 37438 68180 37490
rect 68124 37426 68180 37438
rect 68684 37490 68740 37772
rect 68684 37438 68686 37490
rect 68738 37438 68740 37490
rect 68684 37426 68740 37438
rect 67788 26852 67956 26908
rect 68012 32900 68068 32910
rect 67788 23380 67844 26852
rect 67788 23314 67844 23324
rect 66556 20850 66612 20860
rect 67116 22260 67172 22270
rect 65916 19628 66180 19638
rect 65972 19572 66020 19628
rect 66076 19572 66124 19628
rect 65916 19562 66180 19572
rect 67116 19012 67172 22204
rect 68012 21588 68068 32844
rect 68908 28196 68964 58156
rect 69244 50428 69300 76524
rect 69468 76514 69524 76524
rect 69692 76580 69748 79200
rect 70252 77250 70308 77262
rect 70252 77198 70254 77250
rect 70306 77198 70308 77250
rect 70252 76580 70308 77198
rect 70364 77028 70420 79200
rect 70364 76962 70420 76972
rect 71036 77026 71092 79200
rect 71036 76974 71038 77026
rect 71090 76974 71092 77026
rect 71036 76962 71092 76974
rect 69692 76514 69748 76524
rect 70028 76578 70308 76580
rect 70028 76526 70254 76578
rect 70306 76526 70308 76578
rect 70028 76524 70308 76526
rect 69356 76020 69412 76030
rect 69356 67228 69412 75964
rect 70028 75794 70084 76524
rect 70252 76514 70308 76524
rect 70588 76748 71540 76804
rect 70588 76578 70644 76748
rect 70924 76580 70980 76590
rect 70588 76526 70590 76578
rect 70642 76526 70644 76578
rect 70588 76514 70644 76526
rect 70700 76524 70924 76580
rect 70028 75742 70030 75794
rect 70082 75742 70084 75794
rect 70028 75730 70084 75742
rect 70476 76132 70532 76142
rect 69356 67172 69524 67228
rect 69244 50372 69412 50428
rect 69020 40964 69076 40974
rect 69244 40964 69300 40974
rect 69020 40962 69300 40964
rect 69020 40910 69022 40962
rect 69074 40910 69246 40962
rect 69298 40910 69300 40962
rect 69020 40908 69300 40910
rect 69020 40404 69076 40908
rect 69244 40898 69300 40908
rect 69356 40628 69412 50372
rect 69468 40740 69524 67172
rect 70028 66276 70084 66286
rect 70028 50428 70084 66220
rect 69916 50372 70084 50428
rect 69804 41858 69860 41870
rect 69804 41806 69806 41858
rect 69858 41806 69860 41858
rect 69804 41746 69860 41806
rect 69804 41694 69806 41746
rect 69858 41694 69860 41746
rect 69804 41682 69860 41694
rect 69580 41412 69636 41422
rect 69580 41074 69636 41356
rect 69580 41022 69582 41074
rect 69634 41022 69636 41074
rect 69580 41010 69636 41022
rect 69468 40684 69636 40740
rect 69356 40514 69412 40572
rect 69356 40462 69358 40514
rect 69410 40462 69412 40514
rect 69356 40450 69412 40462
rect 69020 40338 69076 40348
rect 69468 40290 69524 40302
rect 69468 40238 69470 40290
rect 69522 40238 69524 40290
rect 69244 39620 69300 39630
rect 69132 39618 69300 39620
rect 69132 39566 69246 39618
rect 69298 39566 69300 39618
rect 69132 39564 69300 39566
rect 69020 39172 69076 39182
rect 69132 39172 69188 39564
rect 69244 39554 69300 39564
rect 69356 39396 69412 39406
rect 69356 39302 69412 39340
rect 69076 39116 69188 39172
rect 69020 39106 69076 39116
rect 69020 38836 69076 38846
rect 69020 37490 69076 38780
rect 69132 38668 69188 39116
rect 69244 39060 69300 39070
rect 69244 38966 69300 39004
rect 69132 38612 69300 38668
rect 69244 38050 69300 38612
rect 69244 37998 69246 38050
rect 69298 37998 69300 38050
rect 69244 37986 69300 37998
rect 69020 37438 69022 37490
rect 69074 37438 69076 37490
rect 69020 37426 69076 37438
rect 69244 37826 69300 37838
rect 69244 37774 69246 37826
rect 69298 37774 69300 37826
rect 69020 36260 69076 36270
rect 69020 36166 69076 36204
rect 68908 28130 68964 28140
rect 68908 23604 68964 23614
rect 68908 22484 68964 23548
rect 68908 22418 68964 22428
rect 69244 22484 69300 37774
rect 69356 37266 69412 37278
rect 69356 37214 69358 37266
rect 69410 37214 69412 37266
rect 69356 36260 69412 37214
rect 69356 36194 69412 36204
rect 69244 22418 69300 22428
rect 69468 22372 69524 40238
rect 69580 38388 69636 40684
rect 69692 40402 69748 40414
rect 69692 40350 69694 40402
rect 69746 40350 69748 40402
rect 69692 39508 69748 40350
rect 69692 39442 69748 39452
rect 69692 38948 69748 38958
rect 69692 38854 69748 38892
rect 69580 38322 69636 38332
rect 69804 38724 69860 38734
rect 69804 38164 69860 38668
rect 69804 38050 69860 38108
rect 69804 37998 69806 38050
rect 69858 37998 69860 38050
rect 69804 37986 69860 37998
rect 69692 37828 69748 37838
rect 69692 37490 69748 37772
rect 69692 37438 69694 37490
rect 69746 37438 69748 37490
rect 69692 37426 69748 37438
rect 69916 32900 69972 50372
rect 70476 42308 70532 76076
rect 70700 75794 70756 76524
rect 70924 76486 70980 76524
rect 71260 76578 71316 76590
rect 71260 76526 71262 76578
rect 71314 76526 71316 76578
rect 70700 75742 70702 75794
rect 70754 75742 70756 75794
rect 70700 75730 70756 75742
rect 70476 42242 70532 42252
rect 70812 53060 70868 53070
rect 70252 41858 70308 41870
rect 70252 41806 70254 41858
rect 70306 41806 70308 41858
rect 70140 41746 70196 41758
rect 70140 41694 70142 41746
rect 70194 41694 70196 41746
rect 70140 41186 70196 41694
rect 70140 41134 70142 41186
rect 70194 41134 70196 41186
rect 70140 40402 70196 41134
rect 70252 40852 70308 41806
rect 70700 41858 70756 41870
rect 70700 41806 70702 41858
rect 70754 41806 70756 41858
rect 70252 40786 70308 40796
rect 70476 41636 70532 41646
rect 70476 41298 70532 41580
rect 70476 41246 70478 41298
rect 70530 41246 70532 41298
rect 70476 40516 70532 41246
rect 70700 41300 70756 41806
rect 70700 40740 70756 41244
rect 70700 40674 70756 40684
rect 70476 40450 70532 40460
rect 70700 40516 70756 40526
rect 70140 40350 70142 40402
rect 70194 40350 70196 40402
rect 70140 40180 70196 40350
rect 70700 40402 70756 40460
rect 70700 40350 70702 40402
rect 70754 40350 70756 40402
rect 70700 40338 70756 40350
rect 70140 40114 70196 40124
rect 70700 39732 70756 39742
rect 70364 39620 70420 39630
rect 70364 39526 70420 39564
rect 70588 39620 70644 39630
rect 70700 39620 70756 39676
rect 70588 39618 70756 39620
rect 70588 39566 70590 39618
rect 70642 39566 70756 39618
rect 70588 39564 70756 39566
rect 70588 39554 70644 39564
rect 70028 39508 70084 39518
rect 70028 38836 70084 39452
rect 70028 38770 70084 38780
rect 70252 39394 70308 39406
rect 70252 39342 70254 39394
rect 70306 39342 70308 39394
rect 70140 38276 70196 38286
rect 70140 37938 70196 38220
rect 70140 37886 70142 37938
rect 70194 37886 70196 37938
rect 70140 37874 70196 37886
rect 69916 32834 69972 32844
rect 70252 27858 70308 39342
rect 70476 39396 70532 39406
rect 70476 39060 70532 39340
rect 70476 39004 70644 39060
rect 70364 38836 70420 38846
rect 70364 38742 70420 38780
rect 70476 38722 70532 38734
rect 70476 38670 70478 38722
rect 70530 38670 70532 38722
rect 70476 38668 70532 38670
rect 70364 38612 70532 38668
rect 70588 38668 70644 39004
rect 70700 38836 70756 38846
rect 70700 38742 70756 38780
rect 70588 38612 70756 38668
rect 70364 28642 70420 38612
rect 70588 38164 70644 38174
rect 70588 38070 70644 38108
rect 70588 37828 70644 37838
rect 70588 37380 70644 37772
rect 70588 37286 70644 37324
rect 70588 35588 70644 35598
rect 70588 32004 70644 35532
rect 70588 31938 70644 31948
rect 70700 30548 70756 38612
rect 70812 34356 70868 53004
rect 71148 41858 71204 41870
rect 71148 41806 71150 41858
rect 71202 41806 71204 41858
rect 71036 41746 71092 41758
rect 71036 41694 71038 41746
rect 71090 41694 71092 41746
rect 71036 41412 71092 41694
rect 71148 41748 71204 41806
rect 71148 41682 71204 41692
rect 71148 41412 71204 41422
rect 71036 41410 71204 41412
rect 71036 41358 71150 41410
rect 71202 41358 71204 41410
rect 71036 41356 71204 41358
rect 71148 41346 71204 41356
rect 70924 41186 70980 41198
rect 70924 41134 70926 41186
rect 70978 41134 70980 41186
rect 70924 40852 70980 41134
rect 70924 40786 70980 40796
rect 70924 40514 70980 40526
rect 70924 40462 70926 40514
rect 70978 40462 70980 40514
rect 70924 39732 70980 40462
rect 71260 40292 71316 76526
rect 71372 75906 71428 75918
rect 71372 75854 71374 75906
rect 71426 75854 71428 75906
rect 71372 75794 71428 75854
rect 71372 75742 71374 75794
rect 71426 75742 71428 75794
rect 71372 75730 71428 75742
rect 71372 41300 71428 41310
rect 71372 41206 71428 41244
rect 71372 40628 71428 40638
rect 71372 40534 71428 40572
rect 71260 40226 71316 40236
rect 71036 39788 71428 39844
rect 71036 39732 71092 39788
rect 70980 39676 71092 39732
rect 70924 39666 70980 39676
rect 70924 39508 70980 39518
rect 70924 39414 70980 39452
rect 70924 38948 70980 38958
rect 71036 38948 71092 39676
rect 71372 39618 71428 39788
rect 71372 39566 71374 39618
rect 71426 39566 71428 39618
rect 71372 39554 71428 39566
rect 71484 39620 71540 76748
rect 71596 76578 71652 76590
rect 71596 76526 71598 76578
rect 71650 76526 71652 76578
rect 71596 67228 71652 76526
rect 71708 76580 71764 79200
rect 71708 76514 71764 76524
rect 71820 77028 71876 77038
rect 71820 76466 71876 76972
rect 71820 76414 71822 76466
rect 71874 76414 71876 76466
rect 71820 75906 71876 76414
rect 71820 75854 71822 75906
rect 71874 75854 71876 75906
rect 71820 75842 71876 75854
rect 71932 77026 71988 77038
rect 71932 76974 71934 77026
rect 71986 76974 71988 77026
rect 71932 75794 71988 76974
rect 72268 76578 72324 76590
rect 72268 76526 72270 76578
rect 72322 76526 72324 76578
rect 72268 76244 72324 76526
rect 72268 76178 72324 76188
rect 71932 75742 71934 75794
rect 71986 75742 71988 75794
rect 71932 75730 71988 75742
rect 72380 75794 72436 79200
rect 72604 77026 72660 77038
rect 72604 76974 72606 77026
rect 72658 76974 72660 77026
rect 72604 76690 72660 76974
rect 72604 76638 72606 76690
rect 72658 76638 72660 76690
rect 72604 76626 72660 76638
rect 73052 76692 73108 79200
rect 73052 76626 73108 76636
rect 72940 76580 72996 76590
rect 72380 75742 72382 75794
rect 72434 75742 72436 75794
rect 72380 75684 72436 75742
rect 72828 76578 72996 76580
rect 72828 76526 72942 76578
rect 72994 76526 72996 76578
rect 72828 76524 72996 76526
rect 72604 75684 72660 75694
rect 72380 75682 72660 75684
rect 72380 75630 72606 75682
rect 72658 75630 72660 75682
rect 72380 75628 72660 75630
rect 72604 75618 72660 75628
rect 72156 68852 72212 68862
rect 71596 67172 72100 67228
rect 72044 50428 72100 67172
rect 71820 50372 72100 50428
rect 71596 41748 71652 41758
rect 71596 41410 71652 41692
rect 71596 41358 71598 41410
rect 71650 41358 71652 41410
rect 71596 41346 71652 41358
rect 71708 41524 71764 41534
rect 71708 41410 71764 41468
rect 71708 41358 71710 41410
rect 71762 41358 71764 41410
rect 71708 41346 71764 41358
rect 71260 39506 71316 39518
rect 71260 39454 71262 39506
rect 71314 39454 71316 39506
rect 70924 38946 71092 38948
rect 70924 38894 70926 38946
rect 70978 38894 71092 38946
rect 70924 38892 71092 38894
rect 70924 38882 70980 38892
rect 71036 38050 71092 38892
rect 71036 37998 71038 38050
rect 71090 37998 71092 38050
rect 71036 37986 71092 37998
rect 71148 39394 71204 39406
rect 71148 39342 71150 39394
rect 71202 39342 71204 39394
rect 70924 37940 70980 37950
rect 70924 37490 70980 37884
rect 70924 37438 70926 37490
rect 70978 37438 70980 37490
rect 70924 37426 70980 37438
rect 71148 35028 71204 39342
rect 71260 39396 71316 39454
rect 71260 39330 71316 39340
rect 71372 39060 71428 39070
rect 71484 39060 71540 39564
rect 71372 39058 71540 39060
rect 71372 39006 71374 39058
rect 71426 39006 71540 39058
rect 71372 39004 71540 39006
rect 71372 38994 71428 39004
rect 71260 38836 71316 38846
rect 71820 38836 71876 50372
rect 72044 45892 72100 45902
rect 71932 39844 71988 39854
rect 71932 39730 71988 39788
rect 71932 39678 71934 39730
rect 71986 39678 71988 39730
rect 71932 39666 71988 39678
rect 71316 38780 71876 38836
rect 71260 38668 71316 38780
rect 71260 38612 71428 38668
rect 71260 38052 71316 38062
rect 71260 37958 71316 37996
rect 71260 37380 71316 37390
rect 71260 37286 71316 37324
rect 71260 36596 71316 36606
rect 71372 36596 71428 38612
rect 71932 38164 71988 38174
rect 71820 38052 71876 38062
rect 71708 37996 71820 38052
rect 71596 37940 71652 37950
rect 71596 37846 71652 37884
rect 71260 36594 71428 36596
rect 71260 36542 71262 36594
rect 71314 36542 71428 36594
rect 71260 36540 71428 36542
rect 71484 37826 71540 37838
rect 71484 37774 71486 37826
rect 71538 37774 71540 37826
rect 71260 36530 71316 36540
rect 71484 35252 71540 37774
rect 71596 37492 71652 37502
rect 71708 37492 71764 37996
rect 71820 37986 71876 37996
rect 71596 37490 71764 37492
rect 71596 37438 71598 37490
rect 71650 37438 71764 37490
rect 71596 37436 71764 37438
rect 71596 37426 71652 37436
rect 71932 36594 71988 38108
rect 71932 36542 71934 36594
rect 71986 36542 71988 36594
rect 71932 36530 71988 36542
rect 71708 35588 71764 35598
rect 71708 35494 71764 35532
rect 72044 35308 72100 45836
rect 72156 41860 72212 68796
rect 72828 67228 72884 76524
rect 72940 76514 72996 76524
rect 73164 76580 73220 76590
rect 73164 76468 73220 76524
rect 73724 76580 73780 79200
rect 74396 77026 74452 79200
rect 75068 77250 75124 79200
rect 75740 77476 75796 79200
rect 76412 77476 76468 79200
rect 75740 77420 76244 77476
rect 76412 77420 76916 77476
rect 75068 77198 75070 77250
rect 75122 77198 75124 77250
rect 75068 77186 75124 77198
rect 75852 77250 75908 77262
rect 75852 77198 75854 77250
rect 75906 77198 75908 77250
rect 74396 76974 74398 77026
rect 74450 76974 74452 77026
rect 74396 76962 74452 76974
rect 75068 77026 75124 77038
rect 75068 76974 75070 77026
rect 75122 76974 75124 77026
rect 73724 76514 73780 76524
rect 74060 76692 74116 76702
rect 73164 76466 73444 76468
rect 73164 76414 73166 76466
rect 73218 76414 73444 76466
rect 73164 76412 73444 76414
rect 73164 76402 73220 76412
rect 73388 75794 73444 76412
rect 73388 75742 73390 75794
rect 73442 75742 73444 75794
rect 73388 75730 73444 75742
rect 73948 75796 74004 75806
rect 74060 75796 74116 76636
rect 73948 75794 74116 75796
rect 73948 75742 73950 75794
rect 74002 75742 74116 75794
rect 73948 75740 74116 75742
rect 74396 76578 74452 76590
rect 74396 76526 74398 76578
rect 74450 76526 74452 76578
rect 73948 75730 74004 75740
rect 73836 75684 73892 75694
rect 72940 75460 72996 75470
rect 72940 75458 73332 75460
rect 72940 75406 72942 75458
rect 72994 75406 73332 75458
rect 72940 75404 73332 75406
rect 72940 75394 72996 75404
rect 73276 67228 73332 75404
rect 73724 74004 73780 74014
rect 72828 67172 72996 67228
rect 73276 67172 73556 67228
rect 72940 50428 72996 67172
rect 72828 50372 72996 50428
rect 72156 41794 72212 41804
rect 72604 48580 72660 48590
rect 72268 40516 72324 40526
rect 72268 38276 72324 40460
rect 72380 40292 72436 40302
rect 72380 39618 72436 40236
rect 72380 39566 72382 39618
rect 72434 39566 72436 39618
rect 72380 39396 72436 39566
rect 72380 39330 72436 39340
rect 72492 40290 72548 40302
rect 72492 40238 72494 40290
rect 72546 40238 72548 40290
rect 72492 38836 72548 40238
rect 72492 38742 72548 38780
rect 72492 38612 72548 38622
rect 72268 38164 72324 38220
rect 72156 38108 72324 38164
rect 72380 38556 72492 38612
rect 72156 38050 72212 38108
rect 72156 37998 72158 38050
rect 72210 37998 72212 38050
rect 72156 37986 72212 37998
rect 72268 37940 72324 37950
rect 72268 37380 72324 37884
rect 72380 37380 72436 38556
rect 72492 38546 72548 38556
rect 72604 38164 72660 48524
rect 72828 39620 72884 50372
rect 73164 45668 73220 45678
rect 73052 45612 73164 45668
rect 72940 40740 72996 40750
rect 72940 40626 72996 40684
rect 72940 40574 72942 40626
rect 72994 40574 72996 40626
rect 72940 40562 72996 40574
rect 72828 39554 72884 39564
rect 72940 39730 72996 39742
rect 72940 39678 72942 39730
rect 72994 39678 72996 39730
rect 72940 39172 72996 39678
rect 73052 39396 73108 45612
rect 73164 45602 73220 45612
rect 73276 41076 73332 41086
rect 73276 40982 73332 41020
rect 73388 40962 73444 40974
rect 73388 40910 73390 40962
rect 73442 40910 73444 40962
rect 73388 40628 73444 40910
rect 73164 40572 73444 40628
rect 73164 39618 73220 40572
rect 73388 40404 73444 40414
rect 73388 40310 73444 40348
rect 73164 39566 73166 39618
rect 73218 39566 73220 39618
rect 73164 39554 73220 39566
rect 73276 39732 73332 39742
rect 73052 39340 73220 39396
rect 72940 39106 72996 39116
rect 72716 38948 72772 38958
rect 73052 38948 73108 38958
rect 72716 38946 73108 38948
rect 72716 38894 72718 38946
rect 72770 38894 73054 38946
rect 73106 38894 73108 38946
rect 72716 38892 73108 38894
rect 72716 38882 72772 38892
rect 72604 38098 72660 38108
rect 72940 38164 72996 38174
rect 72940 38070 72996 38108
rect 72828 37940 72884 37950
rect 72828 37846 72884 37884
rect 72492 37828 72548 37838
rect 72716 37828 72772 37838
rect 73052 37828 73108 38892
rect 73164 38668 73220 39340
rect 73276 38946 73332 39676
rect 73500 39396 73556 67172
rect 73612 41972 73668 41982
rect 73612 41186 73668 41916
rect 73612 41134 73614 41186
rect 73666 41134 73668 41186
rect 73612 41122 73668 41134
rect 73612 40516 73668 40526
rect 73724 40516 73780 73948
rect 73836 45332 73892 75628
rect 74060 75460 74116 75470
rect 74060 75122 74116 75404
rect 74060 75070 74062 75122
rect 74114 75070 74116 75122
rect 74060 75058 74116 75070
rect 73836 45266 73892 45276
rect 74172 74788 74228 74798
rect 74060 41972 74116 41982
rect 74060 41878 74116 41916
rect 74172 41524 74228 74732
rect 74396 67228 74452 76526
rect 74508 76580 74564 76590
rect 74508 75794 74564 76524
rect 74508 75742 74510 75794
rect 74562 75742 74564 75794
rect 74508 75730 74564 75742
rect 74732 76578 74788 76590
rect 74732 76526 74734 76578
rect 74786 76526 74788 76578
rect 74508 75572 74564 75582
rect 74508 75122 74564 75516
rect 74508 75070 74510 75122
rect 74562 75070 74564 75122
rect 74508 75058 74564 75070
rect 74620 74116 74676 74126
rect 74396 67172 74564 67228
rect 74060 41468 74228 41524
rect 74396 41524 74452 41534
rect 73836 41076 73892 41086
rect 73836 40628 73892 41020
rect 73948 40628 74004 40638
rect 73836 40626 74004 40628
rect 73836 40574 73950 40626
rect 74002 40574 74004 40626
rect 73836 40572 74004 40574
rect 73948 40562 74004 40572
rect 73724 40460 73892 40516
rect 73612 40422 73668 40460
rect 73276 38894 73278 38946
rect 73330 38894 73332 38946
rect 73276 38882 73332 38894
rect 73388 39340 73556 39396
rect 73612 39618 73668 39630
rect 73612 39566 73614 39618
rect 73666 39566 73668 39618
rect 73164 38612 73332 38668
rect 73276 38276 73332 38612
rect 73388 38612 73444 39340
rect 73500 39060 73556 39070
rect 73612 39060 73668 39566
rect 73500 39058 73668 39060
rect 73500 39006 73502 39058
rect 73554 39006 73668 39058
rect 73500 39004 73668 39006
rect 73500 38994 73556 39004
rect 73724 38836 73780 38846
rect 73724 38742 73780 38780
rect 73836 38612 73892 40460
rect 73948 40404 74004 40414
rect 74060 40404 74116 41468
rect 74396 41410 74452 41468
rect 74396 41358 74398 41410
rect 74450 41358 74452 41410
rect 74396 41346 74452 41358
rect 74004 40348 74116 40404
rect 74172 41300 74228 41310
rect 73948 40338 74004 40348
rect 74060 40180 74116 40190
rect 74060 39618 74116 40124
rect 74172 39956 74228 41244
rect 74284 40516 74340 40526
rect 74284 40422 74340 40460
rect 74172 39900 74452 39956
rect 74060 39566 74062 39618
rect 74114 39566 74116 39618
rect 74060 39554 74116 39566
rect 74172 39620 74228 39630
rect 74172 38948 74228 39564
rect 74172 38834 74228 38892
rect 74172 38782 74174 38834
rect 74226 38782 74228 38834
rect 74172 38770 74228 38782
rect 74396 39058 74452 39900
rect 74396 39006 74398 39058
rect 74450 39006 74452 39058
rect 73836 38556 74004 38612
rect 73388 38546 73444 38556
rect 73276 38220 73892 38276
rect 73164 38164 73220 38174
rect 73164 38050 73220 38108
rect 73164 37998 73166 38050
rect 73218 37998 73220 38050
rect 73164 37986 73220 37998
rect 73276 38050 73332 38062
rect 73276 37998 73278 38050
rect 73330 37998 73332 38050
rect 72492 37826 72716 37828
rect 72492 37774 72494 37826
rect 72546 37774 72716 37826
rect 72492 37772 72716 37774
rect 72492 37762 72548 37772
rect 72380 37324 72548 37380
rect 72268 37286 72324 37324
rect 72492 37266 72548 37324
rect 72492 37214 72494 37266
rect 72546 37214 72548 37266
rect 72380 37156 72436 37166
rect 71484 35186 71540 35196
rect 71932 35252 72100 35308
rect 71036 34972 71204 35028
rect 71260 35028 71316 35038
rect 70924 34804 70980 34814
rect 70924 34710 70980 34748
rect 70812 34290 70868 34300
rect 70700 30482 70756 30492
rect 70700 30324 70756 30334
rect 70364 28590 70366 28642
rect 70418 28590 70420 28642
rect 70364 28578 70420 28590
rect 70588 28754 70644 28766
rect 70588 28702 70590 28754
rect 70642 28702 70644 28754
rect 70252 27806 70254 27858
rect 70306 27806 70308 27858
rect 70252 27794 70308 27806
rect 70140 27746 70196 27758
rect 70140 27694 70142 27746
rect 70194 27694 70196 27746
rect 70140 27412 70196 27694
rect 70140 27346 70196 27356
rect 70588 27188 70644 28702
rect 70700 28642 70756 30268
rect 70924 29314 70980 29326
rect 70924 29262 70926 29314
rect 70978 29262 70980 29314
rect 70924 29092 70980 29262
rect 70924 29026 70980 29036
rect 70700 28590 70702 28642
rect 70754 28590 70756 28642
rect 70700 28578 70756 28590
rect 70812 28866 70868 28878
rect 70812 28814 70814 28866
rect 70866 28814 70868 28866
rect 70812 28644 70868 28814
rect 70812 28578 70868 28588
rect 70700 27860 70756 27870
rect 70700 27766 70756 27804
rect 70924 27858 70980 27870
rect 70924 27806 70926 27858
rect 70978 27806 70980 27858
rect 70812 27746 70868 27758
rect 70812 27694 70814 27746
rect 70866 27694 70868 27746
rect 70252 27132 70644 27188
rect 70700 27524 70756 27534
rect 70252 25060 70308 27132
rect 70700 27074 70756 27468
rect 70700 27022 70702 27074
rect 70754 27022 70756 27074
rect 70700 27010 70756 27022
rect 70588 26962 70644 26974
rect 70588 26910 70590 26962
rect 70642 26910 70644 26962
rect 70476 26852 70532 26862
rect 70252 24994 70308 25004
rect 70364 26850 70532 26852
rect 70364 26798 70478 26850
rect 70530 26798 70532 26850
rect 70364 26796 70532 26798
rect 70364 24388 70420 26796
rect 70476 26786 70532 26796
rect 70476 25396 70532 25406
rect 70476 25302 70532 25340
rect 70476 24388 70532 24398
rect 70364 24332 70476 24388
rect 70476 24322 70532 24332
rect 70588 23828 70644 26910
rect 70812 25844 70868 27694
rect 70924 26292 70980 27806
rect 71036 27074 71092 34972
rect 71260 34914 71316 34972
rect 71932 35028 71988 35252
rect 71932 34962 71988 34972
rect 71260 34862 71262 34914
rect 71314 34862 71316 34914
rect 71260 34850 71316 34862
rect 71596 34916 71652 34926
rect 71596 34822 71652 34860
rect 71820 34916 71876 34926
rect 71820 34822 71876 34860
rect 71372 34690 71428 34702
rect 71372 34638 71374 34690
rect 71426 34638 71428 34690
rect 71372 34468 71428 34638
rect 71932 34692 71988 34702
rect 71932 34598 71988 34636
rect 71372 34412 71540 34468
rect 71260 34356 71316 34366
rect 71260 34020 71316 34300
rect 71372 34244 71428 34254
rect 71372 34150 71428 34188
rect 71260 33964 71428 34020
rect 71372 32674 71428 33964
rect 71372 32622 71374 32674
rect 71426 32622 71428 32674
rect 71260 32564 71316 32574
rect 71260 32470 71316 32508
rect 71372 31892 71428 32622
rect 71372 31826 71428 31836
rect 71372 30996 71428 31006
rect 71372 30660 71428 30940
rect 71484 30772 71540 34412
rect 71820 34356 71876 34366
rect 72044 34356 72100 35252
rect 72268 37154 72436 37156
rect 72268 37102 72382 37154
rect 72434 37102 72436 37154
rect 72268 37100 72436 37102
rect 72156 35028 72212 35038
rect 72156 34914 72212 34972
rect 72156 34862 72158 34914
rect 72210 34862 72212 34914
rect 72156 34850 72212 34862
rect 72268 34692 72324 37100
rect 72380 37090 72436 37100
rect 72492 36706 72548 37214
rect 72716 37266 72772 37772
rect 72940 37772 73108 37828
rect 73164 37828 73220 37838
rect 73276 37828 73332 37998
rect 73724 37938 73780 37950
rect 73724 37886 73726 37938
rect 73778 37886 73780 37938
rect 73220 37772 73332 37828
rect 73612 37828 73668 37838
rect 73724 37828 73780 37886
rect 73668 37772 73780 37828
rect 72940 37716 72996 37772
rect 73164 37762 73220 37772
rect 72716 37214 72718 37266
rect 72770 37214 72772 37266
rect 72716 37202 72772 37214
rect 72828 37660 72996 37716
rect 72492 36654 72494 36706
rect 72546 36654 72548 36706
rect 72492 36642 72548 36654
rect 72604 37156 72660 37166
rect 72492 36484 72548 36494
rect 72492 36390 72548 36428
rect 72604 35924 72660 37100
rect 72828 37044 72884 37660
rect 73052 37380 73108 37390
rect 73052 37266 73108 37324
rect 73052 37214 73054 37266
rect 73106 37214 73108 37266
rect 73052 37202 73108 37214
rect 73388 37380 73444 37390
rect 73388 37266 73444 37324
rect 73388 37214 73390 37266
rect 73442 37214 73444 37266
rect 73276 37156 73332 37166
rect 73276 37062 73332 37100
rect 72492 35868 72660 35924
rect 72716 36988 72884 37044
rect 72268 34626 72324 34636
rect 72380 34804 72436 34814
rect 72380 34356 72436 34748
rect 72492 34580 72548 35868
rect 72604 35698 72660 35710
rect 72604 35646 72606 35698
rect 72658 35646 72660 35698
rect 72604 35588 72660 35646
rect 72604 35522 72660 35532
rect 72492 34524 72660 34580
rect 72492 34356 72548 34366
rect 71820 34354 72100 34356
rect 71820 34302 71822 34354
rect 71874 34302 72100 34354
rect 71820 34300 72100 34302
rect 72156 34354 72548 34356
rect 72156 34302 72494 34354
rect 72546 34302 72548 34354
rect 72156 34300 72548 34302
rect 71820 34290 71876 34300
rect 72044 33460 72100 33470
rect 71708 33292 71988 33348
rect 71708 33234 71764 33292
rect 71708 33182 71710 33234
rect 71762 33182 71764 33234
rect 71708 32562 71764 33182
rect 71708 32510 71710 32562
rect 71762 32510 71764 32562
rect 71596 32452 71652 32462
rect 71596 32358 71652 32396
rect 71708 30996 71764 32510
rect 71708 30930 71764 30940
rect 71820 33122 71876 33134
rect 71820 33070 71822 33122
rect 71874 33070 71876 33122
rect 71484 30716 71652 30772
rect 71372 30604 71540 30660
rect 71372 30212 71428 30222
rect 71148 29988 71204 29998
rect 71148 29894 71204 29932
rect 71372 29650 71428 30156
rect 71484 30098 71540 30604
rect 71484 30046 71486 30098
rect 71538 30046 71540 30098
rect 71484 30034 71540 30046
rect 71372 29598 71374 29650
rect 71426 29598 71428 29650
rect 71372 29586 71428 29598
rect 71036 27022 71038 27074
rect 71090 27022 71092 27074
rect 71036 27010 71092 27022
rect 71484 28532 71540 28542
rect 71484 27746 71540 28476
rect 71484 27694 71486 27746
rect 71538 27694 71540 27746
rect 71484 26740 71540 27694
rect 70924 26226 70980 26236
rect 71148 26684 71540 26740
rect 70588 23762 70644 23772
rect 70700 25788 70868 25844
rect 70700 22932 70756 25788
rect 70924 25508 70980 25518
rect 71036 25508 71092 25518
rect 70980 25506 71092 25508
rect 70980 25454 71038 25506
rect 71090 25454 71092 25506
rect 70980 25452 71092 25454
rect 70924 25414 70980 25452
rect 71036 25442 71092 25452
rect 71036 25060 71092 25070
rect 71036 23716 71092 25004
rect 71036 23650 71092 23660
rect 70700 22866 70756 22876
rect 71036 22932 71092 22942
rect 69468 22306 69524 22316
rect 68012 21522 68068 21532
rect 70252 22260 70308 22270
rect 67116 18946 67172 18956
rect 68572 18900 68628 18910
rect 65916 18060 66180 18070
rect 65972 18004 66020 18060
rect 66076 18004 66124 18060
rect 65916 17994 66180 18004
rect 65916 16492 66180 16502
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 65916 16426 66180 16436
rect 65916 14924 66180 14934
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 65916 14858 66180 14868
rect 65916 13356 66180 13366
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 65916 13290 66180 13300
rect 65916 11788 66180 11798
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 65916 11722 66180 11732
rect 67452 11284 67508 11294
rect 65916 10220 66180 10230
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 65916 10154 66180 10164
rect 64764 9762 64820 9772
rect 67116 9268 67172 9278
rect 65916 8652 66180 8662
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 65916 8586 66180 8596
rect 66668 7588 66724 7598
rect 66724 7532 67060 7588
rect 66668 7494 66724 7532
rect 67004 7474 67060 7532
rect 67004 7422 67006 7474
rect 67058 7422 67060 7474
rect 67004 7410 67060 7422
rect 65916 7084 66180 7094
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 65916 7018 66180 7028
rect 67116 5908 67172 9212
rect 67340 6466 67396 6478
rect 67340 6414 67342 6466
rect 67394 6414 67396 6466
rect 67340 6244 67396 6414
rect 67340 6178 67396 6188
rect 67340 5908 67396 5918
rect 67116 5906 67396 5908
rect 67116 5854 67342 5906
rect 67394 5854 67396 5906
rect 67116 5852 67396 5854
rect 64652 5170 64708 5180
rect 65548 5794 65604 5806
rect 65548 5742 65550 5794
rect 65602 5742 65604 5794
rect 65548 5124 65604 5742
rect 65916 5516 66180 5526
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 65916 5450 66180 5460
rect 65548 5058 65604 5068
rect 66332 5348 66388 5358
rect 64540 4246 64596 4284
rect 65660 4340 65716 4350
rect 65548 4226 65604 4238
rect 65548 4174 65550 4226
rect 65602 4174 65604 4226
rect 64092 4116 64148 4126
rect 63868 3666 63924 3678
rect 63868 3614 63870 3666
rect 63922 3614 63924 3666
rect 63868 3444 63924 3614
rect 63868 3378 63924 3388
rect 63420 924 63700 980
rect 63420 800 63476 924
rect 64092 800 64148 4060
rect 65548 3892 65604 4174
rect 65548 3826 65604 3836
rect 65660 3666 65716 4284
rect 65916 3948 66180 3958
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 65916 3882 66180 3892
rect 65660 3614 65662 3666
rect 65714 3614 65716 3666
rect 65660 3602 65716 3614
rect 65436 3556 65492 3566
rect 64764 3444 64820 3454
rect 64764 800 64820 3388
rect 65436 800 65492 3500
rect 66332 2660 66388 5292
rect 66444 5236 66500 5246
rect 66444 3554 66500 5180
rect 67116 5234 67172 5852
rect 67340 5842 67396 5852
rect 67116 5182 67118 5234
rect 67170 5182 67172 5234
rect 67116 5170 67172 5182
rect 67452 5234 67508 11228
rect 68012 7252 68068 7262
rect 67788 7250 68068 7252
rect 67788 7198 68014 7250
rect 68066 7198 68068 7250
rect 67788 7196 68068 7198
rect 67452 5182 67454 5234
rect 67506 5182 67508 5234
rect 66444 3502 66446 3554
rect 66498 3502 66500 3554
rect 66444 3490 66500 3502
rect 66780 5124 66836 5134
rect 66108 2604 66388 2660
rect 66108 800 66164 2604
rect 66780 800 66836 5068
rect 67452 4338 67508 5182
rect 67452 4286 67454 4338
rect 67506 4286 67508 4338
rect 67452 4274 67508 4286
rect 67564 6468 67620 6478
rect 67452 3780 67508 3790
rect 67452 3686 67508 3724
rect 67564 3220 67620 6412
rect 67788 5124 67844 7196
rect 68012 7186 68068 7196
rect 67900 6692 67956 6702
rect 68348 6692 68404 6702
rect 67900 6690 68404 6692
rect 67900 6638 67902 6690
rect 67954 6638 68350 6690
rect 68402 6638 68404 6690
rect 67900 6636 68404 6638
rect 67900 6356 67956 6636
rect 68348 6626 68404 6636
rect 67900 6290 67956 6300
rect 68460 6244 68516 6254
rect 67788 5058 67844 5068
rect 68124 5236 68180 5246
rect 67452 3164 67620 3220
rect 67452 800 67508 3164
rect 68124 800 68180 5180
rect 68460 5122 68516 6188
rect 68572 6132 68628 18844
rect 70252 16212 70308 22204
rect 70476 20692 70532 20702
rect 70476 19460 70532 20636
rect 70476 19394 70532 19404
rect 70924 18450 70980 18462
rect 70924 18398 70926 18450
rect 70978 18398 70980 18450
rect 70588 18340 70644 18350
rect 70924 18340 70980 18398
rect 70588 18338 70980 18340
rect 70588 18286 70590 18338
rect 70642 18286 70980 18338
rect 70588 18284 70980 18286
rect 70588 17892 70644 18284
rect 70588 17826 70644 17836
rect 71036 16324 71092 22876
rect 71148 18676 71204 26684
rect 71372 26178 71428 26190
rect 71372 26126 71374 26178
rect 71426 26126 71428 26178
rect 71372 25844 71428 26126
rect 71372 25778 71428 25788
rect 71260 25732 71316 25742
rect 71260 25638 71316 25676
rect 71596 25284 71652 30716
rect 71820 30212 71876 33070
rect 71932 32788 71988 33292
rect 72044 33346 72100 33404
rect 72044 33294 72046 33346
rect 72098 33294 72100 33346
rect 72044 33282 72100 33294
rect 72156 33346 72212 34300
rect 72492 34290 72548 34300
rect 72604 33684 72660 34524
rect 72716 34132 72772 36988
rect 73388 36932 73444 37214
rect 73612 37266 73668 37772
rect 73612 37214 73614 37266
rect 73666 37214 73668 37266
rect 73612 37202 73668 37214
rect 73724 37268 73780 37278
rect 73164 36876 73444 36932
rect 72940 36820 72996 36830
rect 72828 36764 72940 36820
rect 72828 35308 72884 36764
rect 72940 36754 72996 36764
rect 72940 36596 72996 36606
rect 73164 36596 73220 36876
rect 72940 36594 73220 36596
rect 72940 36542 72942 36594
rect 72994 36542 73220 36594
rect 72940 36540 73220 36542
rect 73276 36706 73332 36718
rect 73276 36654 73278 36706
rect 73330 36654 73332 36706
rect 73276 36594 73332 36654
rect 73276 36542 73278 36594
rect 73330 36542 73332 36594
rect 72940 36530 72996 36540
rect 73276 36530 73332 36542
rect 72940 35980 73444 36036
rect 72940 35922 72996 35980
rect 72940 35870 72942 35922
rect 72994 35870 72996 35922
rect 72940 35858 72996 35870
rect 73276 35810 73332 35822
rect 73276 35758 73278 35810
rect 73330 35758 73332 35810
rect 72828 35252 72996 35308
rect 72940 35140 72996 35252
rect 72940 35074 72996 35084
rect 72828 34914 72884 34926
rect 72828 34862 72830 34914
rect 72882 34862 72884 34914
rect 72828 34804 72884 34862
rect 73052 34916 73108 34926
rect 73276 34916 73332 35758
rect 73388 35812 73444 35980
rect 73612 35812 73668 35822
rect 73724 35812 73780 37212
rect 73388 35810 73780 35812
rect 73388 35758 73614 35810
rect 73666 35758 73780 35810
rect 73388 35756 73780 35758
rect 73612 35746 73668 35756
rect 73724 35364 73780 35374
rect 73612 35308 73724 35364
rect 73052 34914 73220 34916
rect 73052 34862 73054 34914
rect 73106 34862 73220 34914
rect 73052 34860 73220 34862
rect 73052 34850 73108 34860
rect 72828 34738 72884 34748
rect 73052 34692 73108 34702
rect 72940 34690 73108 34692
rect 72940 34638 73054 34690
rect 73106 34638 73108 34690
rect 72940 34636 73108 34638
rect 73164 34692 73220 34860
rect 73276 34822 73332 34860
rect 73500 34916 73556 34954
rect 73500 34850 73556 34860
rect 73388 34692 73444 34702
rect 73164 34636 73332 34692
rect 72940 34468 72996 34636
rect 73052 34626 73108 34636
rect 72940 34402 72996 34412
rect 73276 34356 73332 34636
rect 73276 34290 73332 34300
rect 73388 34354 73444 34636
rect 73388 34302 73390 34354
rect 73442 34302 73444 34354
rect 73388 34290 73444 34302
rect 73052 34132 73108 34142
rect 72716 34130 73108 34132
rect 72716 34078 72718 34130
rect 72770 34078 73054 34130
rect 73106 34078 73108 34130
rect 72716 34076 73108 34078
rect 72716 34066 72772 34076
rect 73052 34066 73108 34076
rect 73388 34132 73444 34142
rect 73612 34132 73668 35308
rect 73724 35298 73780 35308
rect 73836 34914 73892 38220
rect 73948 37938 74004 38556
rect 74284 38052 74340 38062
rect 74284 37958 74340 37996
rect 73948 37886 73950 37938
rect 74002 37886 74004 37938
rect 73948 37492 74004 37886
rect 73948 37426 74004 37436
rect 74060 37826 74116 37838
rect 74060 37774 74062 37826
rect 74114 37774 74116 37826
rect 73948 36372 74004 36382
rect 73948 36278 74004 36316
rect 73836 34862 73838 34914
rect 73890 34862 73892 34914
rect 73836 34850 73892 34862
rect 73948 35812 74004 35822
rect 73948 35698 74004 35756
rect 73948 35646 73950 35698
rect 74002 35646 74004 35698
rect 73948 34916 74004 35646
rect 74060 35364 74116 37774
rect 74284 37266 74340 37278
rect 74284 37214 74286 37266
rect 74338 37214 74340 37266
rect 74284 37044 74340 37214
rect 74284 36978 74340 36988
rect 74284 36820 74340 36830
rect 74172 36764 74284 36820
rect 74172 35810 74228 36764
rect 74284 36754 74340 36764
rect 74396 36596 74452 39006
rect 74508 39060 74564 67172
rect 74620 40852 74676 74060
rect 74732 74004 74788 76526
rect 74956 76580 75012 76590
rect 74956 76466 75012 76524
rect 74956 76414 74958 76466
rect 75010 76414 75012 76466
rect 74956 76402 75012 76414
rect 74732 73938 74788 73948
rect 74844 75796 74900 75806
rect 74844 50428 74900 75740
rect 75068 75794 75124 76974
rect 75740 77026 75796 77038
rect 75740 76974 75742 77026
rect 75794 76974 75796 77026
rect 75404 76804 75460 76814
rect 75404 76690 75460 76748
rect 75404 76638 75406 76690
rect 75458 76638 75460 76690
rect 75404 76626 75460 76638
rect 75740 76578 75796 76974
rect 75740 76526 75742 76578
rect 75794 76526 75796 76578
rect 75740 76514 75796 76526
rect 75068 75742 75070 75794
rect 75122 75742 75124 75794
rect 75068 75730 75124 75742
rect 75404 75908 75460 75918
rect 75404 75682 75460 75852
rect 75404 75630 75406 75682
rect 75458 75630 75460 75682
rect 75404 75618 75460 75630
rect 75628 75684 75684 75694
rect 75628 75570 75684 75628
rect 75628 75518 75630 75570
rect 75682 75518 75684 75570
rect 75628 75506 75684 75518
rect 75404 75236 75460 75246
rect 74956 75124 75012 75134
rect 74956 75030 75012 75068
rect 75404 75122 75460 75180
rect 75404 75070 75406 75122
rect 75458 75070 75460 75122
rect 75404 75058 75460 75070
rect 75628 75010 75684 75022
rect 75628 74958 75630 75010
rect 75682 74958 75684 75010
rect 75292 74228 75348 74238
rect 75292 74134 75348 74172
rect 75628 61348 75684 74958
rect 75740 74228 75796 74238
rect 75852 74228 75908 77198
rect 76076 76580 76132 76590
rect 76076 76486 76132 76524
rect 76188 75682 76244 77420
rect 76412 77250 76468 77262
rect 76412 77198 76414 77250
rect 76466 77198 76468 77250
rect 76412 76690 76468 77198
rect 76412 76638 76414 76690
rect 76466 76638 76468 76690
rect 76412 76626 76468 76638
rect 76636 77026 76692 77038
rect 76636 76974 76638 77026
rect 76690 76974 76692 77026
rect 76188 75630 76190 75682
rect 76242 75630 76244 75682
rect 76076 75348 76132 75358
rect 75964 75236 76020 75246
rect 75964 75010 76020 75180
rect 75964 74958 75966 75010
rect 76018 74958 76020 75010
rect 75964 74946 76020 74958
rect 75740 74226 75908 74228
rect 75740 74174 75742 74226
rect 75794 74174 75908 74226
rect 75740 74172 75908 74174
rect 75740 74162 75796 74172
rect 76076 73554 76132 75292
rect 76188 75124 76244 75630
rect 76188 75058 76244 75068
rect 76412 75908 76468 75918
rect 76300 74788 76356 74798
rect 76300 74694 76356 74732
rect 76412 74226 76468 75852
rect 76524 75796 76580 75806
rect 76524 75570 76580 75740
rect 76524 75518 76526 75570
rect 76578 75518 76580 75570
rect 76524 75506 76580 75518
rect 76412 74174 76414 74226
rect 76466 74174 76468 74226
rect 76412 74162 76468 74174
rect 76524 74788 76580 74798
rect 76076 73502 76078 73554
rect 76130 73502 76132 73554
rect 76076 73490 76132 73502
rect 76524 73554 76580 74732
rect 76524 73502 76526 73554
rect 76578 73502 76580 73554
rect 76524 73490 76580 73502
rect 76636 73106 76692 76974
rect 76748 76356 76804 76366
rect 76748 76262 76804 76300
rect 76860 75682 76916 77420
rect 76860 75630 76862 75682
rect 76914 75630 76916 75682
rect 76860 75572 76916 75630
rect 76860 75506 76916 75516
rect 76972 76916 77028 76926
rect 76860 75124 76916 75134
rect 76972 75124 77028 76860
rect 77084 75348 77140 79200
rect 77196 79044 77252 79054
rect 77196 77026 77252 78988
rect 77196 76974 77198 77026
rect 77250 76974 77252 77026
rect 77196 76466 77252 76974
rect 77756 76580 77812 79200
rect 77196 76414 77198 76466
rect 77250 76414 77252 76466
rect 77196 76402 77252 76414
rect 77420 76524 77812 76580
rect 77980 78036 78036 78046
rect 77084 75282 77140 75292
rect 77196 75458 77252 75470
rect 77196 75406 77198 75458
rect 77250 75406 77252 75458
rect 77196 75124 77252 75406
rect 76860 75122 77028 75124
rect 76860 75070 76862 75122
rect 76914 75070 77028 75122
rect 76860 75068 77028 75070
rect 77084 75068 77252 75124
rect 76860 73556 76916 75068
rect 76972 74116 77028 74126
rect 76972 74022 77028 74060
rect 76972 73556 77028 73566
rect 76860 73554 77028 73556
rect 76860 73502 76974 73554
rect 77026 73502 77028 73554
rect 76860 73500 77028 73502
rect 76972 73490 77028 73500
rect 76636 73054 76638 73106
rect 76690 73054 76692 73106
rect 76636 73042 76692 73054
rect 75068 61292 75684 61348
rect 76412 72548 76468 72558
rect 74844 50372 75012 50428
rect 74956 42196 75012 50372
rect 74956 42130 75012 42140
rect 74956 41972 75012 41982
rect 74844 41970 75012 41972
rect 74844 41918 74958 41970
rect 75010 41918 75012 41970
rect 74844 41916 75012 41918
rect 74732 41858 74788 41870
rect 74732 41806 74734 41858
rect 74786 41806 74788 41858
rect 74732 41636 74788 41806
rect 74732 41570 74788 41580
rect 74732 41412 74788 41422
rect 74844 41412 74900 41916
rect 74956 41906 75012 41916
rect 75068 41972 75124 61292
rect 75852 59108 75908 59118
rect 75740 45332 75796 45342
rect 75740 42866 75796 45276
rect 75740 42814 75742 42866
rect 75794 42814 75796 42866
rect 75740 42644 75796 42814
rect 75740 42578 75796 42588
rect 75292 42532 75348 42542
rect 75068 41906 75124 41916
rect 75180 42476 75292 42532
rect 74732 41410 74900 41412
rect 74732 41358 74734 41410
rect 74786 41358 74900 41410
rect 74732 41356 74900 41358
rect 75068 41636 75124 41646
rect 74732 41346 74788 41356
rect 75068 41298 75124 41580
rect 75068 41246 75070 41298
rect 75122 41246 75124 41298
rect 75068 41234 75124 41246
rect 74620 40796 74788 40852
rect 74620 40628 74676 40638
rect 74620 40534 74676 40572
rect 74620 39732 74676 39742
rect 74732 39732 74788 40796
rect 75068 40740 75124 40750
rect 75068 40404 75124 40684
rect 75180 40626 75236 42476
rect 75292 42466 75348 42476
rect 75292 42082 75348 42094
rect 75292 42030 75294 42082
rect 75346 42030 75348 42082
rect 75292 41972 75348 42030
rect 75628 41972 75684 41982
rect 75292 41970 75684 41972
rect 75292 41918 75630 41970
rect 75682 41918 75684 41970
rect 75292 41916 75684 41918
rect 75628 41906 75684 41916
rect 75292 41300 75348 41310
rect 75292 41206 75348 41244
rect 75180 40574 75182 40626
rect 75234 40574 75236 40626
rect 75180 40562 75236 40574
rect 75628 40962 75684 40974
rect 75628 40910 75630 40962
rect 75682 40910 75684 40962
rect 75292 40404 75348 40414
rect 75068 40348 75236 40404
rect 74676 39676 74788 39732
rect 74956 40178 75012 40190
rect 74956 40126 74958 40178
rect 75010 40126 75012 40178
rect 74620 39638 74676 39676
rect 74956 39508 75012 40126
rect 75068 39620 75124 39630
rect 75068 39526 75124 39564
rect 74508 38994 74564 39004
rect 74620 39452 75012 39508
rect 74620 38668 74676 39452
rect 75068 39396 75124 39406
rect 74508 38612 74676 38668
rect 74844 38834 74900 38846
rect 74844 38782 74846 38834
rect 74898 38782 74900 38834
rect 74844 38724 74900 38782
rect 74844 38658 74900 38668
rect 74508 37604 74564 38612
rect 74620 38052 74676 38062
rect 74676 37996 74900 38052
rect 74620 37958 74676 37996
rect 74732 37826 74788 37838
rect 74732 37774 74734 37826
rect 74786 37774 74788 37826
rect 74508 37548 74676 37604
rect 74284 36540 74452 36596
rect 74508 37378 74564 37390
rect 74508 37326 74510 37378
rect 74562 37326 74564 37378
rect 74284 36036 74340 36540
rect 74508 36484 74564 37326
rect 74620 36932 74676 37548
rect 74620 36866 74676 36876
rect 74620 36484 74676 36494
rect 74508 36482 74676 36484
rect 74508 36430 74622 36482
rect 74674 36430 74676 36482
rect 74508 36428 74676 36430
rect 74620 36418 74676 36428
rect 74396 36372 74452 36382
rect 74396 36278 74452 36316
rect 74284 35980 74564 36036
rect 74172 35758 74174 35810
rect 74226 35758 74228 35810
rect 74172 35746 74228 35758
rect 74508 35810 74564 35980
rect 74732 35924 74788 37774
rect 74844 37378 74900 37996
rect 75068 38050 75124 39340
rect 75180 39172 75236 40348
rect 75348 40348 75460 40404
rect 75292 40338 75348 40348
rect 75292 40180 75348 40190
rect 75292 40086 75348 40124
rect 75292 39620 75348 39630
rect 75292 39394 75348 39564
rect 75404 39618 75460 40348
rect 75628 40180 75684 40910
rect 75852 40404 75908 59052
rect 76412 50428 76468 72492
rect 77084 68852 77140 75068
rect 77308 74900 77364 74910
rect 77420 74900 77476 76524
rect 77868 76468 77924 76478
rect 77756 76466 77924 76468
rect 77756 76414 77870 76466
rect 77922 76414 77924 76466
rect 77756 76412 77924 76414
rect 77756 75348 77812 76412
rect 77868 76402 77924 76412
rect 77868 76020 77924 76030
rect 77868 75570 77924 75964
rect 77868 75518 77870 75570
rect 77922 75518 77924 75570
rect 77868 75506 77924 75518
rect 77756 75282 77812 75292
rect 77532 75012 77588 75022
rect 77532 74918 77588 74956
rect 77868 75010 77924 75022
rect 77868 74958 77870 75010
rect 77922 74958 77924 75010
rect 77308 74898 77476 74900
rect 77308 74846 77310 74898
rect 77362 74846 77476 74898
rect 77308 74844 77476 74846
rect 77308 74788 77364 74844
rect 77308 74722 77364 74732
rect 77756 74340 77812 74350
rect 77532 74338 77812 74340
rect 77532 74286 77758 74338
rect 77810 74286 77812 74338
rect 77532 74284 77812 74286
rect 77532 74114 77588 74284
rect 77756 74274 77812 74284
rect 77532 74062 77534 74114
rect 77586 74062 77588 74114
rect 77532 74050 77588 74062
rect 77420 73556 77476 73566
rect 77420 73462 77476 73500
rect 77644 73220 77700 73230
rect 77644 73126 77700 73164
rect 77196 73106 77252 73118
rect 77196 73054 77198 73106
rect 77250 73054 77252 73106
rect 77196 72658 77252 73054
rect 77196 72606 77198 72658
rect 77250 72606 77252 72658
rect 77196 72594 77252 72606
rect 77868 72548 77924 74958
rect 77980 74338 78036 77980
rect 78204 76578 78260 76590
rect 78204 76526 78206 76578
rect 78258 76526 78260 76578
rect 78204 76132 78260 76526
rect 78204 76066 78260 76076
rect 78092 75684 78148 75694
rect 78092 75460 78148 75628
rect 78428 75572 78484 79200
rect 78428 75506 78484 75516
rect 78092 75394 78148 75404
rect 79100 75236 79156 79200
rect 79100 75170 79156 75180
rect 77980 74286 77982 74338
rect 78034 74286 78036 74338
rect 77980 74226 78036 74286
rect 77980 74174 77982 74226
rect 78034 74174 78036 74226
rect 77980 74162 78036 74174
rect 78092 74898 78148 74910
rect 78092 74846 78094 74898
rect 78146 74846 78148 74898
rect 78092 74676 78148 74846
rect 78092 74228 78148 74620
rect 78092 74162 78148 74172
rect 78204 73556 78260 73566
rect 78204 73462 78260 73500
rect 77868 72482 77924 72492
rect 77644 72436 77700 72446
rect 77644 72342 77700 72380
rect 78204 72436 78260 72446
rect 78204 72342 78260 72380
rect 77868 72324 77924 72334
rect 77868 72322 78148 72324
rect 77868 72270 77870 72322
rect 77922 72270 78148 72322
rect 77868 72268 78148 72270
rect 77868 72258 77924 72268
rect 77868 71876 77924 71886
rect 77868 71782 77924 71820
rect 77644 71764 77700 71774
rect 77644 71670 77700 71708
rect 77756 71092 77812 71102
rect 77756 70998 77812 71036
rect 77420 70756 77476 70766
rect 77420 70662 77476 70700
rect 77644 69186 77700 69198
rect 77868 69188 77924 69198
rect 77644 69134 77646 69186
rect 77698 69134 77700 69186
rect 77644 69076 77700 69134
rect 77644 69010 77700 69020
rect 77756 69186 77924 69188
rect 77756 69134 77870 69186
rect 77922 69134 77924 69186
rect 77756 69132 77924 69134
rect 77084 68786 77140 68796
rect 77420 68516 77476 68526
rect 77420 68422 77476 68460
rect 77644 68514 77700 68526
rect 77644 68462 77646 68514
rect 77698 68462 77700 68514
rect 77644 67844 77700 68462
rect 77644 67778 77700 67788
rect 77644 66946 77700 66958
rect 77644 66894 77646 66946
rect 77698 66894 77700 66946
rect 77644 66836 77700 66894
rect 77644 66770 77700 66780
rect 77644 66276 77700 66286
rect 77644 66182 77700 66220
rect 77420 66050 77476 66062
rect 77420 65998 77422 66050
rect 77474 65998 77476 66050
rect 77420 65716 77476 65998
rect 77420 65650 77476 65660
rect 77644 64708 77700 64718
rect 77644 64614 77700 64652
rect 77420 64596 77476 64606
rect 77420 64502 77476 64540
rect 77644 63924 77700 63934
rect 77644 63830 77700 63868
rect 77644 63140 77700 63150
rect 76972 63138 77700 63140
rect 76972 63086 77646 63138
rect 77698 63086 77700 63138
rect 76972 63084 77700 63086
rect 76972 50428 77028 63084
rect 77644 63074 77700 63084
rect 77420 62916 77476 62926
rect 77420 62822 77476 62860
rect 77644 61346 77700 61358
rect 77644 61294 77646 61346
rect 77698 61294 77700 61346
rect 77644 61236 77700 61294
rect 77644 61170 77700 61180
rect 77644 60788 77700 60798
rect 77644 60694 77700 60732
rect 77420 59106 77476 59118
rect 77420 59054 77422 59106
rect 77474 59054 77476 59106
rect 77420 58996 77476 59054
rect 77644 59108 77700 59118
rect 77644 59014 77700 59052
rect 77420 58930 77476 58940
rect 77644 58210 77700 58222
rect 77644 58158 77646 58210
rect 77698 58158 77700 58210
rect 77644 57876 77700 58158
rect 77644 57810 77700 57820
rect 77644 56756 77700 56766
rect 77644 56662 77700 56700
rect 77420 55970 77476 55982
rect 77420 55918 77422 55970
rect 77474 55918 77476 55970
rect 77420 55636 77476 55918
rect 77644 55972 77700 55982
rect 77644 55878 77700 55916
rect 77420 55570 77476 55580
rect 77756 55468 77812 69132
rect 77868 69122 77924 69132
rect 78092 67228 78148 72268
rect 78540 71876 78596 71886
rect 78596 71820 78820 71876
rect 78540 71810 78596 71820
rect 78204 71764 78260 71774
rect 78204 71316 78260 71708
rect 78204 71250 78260 71260
rect 78204 70756 78260 70766
rect 78204 70196 78260 70700
rect 78204 70130 78260 70140
rect 78204 69186 78260 69198
rect 78204 69134 78206 69186
rect 78258 69134 78260 69186
rect 78204 69076 78260 69134
rect 78204 69010 78260 69020
rect 78204 68626 78260 68638
rect 78204 68574 78206 68626
rect 78258 68574 78260 68626
rect 78204 68516 78260 68574
rect 78204 67956 78260 68460
rect 78204 67890 78260 67900
rect 77868 67172 77924 67182
rect 78092 67172 78708 67228
rect 77868 67078 77924 67116
rect 78204 67058 78260 67070
rect 78204 67006 78206 67058
rect 78258 67006 78260 67058
rect 78204 66836 78260 67006
rect 78204 66770 78260 66780
rect 78204 66050 78260 66062
rect 78204 65998 78206 66050
rect 78258 65998 78260 66050
rect 78204 65716 78260 65998
rect 78204 65650 78260 65660
rect 78204 64596 78260 64606
rect 78204 64502 78260 64540
rect 77868 64034 77924 64046
rect 77868 63982 77870 64034
rect 77922 63982 77924 64034
rect 77868 62244 77924 63982
rect 78204 63924 78260 63934
rect 78204 63476 78260 63868
rect 78204 63410 78260 63420
rect 78204 62916 78260 62926
rect 78204 62356 78260 62860
rect 78204 62290 78260 62300
rect 77868 62178 77924 62188
rect 77868 61348 77924 61358
rect 77868 61254 77924 61292
rect 78204 61346 78260 61358
rect 78204 61294 78206 61346
rect 78258 61294 78260 61346
rect 78204 61236 78260 61294
rect 78204 61170 78260 61180
rect 77868 60900 77924 60910
rect 77868 60898 78148 60900
rect 77868 60846 77870 60898
rect 77922 60846 78148 60898
rect 77868 60844 78148 60846
rect 77868 60834 77924 60844
rect 78092 58436 78148 60844
rect 78204 60788 78260 60798
rect 78204 60116 78260 60732
rect 78204 60050 78260 60060
rect 78204 59218 78260 59230
rect 78204 59166 78206 59218
rect 78258 59166 78260 59218
rect 78204 58996 78260 59166
rect 78204 58930 78260 58940
rect 78092 58380 78596 58436
rect 77868 58212 77924 58222
rect 77868 58118 77924 58156
rect 78204 58210 78260 58222
rect 78204 58158 78206 58210
rect 78258 58158 78260 58210
rect 78204 57876 78260 58158
rect 78204 57810 78260 57820
rect 78204 56756 78260 56766
rect 78204 56662 78260 56700
rect 77868 56644 77924 56654
rect 77868 56550 77924 56588
rect 78204 56082 78260 56094
rect 78204 56030 78206 56082
rect 78258 56030 78260 56082
rect 78204 55636 78260 56030
rect 78204 55570 78260 55580
rect 77756 55412 78484 55468
rect 77644 55188 77700 55198
rect 77644 55094 77700 55132
rect 78204 55188 78260 55198
rect 77868 55076 77924 55086
rect 77868 54982 77924 55020
rect 78204 54516 78260 55132
rect 78204 54450 78260 54460
rect 78204 53618 78260 53630
rect 78204 53566 78206 53618
rect 78258 53566 78260 53618
rect 77644 53506 77700 53518
rect 77868 53508 77924 53518
rect 77644 53454 77646 53506
rect 77698 53454 77700 53506
rect 77644 53396 77700 53454
rect 77644 53330 77700 53340
rect 77756 53506 77924 53508
rect 77756 53454 77870 53506
rect 77922 53454 77924 53506
rect 77756 53452 77924 53454
rect 77756 53060 77812 53452
rect 77868 53442 77924 53452
rect 78204 53396 78260 53566
rect 78204 53330 78260 53340
rect 76188 50372 76468 50428
rect 76860 50372 77028 50428
rect 77420 53004 77812 53060
rect 77868 53060 77924 53070
rect 76076 41412 76132 41422
rect 76076 41186 76132 41356
rect 76076 41134 76078 41186
rect 76130 41134 76132 41186
rect 76076 41122 76132 41134
rect 75628 40114 75684 40124
rect 75740 40348 75908 40404
rect 76188 40852 76244 50372
rect 76636 43314 76692 43326
rect 76636 43262 76638 43314
rect 76690 43262 76692 43314
rect 76524 42756 76580 42766
rect 76636 42756 76692 43262
rect 76412 42754 76692 42756
rect 76412 42702 76526 42754
rect 76578 42702 76692 42754
rect 76412 42700 76692 42702
rect 76300 42532 76356 42542
rect 76300 42438 76356 42476
rect 75404 39566 75406 39618
rect 75458 39566 75460 39618
rect 75404 39554 75460 39566
rect 75516 39618 75572 39630
rect 75516 39566 75518 39618
rect 75570 39566 75572 39618
rect 75292 39342 75294 39394
rect 75346 39342 75348 39394
rect 75292 39330 75348 39342
rect 75516 39284 75572 39566
rect 75404 39228 75572 39284
rect 75180 39116 75348 39172
rect 75180 38946 75236 38958
rect 75180 38894 75182 38946
rect 75234 38894 75236 38946
rect 75180 38724 75236 38894
rect 75180 38658 75236 38668
rect 75068 37998 75070 38050
rect 75122 37998 75124 38050
rect 74956 37940 75012 37950
rect 74956 37846 75012 37884
rect 75068 37828 75124 37998
rect 75068 37762 75124 37772
rect 74844 37326 74846 37378
rect 74898 37326 74900 37378
rect 74844 37314 74900 37326
rect 75068 37490 75124 37502
rect 75068 37438 75070 37490
rect 75122 37438 75124 37490
rect 74956 36932 75012 36942
rect 74844 36708 74900 36718
rect 74844 36594 74900 36652
rect 74956 36706 75012 36876
rect 74956 36654 74958 36706
rect 75010 36654 75012 36706
rect 74956 36642 75012 36654
rect 74844 36542 74846 36594
rect 74898 36542 74900 36594
rect 74844 36530 74900 36542
rect 74732 35868 74900 35924
rect 74508 35758 74510 35810
rect 74562 35758 74564 35810
rect 74508 35700 74564 35758
rect 74732 35700 74788 35710
rect 74508 35698 74788 35700
rect 74508 35646 74734 35698
rect 74786 35646 74788 35698
rect 74508 35644 74788 35646
rect 74732 35634 74788 35644
rect 74396 35588 74452 35598
rect 74396 35586 74564 35588
rect 74396 35534 74398 35586
rect 74450 35534 74564 35586
rect 74396 35532 74564 35534
rect 74396 35522 74452 35532
rect 74060 35298 74116 35308
rect 74172 35252 74228 35262
rect 74060 34916 74116 34926
rect 73948 34914 74116 34916
rect 73948 34862 74062 34914
rect 74114 34862 74116 34914
rect 73948 34860 74116 34862
rect 72604 33628 72996 33684
rect 72716 33460 72772 33470
rect 72716 33366 72772 33404
rect 72156 33294 72158 33346
rect 72210 33294 72212 33346
rect 72156 33282 72212 33294
rect 72604 33348 72660 33358
rect 71932 32732 72212 32788
rect 72156 32562 72212 32732
rect 72380 32676 72436 32686
rect 72436 32620 72548 32676
rect 72380 32610 72436 32620
rect 72156 32510 72158 32562
rect 72210 32510 72212 32562
rect 72156 32498 72212 32510
rect 72380 32452 72436 32462
rect 72380 32358 72436 32396
rect 71932 31892 71988 31902
rect 71988 31836 72100 31892
rect 71932 31826 71988 31836
rect 72044 31778 72100 31836
rect 72044 31726 72046 31778
rect 72098 31726 72100 31778
rect 72044 31714 72100 31726
rect 72268 30996 72324 31006
rect 72268 30902 72324 30940
rect 72044 30884 72100 30894
rect 71932 30772 71988 30782
rect 71932 30322 71988 30716
rect 71932 30270 71934 30322
rect 71986 30270 71988 30322
rect 71932 30258 71988 30270
rect 71708 30156 71876 30212
rect 72044 30210 72100 30828
rect 72044 30158 72046 30210
rect 72098 30158 72100 30210
rect 71708 25956 71764 30156
rect 72044 30146 72100 30158
rect 72380 30882 72436 30894
rect 72380 30830 72382 30882
rect 72434 30830 72436 30882
rect 71820 29988 71876 29998
rect 72156 29988 72212 29998
rect 71820 29986 71988 29988
rect 71820 29934 71822 29986
rect 71874 29934 71988 29986
rect 71820 29932 71988 29934
rect 71820 29922 71876 29932
rect 71820 29764 71876 29774
rect 71820 29650 71876 29708
rect 71820 29598 71822 29650
rect 71874 29598 71876 29650
rect 71820 29586 71876 29598
rect 71820 28532 71876 28570
rect 71820 28466 71876 28476
rect 71820 28308 71876 28318
rect 71820 27186 71876 28252
rect 71932 27860 71988 29932
rect 72156 29202 72212 29932
rect 72156 29150 72158 29202
rect 72210 29150 72212 29202
rect 72156 28530 72212 29150
rect 72156 28478 72158 28530
rect 72210 28478 72212 28530
rect 72156 28466 72212 28478
rect 71932 27794 71988 27804
rect 71820 27134 71822 27186
rect 71874 27134 71876 27186
rect 71820 27122 71876 27134
rect 72268 27188 72324 27198
rect 72268 27094 72324 27132
rect 71820 26180 71876 26190
rect 71820 26178 71988 26180
rect 71820 26126 71822 26178
rect 71874 26126 71988 26178
rect 71820 26124 71988 26126
rect 71820 26114 71876 26124
rect 71708 25900 71876 25956
rect 71820 25506 71876 25900
rect 71820 25454 71822 25506
rect 71874 25454 71876 25506
rect 71820 25442 71876 25454
rect 71932 25508 71988 26124
rect 72380 25956 72436 30830
rect 72492 30210 72548 32620
rect 72604 32674 72660 33292
rect 72604 32622 72606 32674
rect 72658 32622 72660 32674
rect 72604 32002 72660 32622
rect 72604 31950 72606 32002
rect 72658 31950 72660 32002
rect 72604 31938 72660 31950
rect 72828 32564 72884 32574
rect 72716 31668 72772 31678
rect 72716 31574 72772 31612
rect 72604 31444 72660 31454
rect 72604 31106 72660 31388
rect 72604 31054 72606 31106
rect 72658 31054 72660 31106
rect 72604 31042 72660 31054
rect 72492 30158 72494 30210
rect 72546 30158 72548 30210
rect 72492 30146 72548 30158
rect 72716 30996 72772 31006
rect 72828 30996 72884 32508
rect 72716 30994 72884 30996
rect 72716 30942 72718 30994
rect 72770 30942 72884 30994
rect 72716 30940 72884 30942
rect 72716 29426 72772 30940
rect 72828 30436 72884 30446
rect 72828 30342 72884 30380
rect 72940 30210 72996 33628
rect 73388 33458 73444 34076
rect 73500 34076 73668 34132
rect 73724 34690 73780 34702
rect 73724 34638 73726 34690
rect 73778 34638 73780 34690
rect 73500 33796 73556 34076
rect 73500 33730 73556 33740
rect 73612 33906 73668 33918
rect 73612 33854 73614 33906
rect 73666 33854 73668 33906
rect 73388 33406 73390 33458
rect 73442 33406 73444 33458
rect 73388 33394 73444 33406
rect 73276 33348 73332 33358
rect 73164 32674 73220 32686
rect 73164 32622 73166 32674
rect 73218 32622 73220 32674
rect 73164 32564 73220 32622
rect 73164 32498 73220 32508
rect 73164 32002 73220 32014
rect 73164 31950 73166 32002
rect 73218 31950 73220 32002
rect 73164 31890 73220 31950
rect 73164 31838 73166 31890
rect 73218 31838 73220 31890
rect 73164 31826 73220 31838
rect 73276 31778 73332 33292
rect 73612 33346 73668 33854
rect 73612 33294 73614 33346
rect 73666 33294 73668 33346
rect 73388 32564 73444 32574
rect 73612 32564 73668 33294
rect 73388 32562 73668 32564
rect 73388 32510 73390 32562
rect 73442 32510 73668 32562
rect 73388 32508 73668 32510
rect 73388 32498 73444 32508
rect 73724 32340 73780 34638
rect 73836 34356 73892 34366
rect 73836 34262 73892 34300
rect 73724 32274 73780 32284
rect 73836 33796 73892 33806
rect 73836 32116 73892 33740
rect 73276 31726 73278 31778
rect 73330 31726 73332 31778
rect 73276 31714 73332 31726
rect 73612 32060 73892 32116
rect 73948 33122 74004 34860
rect 74060 34850 74116 34860
rect 74172 34356 74228 35196
rect 74172 34290 74228 34300
rect 74396 34804 74452 34814
rect 74396 34132 74452 34748
rect 74396 34066 74452 34076
rect 74396 33458 74452 33470
rect 74396 33406 74398 33458
rect 74450 33406 74452 33458
rect 74396 33236 74452 33406
rect 74396 33170 74452 33180
rect 73948 33070 73950 33122
rect 74002 33070 74004 33122
rect 73388 31444 73444 31454
rect 73388 31218 73444 31388
rect 73388 31166 73390 31218
rect 73442 31166 73444 31218
rect 73388 31154 73444 31166
rect 73612 30994 73668 32060
rect 73948 32004 74004 33070
rect 74508 33012 74564 35532
rect 74732 34914 74788 34926
rect 74732 34862 74734 34914
rect 74786 34862 74788 34914
rect 74732 34804 74788 34862
rect 74732 34738 74788 34748
rect 74844 34580 74900 35868
rect 74956 35586 75012 35598
rect 74956 35534 74958 35586
rect 75010 35534 75012 35586
rect 74956 34916 75012 35534
rect 74956 34850 75012 34860
rect 74620 34524 74900 34580
rect 74956 34690 75012 34702
rect 74956 34638 74958 34690
rect 75010 34638 75012 34690
rect 74620 33346 74676 34524
rect 74732 34132 74788 34142
rect 74732 34038 74788 34076
rect 74844 34018 74900 34030
rect 74844 33966 74846 34018
rect 74898 33966 74900 34018
rect 74620 33294 74622 33346
rect 74674 33294 74676 33346
rect 74620 33282 74676 33294
rect 74732 33906 74788 33918
rect 74732 33854 74734 33906
rect 74786 33854 74788 33906
rect 74508 32946 74564 32956
rect 74732 32788 74788 33854
rect 74844 33684 74900 33966
rect 74956 33908 75012 34638
rect 75068 34130 75124 37438
rect 75180 37268 75236 37278
rect 75180 37174 75236 37212
rect 75292 37044 75348 39116
rect 75404 38724 75460 39228
rect 75404 38658 75460 38668
rect 75516 39060 75572 39070
rect 75516 38164 75572 39004
rect 75628 38836 75684 38846
rect 75628 38742 75684 38780
rect 75628 38164 75684 38174
rect 75572 38162 75684 38164
rect 75572 38110 75630 38162
rect 75682 38110 75684 38162
rect 75572 38108 75684 38110
rect 75516 38098 75572 38108
rect 75628 38098 75684 38108
rect 75404 37828 75460 37838
rect 75404 37378 75460 37772
rect 75404 37326 75406 37378
rect 75458 37326 75460 37378
rect 75404 37314 75460 37326
rect 75516 37716 75572 37726
rect 75180 36988 75348 37044
rect 75180 35810 75236 36988
rect 75404 36484 75460 36494
rect 75516 36484 75572 37660
rect 75460 36428 75572 36484
rect 75404 36390 75460 36428
rect 75628 36258 75684 36270
rect 75628 36206 75630 36258
rect 75682 36206 75684 36258
rect 75180 35758 75182 35810
rect 75234 35758 75236 35810
rect 75180 35746 75236 35758
rect 75292 35812 75348 35822
rect 75292 35698 75348 35756
rect 75292 35646 75294 35698
rect 75346 35646 75348 35698
rect 75292 35634 75348 35646
rect 75404 35476 75460 35486
rect 75404 35026 75460 35420
rect 75404 34974 75406 35026
rect 75458 34974 75460 35026
rect 75404 34962 75460 34974
rect 75628 34916 75684 36206
rect 75740 35924 75796 40348
rect 76188 38946 76244 40796
rect 76188 38894 76190 38946
rect 76242 38894 76244 38946
rect 76188 38882 76244 38894
rect 76300 40962 76356 40974
rect 76300 40910 76302 40962
rect 76354 40910 76356 40962
rect 75964 38834 76020 38846
rect 75964 38782 75966 38834
rect 76018 38782 76020 38834
rect 75964 38724 76020 38782
rect 76300 38668 76356 40910
rect 76412 39956 76468 42700
rect 76524 42690 76580 42700
rect 76524 41860 76580 41870
rect 76524 41300 76580 41804
rect 76524 41186 76580 41244
rect 76524 41134 76526 41186
rect 76578 41134 76580 41186
rect 76524 41122 76580 41134
rect 76636 41076 76692 41086
rect 76636 40514 76692 41020
rect 76748 41074 76804 41086
rect 76748 41022 76750 41074
rect 76802 41022 76804 41074
rect 76748 40628 76804 41022
rect 76748 40562 76804 40572
rect 76636 40462 76638 40514
rect 76690 40462 76692 40514
rect 76636 40450 76692 40462
rect 76412 39890 76468 39900
rect 76748 39730 76804 39742
rect 76748 39678 76750 39730
rect 76802 39678 76804 39730
rect 76524 39620 76580 39630
rect 76524 39526 76580 39564
rect 76412 39506 76468 39518
rect 76412 39454 76414 39506
rect 76466 39454 76468 39506
rect 76412 39060 76468 39454
rect 76412 39004 76580 39060
rect 75852 38500 75908 38510
rect 75852 36596 75908 38444
rect 75964 37378 76020 38668
rect 75964 37326 75966 37378
rect 76018 37326 76020 37378
rect 75964 37314 76020 37326
rect 76076 38612 76356 38668
rect 76412 38722 76468 38734
rect 76412 38670 76414 38722
rect 76466 38670 76468 38722
rect 76412 38612 76468 38670
rect 75852 36530 75908 36540
rect 76076 36484 76132 38612
rect 76412 38546 76468 38556
rect 76524 38500 76580 39004
rect 76524 38434 76580 38444
rect 76636 38834 76692 38846
rect 76636 38782 76638 38834
rect 76690 38782 76692 38834
rect 76188 38276 76244 38286
rect 76636 38276 76692 38782
rect 76244 38220 76356 38276
rect 76188 38210 76244 38220
rect 76188 38052 76244 38062
rect 76300 38052 76356 38220
rect 76636 38210 76692 38220
rect 76748 38164 76804 39678
rect 76860 39732 76916 50372
rect 77420 48580 77476 53004
rect 77868 52966 77924 53004
rect 78204 52946 78260 52958
rect 78204 52894 78206 52946
rect 78258 52894 78260 52946
rect 77644 52836 77700 52846
rect 78204 52836 78260 52894
rect 77644 52834 78260 52836
rect 77644 52782 77646 52834
rect 77698 52782 78260 52834
rect 77644 52780 78260 52782
rect 77644 52770 77700 52780
rect 78204 52276 78260 52780
rect 78204 52210 78260 52220
rect 77868 51492 77924 51502
rect 77420 48514 77476 48524
rect 77532 51490 77924 51492
rect 77532 51438 77870 51490
rect 77922 51438 77924 51490
rect 77532 51436 77924 51438
rect 77420 45332 77476 45342
rect 77532 45332 77588 51436
rect 77868 51426 77924 51436
rect 78204 51378 78260 51390
rect 78204 51326 78206 51378
rect 78258 51326 78260 51378
rect 77644 51266 77700 51278
rect 77644 51214 77646 51266
rect 77698 51214 77700 51266
rect 77644 51156 77700 51214
rect 77644 51090 77700 51100
rect 78204 51156 78260 51326
rect 78204 51090 78260 51100
rect 77644 50484 77700 50494
rect 77644 50390 77700 50428
rect 78204 50484 78260 50494
rect 77868 50372 77924 50382
rect 77868 50278 77924 50316
rect 78204 50036 78260 50428
rect 78204 49970 78260 49980
rect 77644 48916 77700 48926
rect 77644 48822 77700 48860
rect 78204 48916 78260 48926
rect 78204 48822 78260 48860
rect 77868 48804 77924 48814
rect 77868 48710 77924 48748
rect 77868 48356 77924 48366
rect 77756 48354 77924 48356
rect 77756 48302 77870 48354
rect 77922 48302 77924 48354
rect 77756 48300 77924 48302
rect 77644 48244 77700 48254
rect 77644 48150 77700 48188
rect 77644 47236 77700 47246
rect 77644 47142 77700 47180
rect 77644 45666 77700 45678
rect 77644 45614 77646 45666
rect 77698 45614 77700 45666
rect 77644 45556 77700 45614
rect 77644 45490 77700 45500
rect 77476 45276 77588 45332
rect 77420 45266 77476 45276
rect 77644 44996 77700 45006
rect 77644 44902 77700 44940
rect 77084 43538 77140 43550
rect 77084 43486 77086 43538
rect 77138 43486 77140 43538
rect 76972 43426 77028 43438
rect 76972 43374 76974 43426
rect 77026 43374 77028 43426
rect 76972 43314 77028 43374
rect 76972 43262 76974 43314
rect 77026 43262 77028 43314
rect 76972 43250 77028 43262
rect 77084 42980 77140 43486
rect 77420 43540 77476 43550
rect 77420 43446 77476 43484
rect 77644 43538 77700 43550
rect 77644 43486 77646 43538
rect 77698 43486 77700 43538
rect 77308 43428 77364 43438
rect 76972 42924 77140 42980
rect 77196 43426 77364 43428
rect 77196 43374 77310 43426
rect 77362 43374 77364 43426
rect 77196 43372 77364 43374
rect 76972 42642 77028 42924
rect 77196 42756 77252 43372
rect 77308 43362 77364 43372
rect 76972 42590 76974 42642
rect 77026 42590 77028 42642
rect 76972 41412 77028 42590
rect 76972 41186 77028 41356
rect 76972 41134 76974 41186
rect 77026 41134 77028 41186
rect 76972 41122 77028 41134
rect 77084 42700 77252 42756
rect 77532 42756 77588 42766
rect 77644 42756 77700 43486
rect 77532 42754 77700 42756
rect 77532 42702 77534 42754
rect 77586 42702 77700 42754
rect 77532 42700 77700 42702
rect 76860 39676 77028 39732
rect 76748 38098 76804 38108
rect 76300 37996 76580 38052
rect 76188 37958 76244 37996
rect 76524 37938 76580 37996
rect 76524 37886 76526 37938
rect 76578 37886 76580 37938
rect 76524 37874 76580 37886
rect 76636 38050 76692 38062
rect 76636 37998 76638 38050
rect 76690 37998 76692 38050
rect 76300 37826 76356 37838
rect 76300 37774 76302 37826
rect 76354 37774 76356 37826
rect 76188 37268 76244 37278
rect 76188 37174 76244 37212
rect 76188 36484 76244 36494
rect 76076 36482 76244 36484
rect 76076 36430 76190 36482
rect 76242 36430 76244 36482
rect 76076 36428 76244 36430
rect 76188 36418 76244 36428
rect 76300 36260 76356 37774
rect 76636 37828 76692 37998
rect 76636 37762 76692 37772
rect 76412 37548 76916 37604
rect 76412 37490 76468 37548
rect 76412 37438 76414 37490
rect 76466 37438 76468 37490
rect 76412 37426 76468 37438
rect 76636 37380 76692 37390
rect 76636 37266 76692 37324
rect 76636 37214 76638 37266
rect 76690 37214 76692 37266
rect 75964 36204 76356 36260
rect 76412 36594 76468 36606
rect 76412 36542 76414 36594
rect 76466 36542 76468 36594
rect 75740 35868 75908 35924
rect 75740 35700 75796 35710
rect 75740 35606 75796 35644
rect 75628 34850 75684 34860
rect 75292 34804 75348 34814
rect 75068 34078 75070 34130
rect 75122 34078 75124 34130
rect 75068 34066 75124 34078
rect 75180 34802 75348 34804
rect 75180 34750 75294 34802
rect 75346 34750 75348 34802
rect 75180 34748 75348 34750
rect 74956 33842 75012 33852
rect 74844 33628 75124 33684
rect 74732 32722 74788 32732
rect 74844 33458 74900 33470
rect 74844 33406 74846 33458
rect 74898 33406 74900 33458
rect 74844 32786 74900 33406
rect 74844 32734 74846 32786
rect 74898 32734 74900 32786
rect 74844 32722 74900 32734
rect 74284 32676 74340 32686
rect 74956 32676 75012 32686
rect 74284 32674 74676 32676
rect 74284 32622 74286 32674
rect 74338 32622 74676 32674
rect 74284 32620 74676 32622
rect 74284 32610 74340 32620
rect 74060 32562 74116 32574
rect 74060 32510 74062 32562
rect 74114 32510 74116 32562
rect 74060 32116 74116 32510
rect 74620 32562 74676 32620
rect 74956 32582 75012 32620
rect 74620 32510 74622 32562
rect 74674 32510 74676 32562
rect 74620 32498 74676 32510
rect 74060 32050 74116 32060
rect 74508 32340 74564 32350
rect 73948 31938 74004 31948
rect 73724 31556 73780 31566
rect 73724 31462 73780 31500
rect 73836 31554 73892 31566
rect 73836 31502 73838 31554
rect 73890 31502 73892 31554
rect 73612 30942 73614 30994
rect 73666 30942 73668 30994
rect 73612 30930 73668 30942
rect 72940 30158 72942 30210
rect 72994 30158 72996 30210
rect 72940 30146 72996 30158
rect 73612 30322 73668 30334
rect 73612 30270 73614 30322
rect 73666 30270 73668 30322
rect 73164 29540 73220 29550
rect 72940 29538 73220 29540
rect 72940 29486 73166 29538
rect 73218 29486 73220 29538
rect 72940 29484 73220 29486
rect 72716 29374 72718 29426
rect 72770 29374 72772 29426
rect 72716 29362 72772 29374
rect 72828 29426 72884 29438
rect 72828 29374 72830 29426
rect 72882 29374 72884 29426
rect 72492 29202 72548 29214
rect 72492 29150 72494 29202
rect 72546 29150 72548 29202
rect 72492 28868 72548 29150
rect 72492 28642 72548 28812
rect 72828 28756 72884 29374
rect 72828 28690 72884 28700
rect 72492 28590 72494 28642
rect 72546 28590 72548 28642
rect 72492 28578 72548 28590
rect 72604 28644 72660 28654
rect 72492 28420 72548 28430
rect 72492 27188 72548 28364
rect 72604 28082 72660 28588
rect 72604 28030 72606 28082
rect 72658 28030 72660 28082
rect 72604 28018 72660 28030
rect 72716 28532 72772 28542
rect 72716 27636 72772 28476
rect 72828 28532 72884 28542
rect 72940 28532 72996 29484
rect 73164 29474 73220 29484
rect 73500 29428 73556 29438
rect 73500 29334 73556 29372
rect 72828 28530 72996 28532
rect 72828 28478 72830 28530
rect 72882 28478 72996 28530
rect 72828 28476 72996 28478
rect 73052 29314 73108 29326
rect 73052 29262 73054 29314
rect 73106 29262 73108 29314
rect 72828 28084 72884 28476
rect 73052 28084 73108 29262
rect 73500 28756 73556 28766
rect 73500 28662 73556 28700
rect 73052 28028 73332 28084
rect 72828 27972 72884 28028
rect 72828 27970 73108 27972
rect 72828 27918 72830 27970
rect 72882 27918 73108 27970
rect 72828 27916 73108 27918
rect 72828 27906 72884 27916
rect 72716 27570 72772 27580
rect 72940 27746 72996 27758
rect 72940 27694 72942 27746
rect 72994 27694 72996 27746
rect 72716 27188 72772 27198
rect 72940 27188 72996 27694
rect 72492 27186 72772 27188
rect 72492 27134 72718 27186
rect 72770 27134 72772 27186
rect 72492 27132 72772 27134
rect 72716 27076 72772 27132
rect 72716 27010 72772 27020
rect 72828 27132 72996 27188
rect 72492 26516 72548 26526
rect 72548 26460 72772 26516
rect 72492 26422 72548 26460
rect 72604 25956 72660 25966
rect 72380 25900 72604 25956
rect 72604 25890 72660 25900
rect 72604 25732 72660 25742
rect 71932 25442 71988 25452
rect 72044 25618 72100 25630
rect 72044 25566 72046 25618
rect 72098 25566 72100 25618
rect 71596 25218 71652 25228
rect 71708 25172 71764 25182
rect 71708 24946 71764 25116
rect 71708 24894 71710 24946
rect 71762 24894 71764 24946
rect 71708 24882 71764 24894
rect 71820 25060 71876 25070
rect 71372 24612 71428 24622
rect 71372 24518 71428 24556
rect 71820 23940 71876 25004
rect 71708 23380 71764 23390
rect 71708 23286 71764 23324
rect 71820 23268 71876 23884
rect 71820 23202 71876 23212
rect 72044 23156 72100 25566
rect 72156 25172 72212 25182
rect 72156 24722 72212 25116
rect 72156 24670 72158 24722
rect 72210 24670 72212 24722
rect 72156 24658 72212 24670
rect 72268 25060 72324 25070
rect 72156 23940 72212 23950
rect 72156 23846 72212 23884
rect 72044 23090 72100 23100
rect 72156 23380 72212 23390
rect 72156 23154 72212 23324
rect 72156 23102 72158 23154
rect 72210 23102 72212 23154
rect 72156 23090 72212 23102
rect 72268 23044 72324 25004
rect 72380 24498 72436 24510
rect 72380 24446 72382 24498
rect 72434 24446 72436 24498
rect 72380 23604 72436 24446
rect 72380 23538 72436 23548
rect 72492 23828 72548 23838
rect 72380 23044 72436 23054
rect 72268 23042 72436 23044
rect 72268 22990 72382 23042
rect 72434 22990 72436 23042
rect 72268 22988 72436 22990
rect 72380 22978 72436 22988
rect 71932 22484 71988 22494
rect 71988 22428 72100 22484
rect 71932 22390 71988 22428
rect 72044 22370 72100 22428
rect 72044 22318 72046 22370
rect 72098 22318 72100 22370
rect 72044 22306 72100 22318
rect 72268 22482 72324 22494
rect 72268 22430 72270 22482
rect 72322 22430 72324 22482
rect 72268 22260 72324 22430
rect 72268 22194 72324 22204
rect 71708 21700 71764 21710
rect 71708 21606 71764 21644
rect 72156 21700 72212 21710
rect 72156 21586 72212 21644
rect 72156 21534 72158 21586
rect 72210 21534 72212 21586
rect 72156 21522 72212 21534
rect 72380 21362 72436 21374
rect 72380 21310 72382 21362
rect 72434 21310 72436 21362
rect 71260 20916 71316 20926
rect 71316 20860 71428 20916
rect 71260 20822 71316 20860
rect 71372 20802 71428 20860
rect 71372 20750 71374 20802
rect 71426 20750 71428 20802
rect 71372 20738 71428 20750
rect 72268 20692 72324 20702
rect 72268 20598 72324 20636
rect 72380 20188 72436 21310
rect 72492 20802 72548 23772
rect 72604 21588 72660 25676
rect 72716 25506 72772 26460
rect 72716 25454 72718 25506
rect 72770 25454 72772 25506
rect 72716 25442 72772 25454
rect 72716 24724 72772 24734
rect 72716 24388 72772 24668
rect 72828 24500 72884 27132
rect 72940 26964 72996 26974
rect 73052 26964 73108 27916
rect 73164 27860 73220 27870
rect 73164 27766 73220 27804
rect 73276 27188 73332 28028
rect 73388 27860 73444 27870
rect 73388 27858 73556 27860
rect 73388 27806 73390 27858
rect 73442 27806 73556 27858
rect 73388 27804 73556 27806
rect 73388 27794 73444 27804
rect 73276 27132 73444 27188
rect 73164 27076 73220 27114
rect 73164 27010 73220 27020
rect 72940 26962 73108 26964
rect 72940 26910 72942 26962
rect 72994 26910 73108 26962
rect 72940 26908 73108 26910
rect 73388 26908 73444 27132
rect 73500 27076 73556 27804
rect 73612 27748 73668 30270
rect 73724 30210 73780 30222
rect 73724 30158 73726 30210
rect 73778 30158 73780 30210
rect 73724 29428 73780 30158
rect 73724 29362 73780 29372
rect 73724 28644 73780 28654
rect 73724 28550 73780 28588
rect 73836 28532 73892 31502
rect 73948 31554 74004 31566
rect 73948 31502 73950 31554
rect 74002 31502 74004 31554
rect 73948 30548 74004 31502
rect 74060 31220 74116 31230
rect 74060 31126 74116 31164
rect 74172 31108 74228 31118
rect 74172 31014 74228 31052
rect 73948 30482 74004 30492
rect 74284 30994 74340 31006
rect 74284 30942 74286 30994
rect 74338 30942 74340 30994
rect 74284 30436 74340 30942
rect 74284 30370 74340 30380
rect 74396 29988 74452 29998
rect 74396 29426 74452 29932
rect 74396 29374 74398 29426
rect 74450 29374 74452 29426
rect 74396 29362 74452 29374
rect 74060 29204 74116 29214
rect 74060 29110 74116 29148
rect 74396 28868 74452 28878
rect 74396 28642 74452 28812
rect 74396 28590 74398 28642
rect 74450 28590 74452 28642
rect 74396 28578 74452 28590
rect 73836 28466 73892 28476
rect 74060 28420 74116 28430
rect 74060 28418 74228 28420
rect 74060 28366 74062 28418
rect 74114 28366 74228 28418
rect 74060 28364 74228 28366
rect 74060 28354 74116 28364
rect 73948 28196 74004 28206
rect 73724 28084 73780 28094
rect 73724 27970 73780 28028
rect 73724 27918 73726 27970
rect 73778 27918 73780 27970
rect 73724 27906 73780 27918
rect 73948 27858 74004 28140
rect 73948 27806 73950 27858
rect 74002 27806 74004 27858
rect 73948 27794 74004 27806
rect 73724 27748 73780 27758
rect 73612 27692 73724 27748
rect 73724 27682 73780 27692
rect 73836 27746 73892 27758
rect 73836 27694 73838 27746
rect 73890 27694 73892 27746
rect 73836 27300 73892 27694
rect 73500 26982 73556 27020
rect 73724 27244 73892 27300
rect 73724 26908 73780 27244
rect 74060 27076 74116 27086
rect 74060 26982 74116 27020
rect 72940 26898 72996 26908
rect 73164 26852 73220 26862
rect 73052 26850 73220 26852
rect 73052 26798 73166 26850
rect 73218 26798 73220 26850
rect 73052 26796 73220 26798
rect 72940 26740 72996 26750
rect 72940 25844 72996 26684
rect 73052 25956 73108 26796
rect 73164 26786 73220 26796
rect 73276 26852 73444 26908
rect 73612 26852 73780 26908
rect 74060 26852 74116 26862
rect 73276 26516 73332 26852
rect 73276 26450 73332 26460
rect 73388 26290 73444 26302
rect 73388 26238 73390 26290
rect 73442 26238 73444 26290
rect 73164 26180 73220 26190
rect 73388 26180 73444 26238
rect 73220 26124 73444 26180
rect 73164 26086 73220 26124
rect 73500 25956 73556 25966
rect 73052 25900 73332 25956
rect 72940 25788 73108 25844
rect 72940 25620 72996 25630
rect 72940 25526 72996 25564
rect 72940 25284 72996 25294
rect 72940 24722 72996 25228
rect 72940 24670 72942 24722
rect 72994 24670 72996 24722
rect 72940 24658 72996 24670
rect 72828 24444 72996 24500
rect 72716 24332 72884 24388
rect 72716 23940 72772 23950
rect 72716 23846 72772 23884
rect 72828 22370 72884 24332
rect 72940 23154 72996 24444
rect 72940 23102 72942 23154
rect 72994 23102 72996 23154
rect 72940 23090 72996 23102
rect 72828 22318 72830 22370
rect 72882 22318 72884 22370
rect 72828 22306 72884 22318
rect 72940 21588 72996 21598
rect 72604 21586 72996 21588
rect 72604 21534 72942 21586
rect 72994 21534 72996 21586
rect 72604 21532 72996 21534
rect 72940 21522 72996 21532
rect 72492 20750 72494 20802
rect 72546 20750 72548 20802
rect 72492 20738 72548 20750
rect 72716 20802 72772 20814
rect 73052 20804 73108 25788
rect 73276 24164 73332 25900
rect 73500 25506 73556 25900
rect 73500 25454 73502 25506
rect 73554 25454 73556 25506
rect 73500 25442 73556 25454
rect 73500 24722 73556 24734
rect 73500 24670 73502 24722
rect 73554 24670 73556 24722
rect 73500 24612 73556 24670
rect 73612 24724 73668 26852
rect 73836 26516 73892 26526
rect 73724 25618 73780 25630
rect 73724 25566 73726 25618
rect 73778 25566 73780 25618
rect 73724 24836 73780 25566
rect 73836 25396 73892 26460
rect 74060 26292 74116 26796
rect 74172 26740 74228 28364
rect 74396 28196 74452 28206
rect 74284 27858 74340 27870
rect 74284 27806 74286 27858
rect 74338 27806 74340 27858
rect 74284 27748 74340 27806
rect 74284 27682 74340 27692
rect 74284 26740 74340 26750
rect 74172 26684 74284 26740
rect 74284 26674 74340 26684
rect 74172 26292 74228 26302
rect 74060 26290 74228 26292
rect 74060 26238 74174 26290
rect 74226 26238 74228 26290
rect 74060 26236 74228 26238
rect 74172 26226 74228 26236
rect 74396 25730 74452 28140
rect 74396 25678 74398 25730
rect 74450 25678 74452 25730
rect 74396 25666 74452 25678
rect 73836 25340 74116 25396
rect 74060 25284 74116 25340
rect 74060 25228 74228 25284
rect 73724 24770 73780 24780
rect 74060 24948 74116 24958
rect 73612 24658 73668 24668
rect 73836 24722 73892 24734
rect 73836 24670 73838 24722
rect 73890 24670 73892 24722
rect 73500 24546 73556 24556
rect 73276 24108 73780 24164
rect 73164 24052 73220 24062
rect 73164 23958 73220 23996
rect 73276 23940 73332 23950
rect 73276 23846 73332 23884
rect 73276 23042 73332 23054
rect 73276 22990 73278 23042
rect 73330 22990 73332 23042
rect 73276 21028 73332 22990
rect 73388 22370 73444 22382
rect 73388 22318 73390 22370
rect 73442 22318 73444 22370
rect 73388 21924 73444 22318
rect 73724 21924 73780 24108
rect 73836 24052 73892 24670
rect 74060 24610 74116 24892
rect 74060 24558 74062 24610
rect 74114 24558 74116 24610
rect 74060 24546 74116 24558
rect 74060 24164 74116 24202
rect 74060 24098 74116 24108
rect 73836 23986 73892 23996
rect 73948 23268 74004 23278
rect 73948 23154 74004 23212
rect 73948 23102 73950 23154
rect 74002 23102 74004 23154
rect 73948 23090 74004 23102
rect 74060 22932 74116 22942
rect 74060 22838 74116 22876
rect 74060 22372 74116 22382
rect 74172 22372 74228 25228
rect 74508 24724 74564 32284
rect 75068 32228 75124 33628
rect 75180 33236 75236 34748
rect 75292 34738 75348 34748
rect 75516 34692 75572 34702
rect 75740 34692 75796 34702
rect 75516 34690 75684 34692
rect 75516 34638 75518 34690
rect 75570 34638 75684 34690
rect 75516 34636 75684 34638
rect 75516 34626 75572 34636
rect 75292 34020 75348 34030
rect 75292 33346 75348 33964
rect 75628 33572 75684 34636
rect 75740 34356 75796 34636
rect 75740 34290 75796 34300
rect 75628 33506 75684 33516
rect 75292 33294 75294 33346
rect 75346 33294 75348 33346
rect 75292 33282 75348 33294
rect 75180 32676 75236 33180
rect 75852 33124 75908 35868
rect 75964 34916 76020 36204
rect 76412 36036 76468 36542
rect 76412 35970 76468 35980
rect 76076 35812 76132 35822
rect 76524 35812 76580 35822
rect 76636 35812 76692 37214
rect 76076 35810 76692 35812
rect 76076 35758 76078 35810
rect 76130 35758 76526 35810
rect 76578 35758 76692 35810
rect 76076 35756 76692 35758
rect 76748 36594 76804 36606
rect 76748 36542 76750 36594
rect 76802 36542 76804 36594
rect 76076 35746 76132 35756
rect 76524 35746 76580 35756
rect 76636 35586 76692 35598
rect 76636 35534 76638 35586
rect 76690 35534 76692 35586
rect 76636 35252 76692 35534
rect 76748 35476 76804 36542
rect 76860 36482 76916 37548
rect 76860 36430 76862 36482
rect 76914 36430 76916 36482
rect 76860 36418 76916 36430
rect 76972 35924 77028 39676
rect 77084 38834 77140 42700
rect 77308 42644 77364 42654
rect 77308 42550 77364 42588
rect 77196 42530 77252 42542
rect 77196 42478 77198 42530
rect 77250 42478 77252 42530
rect 77196 41188 77252 42478
rect 77308 42308 77364 42318
rect 77308 41300 77364 42252
rect 77308 41244 77476 41300
rect 77196 41132 77364 41188
rect 77196 40962 77252 40974
rect 77196 40910 77198 40962
rect 77250 40910 77252 40962
rect 77196 39844 77252 40910
rect 77196 39778 77252 39788
rect 77308 39618 77364 41132
rect 77420 41074 77476 41244
rect 77532 41188 77588 42700
rect 77532 41094 77588 41132
rect 77420 41022 77422 41074
rect 77474 41022 77476 41074
rect 77420 40628 77476 41022
rect 77420 40562 77476 40572
rect 77756 40404 77812 48300
rect 77868 48290 77924 48300
rect 78204 48244 78260 48254
rect 78204 47796 78260 48188
rect 78204 47730 78260 47740
rect 78204 47346 78260 47358
rect 78204 47294 78206 47346
rect 78258 47294 78260 47346
rect 77868 47234 77924 47246
rect 77868 47182 77870 47234
rect 77922 47182 77924 47234
rect 77868 45892 77924 47182
rect 78204 47236 78260 47294
rect 78204 46676 78260 47180
rect 78204 46610 78260 46620
rect 77868 45826 77924 45836
rect 78204 45778 78260 45790
rect 78204 45726 78206 45778
rect 78258 45726 78260 45778
rect 77868 45668 77924 45678
rect 77868 45574 77924 45612
rect 78204 45556 78260 45726
rect 78204 45490 78260 45500
rect 77868 45218 77924 45230
rect 77868 45166 77870 45218
rect 77922 45166 77924 45218
rect 77868 42756 77924 45166
rect 78204 45106 78260 45118
rect 78204 45054 78206 45106
rect 78258 45054 78260 45106
rect 78204 44996 78260 45054
rect 78204 44436 78260 44940
rect 78204 44370 78260 44380
rect 78316 44098 78372 44110
rect 78316 44046 78318 44098
rect 78370 44046 78372 44098
rect 78316 43652 78372 44046
rect 78092 43596 78372 43652
rect 78092 43316 78148 43596
rect 78204 43428 78260 43438
rect 78204 43334 78260 43372
rect 77868 42700 78036 42756
rect 77868 42530 77924 42542
rect 77868 42478 77870 42530
rect 77922 42478 77924 42530
rect 77868 40740 77924 42478
rect 77980 42420 78036 42700
rect 78092 42754 78148 43260
rect 78092 42702 78094 42754
rect 78146 42702 78148 42754
rect 78092 42690 78148 42702
rect 77980 42364 78372 42420
rect 77980 42196 78036 42206
rect 77980 41858 78036 42140
rect 77980 41806 77982 41858
rect 78034 41806 78036 41858
rect 77980 41794 78036 41806
rect 78092 41300 78148 41310
rect 78092 41206 78148 41244
rect 77868 40674 77924 40684
rect 77980 40628 78036 40638
rect 78036 40572 78260 40628
rect 77980 40562 78036 40572
rect 77308 39566 77310 39618
rect 77362 39566 77364 39618
rect 77308 39554 77364 39566
rect 77420 40348 77812 40404
rect 77868 40402 77924 40414
rect 77868 40350 77870 40402
rect 77922 40350 77924 40402
rect 77084 38782 77086 38834
rect 77138 38782 77140 38834
rect 77084 38770 77140 38782
rect 77196 38724 77252 38734
rect 77084 38612 77252 38668
rect 77084 38050 77140 38612
rect 77084 37998 77086 38050
rect 77138 37998 77140 38050
rect 77084 37986 77140 37998
rect 77196 38500 77252 38510
rect 77196 37266 77252 38444
rect 77308 38388 77364 38398
rect 77308 37938 77364 38332
rect 77308 37886 77310 37938
rect 77362 37886 77364 37938
rect 77308 37492 77364 37886
rect 77308 37426 77364 37436
rect 77196 37214 77198 37266
rect 77250 37214 77252 37266
rect 77196 37202 77252 37214
rect 77420 37268 77476 40348
rect 77644 39844 77700 39854
rect 77700 39788 77812 39844
rect 77644 39778 77700 39788
rect 77756 39284 77812 39788
rect 77868 39506 77924 40350
rect 78092 40180 78148 40190
rect 78092 39618 78148 40124
rect 78092 39566 78094 39618
rect 78146 39566 78148 39618
rect 78092 39554 78148 39566
rect 77868 39454 77870 39506
rect 77922 39454 77924 39506
rect 77868 39442 77924 39454
rect 77756 39228 77924 39284
rect 77644 38948 77700 38958
rect 77644 38854 77700 38892
rect 77532 38834 77588 38846
rect 77532 38782 77534 38834
rect 77586 38782 77588 38834
rect 77532 38162 77588 38782
rect 77756 38836 77812 38846
rect 77532 38110 77534 38162
rect 77586 38110 77588 38162
rect 77532 38098 77588 38110
rect 77644 38276 77700 38286
rect 77644 37938 77700 38220
rect 77644 37886 77646 37938
rect 77698 37886 77700 37938
rect 77644 37380 77700 37886
rect 77644 37314 77700 37324
rect 77420 37212 77588 37268
rect 77308 37154 77364 37166
rect 77308 37102 77310 37154
rect 77362 37102 77364 37154
rect 77308 36708 77364 37102
rect 77308 36642 77364 36652
rect 77420 37042 77476 37054
rect 77420 36990 77422 37042
rect 77474 36990 77476 37042
rect 77420 36148 77476 36990
rect 77420 36082 77476 36092
rect 76972 35868 77252 35924
rect 76860 35812 76916 35822
rect 76860 35718 76916 35756
rect 76748 35410 76804 35420
rect 76972 35698 77028 35710
rect 76972 35646 76974 35698
rect 77026 35646 77028 35698
rect 76636 35196 76916 35252
rect 76524 35026 76580 35038
rect 76524 34974 76526 35026
rect 76578 34974 76580 35026
rect 76076 34916 76132 34926
rect 75964 34914 76132 34916
rect 75964 34862 76078 34914
rect 76130 34862 76132 34914
rect 75964 34860 76132 34862
rect 76076 34850 76132 34860
rect 76524 34580 76580 34974
rect 76524 34514 76580 34524
rect 76748 35026 76804 35038
rect 76748 34974 76750 35026
rect 76802 34974 76804 35026
rect 76636 34468 76692 34478
rect 75964 34356 76020 34366
rect 75964 34262 76020 34300
rect 75852 33058 75908 33068
rect 76300 34244 76356 34254
rect 76300 32900 76356 34188
rect 76636 34242 76692 34412
rect 76636 34190 76638 34242
rect 76690 34190 76692 34242
rect 76636 34178 76692 34190
rect 76412 34132 76468 34142
rect 76412 34038 76468 34076
rect 76748 33570 76804 34974
rect 76860 34914 76916 35196
rect 76860 34862 76862 34914
rect 76914 34862 76916 34914
rect 76860 34850 76916 34862
rect 76860 34132 76916 34142
rect 76972 34132 77028 35646
rect 76860 34130 76972 34132
rect 76860 34078 76862 34130
rect 76914 34078 76972 34130
rect 76860 34076 76972 34078
rect 76860 34066 76916 34076
rect 76748 33518 76750 33570
rect 76802 33518 76804 33570
rect 76748 33506 76804 33518
rect 76860 33908 76916 33918
rect 76524 33460 76580 33470
rect 76524 33366 76580 33404
rect 76860 33234 76916 33852
rect 76860 33182 76862 33234
rect 76914 33182 76916 33234
rect 76860 33170 76916 33182
rect 75628 32844 76356 32900
rect 75628 32786 75684 32844
rect 75628 32734 75630 32786
rect 75682 32734 75684 32786
rect 75628 32722 75684 32734
rect 75180 32610 75236 32620
rect 75740 32676 75796 32686
rect 75796 32620 75908 32676
rect 75740 32610 75796 32620
rect 75068 32162 75124 32172
rect 75292 32562 75348 32574
rect 75292 32510 75294 32562
rect 75346 32510 75348 32562
rect 75292 32452 75348 32510
rect 74844 32116 74900 32126
rect 74732 31892 74788 31902
rect 74732 31798 74788 31836
rect 74844 31218 74900 32060
rect 75180 32004 75236 32014
rect 74844 31166 74846 31218
rect 74898 31166 74900 31218
rect 74844 31154 74900 31166
rect 75068 31780 75124 31790
rect 75068 31220 75124 31724
rect 75180 31668 75236 31948
rect 75292 31892 75348 32396
rect 75292 31826 75348 31836
rect 75180 31612 75348 31668
rect 75180 31220 75236 31230
rect 75068 31218 75236 31220
rect 75068 31166 75182 31218
rect 75234 31166 75236 31218
rect 75068 31164 75236 31166
rect 75180 31154 75236 31164
rect 75180 30996 75236 31006
rect 75068 30940 75180 30996
rect 74620 30772 74676 30782
rect 74620 30322 74676 30716
rect 74620 30270 74622 30322
rect 74674 30270 74676 30322
rect 74620 30258 74676 30270
rect 75068 30210 75124 30940
rect 75180 30930 75236 30940
rect 75068 30158 75070 30210
rect 75122 30158 75124 30210
rect 75068 30146 75124 30158
rect 75292 29988 75348 31612
rect 75404 31554 75460 31566
rect 75404 31502 75406 31554
rect 75458 31502 75460 31554
rect 75404 31332 75460 31502
rect 75404 31266 75460 31276
rect 75740 31332 75796 31342
rect 75404 30996 75460 31006
rect 75404 30210 75460 30940
rect 75404 30158 75406 30210
rect 75458 30158 75460 30210
rect 75404 30146 75460 30158
rect 75516 30994 75572 31006
rect 75516 30942 75518 30994
rect 75570 30942 75572 30994
rect 75516 30100 75572 30942
rect 75628 30884 75684 30894
rect 75628 30790 75684 30828
rect 75292 29932 75460 29988
rect 74844 29428 74900 29438
rect 74844 29426 75348 29428
rect 74844 29374 74846 29426
rect 74898 29374 75348 29426
rect 74844 29372 75348 29374
rect 74844 29362 74900 29372
rect 74732 28980 74788 28990
rect 74732 28644 74788 28924
rect 74732 28530 74788 28588
rect 75068 28868 75124 28878
rect 75068 28642 75124 28812
rect 75068 28590 75070 28642
rect 75122 28590 75124 28642
rect 75068 28578 75124 28590
rect 74732 28478 74734 28530
rect 74786 28478 74788 28530
rect 74732 28466 74788 28478
rect 75180 28420 75236 28430
rect 74956 27972 75012 27982
rect 74732 27858 74788 27870
rect 74732 27806 74734 27858
rect 74786 27806 74788 27858
rect 74732 27748 74788 27806
rect 74956 27858 75012 27916
rect 75180 27970 75236 28364
rect 75180 27918 75182 27970
rect 75234 27918 75236 27970
rect 75180 27906 75236 27918
rect 74956 27806 74958 27858
rect 75010 27806 75012 27858
rect 74956 27794 75012 27806
rect 74620 27188 74676 27198
rect 74620 26962 74676 27132
rect 74620 26910 74622 26962
rect 74674 26910 74676 26962
rect 74620 26628 74676 26910
rect 74732 26964 74788 27692
rect 75068 27746 75124 27758
rect 75068 27694 75070 27746
rect 75122 27694 75124 27746
rect 74732 26898 74788 26908
rect 74956 27076 75012 27086
rect 74956 26962 75012 27020
rect 74956 26910 74958 26962
rect 75010 26910 75012 26962
rect 74956 26898 75012 26910
rect 74620 26562 74676 26572
rect 74620 26404 74676 26414
rect 74620 26310 74676 26348
rect 74732 26290 74788 26302
rect 74732 26238 74734 26290
rect 74786 26238 74788 26290
rect 74732 26180 74788 26238
rect 74732 26114 74788 26124
rect 74732 25730 74788 25742
rect 74732 25678 74734 25730
rect 74786 25678 74788 25730
rect 74732 25618 74788 25678
rect 74732 25566 74734 25618
rect 74786 25566 74788 25618
rect 74732 25554 74788 25566
rect 74620 24724 74676 24734
rect 74508 24722 74676 24724
rect 74508 24670 74622 24722
rect 74674 24670 74676 24722
rect 74508 24668 74676 24670
rect 74620 24658 74676 24668
rect 74508 24052 74564 24062
rect 74508 23958 74564 23996
rect 74396 23940 74452 23950
rect 74396 23846 74452 23884
rect 74956 23604 75012 23614
rect 74844 23548 74956 23604
rect 74732 23042 74788 23054
rect 74732 22990 74734 23042
rect 74786 22990 74788 23042
rect 74284 22596 74340 22606
rect 74284 22502 74340 22540
rect 74172 22316 74340 22372
rect 74060 22148 74116 22316
rect 74060 22092 74228 22148
rect 73724 21868 74116 21924
rect 73388 21858 73444 21868
rect 73948 21700 74004 21710
rect 73836 21698 74004 21700
rect 73836 21646 73950 21698
rect 74002 21646 74004 21698
rect 73836 21644 74004 21646
rect 73500 21586 73556 21598
rect 73500 21534 73502 21586
rect 73554 21534 73556 21586
rect 73500 21476 73556 21534
rect 73500 21410 73556 21420
rect 73276 20962 73332 20972
rect 72716 20750 72718 20802
rect 72770 20750 72772 20802
rect 72156 20132 72436 20188
rect 72716 20132 72772 20750
rect 72940 20802 73108 20804
rect 72940 20750 73054 20802
rect 73106 20750 73108 20802
rect 72940 20748 73108 20750
rect 72940 20242 72996 20748
rect 73052 20738 73108 20748
rect 72940 20190 72942 20242
rect 72994 20190 72996 20242
rect 72940 20178 72996 20190
rect 71260 18676 71316 18686
rect 71148 18674 71316 18676
rect 71148 18622 71262 18674
rect 71314 18622 71316 18674
rect 71148 18620 71316 18622
rect 71260 18610 71316 18620
rect 72156 16996 72212 20132
rect 72716 20066 72772 20076
rect 73836 19348 73892 21644
rect 73948 21634 74004 21644
rect 74060 21476 74116 21868
rect 73948 21420 74116 21476
rect 73948 20802 74004 21420
rect 73948 20750 73950 20802
rect 74002 20750 74004 20802
rect 73948 20738 74004 20750
rect 74060 20692 74116 20702
rect 74060 20598 74116 20636
rect 73948 20244 74004 20254
rect 74172 20244 74228 22092
rect 74284 21586 74340 22316
rect 74284 21534 74286 21586
rect 74338 21534 74340 21586
rect 74284 21522 74340 21534
rect 74620 21474 74676 21486
rect 74620 21422 74622 21474
rect 74674 21422 74676 21474
rect 73948 20242 74228 20244
rect 73948 20190 73950 20242
rect 74002 20190 74228 20242
rect 73948 20188 74228 20190
rect 74284 20914 74340 20926
rect 74284 20862 74286 20914
rect 74338 20862 74340 20914
rect 73948 20178 74004 20188
rect 73836 19282 73892 19292
rect 74284 18900 74340 20862
rect 74284 18834 74340 18844
rect 74620 18116 74676 21422
rect 74732 20244 74788 22990
rect 74844 22370 74900 23548
rect 74956 23538 75012 23548
rect 74956 23156 75012 23166
rect 75068 23156 75124 27694
rect 75292 27412 75348 29372
rect 75404 28644 75460 29932
rect 75516 29426 75572 30044
rect 75628 29986 75684 29998
rect 75628 29934 75630 29986
rect 75682 29934 75684 29986
rect 75628 29652 75684 29934
rect 75628 29586 75684 29596
rect 75516 29374 75518 29426
rect 75570 29374 75572 29426
rect 75516 28980 75572 29374
rect 75628 29428 75684 29438
rect 75628 29334 75684 29372
rect 75516 28914 75572 28924
rect 75404 28588 75572 28644
rect 75404 28420 75460 28458
rect 75404 28354 75460 28364
rect 75292 27356 75460 27412
rect 75404 27186 75460 27356
rect 75404 27134 75406 27186
rect 75458 27134 75460 27186
rect 75404 27122 75460 27134
rect 75292 27076 75348 27086
rect 75292 26982 75348 27020
rect 75516 26908 75572 28588
rect 75628 28532 75684 28542
rect 75628 27858 75684 28476
rect 75628 27806 75630 27858
rect 75682 27806 75684 27858
rect 75628 27794 75684 27806
rect 75740 27412 75796 31276
rect 75852 31106 75908 32620
rect 76300 32564 76356 32844
rect 76748 32786 76804 32798
rect 76748 32734 76750 32786
rect 76802 32734 76804 32786
rect 76412 32564 76468 32574
rect 76300 32562 76468 32564
rect 76300 32510 76414 32562
rect 76466 32510 76468 32562
rect 76300 32508 76468 32510
rect 76076 32452 76132 32462
rect 76076 32358 76132 32396
rect 76188 31780 76244 31790
rect 76300 31780 76356 32508
rect 76412 32498 76468 32508
rect 76188 31778 76356 31780
rect 76188 31726 76190 31778
rect 76242 31726 76356 31778
rect 76188 31724 76356 31726
rect 76412 31780 76468 31790
rect 76188 31714 76244 31724
rect 76412 31686 76468 31724
rect 76636 31778 76692 31790
rect 76636 31726 76638 31778
rect 76690 31726 76692 31778
rect 76300 31556 76356 31566
rect 76300 31462 76356 31500
rect 75852 31054 75854 31106
rect 75906 31054 75908 31106
rect 75852 29764 75908 31054
rect 76412 31106 76468 31118
rect 76412 31054 76414 31106
rect 76466 31054 76468 31106
rect 76076 30996 76132 31006
rect 76412 30996 76468 31054
rect 76076 30994 76468 30996
rect 76076 30942 76078 30994
rect 76130 30942 76468 30994
rect 76076 30940 76468 30942
rect 76076 30930 76132 30940
rect 76412 30660 76468 30940
rect 76636 30660 76692 31726
rect 76748 31220 76804 32734
rect 76860 32676 76916 32686
rect 76860 32582 76916 32620
rect 76972 32562 77028 34076
rect 77084 34244 77140 34254
rect 77084 34130 77140 34188
rect 77084 34078 77086 34130
rect 77138 34078 77140 34130
rect 77084 34066 77140 34078
rect 77084 33236 77140 33246
rect 77084 33142 77140 33180
rect 77196 32788 77252 35868
rect 77532 35476 77588 37212
rect 77644 37044 77700 37054
rect 77644 36596 77700 36988
rect 77644 35922 77700 36540
rect 77644 35870 77646 35922
rect 77698 35870 77700 35922
rect 77644 35858 77700 35870
rect 77308 35420 77588 35476
rect 77308 35028 77364 35420
rect 77756 35364 77812 38780
rect 77868 37266 77924 39228
rect 78092 38834 78148 38846
rect 78092 38782 78094 38834
rect 78146 38782 78148 38834
rect 77868 37214 77870 37266
rect 77922 37214 77924 37266
rect 77868 37202 77924 37214
rect 77980 38164 78036 38174
rect 77868 36932 77924 36942
rect 77868 36706 77924 36876
rect 77868 36654 77870 36706
rect 77922 36654 77924 36706
rect 77868 35924 77924 36654
rect 77980 36594 78036 38108
rect 77980 36542 77982 36594
rect 78034 36542 78036 36594
rect 77980 36530 78036 36542
rect 77868 35858 77924 35868
rect 77980 35812 78036 35822
rect 77868 35698 77924 35710
rect 77868 35646 77870 35698
rect 77922 35646 77924 35698
rect 77868 35364 77924 35646
rect 77308 34962 77364 34972
rect 77420 35308 77924 35364
rect 77308 34020 77364 34030
rect 77308 33926 77364 33964
rect 76972 32510 76974 32562
rect 77026 32510 77028 32562
rect 76972 32002 77028 32510
rect 76972 31950 76974 32002
rect 77026 31950 77028 32002
rect 76972 31938 77028 31950
rect 77084 32732 77252 32788
rect 76748 31154 76804 31164
rect 76860 31332 76916 31342
rect 76748 30996 76804 31006
rect 76860 30996 76916 31276
rect 77084 31108 77140 32732
rect 77196 32002 77252 32014
rect 77196 31950 77198 32002
rect 77250 31950 77252 32002
rect 77196 31668 77252 31950
rect 77308 31892 77364 31902
rect 77420 31892 77476 35308
rect 77868 35140 77924 35150
rect 77756 35084 77868 35140
rect 77532 35028 77588 35038
rect 77532 34580 77588 34972
rect 77532 34242 77588 34524
rect 77532 34190 77534 34242
rect 77586 34190 77588 34242
rect 77532 34178 77588 34190
rect 77644 34132 77700 34142
rect 77644 34038 77700 34076
rect 77532 33346 77588 33358
rect 77532 33294 77534 33346
rect 77586 33294 77588 33346
rect 77532 32228 77588 33294
rect 77756 33234 77812 35084
rect 77868 35046 77924 35084
rect 77756 33182 77758 33234
rect 77810 33182 77812 33234
rect 77756 33170 77812 33182
rect 77868 33572 77924 33582
rect 77868 32786 77924 33516
rect 77868 32734 77870 32786
rect 77922 32734 77924 32786
rect 77868 32722 77924 32734
rect 77644 32564 77700 32574
rect 77980 32564 78036 35756
rect 78092 35026 78148 38782
rect 78204 38162 78260 40572
rect 78204 38110 78206 38162
rect 78258 38110 78260 38162
rect 78204 38098 78260 38110
rect 78316 36820 78372 42364
rect 78316 36754 78372 36764
rect 78204 36482 78260 36494
rect 78204 36430 78206 36482
rect 78258 36430 78260 36482
rect 78204 35922 78260 36430
rect 78204 35870 78206 35922
rect 78258 35870 78260 35922
rect 78204 35858 78260 35870
rect 78092 34974 78094 35026
rect 78146 34974 78148 35026
rect 78092 34962 78148 34974
rect 78316 35476 78372 35486
rect 78204 34916 78260 34926
rect 78204 34822 78260 34860
rect 77644 32562 78036 32564
rect 77644 32510 77646 32562
rect 77698 32510 78036 32562
rect 77644 32508 78036 32510
rect 78092 34468 78148 34478
rect 77644 32498 77700 32508
rect 77868 32228 77924 32238
rect 77532 32172 77812 32228
rect 77532 32004 77588 32042
rect 77532 31938 77588 31948
rect 77308 31890 77476 31892
rect 77308 31838 77310 31890
rect 77362 31838 77476 31890
rect 77308 31836 77476 31838
rect 77308 31826 77364 31836
rect 77532 31780 77588 31790
rect 77756 31780 77812 32172
rect 77868 32002 77924 32172
rect 77868 31950 77870 32002
rect 77922 31950 77924 32002
rect 77868 31938 77924 31950
rect 77756 31724 77924 31780
rect 77196 31612 77476 31668
rect 77308 31220 77364 31230
rect 77308 31126 77364 31164
rect 77084 31052 77252 31108
rect 76748 30994 77140 30996
rect 76748 30942 76750 30994
rect 76802 30942 77140 30994
rect 76748 30940 77140 30942
rect 76748 30930 76804 30940
rect 76412 30604 76692 30660
rect 76412 30324 76468 30334
rect 76076 30210 76132 30222
rect 76076 30158 76078 30210
rect 76130 30158 76132 30210
rect 76076 30100 76132 30158
rect 76076 30034 76132 30044
rect 76300 29988 76356 29998
rect 76300 29894 76356 29932
rect 75852 29708 76244 29764
rect 75852 29540 75908 29550
rect 76076 29540 76132 29578
rect 75852 29538 76020 29540
rect 75852 29486 75854 29538
rect 75906 29486 76020 29538
rect 75852 29484 76020 29486
rect 75852 29474 75908 29484
rect 75964 29428 76020 29484
rect 76076 29474 76132 29484
rect 75964 29362 76020 29372
rect 76076 28644 76132 28654
rect 76076 28550 76132 28588
rect 75852 27972 75908 27982
rect 76188 27972 76244 29708
rect 76300 29652 76356 29662
rect 76412 29652 76468 30268
rect 76636 30210 76692 30604
rect 76636 30158 76638 30210
rect 76690 30158 76692 30210
rect 76524 30100 76580 30110
rect 76524 30006 76580 30044
rect 76636 29876 76692 30158
rect 77084 30210 77140 30940
rect 77084 30158 77086 30210
rect 77138 30158 77140 30210
rect 77084 30146 77140 30158
rect 77196 29988 77252 31052
rect 76300 29650 76468 29652
rect 76300 29598 76302 29650
rect 76354 29598 76468 29650
rect 76300 29596 76468 29598
rect 76524 29820 76692 29876
rect 76972 29932 77252 29988
rect 77308 30100 77364 30110
rect 76300 29586 76356 29596
rect 76524 29540 76580 29820
rect 76972 29764 77028 29932
rect 76524 29474 76580 29484
rect 76636 29540 76692 29550
rect 76636 29538 76916 29540
rect 76636 29486 76638 29538
rect 76690 29486 76916 29538
rect 76636 29484 76916 29486
rect 76636 29474 76692 29484
rect 76748 29316 76804 29326
rect 76412 29314 76804 29316
rect 76412 29262 76750 29314
rect 76802 29262 76804 29314
rect 76412 29260 76804 29262
rect 76300 29202 76356 29214
rect 76300 29150 76302 29202
rect 76354 29150 76356 29202
rect 76300 28754 76356 29150
rect 76300 28702 76302 28754
rect 76354 28702 76356 28754
rect 76300 28690 76356 28702
rect 76412 28196 76468 29260
rect 76748 29250 76804 29260
rect 76860 28756 76916 29484
rect 76972 29538 77028 29708
rect 76972 29486 76974 29538
rect 77026 29486 77028 29538
rect 76972 29474 77028 29486
rect 76636 28700 76916 28756
rect 76524 28644 76580 28654
rect 76524 28550 76580 28588
rect 76636 28420 76692 28700
rect 76860 28644 76916 28700
rect 77084 29426 77140 29438
rect 77084 29374 77086 29426
rect 77138 29374 77140 29426
rect 76972 28644 77028 28654
rect 76860 28642 77028 28644
rect 76860 28590 76974 28642
rect 77026 28590 77028 28642
rect 76860 28588 77028 28590
rect 76972 28578 77028 28588
rect 77084 28644 77140 29374
rect 76412 28140 76580 28196
rect 76412 27972 76468 27982
rect 76188 27970 76468 27972
rect 76188 27918 76414 27970
rect 76466 27918 76468 27970
rect 76188 27916 76468 27918
rect 75852 27878 75908 27916
rect 76412 27906 76468 27916
rect 76524 27524 76580 28140
rect 76636 27970 76692 28364
rect 76748 28530 76804 28542
rect 76748 28478 76750 28530
rect 76802 28478 76804 28530
rect 76748 28196 76804 28478
rect 77084 28196 77140 28588
rect 76748 28140 77140 28196
rect 76636 27918 76638 27970
rect 76690 27918 76692 27970
rect 76636 27906 76692 27918
rect 76748 27970 76804 27982
rect 76748 27918 76750 27970
rect 76802 27918 76804 27970
rect 76748 27860 76804 27918
rect 76748 27794 76804 27804
rect 76860 27858 76916 27870
rect 76860 27806 76862 27858
rect 76914 27806 76916 27858
rect 76860 27636 76916 27806
rect 77084 27858 77140 28140
rect 77084 27806 77086 27858
rect 77138 27806 77140 27858
rect 77084 27748 77140 27806
rect 76860 27570 76916 27580
rect 76972 27692 77140 27748
rect 77196 28418 77252 28430
rect 77196 28366 77198 28418
rect 77250 28366 77252 28418
rect 76524 27458 76580 27468
rect 75740 27356 76244 27412
rect 76188 27300 76244 27356
rect 76860 27300 76916 27310
rect 76188 27244 76468 27300
rect 76412 27076 76468 27244
rect 76860 27206 76916 27244
rect 76972 27076 77028 27692
rect 77196 27524 77252 28366
rect 76412 27074 76580 27076
rect 76412 27022 76414 27074
rect 76466 27022 76580 27074
rect 76412 27020 76580 27022
rect 76412 27010 76468 27020
rect 75404 26852 75572 26908
rect 75628 26962 75684 26974
rect 75628 26910 75630 26962
rect 75682 26910 75684 26962
rect 75628 26908 75684 26910
rect 76188 26964 76244 27002
rect 75628 26852 75796 26908
rect 76188 26898 76244 26908
rect 75292 26292 75348 26302
rect 75404 26292 75460 26852
rect 75292 26290 75460 26292
rect 75292 26238 75294 26290
rect 75346 26238 75460 26290
rect 75292 26236 75460 26238
rect 75516 26402 75572 26414
rect 75516 26350 75518 26402
rect 75570 26350 75572 26402
rect 75292 26226 75348 26236
rect 75404 25506 75460 25518
rect 75404 25454 75406 25506
rect 75458 25454 75460 25506
rect 75404 25396 75460 25454
rect 75404 25330 75460 25340
rect 75180 24724 75236 24734
rect 75180 24630 75236 24668
rect 75292 24052 75348 24062
rect 75292 23958 75348 23996
rect 75404 23716 75460 23726
rect 74956 23154 75124 23156
rect 74956 23102 74958 23154
rect 75010 23102 75124 23154
rect 74956 23100 75124 23102
rect 75180 23714 75460 23716
rect 75180 23662 75406 23714
rect 75458 23662 75460 23714
rect 75180 23660 75460 23662
rect 74956 23090 75012 23100
rect 74844 22318 74846 22370
rect 74898 22318 74900 22370
rect 74844 22306 74900 22318
rect 74956 21588 75012 21598
rect 75012 21532 75124 21588
rect 74956 21494 75012 21532
rect 75068 20914 75124 21532
rect 75068 20862 75070 20914
rect 75122 20862 75124 20914
rect 75068 20850 75124 20862
rect 74732 20178 74788 20188
rect 75068 20132 75124 20142
rect 75068 20038 75124 20076
rect 74844 20018 74900 20030
rect 74844 19966 74846 20018
rect 74898 19966 74900 20018
rect 74844 19796 74900 19966
rect 74900 19740 75124 19796
rect 74844 19730 74900 19740
rect 75068 19346 75124 19740
rect 75068 19294 75070 19346
rect 75122 19294 75124 19346
rect 75068 19282 75124 19294
rect 74620 18050 74676 18060
rect 72156 16930 72212 16940
rect 75180 16884 75236 23660
rect 75404 23650 75460 23660
rect 75404 22370 75460 22382
rect 75404 22318 75406 22370
rect 75458 22318 75460 22370
rect 75292 21476 75348 21486
rect 75292 21026 75348 21420
rect 75292 20974 75294 21026
rect 75346 20974 75348 21026
rect 75292 20962 75348 20974
rect 75404 21028 75460 22318
rect 75404 20962 75460 20972
rect 75292 20802 75348 20814
rect 75292 20750 75294 20802
rect 75346 20750 75348 20802
rect 75292 17444 75348 20750
rect 75404 19908 75460 19918
rect 75404 19814 75460 19852
rect 75404 19012 75460 19022
rect 75404 18918 75460 18956
rect 75292 17378 75348 17388
rect 71036 16258 71092 16268
rect 74284 16828 75236 16884
rect 70252 16146 70308 16156
rect 69692 15204 69748 15214
rect 69692 6692 69748 15148
rect 71372 14420 71428 14430
rect 69692 6626 69748 6636
rect 69804 9380 69860 9390
rect 69244 6580 69300 6590
rect 69244 6356 69300 6524
rect 69356 6468 69412 6478
rect 69356 6374 69412 6412
rect 69244 6290 69300 6300
rect 68572 6066 68628 6076
rect 68460 5070 68462 5122
rect 68514 5070 68516 5122
rect 68460 5058 68516 5070
rect 68908 5794 68964 5806
rect 68908 5742 68910 5794
rect 68962 5742 68964 5794
rect 68348 4116 68404 4126
rect 68348 4022 68404 4060
rect 68796 3892 68852 3902
rect 68796 800 68852 3836
rect 68908 3556 68964 5742
rect 69356 5348 69412 5358
rect 69356 5254 69412 5292
rect 68908 3490 68964 3500
rect 69468 3780 69524 3790
rect 69468 800 69524 3724
rect 69804 3668 69860 9324
rect 71260 6692 71316 6702
rect 71036 6636 71260 6692
rect 70476 6468 70532 6478
rect 70364 6412 70476 6468
rect 69804 3666 70308 3668
rect 69804 3614 69806 3666
rect 69858 3614 70308 3666
rect 69804 3612 70308 3614
rect 69804 3602 69860 3612
rect 70252 3554 70308 3612
rect 70252 3502 70254 3554
rect 70306 3502 70308 3554
rect 70252 3490 70308 3502
rect 70364 3220 70420 6412
rect 70476 6402 70532 6412
rect 71036 6130 71092 6636
rect 71260 6598 71316 6636
rect 71036 6078 71038 6130
rect 71090 6078 71092 6130
rect 71036 6066 71092 6078
rect 70476 5796 70532 5806
rect 70476 5348 70532 5740
rect 70476 5282 70532 5292
rect 70812 5684 70868 5694
rect 70476 4226 70532 4238
rect 70476 4174 70478 4226
rect 70530 4174 70532 4226
rect 70476 4004 70532 4174
rect 70476 3938 70532 3948
rect 70140 3164 70420 3220
rect 70140 800 70196 3164
rect 70812 800 70868 5628
rect 71372 5124 71428 14364
rect 73052 12740 73108 12750
rect 71708 7812 71764 7822
rect 71708 7698 71764 7756
rect 71708 7646 71710 7698
rect 71762 7646 71764 7698
rect 71708 7634 71764 7646
rect 72380 7812 72436 7822
rect 72380 7474 72436 7756
rect 72380 7422 72382 7474
rect 72434 7422 72436 7474
rect 72380 7410 72436 7422
rect 72268 6468 72324 6478
rect 72268 6374 72324 6412
rect 71708 5908 71764 5918
rect 71708 5814 71764 5852
rect 72268 5908 72324 5918
rect 72268 5814 72324 5852
rect 72828 5796 72884 5806
rect 72268 5236 72324 5246
rect 72268 5142 72324 5180
rect 71036 5122 71428 5124
rect 71036 5070 71374 5122
rect 71426 5070 71428 5122
rect 71036 5068 71428 5070
rect 71036 4562 71092 5068
rect 71372 5058 71428 5068
rect 72156 5124 72212 5134
rect 71036 4510 71038 4562
rect 71090 4510 71092 4562
rect 71036 4498 71092 4510
rect 71708 4564 71764 4574
rect 71708 4470 71764 4508
rect 71484 4116 71540 4126
rect 71260 3668 71316 3678
rect 71260 3574 71316 3612
rect 71484 800 71540 4060
rect 72156 800 72212 5068
rect 72268 4564 72324 4574
rect 72268 4338 72324 4508
rect 72268 4286 72270 4338
rect 72322 4286 72324 4338
rect 72268 4274 72324 4286
rect 72828 800 72884 5740
rect 73052 4228 73108 12684
rect 73836 8818 73892 8830
rect 73836 8766 73838 8818
rect 73890 8766 73892 8818
rect 73612 8372 73668 8382
rect 73612 6244 73668 8316
rect 73612 6178 73668 6188
rect 73276 5684 73332 5694
rect 73276 5590 73332 5628
rect 73052 4162 73108 4172
rect 73500 5236 73556 5246
rect 73276 4114 73332 4126
rect 73276 4062 73278 4114
rect 73330 4062 73332 4114
rect 73276 3892 73332 4062
rect 73276 3826 73332 3836
rect 73500 800 73556 5180
rect 73836 4900 73892 8766
rect 74284 8428 74340 16828
rect 75516 15148 75572 26350
rect 75628 25282 75684 25294
rect 75628 25230 75630 25282
rect 75682 25230 75684 25282
rect 75628 24948 75684 25230
rect 75740 25172 75796 26852
rect 76188 26516 76244 26526
rect 76188 26422 76244 26460
rect 76524 26290 76580 27020
rect 76860 27020 77028 27076
rect 77084 27468 77252 27524
rect 76748 26516 76804 26526
rect 76860 26516 76916 27020
rect 76748 26514 76916 26516
rect 76748 26462 76750 26514
rect 76802 26462 76916 26514
rect 76748 26460 76916 26462
rect 76972 26850 77028 26862
rect 76972 26798 76974 26850
rect 77026 26798 77028 26850
rect 76748 26450 76804 26460
rect 76524 26238 76526 26290
rect 76578 26238 76580 26290
rect 76524 26226 76580 26238
rect 75740 25106 75796 25116
rect 75852 26180 75908 26190
rect 75628 24882 75684 24892
rect 75852 24946 75908 26124
rect 76972 25844 77028 26798
rect 76972 25778 77028 25788
rect 76524 25508 76580 25518
rect 77084 25508 77140 27468
rect 77196 27300 77252 27310
rect 77196 27206 77252 27244
rect 77308 26514 77364 30044
rect 77420 30098 77476 31612
rect 77532 31218 77588 31724
rect 77532 31166 77534 31218
rect 77586 31166 77588 31218
rect 77532 31154 77588 31166
rect 77756 31554 77812 31566
rect 77756 31502 77758 31554
rect 77810 31502 77812 31554
rect 77420 30046 77422 30098
rect 77474 30046 77476 30098
rect 77420 30034 77476 30046
rect 77532 30548 77588 30558
rect 77532 29428 77588 30492
rect 77644 30436 77700 30446
rect 77644 29650 77700 30380
rect 77756 30324 77812 31502
rect 77868 31108 77924 31724
rect 78092 31220 78148 34412
rect 78204 34356 78260 34366
rect 78204 34262 78260 34300
rect 78204 33460 78260 33470
rect 78204 33366 78260 33404
rect 78316 32788 78372 35420
rect 78092 31154 78148 31164
rect 78204 32732 78372 32788
rect 78204 32562 78260 32732
rect 78428 32676 78484 55412
rect 78540 38388 78596 58380
rect 78540 38322 78596 38332
rect 78540 37492 78596 37502
rect 78540 33460 78596 37436
rect 78652 35812 78708 67172
rect 78652 35746 78708 35756
rect 78764 34468 78820 71820
rect 78876 71092 78932 71102
rect 78876 67228 78932 71036
rect 78876 67172 79492 67228
rect 78764 34402 78820 34412
rect 78876 64708 78932 64718
rect 78540 33394 78596 33404
rect 78204 32510 78206 32562
rect 78258 32510 78260 32562
rect 77868 31106 78036 31108
rect 77868 31054 77870 31106
rect 77922 31054 78036 31106
rect 77868 31052 78036 31054
rect 77868 31042 77924 31052
rect 77756 30268 77924 30324
rect 77868 30098 77924 30268
rect 77868 30046 77870 30098
rect 77922 30046 77924 30098
rect 77868 30034 77924 30046
rect 77868 29876 77924 29886
rect 77644 29598 77646 29650
rect 77698 29598 77700 29650
rect 77644 29586 77700 29598
rect 77756 29652 77812 29662
rect 77756 29558 77812 29596
rect 77532 29372 77812 29428
rect 77532 29202 77588 29214
rect 77532 29150 77534 29202
rect 77586 29150 77588 29202
rect 77420 28980 77476 28990
rect 77420 28642 77476 28924
rect 77420 28590 77422 28642
rect 77474 28590 77476 28642
rect 77420 28308 77476 28590
rect 77420 28242 77476 28252
rect 77532 27970 77588 29150
rect 77644 28644 77700 28654
rect 77644 28550 77700 28588
rect 77756 28420 77812 29372
rect 77868 28532 77924 29820
rect 77868 28466 77924 28476
rect 77644 28364 77812 28420
rect 77644 28082 77700 28364
rect 77644 28030 77646 28082
rect 77698 28030 77700 28082
rect 77644 28018 77700 28030
rect 77532 27918 77534 27970
rect 77586 27918 77588 27970
rect 77532 27300 77588 27918
rect 77756 27972 77812 27982
rect 77756 27878 77812 27916
rect 77308 26462 77310 26514
rect 77362 26462 77364 26514
rect 77308 26450 77364 26462
rect 77420 27076 77476 27086
rect 75852 24894 75854 24946
rect 75906 24894 75908 24946
rect 75852 24882 75908 24894
rect 76188 25394 76244 25406
rect 76188 25342 76190 25394
rect 76242 25342 76244 25394
rect 76188 25284 76244 25342
rect 76524 25394 76580 25452
rect 76524 25342 76526 25394
rect 76578 25342 76580 25394
rect 76524 25330 76580 25342
rect 76972 25452 77140 25508
rect 77420 25508 77476 27020
rect 77532 26962 77588 27244
rect 77868 27076 77924 27086
rect 77980 27076 78036 31052
rect 78092 30772 78148 30782
rect 78204 30772 78260 32510
rect 78148 30716 78260 30772
rect 78316 32620 78428 32676
rect 78092 30706 78148 30716
rect 78204 30212 78260 30222
rect 78204 29092 78260 30156
rect 78204 29026 78260 29036
rect 78204 28756 78260 28766
rect 78316 28756 78372 32620
rect 78428 32610 78484 32620
rect 78540 33236 78596 33246
rect 78540 30212 78596 33180
rect 78540 30146 78596 30156
rect 78876 30100 78932 64652
rect 78988 50372 79044 50382
rect 79044 50316 79268 50372
rect 78988 50306 79044 50316
rect 78988 48804 79044 48814
rect 78988 35252 79044 48748
rect 78988 35186 79044 35196
rect 79100 33572 79156 33582
rect 79212 33572 79268 50316
rect 79436 38668 79492 67172
rect 79324 38612 79492 38668
rect 79324 35028 79380 38612
rect 79324 34962 79380 34972
rect 79436 38388 79492 38398
rect 79156 33516 79268 33572
rect 79100 33506 79156 33516
rect 78876 30034 78932 30044
rect 79436 29764 79492 38332
rect 79100 29708 79492 29764
rect 79100 28980 79156 29708
rect 79100 28914 79156 28924
rect 78204 28754 78372 28756
rect 78204 28702 78206 28754
rect 78258 28702 78372 28754
rect 78204 28700 78372 28702
rect 78204 28690 78260 28700
rect 77924 27020 78036 27076
rect 78204 27636 78260 27646
rect 77868 26982 77924 27020
rect 77532 26910 77534 26962
rect 77586 26910 77588 26962
rect 77532 26290 77588 26910
rect 77756 26740 77812 26750
rect 77756 26514 77812 26684
rect 77756 26462 77758 26514
rect 77810 26462 77812 26514
rect 77756 26450 77812 26462
rect 77532 26238 77534 26290
rect 77586 26238 77588 26290
rect 77532 26226 77588 26238
rect 77644 26292 77700 26302
rect 77644 26198 77700 26236
rect 75740 24834 75796 24846
rect 75740 24782 75742 24834
rect 75794 24782 75796 24834
rect 75628 24724 75684 24734
rect 75628 24052 75684 24668
rect 75740 24500 75796 24782
rect 75740 24276 75796 24444
rect 75740 24210 75796 24220
rect 75964 24498 76020 24510
rect 75964 24446 75966 24498
rect 76018 24446 76020 24498
rect 75628 23996 75796 24052
rect 75628 23826 75684 23838
rect 75628 23774 75630 23826
rect 75682 23774 75684 23826
rect 75628 23266 75684 23774
rect 75740 23378 75796 23996
rect 75964 23716 76020 24446
rect 76188 24052 76244 25228
rect 76524 25060 76580 25070
rect 76524 24946 76580 25004
rect 76524 24894 76526 24946
rect 76578 24894 76580 24946
rect 76524 24882 76580 24894
rect 76524 24724 76580 24734
rect 76860 24724 76916 24734
rect 76412 24500 76468 24510
rect 76188 23996 76356 24052
rect 76188 23828 76244 23838
rect 76188 23716 76244 23772
rect 75740 23326 75742 23378
rect 75794 23326 75796 23378
rect 75740 23314 75796 23326
rect 75852 23660 76244 23716
rect 75628 23214 75630 23266
rect 75682 23214 75684 23266
rect 75628 23156 75684 23214
rect 75852 23156 75908 23660
rect 76188 23492 76244 23502
rect 75628 23100 75908 23156
rect 75964 23156 76020 23166
rect 75964 23154 76132 23156
rect 75964 23102 75966 23154
rect 76018 23102 76132 23154
rect 75964 23100 76132 23102
rect 75964 23090 76020 23100
rect 75740 22036 75796 22046
rect 75740 21588 75796 21980
rect 76076 21924 76132 23100
rect 76188 22370 76244 23436
rect 76188 22318 76190 22370
rect 76242 22318 76244 22370
rect 76188 22306 76244 22318
rect 76300 22036 76356 23996
rect 76412 24050 76468 24444
rect 76412 23998 76414 24050
rect 76466 23998 76468 24050
rect 76412 23986 76468 23998
rect 76300 21970 76356 21980
rect 76412 23714 76468 23726
rect 76412 23662 76414 23714
rect 76466 23662 76468 23714
rect 76076 21868 76244 21924
rect 76076 21700 76132 21710
rect 76076 21606 76132 21644
rect 75740 21494 75796 21532
rect 75628 20690 75684 20702
rect 75628 20638 75630 20690
rect 75682 20638 75684 20690
rect 75628 20356 75684 20638
rect 75628 20300 76020 20356
rect 75628 20130 75684 20142
rect 75628 20078 75630 20130
rect 75682 20078 75684 20130
rect 75628 16996 75684 20078
rect 75964 20132 76020 20300
rect 76076 20132 76132 20142
rect 75964 20130 76132 20132
rect 75964 20078 76078 20130
rect 76130 20078 76132 20130
rect 75964 20076 76132 20078
rect 75740 20020 75796 20030
rect 75740 19906 75796 19964
rect 75740 19854 75742 19906
rect 75794 19854 75796 19906
rect 75740 19842 75796 19854
rect 75964 19908 76020 20076
rect 76076 20066 76132 20076
rect 75964 19124 76020 19852
rect 75964 19058 76020 19068
rect 76076 19348 76132 19358
rect 75628 16930 75684 16940
rect 75180 15092 75572 15148
rect 74620 14756 74676 14766
rect 74620 12404 74676 14700
rect 75180 12404 75236 15092
rect 76076 13524 76132 19292
rect 76188 13972 76244 21868
rect 76300 21700 76356 21710
rect 76300 20018 76356 21644
rect 76412 20468 76468 23662
rect 76524 23378 76580 24668
rect 76524 23326 76526 23378
rect 76578 23326 76580 23378
rect 76524 23314 76580 23326
rect 76636 24722 76916 24724
rect 76636 24670 76862 24722
rect 76914 24670 76916 24722
rect 76636 24668 76916 24670
rect 76524 22260 76580 22270
rect 76636 22260 76692 24668
rect 76860 24658 76916 24668
rect 76860 24500 76916 24510
rect 76860 24406 76916 24444
rect 76972 24164 77028 25452
rect 77420 25414 77476 25452
rect 77644 26068 77700 26078
rect 77084 25282 77140 25294
rect 77084 25230 77086 25282
rect 77138 25230 77140 25282
rect 77084 25172 77140 25230
rect 77140 25116 77252 25172
rect 77084 25106 77140 25116
rect 77196 24836 77252 25116
rect 77644 24946 77700 26012
rect 77868 25844 77924 25854
rect 77868 25394 77924 25788
rect 78204 25732 78260 27580
rect 78204 25506 78260 25676
rect 78204 25454 78206 25506
rect 78258 25454 78260 25506
rect 78204 25442 78260 25454
rect 77868 25342 77870 25394
rect 77922 25342 77924 25394
rect 77868 25330 77924 25342
rect 77644 24894 77646 24946
rect 77698 24894 77700 24946
rect 77644 24882 77700 24894
rect 77756 24948 77812 24958
rect 77532 24836 77588 24846
rect 77196 24834 77588 24836
rect 77196 24782 77198 24834
rect 77250 24782 77534 24834
rect 77586 24782 77588 24834
rect 77196 24780 77588 24782
rect 77196 24770 77252 24780
rect 76972 24108 77252 24164
rect 77084 23940 77140 23950
rect 76972 23938 77140 23940
rect 76972 23886 77086 23938
rect 77138 23886 77140 23938
rect 76972 23884 77140 23886
rect 76748 23828 76804 23838
rect 76804 23772 76916 23828
rect 76748 23762 76804 23772
rect 76860 23714 76916 23772
rect 76860 23662 76862 23714
rect 76914 23662 76916 23714
rect 76860 23650 76916 23662
rect 76524 22258 76692 22260
rect 76524 22206 76526 22258
rect 76578 22206 76692 22258
rect 76524 22204 76692 22206
rect 76748 23268 76804 23278
rect 76972 23268 77028 23884
rect 77084 23874 77140 23884
rect 77196 23604 77252 24108
rect 77532 24162 77588 24780
rect 77532 24110 77534 24162
rect 77586 24110 77588 24162
rect 77532 24098 77588 24110
rect 77644 24724 77700 24734
rect 77644 23940 77700 24668
rect 77196 23538 77252 23548
rect 77532 23884 77700 23940
rect 77532 23492 77588 23884
rect 77756 23826 77812 24892
rect 77868 24724 77924 24734
rect 77868 24722 78036 24724
rect 77868 24670 77870 24722
rect 77922 24670 78036 24722
rect 77868 24668 78036 24670
rect 77868 24658 77924 24668
rect 77756 23774 77758 23826
rect 77810 23774 77812 23826
rect 77756 23762 77812 23774
rect 77644 23716 77700 23726
rect 77644 23622 77700 23660
rect 77532 23436 77700 23492
rect 77644 23378 77700 23436
rect 77644 23326 77646 23378
rect 77698 23326 77700 23378
rect 77644 23314 77700 23326
rect 76748 23266 77028 23268
rect 76748 23214 76750 23266
rect 76802 23214 77028 23266
rect 76748 23212 77028 23214
rect 77084 23268 77140 23278
rect 77532 23268 77588 23278
rect 77084 23266 77588 23268
rect 77084 23214 77086 23266
rect 77138 23214 77534 23266
rect 77586 23214 77588 23266
rect 77084 23212 77588 23214
rect 76524 22194 76580 22204
rect 76748 22036 76804 23212
rect 77084 23202 77140 23212
rect 76860 23044 76916 23054
rect 76860 22594 76916 22988
rect 76860 22542 76862 22594
rect 76914 22542 76916 22594
rect 76860 22530 76916 22542
rect 77196 22594 77252 23212
rect 77196 22542 77198 22594
rect 77250 22542 77252 22594
rect 77196 22530 77252 22542
rect 77532 22594 77588 23212
rect 77532 22542 77534 22594
rect 77586 22542 77588 22594
rect 76972 22148 77028 22158
rect 76636 21980 76804 22036
rect 76860 22146 77028 22148
rect 76860 22094 76974 22146
rect 77026 22094 77028 22146
rect 76860 22092 77028 22094
rect 76636 21700 76692 21980
rect 76860 21812 76916 22092
rect 76972 22082 77028 22092
rect 76636 21606 76692 21644
rect 76748 21756 76916 21812
rect 76524 21028 76580 21038
rect 76524 20934 76580 20972
rect 76748 20804 76804 21756
rect 76972 21700 77028 21710
rect 76412 20402 76468 20412
rect 76524 20748 76804 20804
rect 76860 21698 77028 21700
rect 76860 21646 76974 21698
rect 77026 21646 77028 21698
rect 76860 21644 77028 21646
rect 76860 21028 76916 21644
rect 76972 21634 77028 21644
rect 77532 21698 77588 22542
rect 77644 23156 77700 23166
rect 77644 22482 77700 23100
rect 77644 22430 77646 22482
rect 77698 22430 77700 22482
rect 77644 22418 77700 22430
rect 77868 23154 77924 23166
rect 77868 23102 77870 23154
rect 77922 23102 77924 23154
rect 77756 22148 77812 22158
rect 77532 21646 77534 21698
rect 77586 21646 77588 21698
rect 77532 21634 77588 21646
rect 77644 22146 77812 22148
rect 77644 22094 77758 22146
rect 77810 22094 77812 22146
rect 77644 22092 77812 22094
rect 77196 21028 77252 21038
rect 77644 21028 77700 22092
rect 77756 22082 77812 22092
rect 77868 22148 77924 23102
rect 77868 22082 77924 22092
rect 77868 21812 77924 21822
rect 77756 21700 77812 21710
rect 77756 21606 77812 21644
rect 77868 21474 77924 21756
rect 77868 21422 77870 21474
rect 77922 21422 77924 21474
rect 77868 21410 77924 21422
rect 77980 21252 78036 24668
rect 78540 24276 78596 24286
rect 78316 23492 78372 23502
rect 76860 21026 77252 21028
rect 76860 20974 76862 21026
rect 76914 20974 77198 21026
rect 77250 20974 77252 21026
rect 76860 20972 77252 20974
rect 76300 19966 76302 20018
rect 76354 19966 76356 20018
rect 76300 19954 76356 19966
rect 76412 20020 76468 20030
rect 76412 15148 76468 19964
rect 76524 19348 76580 20748
rect 76524 19282 76580 19292
rect 76636 20578 76692 20590
rect 76636 20526 76638 20578
rect 76690 20526 76692 20578
rect 76636 19236 76692 20526
rect 76748 20132 76804 20142
rect 76860 20132 76916 20972
rect 77196 20962 77252 20972
rect 77420 20972 77700 21028
rect 77868 21196 78036 21252
rect 78204 23156 78260 23166
rect 77308 20916 77364 20926
rect 77308 20822 77364 20860
rect 76748 20130 76916 20132
rect 76748 20078 76750 20130
rect 76802 20078 76916 20130
rect 76748 20076 76916 20078
rect 76748 20066 76804 20076
rect 76860 20020 76916 20076
rect 76860 19954 76916 19964
rect 76972 20244 77028 20254
rect 77420 20244 77476 20972
rect 77532 20804 77588 20814
rect 77532 20710 77588 20748
rect 77868 20690 77924 21196
rect 77868 20638 77870 20690
rect 77922 20638 77924 20690
rect 77868 20626 77924 20638
rect 77980 20916 78036 20926
rect 76972 19906 77028 20188
rect 77308 20188 77476 20244
rect 77084 20020 77140 20030
rect 77084 20018 77252 20020
rect 77084 19966 77086 20018
rect 77138 19966 77252 20018
rect 77084 19964 77252 19966
rect 77084 19954 77140 19964
rect 76972 19854 76974 19906
rect 77026 19854 77028 19906
rect 76972 19842 77028 19854
rect 76860 19236 76916 19246
rect 76636 19180 76804 19236
rect 76524 19124 76580 19134
rect 76524 18564 76580 19068
rect 76636 19010 76692 19022
rect 76636 18958 76638 19010
rect 76690 18958 76692 19010
rect 76636 18900 76692 18958
rect 76748 19012 76804 19180
rect 76860 19234 77140 19236
rect 76860 19182 76862 19234
rect 76914 19182 77140 19234
rect 76860 19180 77140 19182
rect 76860 19170 76916 19180
rect 76748 18946 76804 18956
rect 76636 18834 76692 18844
rect 76748 18676 76804 18686
rect 76748 18582 76804 18620
rect 76524 18498 76580 18508
rect 76972 17556 77028 17566
rect 77084 17556 77140 19180
rect 77196 19122 77252 19964
rect 77196 19070 77198 19122
rect 77250 19070 77252 19122
rect 77196 19058 77252 19070
rect 77196 18900 77252 18910
rect 77196 18450 77252 18844
rect 77196 18398 77198 18450
rect 77250 18398 77252 18450
rect 77196 18386 77252 18398
rect 77196 17556 77252 17566
rect 77084 17554 77252 17556
rect 77084 17502 77198 17554
rect 77250 17502 77252 17554
rect 77084 17500 77252 17502
rect 76972 17462 77028 17500
rect 77196 17490 77252 17500
rect 77308 17332 77364 20188
rect 77644 20132 77700 20142
rect 77644 20038 77700 20076
rect 77420 20020 77476 20030
rect 77420 19926 77476 19964
rect 77644 19908 77700 19918
rect 77644 19814 77700 19852
rect 77532 19124 77588 19134
rect 77532 18676 77588 19068
rect 77980 19124 78036 20860
rect 77980 19058 78036 19068
rect 78092 20804 78148 20814
rect 77868 19012 77924 19022
rect 77868 18918 77924 18956
rect 78092 18676 78148 20748
rect 78204 20802 78260 23100
rect 78204 20750 78206 20802
rect 78258 20750 78260 20802
rect 78204 19684 78260 20750
rect 78316 20130 78372 23436
rect 78316 20078 78318 20130
rect 78370 20078 78372 20130
rect 78316 20066 78372 20078
rect 78428 22036 78484 22046
rect 78204 19628 78372 19684
rect 78204 19236 78260 19246
rect 78204 18900 78260 19180
rect 78204 18834 78260 18844
rect 77532 18610 77588 18620
rect 77868 18620 78148 18676
rect 78204 18676 78260 18686
rect 77420 18564 77476 18574
rect 77420 18470 77476 18508
rect 77756 18452 77812 18490
rect 77756 18386 77812 18396
rect 77756 18228 77812 18238
rect 77756 18134 77812 18172
rect 77644 17668 77700 17678
rect 77532 17556 77588 17566
rect 77532 17462 77588 17500
rect 77308 17266 77364 17276
rect 77532 17220 77588 17230
rect 77308 16996 77364 17006
rect 77196 16884 77252 16894
rect 77196 16790 77252 16828
rect 76300 15092 76468 15148
rect 76300 14308 76356 15092
rect 77308 14420 77364 16940
rect 77308 14354 77364 14364
rect 77420 16772 77476 16782
rect 76300 14252 76580 14308
rect 76300 13972 76356 13982
rect 76188 13916 76300 13972
rect 76300 13906 76356 13916
rect 76076 13458 76132 13468
rect 74620 12402 75012 12404
rect 74620 12350 74622 12402
rect 74674 12350 75012 12402
rect 74620 12348 75012 12350
rect 74620 12338 74676 12348
rect 74956 12178 75012 12348
rect 74956 12126 74958 12178
rect 75010 12126 75012 12178
rect 74956 12114 75012 12126
rect 75180 12178 75236 12348
rect 75964 12404 76020 12414
rect 76020 12348 76356 12404
rect 75964 12310 76020 12348
rect 75180 12126 75182 12178
rect 75234 12126 75236 12178
rect 75180 12114 75236 12126
rect 75516 11954 75572 11966
rect 75516 11902 75518 11954
rect 75570 11902 75572 11954
rect 75516 11396 75572 11902
rect 75516 11330 75572 11340
rect 76188 11170 76244 11182
rect 76188 11118 76190 11170
rect 76242 11118 76244 11170
rect 75852 10386 75908 10398
rect 75852 10334 75854 10386
rect 75906 10334 75908 10386
rect 74060 8372 74340 8428
rect 74844 9602 74900 9614
rect 74844 9550 74846 9602
rect 74898 9550 74900 9602
rect 74844 8428 74900 9550
rect 75292 9604 75348 9642
rect 75292 9538 75348 9548
rect 75628 9604 75684 9614
rect 75628 9602 75796 9604
rect 75628 9550 75630 9602
rect 75682 9550 75796 9602
rect 75628 9548 75796 9550
rect 75628 9538 75684 9548
rect 75292 9380 75348 9390
rect 75180 9042 75236 9054
rect 75180 8990 75182 9042
rect 75234 8990 75236 9042
rect 74844 8372 75124 8428
rect 74060 8148 74116 8372
rect 74060 8082 74116 8092
rect 74620 8034 74676 8046
rect 74620 7982 74622 8034
rect 74674 7982 74676 8034
rect 73948 7362 74004 7374
rect 73948 7310 73950 7362
rect 74002 7310 74004 7362
rect 73948 5124 74004 7310
rect 73948 5058 74004 5068
rect 73836 4844 74004 4900
rect 73612 3444 73668 3454
rect 73612 3350 73668 3388
rect 73948 2996 74004 4844
rect 74172 4228 74228 4238
rect 74060 4004 74116 4014
rect 74060 3554 74116 3948
rect 74060 3502 74062 3554
rect 74114 3502 74116 3554
rect 74060 3490 74116 3502
rect 74060 2996 74116 3006
rect 73948 2940 74060 2996
rect 74060 2930 74116 2940
rect 74172 800 74228 4172
rect 74620 980 74676 7982
rect 74732 7700 74788 7710
rect 74732 6802 74788 7644
rect 74732 6750 74734 6802
rect 74786 6750 74788 6802
rect 74732 6738 74788 6750
rect 74956 6690 75012 6702
rect 74956 6638 74958 6690
rect 75010 6638 75012 6690
rect 74956 6580 75012 6638
rect 74732 6524 74956 6580
rect 74732 5234 74788 6524
rect 74956 6514 75012 6524
rect 75068 5460 75124 8372
rect 75180 6916 75236 8990
rect 75292 8258 75348 9324
rect 75740 8428 75796 9548
rect 75292 8206 75294 8258
rect 75346 8206 75348 8258
rect 75292 8194 75348 8206
rect 75628 8372 75796 8428
rect 75628 8260 75684 8372
rect 75628 8194 75684 8204
rect 75292 7700 75348 7710
rect 75292 7474 75348 7644
rect 75292 7422 75294 7474
rect 75346 7422 75348 7474
rect 75292 7410 75348 7422
rect 75180 6850 75236 6860
rect 75292 6804 75348 6814
rect 75852 6804 75908 10334
rect 76188 9380 76244 11118
rect 76188 9314 76244 9324
rect 76300 9938 76356 12348
rect 76412 11396 76468 11406
rect 76412 11302 76468 11340
rect 76300 9886 76302 9938
rect 76354 9886 76356 9938
rect 75180 6692 75236 6702
rect 75292 6692 75348 6748
rect 75180 6690 75348 6692
rect 75180 6638 75182 6690
rect 75234 6638 75348 6690
rect 75180 6636 75348 6638
rect 75404 6748 75908 6804
rect 76076 9042 76132 9054
rect 76076 8990 76078 9042
rect 76130 8990 76132 9042
rect 75180 6626 75236 6636
rect 75068 5394 75124 5404
rect 74732 5182 74734 5234
rect 74786 5182 74788 5234
rect 74732 5170 74788 5182
rect 75180 5348 75236 5358
rect 75068 5124 75124 5134
rect 74956 5122 75124 5124
rect 74956 5070 75070 5122
rect 75122 5070 75124 5122
rect 74956 5068 75124 5070
rect 74620 914 74676 924
rect 74844 3444 74900 3454
rect 74956 3444 75012 5068
rect 75068 5058 75124 5068
rect 75180 4338 75236 5292
rect 75180 4286 75182 4338
rect 75234 4286 75236 4338
rect 75180 4274 75236 4286
rect 75068 3780 75124 3790
rect 75068 3686 75124 3724
rect 74900 3388 75012 3444
rect 74844 800 74900 3388
rect 75404 1876 75460 6748
rect 75516 6468 75572 6478
rect 75516 6374 75572 6412
rect 75516 6244 75572 6254
rect 75516 5234 75572 6188
rect 76076 6132 76132 8990
rect 76188 8260 76244 8270
rect 76188 6690 76244 8204
rect 76300 7476 76356 9886
rect 76524 8260 76580 14252
rect 77084 13972 77140 13982
rect 76524 8194 76580 8204
rect 76860 8372 76916 8382
rect 76412 8148 76468 8158
rect 76412 8036 76468 8092
rect 76860 8146 76916 8316
rect 76860 8094 76862 8146
rect 76914 8094 76916 8146
rect 76524 8036 76580 8046
rect 76412 8034 76580 8036
rect 76412 7982 76526 8034
rect 76578 7982 76580 8034
rect 76412 7980 76580 7982
rect 76524 7970 76580 7980
rect 76300 7420 76468 7476
rect 76188 6638 76190 6690
rect 76242 6638 76244 6690
rect 76188 6626 76244 6638
rect 76300 7250 76356 7262
rect 76300 7198 76302 7250
rect 76354 7198 76356 7250
rect 76076 6076 76244 6132
rect 75628 5796 75684 5806
rect 75628 5702 75684 5740
rect 75516 5182 75518 5234
rect 75570 5182 75572 5234
rect 75516 5170 75572 5182
rect 76188 5010 76244 6076
rect 76300 5236 76356 7198
rect 76412 6804 76468 7420
rect 76412 6710 76468 6748
rect 76860 6580 76916 8094
rect 77084 8148 77140 13916
rect 77196 11170 77252 11182
rect 77196 11118 77198 11170
rect 77250 11118 77252 11170
rect 77196 9828 77252 11118
rect 77420 10612 77476 16716
rect 77532 13412 77588 17164
rect 77644 17106 77700 17612
rect 77868 17554 77924 18620
rect 77868 17502 77870 17554
rect 77922 17502 77924 17554
rect 77868 17490 77924 17502
rect 77980 18452 78036 18462
rect 77868 17332 77924 17342
rect 77644 17054 77646 17106
rect 77698 17054 77700 17106
rect 77644 17042 77700 17054
rect 77756 17276 77868 17332
rect 77644 15876 77700 15886
rect 77644 15782 77700 15820
rect 77644 14306 77700 14318
rect 77644 14254 77646 14306
rect 77698 14254 77700 14306
rect 77644 14196 77700 14254
rect 77644 14130 77700 14140
rect 77756 13972 77812 17276
rect 77868 17266 77924 17276
rect 77868 17108 77924 17118
rect 77980 17108 78036 18396
rect 78204 17668 78260 18620
rect 78316 18450 78372 19628
rect 78428 19236 78484 21980
rect 78428 19170 78484 19180
rect 78316 18398 78318 18450
rect 78370 18398 78372 18450
rect 78316 18386 78372 18398
rect 78204 17574 78260 17612
rect 77868 17106 78036 17108
rect 77868 17054 77870 17106
rect 77922 17054 78036 17106
rect 77868 17052 78036 17054
rect 78204 17444 78260 17454
rect 77868 17042 77924 17052
rect 78092 16884 78148 16894
rect 78092 16790 78148 16828
rect 78204 16660 78260 17388
rect 77868 16604 78260 16660
rect 77868 15986 77924 16604
rect 77868 15934 77870 15986
rect 77922 15934 77924 15986
rect 77868 15922 77924 15934
rect 78204 15986 78260 15998
rect 78204 15934 78206 15986
rect 78258 15934 78260 15986
rect 78204 15876 78260 15934
rect 78204 15316 78260 15820
rect 78204 15250 78260 15260
rect 78540 15148 78596 24220
rect 78652 22148 78708 22158
rect 78652 17332 78708 22092
rect 78652 17266 78708 17276
rect 78316 15092 78596 15148
rect 77868 14420 77924 14430
rect 77868 14326 77924 14364
rect 78204 14418 78260 14430
rect 78204 14366 78206 14418
rect 78258 14366 78260 14418
rect 78204 14196 78260 14366
rect 78204 14130 78260 14140
rect 77868 13972 77924 13982
rect 77756 13970 77924 13972
rect 77756 13918 77870 13970
rect 77922 13918 77924 13970
rect 77756 13916 77924 13918
rect 77868 13906 77924 13916
rect 78092 13746 78148 13758
rect 78092 13694 78094 13746
rect 78146 13694 78148 13746
rect 77644 13636 77700 13646
rect 78092 13636 78148 13694
rect 77644 13634 78148 13636
rect 77644 13582 77646 13634
rect 77698 13582 78148 13634
rect 77644 13580 78148 13582
rect 77644 13570 77700 13580
rect 78092 13524 78148 13580
rect 78092 13458 78148 13468
rect 77532 13356 77924 13412
rect 77756 13188 77812 13198
rect 77756 12180 77812 13132
rect 77868 12402 77924 13356
rect 78316 13300 78372 15092
rect 77868 12350 77870 12402
rect 77922 12350 77924 12402
rect 77868 12338 77924 12350
rect 77980 13244 78372 13300
rect 77756 12124 77924 12180
rect 77644 12066 77700 12078
rect 77644 12014 77646 12066
rect 77698 12014 77700 12066
rect 77644 11956 77700 12014
rect 77644 11890 77700 11900
rect 77868 11282 77924 12124
rect 77868 11230 77870 11282
rect 77922 11230 77924 11282
rect 77868 11218 77924 11230
rect 77644 11170 77700 11182
rect 77644 11118 77646 11170
rect 77698 11118 77700 11170
rect 77644 10836 77700 11118
rect 77644 10770 77700 10780
rect 77420 10556 77924 10612
rect 77196 9772 77588 9828
rect 77196 9602 77252 9614
rect 77196 9550 77198 9602
rect 77250 9550 77252 9602
rect 77196 8372 77252 9550
rect 77196 8306 77252 8316
rect 77196 8148 77252 8158
rect 77084 8146 77252 8148
rect 77084 8094 77198 8146
rect 77250 8094 77252 8146
rect 77084 8092 77252 8094
rect 77196 8082 77252 8092
rect 77532 8146 77588 9772
rect 77644 9716 77700 9726
rect 77644 9622 77700 9660
rect 77868 9714 77924 10556
rect 77868 9662 77870 9714
rect 77922 9662 77924 9714
rect 77868 9650 77924 9662
rect 77868 8932 77924 8942
rect 77868 8838 77924 8876
rect 77532 8094 77534 8146
rect 77586 8094 77588 8146
rect 77532 7476 77588 8094
rect 77868 8260 77924 8270
rect 77868 8146 77924 8204
rect 77868 8094 77870 8146
rect 77922 8094 77924 8146
rect 77868 8082 77924 8094
rect 77532 7410 77588 7420
rect 77196 6916 77252 6926
rect 77084 6692 77140 6702
rect 76860 6514 76916 6524
rect 76972 6690 77140 6692
rect 76972 6638 77086 6690
rect 77138 6638 77140 6690
rect 76972 6636 77140 6638
rect 76748 6468 76804 6478
rect 76300 5170 76356 5180
rect 76524 6466 76804 6468
rect 76524 6414 76750 6466
rect 76802 6414 76804 6466
rect 76524 6412 76804 6414
rect 76524 5122 76580 6412
rect 76748 6402 76804 6412
rect 76860 6356 76916 6366
rect 76972 6356 77028 6636
rect 77084 6626 77140 6636
rect 76916 6300 77028 6356
rect 76860 6290 76916 6300
rect 76524 5070 76526 5122
rect 76578 5070 76580 5122
rect 76524 5058 76580 5070
rect 76972 5124 77028 6300
rect 76972 5058 77028 5068
rect 76188 4958 76190 5010
rect 76242 4958 76244 5010
rect 76188 4946 76244 4958
rect 77196 5010 77252 6860
rect 77532 6804 77588 6814
rect 77308 6692 77364 6702
rect 77532 6692 77588 6748
rect 77308 6690 77588 6692
rect 77308 6638 77310 6690
rect 77362 6638 77588 6690
rect 77308 6636 77588 6638
rect 77308 6626 77364 6636
rect 77420 6468 77476 6478
rect 77308 6132 77364 6142
rect 77308 5906 77364 6076
rect 77308 5854 77310 5906
rect 77362 5854 77364 5906
rect 77308 5842 77364 5854
rect 77420 5122 77476 6412
rect 77420 5070 77422 5122
rect 77474 5070 77476 5122
rect 77420 5058 77476 5070
rect 77196 4958 77198 5010
rect 77250 4958 77252 5010
rect 77196 4946 77252 4958
rect 77532 4788 77588 6636
rect 77644 6468 77700 6478
rect 77644 6466 77924 6468
rect 77644 6414 77646 6466
rect 77698 6414 77924 6466
rect 77644 6412 77924 6414
rect 77644 6402 77700 6412
rect 77868 5122 77924 6412
rect 77868 5070 77870 5122
rect 77922 5070 77924 5122
rect 77868 5058 77924 5070
rect 77196 4732 77588 4788
rect 76188 4116 76244 4126
rect 76188 4022 76244 4060
rect 77196 3666 77252 4732
rect 77196 3614 77198 3666
rect 77250 3614 77252 3666
rect 77196 3602 77252 3614
rect 77868 3444 77924 3454
rect 77980 3444 78036 13244
rect 78204 12178 78260 12190
rect 78204 12126 78206 12178
rect 78258 12126 78260 12178
rect 78204 11956 78260 12126
rect 78204 11890 78260 11900
rect 78204 11282 78260 11294
rect 78204 11230 78206 11282
rect 78258 11230 78260 11282
rect 78204 10836 78260 11230
rect 78204 10770 78260 10780
rect 78204 10612 78260 10622
rect 78204 10610 78372 10612
rect 78204 10558 78206 10610
rect 78258 10558 78372 10610
rect 78204 10556 78372 10558
rect 78204 10546 78260 10556
rect 78204 9716 78260 9726
rect 78204 9622 78260 9660
rect 78092 9604 78148 9614
rect 78092 8596 78148 9548
rect 78092 8428 78148 8540
rect 78092 8372 78260 8428
rect 78204 8258 78260 8372
rect 78204 8206 78206 8258
rect 78258 8206 78260 8258
rect 78204 8194 78260 8206
rect 78092 6804 78148 6814
rect 78092 6710 78148 6748
rect 78204 6132 78260 6142
rect 78204 6038 78260 6076
rect 78316 5572 78372 10556
rect 78204 5516 78372 5572
rect 78428 8932 78484 8942
rect 78092 5236 78148 5246
rect 78092 3554 78148 5180
rect 78204 5010 78260 5516
rect 78204 4958 78206 5010
rect 78258 4958 78260 5010
rect 78204 4946 78260 4958
rect 78316 5124 78372 5134
rect 78204 4564 78260 4574
rect 78316 4564 78372 5068
rect 78204 4562 78372 4564
rect 78204 4510 78206 4562
rect 78258 4510 78372 4562
rect 78204 4508 78372 4510
rect 78204 4498 78260 4508
rect 78428 4116 78484 8876
rect 78428 4050 78484 4060
rect 78092 3502 78094 3554
rect 78146 3502 78148 3554
rect 78092 3490 78148 3502
rect 77868 3442 78036 3444
rect 77868 3390 77870 3442
rect 77922 3390 78036 3442
rect 77868 3388 78036 3390
rect 77868 3378 77924 3388
rect 75516 1876 75572 1886
rect 75404 1820 75516 1876
rect 75516 1810 75572 1820
rect 4060 700 4676 756
rect 4928 0 5040 800
rect 5600 0 5712 800
rect 6272 0 6384 800
rect 6944 0 7056 800
rect 7616 0 7728 800
rect 8288 0 8400 800
rect 8960 0 9072 800
rect 9632 0 9744 800
rect 10304 0 10416 800
rect 10976 0 11088 800
rect 11648 0 11760 800
rect 12320 0 12432 800
rect 12992 0 13104 800
rect 13664 0 13776 800
rect 14336 0 14448 800
rect 15008 0 15120 800
rect 15680 0 15792 800
rect 16352 0 16464 800
rect 17024 0 17136 800
rect 17696 0 17808 800
rect 18368 0 18480 800
rect 19040 0 19152 800
rect 19712 0 19824 800
rect 20384 0 20496 800
rect 21056 0 21168 800
rect 21728 0 21840 800
rect 22400 0 22512 800
rect 23072 0 23184 800
rect 23744 0 23856 800
rect 24416 0 24528 800
rect 25088 0 25200 800
rect 25760 0 25872 800
rect 26432 0 26544 800
rect 27104 0 27216 800
rect 27776 0 27888 800
rect 28448 0 28560 800
rect 29120 0 29232 800
rect 29792 0 29904 800
rect 30464 0 30576 800
rect 31136 0 31248 800
rect 31808 0 31920 800
rect 32480 0 32592 800
rect 33152 0 33264 800
rect 33824 0 33936 800
rect 34496 0 34608 800
rect 35168 0 35280 800
rect 35840 0 35952 800
rect 36512 0 36624 800
rect 37184 0 37296 800
rect 37856 0 37968 800
rect 38528 0 38640 800
rect 39200 0 39312 800
rect 39872 0 39984 800
rect 40544 0 40656 800
rect 41216 0 41328 800
rect 41888 0 42000 800
rect 42560 0 42672 800
rect 43232 0 43344 800
rect 43904 0 44016 800
rect 44576 0 44688 800
rect 45248 0 45360 800
rect 45920 0 46032 800
rect 46592 0 46704 800
rect 47264 0 47376 800
rect 47936 0 48048 800
rect 48608 0 48720 800
rect 49280 0 49392 800
rect 49952 0 50064 800
rect 50624 0 50736 800
rect 51296 0 51408 800
rect 51968 0 52080 800
rect 52640 0 52752 800
rect 53312 0 53424 800
rect 53984 0 54096 800
rect 54656 0 54768 800
rect 55328 0 55440 800
rect 56000 0 56112 800
rect 56672 0 56784 800
rect 57344 0 57456 800
rect 58016 0 58128 800
rect 58688 0 58800 800
rect 59360 0 59472 800
rect 60032 0 60144 800
rect 60704 0 60816 800
rect 61376 0 61488 800
rect 62048 0 62160 800
rect 62720 0 62832 800
rect 63392 0 63504 800
rect 64064 0 64176 800
rect 64736 0 64848 800
rect 65408 0 65520 800
rect 66080 0 66192 800
rect 66752 0 66864 800
rect 67424 0 67536 800
rect 68096 0 68208 800
rect 68768 0 68880 800
rect 69440 0 69552 800
rect 70112 0 70224 800
rect 70784 0 70896 800
rect 71456 0 71568 800
rect 72128 0 72240 800
rect 72800 0 72912 800
rect 73472 0 73584 800
rect 74144 0 74256 800
rect 74816 0 74928 800
<< via2 >>
rect 2156 77308 2212 77364
rect 1932 76242 1988 76244
rect 1932 76190 1934 76242
rect 1934 76190 1986 76242
rect 1986 76190 1988 76242
rect 1932 76188 1988 76190
rect 1932 75292 1988 75348
rect 4476 76074 4532 76076
rect 4476 76022 4478 76074
rect 4478 76022 4530 76074
rect 4530 76022 4532 76074
rect 4476 76020 4532 76022
rect 4580 76074 4636 76076
rect 4580 76022 4582 76074
rect 4582 76022 4634 76074
rect 4634 76022 4636 76074
rect 4580 76020 4636 76022
rect 4684 76074 4740 76076
rect 4684 76022 4686 76074
rect 4686 76022 4738 76074
rect 4738 76022 4740 76074
rect 4684 76020 4740 76022
rect 4476 74506 4532 74508
rect 4476 74454 4478 74506
rect 4478 74454 4530 74506
rect 4530 74454 4532 74506
rect 4476 74452 4532 74454
rect 4580 74506 4636 74508
rect 4580 74454 4582 74506
rect 4582 74454 4634 74506
rect 4634 74454 4636 74506
rect 4580 74452 4636 74454
rect 4684 74506 4740 74508
rect 4684 74454 4686 74506
rect 4686 74454 4738 74506
rect 4738 74454 4740 74506
rect 4684 74452 4740 74454
rect 1932 74226 1988 74228
rect 1932 74174 1934 74226
rect 1934 74174 1986 74226
rect 1986 74174 1988 74226
rect 1932 74172 1988 74174
rect 1932 73106 1988 73108
rect 1932 73054 1934 73106
rect 1934 73054 1986 73106
rect 1986 73054 1988 73106
rect 1932 73052 1988 73054
rect 4476 72938 4532 72940
rect 4476 72886 4478 72938
rect 4478 72886 4530 72938
rect 4530 72886 4532 72938
rect 4476 72884 4532 72886
rect 4580 72938 4636 72940
rect 4580 72886 4582 72938
rect 4582 72886 4634 72938
rect 4634 72886 4636 72938
rect 4580 72884 4636 72886
rect 4684 72938 4740 72940
rect 4684 72886 4686 72938
rect 4686 72886 4738 72938
rect 4738 72886 4740 72938
rect 4684 72884 4740 72886
rect 2940 72492 2996 72548
rect 1932 71932 1988 71988
rect 3164 71986 3220 71988
rect 3164 71934 3166 71986
rect 3166 71934 3218 71986
rect 3218 71934 3220 71986
rect 3164 71932 3220 71934
rect 4956 72546 5012 72548
rect 4956 72494 4958 72546
rect 4958 72494 5010 72546
rect 5010 72494 5012 72546
rect 4956 72492 5012 72494
rect 5740 72492 5796 72548
rect 8316 76300 8372 76356
rect 3948 71932 4004 71988
rect 1932 70588 1988 70644
rect 2716 70140 2772 70196
rect 1932 69468 1988 69524
rect 1932 67228 1988 67284
rect 4476 71370 4532 71372
rect 4476 71318 4478 71370
rect 4478 71318 4530 71370
rect 4530 71318 4532 71370
rect 4476 71316 4532 71318
rect 4580 71370 4636 71372
rect 4580 71318 4582 71370
rect 4582 71318 4634 71370
rect 4634 71318 4636 71370
rect 4580 71316 4636 71318
rect 4684 71370 4740 71372
rect 4684 71318 4686 71370
rect 4686 71318 4738 71370
rect 4738 71318 4740 71370
rect 4684 71316 4740 71318
rect 3836 70194 3892 70196
rect 3836 70142 3838 70194
rect 3838 70142 3890 70194
rect 3890 70142 3892 70194
rect 3836 70140 3892 70142
rect 4476 69802 4532 69804
rect 4476 69750 4478 69802
rect 4478 69750 4530 69802
rect 4530 69750 4532 69802
rect 4476 69748 4532 69750
rect 4580 69802 4636 69804
rect 4580 69750 4582 69802
rect 4582 69750 4634 69802
rect 4634 69750 4636 69802
rect 4580 69748 4636 69750
rect 4684 69802 4740 69804
rect 4684 69750 4686 69802
rect 4686 69750 4738 69802
rect 4738 69750 4740 69802
rect 4684 69748 4740 69750
rect 2716 68402 2772 68404
rect 2716 68350 2718 68402
rect 2718 68350 2770 68402
rect 2770 68350 2772 68402
rect 2716 68348 2772 68350
rect 4476 68234 4532 68236
rect 4476 68182 4478 68234
rect 4478 68182 4530 68234
rect 4530 68182 4532 68234
rect 4476 68180 4532 68182
rect 4580 68234 4636 68236
rect 4580 68182 4582 68234
rect 4582 68182 4634 68234
rect 4634 68182 4636 68234
rect 4580 68180 4636 68182
rect 4684 68234 4740 68236
rect 4684 68182 4686 68234
rect 4686 68182 4738 68234
rect 4738 68182 4740 68234
rect 4684 68180 4740 68182
rect 1932 66386 1988 66388
rect 1932 66334 1934 66386
rect 1934 66334 1986 66386
rect 1986 66334 1988 66386
rect 1932 66332 1988 66334
rect 2716 67170 2772 67172
rect 2716 67118 2718 67170
rect 2718 67118 2770 67170
rect 2770 67118 2772 67170
rect 2716 67116 2772 67118
rect 2268 67004 2324 67060
rect 1932 63868 1988 63924
rect 3724 67170 3780 67172
rect 3724 67118 3726 67170
rect 3726 67118 3778 67170
rect 3778 67118 3780 67170
rect 3724 67116 3780 67118
rect 4284 67116 4340 67172
rect 3388 67058 3444 67060
rect 3388 67006 3390 67058
rect 3390 67006 3442 67058
rect 3442 67006 3444 67058
rect 3388 67004 3444 67006
rect 4476 66666 4532 66668
rect 4476 66614 4478 66666
rect 4478 66614 4530 66666
rect 4530 66614 4532 66666
rect 4476 66612 4532 66614
rect 4580 66666 4636 66668
rect 4580 66614 4582 66666
rect 4582 66614 4634 66666
rect 4634 66614 4636 66666
rect 4580 66612 4636 66614
rect 4684 66666 4740 66668
rect 4684 66614 4686 66666
rect 4686 66614 4738 66666
rect 4738 66614 4740 66666
rect 4684 66612 4740 66614
rect 3052 66220 3108 66276
rect 3836 66274 3892 66276
rect 3836 66222 3838 66274
rect 3838 66222 3890 66274
rect 3890 66222 3892 66274
rect 3836 66220 3892 66222
rect 2716 65266 2772 65268
rect 2716 65214 2718 65266
rect 2718 65214 2770 65266
rect 2770 65214 2772 65266
rect 2716 65212 2772 65214
rect 4476 65098 4532 65100
rect 4476 65046 4478 65098
rect 4478 65046 4530 65098
rect 4530 65046 4532 65098
rect 4476 65044 4532 65046
rect 4580 65098 4636 65100
rect 4580 65046 4582 65098
rect 4582 65046 4634 65098
rect 4634 65046 4636 65098
rect 4580 65044 4636 65046
rect 4684 65098 4740 65100
rect 4684 65046 4686 65098
rect 4686 65046 4738 65098
rect 4738 65046 4740 65098
rect 4684 65044 4740 65046
rect 1932 62748 1988 62804
rect 1932 61628 1988 61684
rect 2828 64034 2884 64036
rect 2828 63982 2830 64034
rect 2830 63982 2882 64034
rect 2882 63982 2884 64034
rect 2828 63980 2884 63982
rect 3724 63980 3780 64036
rect 4476 63530 4532 63532
rect 4476 63478 4478 63530
rect 4478 63478 4530 63530
rect 4530 63478 4532 63530
rect 4476 63476 4532 63478
rect 4580 63530 4636 63532
rect 4580 63478 4582 63530
rect 4582 63478 4634 63530
rect 4634 63478 4636 63530
rect 4580 63476 4636 63478
rect 4684 63530 4740 63532
rect 4684 63478 4686 63530
rect 4686 63478 4738 63530
rect 4738 63478 4740 63530
rect 4684 63476 4740 63478
rect 2828 62076 2884 62132
rect 3612 62076 3668 62132
rect 4476 61962 4532 61964
rect 4476 61910 4478 61962
rect 4478 61910 4530 61962
rect 4530 61910 4532 61962
rect 4476 61908 4532 61910
rect 4580 61962 4636 61964
rect 4580 61910 4582 61962
rect 4582 61910 4634 61962
rect 4634 61910 4636 61962
rect 4580 61908 4636 61910
rect 4684 61962 4740 61964
rect 4684 61910 4686 61962
rect 4686 61910 4738 61962
rect 4738 61910 4740 61962
rect 4684 61908 4740 61910
rect 2828 61292 2884 61348
rect 4172 61292 4228 61348
rect 2716 60562 2772 60564
rect 2716 60510 2718 60562
rect 2718 60510 2770 60562
rect 2770 60510 2772 60562
rect 2716 60508 2772 60510
rect 1932 59388 1988 59444
rect 2716 59948 2772 60004
rect 3836 60002 3892 60004
rect 3836 59950 3838 60002
rect 3838 59950 3890 60002
rect 3890 59950 3892 60002
rect 3836 59948 3892 59950
rect 2156 59164 2212 59220
rect 1932 57426 1988 57428
rect 1932 57374 1934 57426
rect 1934 57374 1986 57426
rect 1986 57374 1988 57426
rect 1932 57372 1988 57374
rect 1932 56028 1988 56084
rect 1932 53788 1988 53844
rect 2940 59218 2996 59220
rect 2940 59166 2942 59218
rect 2942 59166 2994 59218
rect 2994 59166 2996 59218
rect 2940 59164 2996 59166
rect 3500 59218 3556 59220
rect 3500 59166 3502 59218
rect 3502 59166 3554 59218
rect 3554 59166 3556 59218
rect 3500 59164 3556 59166
rect 2716 58210 2772 58212
rect 2716 58158 2718 58210
rect 2718 58158 2770 58210
rect 2770 58158 2772 58210
rect 2716 58156 2772 58158
rect 2716 56140 2772 56196
rect 3388 56194 3444 56196
rect 3388 56142 3390 56194
rect 3390 56142 3442 56194
rect 3442 56142 3444 56194
rect 3388 56140 3444 56142
rect 2716 55074 2772 55076
rect 2716 55022 2718 55074
rect 2718 55022 2770 55074
rect 2770 55022 2772 55074
rect 2716 55020 2772 55022
rect 1932 52722 1988 52724
rect 1932 52670 1934 52722
rect 1934 52670 1986 52722
rect 1986 52670 1988 52722
rect 1932 52668 1988 52670
rect 1932 51548 1988 51604
rect 1932 50706 1988 50708
rect 1932 50654 1934 50706
rect 1934 50654 1986 50706
rect 1986 50654 1988 50706
rect 1932 50652 1988 50654
rect 1932 49586 1988 49588
rect 1932 49534 1934 49586
rect 1934 49534 1986 49586
rect 1986 49534 1988 49586
rect 1932 49532 1988 49534
rect 1932 48188 1988 48244
rect 1932 45948 1988 46004
rect 2492 53506 2548 53508
rect 2492 53454 2494 53506
rect 2494 53454 2546 53506
rect 2546 53454 2548 53506
rect 2492 53452 2548 53454
rect 3164 53618 3220 53620
rect 3164 53566 3166 53618
rect 3166 53566 3218 53618
rect 3218 53566 3220 53618
rect 3164 53564 3220 53566
rect 2940 53452 2996 53508
rect 3836 53452 3892 53508
rect 3948 53564 4004 53620
rect 2380 48242 2436 48244
rect 2380 48190 2382 48242
rect 2382 48190 2434 48242
rect 2434 48190 2436 48242
rect 2380 48188 2436 48190
rect 2380 45724 2436 45780
rect 2828 50540 2884 50596
rect 3836 50594 3892 50596
rect 3836 50542 3838 50594
rect 3838 50542 3890 50594
rect 3890 50542 3892 50594
rect 3836 50540 3892 50542
rect 3164 49532 3220 49588
rect 2716 48972 2772 49028
rect 3612 49532 3668 49588
rect 2940 48242 2996 48244
rect 2940 48190 2942 48242
rect 2942 48190 2994 48242
rect 2994 48190 2996 48242
rect 2940 48188 2996 48190
rect 3836 49026 3892 49028
rect 3836 48974 3838 49026
rect 3838 48974 3890 49026
rect 3890 48974 3892 49026
rect 3836 48972 3892 48974
rect 2716 47234 2772 47236
rect 2716 47182 2718 47234
rect 2718 47182 2770 47234
rect 2770 47182 2772 47234
rect 2716 47180 2772 47182
rect 2716 45890 2772 45892
rect 2716 45838 2718 45890
rect 2718 45838 2770 45890
rect 2770 45838 2772 45890
rect 2716 45836 2772 45838
rect 3276 45836 3332 45892
rect 3052 45778 3108 45780
rect 3052 45726 3054 45778
rect 3054 45726 3106 45778
rect 3106 45726 3108 45778
rect 3052 45724 3108 45726
rect 2716 44882 2772 44884
rect 2716 44830 2718 44882
rect 2718 44830 2770 44882
rect 2770 44830 2772 44882
rect 2716 44828 2772 44830
rect 2716 44098 2772 44100
rect 2716 44046 2718 44098
rect 2718 44046 2770 44098
rect 2770 44046 2772 44098
rect 2716 44044 2772 44046
rect 1932 42866 1988 42868
rect 1932 42814 1934 42866
rect 1934 42814 1986 42866
rect 1986 42814 1988 42866
rect 1932 42812 1988 42814
rect 1708 41916 1764 41972
rect 1932 41746 1988 41748
rect 1932 41694 1934 41746
rect 1934 41694 1986 41746
rect 1986 41694 1988 41746
rect 1932 41692 1988 41694
rect 1932 40348 1988 40404
rect 1932 39228 1988 39284
rect 2268 43538 2324 43540
rect 2268 43486 2270 43538
rect 2270 43486 2322 43538
rect 2322 43486 2324 43538
rect 2268 43484 2324 43486
rect 2268 40626 2324 40628
rect 2268 40574 2270 40626
rect 2270 40574 2322 40626
rect 2322 40574 2324 40626
rect 2268 40572 2324 40574
rect 2828 43484 2884 43540
rect 2716 42700 2772 42756
rect 3164 40402 3220 40404
rect 3164 40350 3166 40402
rect 3166 40350 3218 40402
rect 3218 40350 3220 40402
rect 3164 40348 3220 40350
rect 2604 39564 2660 39620
rect 2940 39004 2996 39060
rect 3612 45724 3668 45780
rect 3836 42754 3892 42756
rect 3836 42702 3838 42754
rect 3838 42702 3890 42754
rect 3890 42702 3892 42754
rect 3836 42700 3892 42702
rect 3836 41970 3892 41972
rect 3836 41918 3838 41970
rect 3838 41918 3890 41970
rect 3890 41918 3892 41970
rect 3836 41916 3892 41918
rect 4476 60394 4532 60396
rect 4476 60342 4478 60394
rect 4478 60342 4530 60394
rect 4530 60342 4532 60394
rect 4476 60340 4532 60342
rect 4580 60394 4636 60396
rect 4580 60342 4582 60394
rect 4582 60342 4634 60394
rect 4634 60342 4636 60394
rect 4580 60340 4636 60342
rect 4684 60394 4740 60396
rect 4684 60342 4686 60394
rect 4686 60342 4738 60394
rect 4738 60342 4740 60394
rect 4684 60340 4740 60342
rect 4476 58826 4532 58828
rect 4476 58774 4478 58826
rect 4478 58774 4530 58826
rect 4530 58774 4532 58826
rect 4476 58772 4532 58774
rect 4580 58826 4636 58828
rect 4580 58774 4582 58826
rect 4582 58774 4634 58826
rect 4634 58774 4636 58826
rect 4580 58772 4636 58774
rect 4684 58826 4740 58828
rect 4684 58774 4686 58826
rect 4686 58774 4738 58826
rect 4738 58774 4740 58826
rect 4684 58772 4740 58774
rect 4476 57258 4532 57260
rect 4476 57206 4478 57258
rect 4478 57206 4530 57258
rect 4530 57206 4532 57258
rect 4476 57204 4532 57206
rect 4580 57258 4636 57260
rect 4580 57206 4582 57258
rect 4582 57206 4634 57258
rect 4634 57206 4636 57258
rect 4580 57204 4636 57206
rect 4684 57258 4740 57260
rect 4684 57206 4686 57258
rect 4686 57206 4738 57258
rect 4738 57206 4740 57258
rect 4684 57204 4740 57206
rect 4844 56140 4900 56196
rect 4476 55690 4532 55692
rect 4476 55638 4478 55690
rect 4478 55638 4530 55690
rect 4530 55638 4532 55690
rect 4476 55636 4532 55638
rect 4580 55690 4636 55692
rect 4580 55638 4582 55690
rect 4582 55638 4634 55690
rect 4634 55638 4636 55690
rect 4580 55636 4636 55638
rect 4684 55690 4740 55692
rect 4684 55638 4686 55690
rect 4686 55638 4738 55690
rect 4738 55638 4740 55690
rect 4684 55636 4740 55638
rect 4476 54122 4532 54124
rect 4476 54070 4478 54122
rect 4478 54070 4530 54122
rect 4530 54070 4532 54122
rect 4476 54068 4532 54070
rect 4580 54122 4636 54124
rect 4580 54070 4582 54122
rect 4582 54070 4634 54122
rect 4634 54070 4636 54122
rect 4580 54068 4636 54070
rect 4684 54122 4740 54124
rect 4684 54070 4686 54122
rect 4686 54070 4738 54122
rect 4738 54070 4740 54122
rect 4684 54068 4740 54070
rect 4476 52554 4532 52556
rect 4476 52502 4478 52554
rect 4478 52502 4530 52554
rect 4530 52502 4532 52554
rect 4476 52500 4532 52502
rect 4580 52554 4636 52556
rect 4580 52502 4582 52554
rect 4582 52502 4634 52554
rect 4634 52502 4636 52554
rect 4580 52500 4636 52502
rect 4684 52554 4740 52556
rect 4684 52502 4686 52554
rect 4686 52502 4738 52554
rect 4738 52502 4740 52554
rect 4684 52500 4740 52502
rect 4476 50986 4532 50988
rect 4476 50934 4478 50986
rect 4478 50934 4530 50986
rect 4530 50934 4532 50986
rect 4476 50932 4532 50934
rect 4580 50986 4636 50988
rect 4580 50934 4582 50986
rect 4582 50934 4634 50986
rect 4634 50934 4636 50986
rect 4580 50932 4636 50934
rect 4684 50986 4740 50988
rect 4684 50934 4686 50986
rect 4686 50934 4738 50986
rect 4738 50934 4740 50986
rect 4684 50932 4740 50934
rect 4476 49418 4532 49420
rect 4476 49366 4478 49418
rect 4478 49366 4530 49418
rect 4530 49366 4532 49418
rect 4476 49364 4532 49366
rect 4580 49418 4636 49420
rect 4580 49366 4582 49418
rect 4582 49366 4634 49418
rect 4634 49366 4636 49418
rect 4580 49364 4636 49366
rect 4684 49418 4740 49420
rect 4684 49366 4686 49418
rect 4686 49366 4738 49418
rect 4738 49366 4740 49418
rect 4684 49364 4740 49366
rect 4476 47850 4532 47852
rect 4476 47798 4478 47850
rect 4478 47798 4530 47850
rect 4530 47798 4532 47850
rect 4476 47796 4532 47798
rect 4580 47850 4636 47852
rect 4580 47798 4582 47850
rect 4582 47798 4634 47850
rect 4634 47798 4636 47850
rect 4580 47796 4636 47798
rect 4684 47850 4740 47852
rect 4684 47798 4686 47850
rect 4686 47798 4738 47850
rect 4738 47798 4740 47850
rect 4684 47796 4740 47798
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 4284 45890 4340 45892
rect 4284 45838 4286 45890
rect 4286 45838 4338 45890
rect 4338 45838 4340 45890
rect 4284 45836 4340 45838
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 4732 41970 4788 41972
rect 4732 41918 4734 41970
rect 4734 41918 4786 41970
rect 4786 41918 4788 41970
rect 4732 41916 4788 41918
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 5404 40626 5460 40628
rect 5404 40574 5406 40626
rect 5406 40574 5458 40626
rect 5458 40574 5460 40626
rect 5404 40572 5460 40574
rect 4060 40514 4116 40516
rect 4060 40462 4062 40514
rect 4062 40462 4114 40514
rect 4114 40462 4116 40514
rect 4060 40460 4116 40462
rect 4508 40514 4564 40516
rect 4508 40462 4510 40514
rect 4510 40462 4562 40514
rect 4562 40462 4564 40514
rect 4508 40460 4564 40462
rect 5180 40460 5236 40516
rect 4956 40402 5012 40404
rect 4956 40350 4958 40402
rect 4958 40350 5010 40402
rect 5010 40350 5012 40402
rect 4956 40348 5012 40350
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 3836 39618 3892 39620
rect 3836 39566 3838 39618
rect 3838 39566 3890 39618
rect 3890 39566 3892 39618
rect 3836 39564 3892 39566
rect 4732 39618 4788 39620
rect 4732 39566 4734 39618
rect 4734 39566 4786 39618
rect 4786 39566 4788 39618
rect 4732 39564 4788 39566
rect 5180 39340 5236 39396
rect 3276 39004 3332 39060
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 3388 38108 3444 38164
rect 2044 37378 2100 37380
rect 2044 37326 2046 37378
rect 2046 37326 2098 37378
rect 2098 37326 2100 37378
rect 2044 37324 2100 37326
rect 1708 36988 1764 37044
rect 2492 36988 2548 37044
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 2044 36258 2100 36260
rect 2044 36206 2046 36258
rect 2046 36206 2098 36258
rect 2098 36206 2100 36258
rect 2044 36204 2100 36206
rect 1708 35868 1764 35924
rect 2492 35868 2548 35924
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 1708 34802 1764 34804
rect 1708 34750 1710 34802
rect 1710 34750 1762 34802
rect 1762 34750 1764 34802
rect 1708 34748 1764 34750
rect 2492 34802 2548 34804
rect 2492 34750 2494 34802
rect 2494 34750 2546 34802
rect 2546 34750 2548 34802
rect 2492 34748 2548 34750
rect 2044 34690 2100 34692
rect 2044 34638 2046 34690
rect 2046 34638 2098 34690
rect 2098 34638 2100 34690
rect 2044 34636 2100 34638
rect 2044 34242 2100 34244
rect 2044 34190 2046 34242
rect 2046 34190 2098 34242
rect 2098 34190 2100 34242
rect 2044 34188 2100 34190
rect 1708 33628 1764 33684
rect 2492 33628 2548 33684
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 2044 33122 2100 33124
rect 2044 33070 2046 33122
rect 2046 33070 2098 33122
rect 2098 33070 2100 33122
rect 2044 33068 2100 33070
rect 1708 32508 1764 32564
rect 2492 32508 2548 32564
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 2044 31724 2100 31780
rect 1708 31388 1764 31444
rect 2492 31388 2548 31444
rect 2044 31106 2100 31108
rect 2044 31054 2046 31106
rect 2046 31054 2098 31106
rect 2098 31054 2100 31106
rect 2044 31052 2100 31054
rect 1708 30828 1764 30884
rect 2492 30882 2548 30884
rect 2492 30830 2494 30882
rect 2494 30830 2546 30882
rect 2546 30830 2548 30882
rect 2492 30828 2548 30830
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 1708 30268 1764 30324
rect 2044 29538 2100 29540
rect 2044 29486 2046 29538
rect 2046 29486 2098 29538
rect 2098 29486 2100 29538
rect 2044 29484 2100 29486
rect 1708 29148 1764 29204
rect 2492 29148 2548 29204
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 2044 28700 2100 28756
rect 1708 28028 1764 28084
rect 2492 28028 2548 28084
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 2044 27244 2100 27300
rect 1708 26962 1764 26964
rect 1708 26910 1710 26962
rect 1710 26910 1762 26962
rect 1762 26910 1764 26962
rect 1708 26908 1764 26910
rect 2492 26962 2548 26964
rect 2492 26910 2494 26962
rect 2494 26910 2546 26962
rect 2546 26910 2548 26962
rect 2492 26908 2548 26910
rect 2044 26012 2100 26068
rect 1708 25788 1764 25844
rect 2492 25788 2548 25844
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 2044 25564 2100 25620
rect 1708 24668 1764 24724
rect 2492 24668 2548 24724
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 8316 24332 8372 24388
rect 9996 74844 10052 74900
rect 4684 24276 4740 24278
rect 2044 23884 2100 23940
rect 1708 23548 1764 23604
rect 2492 23548 2548 23604
rect 1708 22988 1764 23044
rect 2492 23042 2548 23044
rect 2492 22990 2494 23042
rect 2494 22990 2546 23042
rect 2546 22990 2548 23042
rect 2492 22988 2548 22990
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 2044 22540 2100 22596
rect 1708 22428 1764 22484
rect 11900 75906 11956 75908
rect 11900 75854 11902 75906
rect 11902 75854 11954 75906
rect 11954 75854 11956 75906
rect 11900 75852 11956 75854
rect 11564 75516 11620 75572
rect 11676 74732 11732 74788
rect 9996 21756 10052 21812
rect 11452 22876 11508 22932
rect 2044 21698 2100 21700
rect 2044 21646 2046 21698
rect 2046 21646 2098 21698
rect 2098 21646 2100 21698
rect 2044 21644 2100 21646
rect 1708 21308 1764 21364
rect 2492 21308 2548 21364
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 2044 20860 2100 20916
rect 1708 20188 1764 20244
rect 2044 20300 2100 20356
rect 1708 19122 1764 19124
rect 1708 19070 1710 19122
rect 1710 19070 1762 19122
rect 1762 19070 1764 19122
rect 1708 19068 1764 19070
rect 2492 20188 2548 20244
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 7532 19292 7588 19348
rect 2492 19122 2548 19124
rect 2492 19070 2494 19122
rect 2494 19070 2546 19122
rect 2546 19070 2548 19122
rect 2492 19068 2548 19070
rect 6300 18620 6356 18676
rect 2044 18284 2100 18340
rect 1708 17948 1764 18004
rect 2492 17948 2548 18004
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 2044 17836 2100 17892
rect 1708 17388 1764 17444
rect 2492 17442 2548 17444
rect 2492 17390 2494 17442
rect 2494 17390 2546 17442
rect 2546 17390 2548 17442
rect 2492 17388 2548 17390
rect 1708 16828 1764 16884
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 2044 16268 2100 16324
rect 2156 16044 2212 16100
rect 1708 15708 1764 15764
rect 2044 15426 2100 15428
rect 2044 15374 2046 15426
rect 2046 15374 2098 15426
rect 2098 15374 2100 15426
rect 2044 15372 2100 15374
rect 1708 14588 1764 14644
rect 1596 14364 1652 14420
rect 2044 13970 2100 13972
rect 2044 13918 2046 13970
rect 2046 13918 2098 13970
rect 2098 13918 2100 13970
rect 2044 13916 2100 13918
rect 1708 13468 1764 13524
rect 1932 13020 1988 13076
rect 1708 12348 1764 12404
rect 1708 11282 1764 11284
rect 1708 11230 1710 11282
rect 1710 11230 1762 11282
rect 1762 11230 1764 11282
rect 1708 11228 1764 11230
rect 1708 10108 1764 10164
rect 1708 9548 1764 9604
rect 1708 8988 1764 9044
rect 1708 7868 1764 7924
rect 1708 7308 1764 7364
rect 1708 6748 1764 6804
rect 2044 12850 2100 12852
rect 2044 12798 2046 12850
rect 2046 12798 2098 12850
rect 2098 12798 2100 12850
rect 2044 12796 2100 12798
rect 2044 11282 2100 11284
rect 2044 11230 2046 11282
rect 2046 11230 2098 11282
rect 2098 11230 2100 11282
rect 2044 11228 2100 11230
rect 2044 10722 2100 10724
rect 2044 10670 2046 10722
rect 2046 10670 2098 10722
rect 2098 10670 2100 10722
rect 2044 10668 2100 10670
rect 2492 15708 2548 15764
rect 5852 15148 5908 15204
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 2492 14588 2548 14644
rect 2492 13468 2548 13524
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 2492 12348 2548 12404
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 2492 11170 2548 11172
rect 2492 11118 2494 11170
rect 2494 11118 2546 11170
rect 2546 11118 2548 11170
rect 2492 11116 2548 11118
rect 2380 10332 2436 10388
rect 2492 10108 2548 10164
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 2492 9602 2548 9604
rect 2492 9550 2494 9602
rect 2494 9550 2546 9602
rect 2546 9550 2548 9602
rect 2492 9548 2548 9550
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 2492 7868 2548 7924
rect 2044 7698 2100 7700
rect 2044 7646 2046 7698
rect 2046 7646 2098 7698
rect 2098 7646 2100 7698
rect 2044 7644 2100 7646
rect 5852 7644 5908 7700
rect 2492 7362 2548 7364
rect 2492 7310 2494 7362
rect 2494 7310 2546 7362
rect 2546 7310 2548 7362
rect 2492 7308 2548 7310
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 6076 6972 6132 7028
rect 2156 6748 2212 6804
rect 4284 6524 4340 6580
rect 3612 6076 3668 6132
rect 1708 5628 1764 5684
rect 2380 5964 2436 6020
rect 1596 4956 1652 5012
rect 2492 5628 2548 5684
rect 1708 4508 1764 4564
rect 1820 4172 1876 4228
rect 1820 3554 1876 3556
rect 1820 3502 1822 3554
rect 1822 3502 1874 3554
rect 1874 3502 1876 3554
rect 1820 3500 1876 3502
rect 2492 4508 2548 4564
rect 2716 4956 2772 5012
rect 2492 4226 2548 4228
rect 2492 4174 2494 4226
rect 2494 4174 2546 4226
rect 2546 4174 2548 4226
rect 2492 4172 2548 4174
rect 3388 3554 3444 3556
rect 3388 3502 3390 3554
rect 3390 3502 3442 3554
rect 3442 3502 3444 3554
rect 3388 3500 3444 3502
rect 4956 6412 5012 6468
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 4844 5516 4900 5572
rect 3948 3442 4004 3444
rect 3948 3390 3950 3442
rect 3950 3390 4002 3442
rect 4002 3390 4004 3442
rect 3948 3388 4004 3390
rect 2380 2268 2436 2324
rect 4508 4284 4564 4340
rect 4620 4172 4676 4228
rect 4172 3388 4228 3444
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 4732 3724 4788 3780
rect 5628 5852 5684 5908
rect 5404 3836 5460 3892
rect 5068 3724 5124 3780
rect 5852 3612 5908 3668
rect 5628 3500 5684 3556
rect 9996 15260 10052 15316
rect 8316 14588 8372 14644
rect 8316 12796 8372 12852
rect 8316 12348 8372 12404
rect 9436 12012 9492 12068
rect 8316 11228 8372 11284
rect 8204 10444 8260 10500
rect 8428 9884 8484 9940
rect 8092 9714 8148 9716
rect 8092 9662 8094 9714
rect 8094 9662 8146 9714
rect 8146 9662 8148 9714
rect 8092 9660 8148 9662
rect 7532 6748 7588 6804
rect 9548 11282 9604 11284
rect 9548 11230 9550 11282
rect 9550 11230 9602 11282
rect 9602 11230 9604 11282
rect 9548 11228 9604 11230
rect 10332 12066 10388 12068
rect 10332 12014 10334 12066
rect 10334 12014 10386 12066
rect 10386 12014 10388 12066
rect 10332 12012 10388 12014
rect 11116 10834 11172 10836
rect 11116 10782 11118 10834
rect 11118 10782 11170 10834
rect 11170 10782 11172 10834
rect 11116 10780 11172 10782
rect 9996 10332 10052 10388
rect 12124 76300 12180 76356
rect 13356 76354 13412 76356
rect 13356 76302 13358 76354
rect 13358 76302 13410 76354
rect 13410 76302 13412 76354
rect 13356 76300 13412 76302
rect 12572 75852 12628 75908
rect 12684 75682 12740 75684
rect 12684 75630 12686 75682
rect 12686 75630 12738 75682
rect 12738 75630 12740 75682
rect 12684 75628 12740 75630
rect 13580 75682 13636 75684
rect 13580 75630 13582 75682
rect 13582 75630 13634 75682
rect 13634 75630 13636 75682
rect 13580 75628 13636 75630
rect 13916 75516 13972 75572
rect 13468 74898 13524 74900
rect 13468 74846 13470 74898
rect 13470 74846 13522 74898
rect 13522 74846 13524 74898
rect 13468 74844 13524 74846
rect 14252 74844 14308 74900
rect 14028 74114 14084 74116
rect 14028 74062 14030 74114
rect 14030 74062 14082 74114
rect 14082 74062 14084 74114
rect 14028 74060 14084 74062
rect 12908 73948 12964 74004
rect 14364 74002 14420 74004
rect 14364 73950 14366 74002
rect 14366 73950 14418 74002
rect 14418 73950 14420 74002
rect 14364 73948 14420 73950
rect 12684 23996 12740 24052
rect 13468 23436 13524 23492
rect 14252 24332 14308 24388
rect 11676 13020 11732 13076
rect 12908 22428 12964 22484
rect 11676 11452 11732 11508
rect 12460 11506 12516 11508
rect 12460 11454 12462 11506
rect 12462 11454 12514 11506
rect 12514 11454 12516 11506
rect 12460 11452 12516 11454
rect 15372 76690 15428 76692
rect 15372 76638 15374 76690
rect 15374 76638 15426 76690
rect 15426 76638 15428 76690
rect 15372 76636 15428 76638
rect 14364 22876 14420 22932
rect 16604 76636 16660 76692
rect 16380 76300 16436 76356
rect 17164 76354 17220 76356
rect 17164 76302 17166 76354
rect 17166 76302 17218 76354
rect 17218 76302 17220 76354
rect 17164 76300 17220 76302
rect 16380 74060 16436 74116
rect 19836 76858 19892 76860
rect 19836 76806 19838 76858
rect 19838 76806 19890 76858
rect 19890 76806 19892 76858
rect 19836 76804 19892 76806
rect 19940 76858 19996 76860
rect 19940 76806 19942 76858
rect 19942 76806 19994 76858
rect 19994 76806 19996 76858
rect 19940 76804 19996 76806
rect 20044 76858 20100 76860
rect 20044 76806 20046 76858
rect 20046 76806 20098 76858
rect 20098 76806 20100 76858
rect 20044 76804 20100 76806
rect 17948 75516 18004 75572
rect 19180 75516 19236 75572
rect 16380 24556 16436 24612
rect 14700 22428 14756 22484
rect 14924 23436 14980 23492
rect 14924 23100 14980 23156
rect 11564 11282 11620 11284
rect 11564 11230 11566 11282
rect 11566 11230 11618 11282
rect 11618 11230 11620 11282
rect 11564 11228 11620 11230
rect 11228 9996 11284 10052
rect 9324 9714 9380 9716
rect 9324 9662 9326 9714
rect 9326 9662 9378 9714
rect 9378 9662 9380 9714
rect 9324 9660 9380 9662
rect 8876 8930 8932 8932
rect 8876 8878 8878 8930
rect 8878 8878 8930 8930
rect 8930 8878 8932 8930
rect 8876 8876 8932 8878
rect 6300 5964 6356 6020
rect 6636 6018 6692 6020
rect 6636 5966 6638 6018
rect 6638 5966 6690 6018
rect 6690 5966 6692 6018
rect 6636 5964 6692 5966
rect 6860 5740 6916 5796
rect 6300 5404 6356 5460
rect 6076 5068 6132 5124
rect 6188 4844 6244 4900
rect 6188 4172 6244 4228
rect 6412 4172 6468 4228
rect 6524 4844 6580 4900
rect 6300 4114 6356 4116
rect 6300 4062 6302 4114
rect 6302 4062 6354 4114
rect 6354 4062 6356 4114
rect 6300 4060 6356 4062
rect 6748 5010 6804 5012
rect 6748 4958 6750 5010
rect 6750 4958 6802 5010
rect 6802 4958 6804 5010
rect 6748 4956 6804 4958
rect 6860 4844 6916 4900
rect 6636 4338 6692 4340
rect 6636 4286 6638 4338
rect 6638 4286 6690 4338
rect 6690 4286 6692 4338
rect 6636 4284 6692 4286
rect 7084 4620 7140 4676
rect 6972 4114 7028 4116
rect 6972 4062 6974 4114
rect 6974 4062 7026 4114
rect 7026 4062 7028 4114
rect 6972 4060 7028 4062
rect 6524 3948 6580 4004
rect 6972 3836 7028 3892
rect 6524 3554 6580 3556
rect 6524 3502 6526 3554
rect 6526 3502 6578 3554
rect 6578 3502 6580 3554
rect 6524 3500 6580 3502
rect 6748 3330 6804 3332
rect 6748 3278 6750 3330
rect 6750 3278 6802 3330
rect 6802 3278 6804 3330
rect 6748 3276 6804 3278
rect 7308 4956 7364 5012
rect 7868 6188 7924 6244
rect 7980 6076 8036 6132
rect 8204 6914 8260 6916
rect 8204 6862 8206 6914
rect 8206 6862 8258 6914
rect 8258 6862 8260 6914
rect 8204 6860 8260 6862
rect 8652 6860 8708 6916
rect 8988 8818 9044 8820
rect 8988 8766 8990 8818
rect 8990 8766 9042 8818
rect 9042 8766 9044 8818
rect 8988 8764 9044 8766
rect 8876 6914 8932 6916
rect 8876 6862 8878 6914
rect 8878 6862 8930 6914
rect 8930 6862 8932 6914
rect 8876 6860 8932 6862
rect 8652 6466 8708 6468
rect 8652 6414 8654 6466
rect 8654 6414 8706 6466
rect 8706 6414 8708 6466
rect 8652 6412 8708 6414
rect 9996 9660 10052 9716
rect 9548 7084 9604 7140
rect 9436 6578 9492 6580
rect 9436 6526 9438 6578
rect 9438 6526 9490 6578
rect 9490 6526 9492 6578
rect 9436 6524 9492 6526
rect 8988 6412 9044 6468
rect 8316 6130 8372 6132
rect 8316 6078 8318 6130
rect 8318 6078 8370 6130
rect 8370 6078 8372 6130
rect 8316 6076 8372 6078
rect 8988 6076 9044 6132
rect 8092 5852 8148 5908
rect 8428 5964 8484 6020
rect 7644 5292 7700 5348
rect 7980 5068 8036 5124
rect 7644 4844 7700 4900
rect 7644 4450 7700 4452
rect 7644 4398 7646 4450
rect 7646 4398 7698 4450
rect 7698 4398 7700 4450
rect 7644 4396 7700 4398
rect 7308 4060 7364 4116
rect 7196 3500 7252 3556
rect 7420 3836 7476 3892
rect 8316 5180 8372 5236
rect 8652 5516 8708 5572
rect 8988 5346 9044 5348
rect 8988 5294 8990 5346
rect 8990 5294 9042 5346
rect 9042 5294 9044 5346
rect 8988 5292 9044 5294
rect 8876 5122 8932 5124
rect 8876 5070 8878 5122
rect 8878 5070 8930 5122
rect 8930 5070 8932 5122
rect 8876 5068 8932 5070
rect 9660 6412 9716 6468
rect 11564 10834 11620 10836
rect 11564 10782 11566 10834
rect 11566 10782 11618 10834
rect 11618 10782 11620 10834
rect 11564 10780 11620 10782
rect 11452 10498 11508 10500
rect 11452 10446 11454 10498
rect 11454 10446 11506 10498
rect 11506 10446 11508 10498
rect 11452 10444 11508 10446
rect 12684 10610 12740 10612
rect 12684 10558 12686 10610
rect 12686 10558 12738 10610
rect 12738 10558 12740 10610
rect 12684 10556 12740 10558
rect 11900 9772 11956 9828
rect 12236 9996 12292 10052
rect 11340 9548 11396 9604
rect 12012 9602 12068 9604
rect 12012 9550 12014 9602
rect 12014 9550 12066 9602
rect 12066 9550 12068 9602
rect 12012 9548 12068 9550
rect 10332 8930 10388 8932
rect 10332 8878 10334 8930
rect 10334 8878 10386 8930
rect 10386 8878 10388 8930
rect 10332 8876 10388 8878
rect 12572 9826 12628 9828
rect 12572 9774 12574 9826
rect 12574 9774 12626 9826
rect 12626 9774 12628 9826
rect 12572 9772 12628 9774
rect 12460 8930 12516 8932
rect 12460 8878 12462 8930
rect 12462 8878 12514 8930
rect 12514 8878 12516 8930
rect 12460 8876 12516 8878
rect 12124 8764 12180 8820
rect 13468 9884 13524 9940
rect 13916 9884 13972 9940
rect 13244 9772 13300 9828
rect 14028 9826 14084 9828
rect 14028 9774 14030 9826
rect 14030 9774 14082 9826
rect 14082 9774 14084 9826
rect 14028 9772 14084 9774
rect 13468 9602 13524 9604
rect 13468 9550 13470 9602
rect 13470 9550 13522 9602
rect 13522 9550 13524 9602
rect 13468 9548 13524 9550
rect 14140 9548 14196 9604
rect 13804 9266 13860 9268
rect 13804 9214 13806 9266
rect 13806 9214 13858 9266
rect 13858 9214 13860 9266
rect 13804 9212 13860 9214
rect 14252 9212 14308 9268
rect 13244 8930 13300 8932
rect 13244 8878 13246 8930
rect 13246 8878 13298 8930
rect 13298 8878 13300 8930
rect 13244 8876 13300 8878
rect 9996 6412 10052 6468
rect 10780 6748 10836 6804
rect 10220 5852 10276 5908
rect 8540 4620 8596 4676
rect 8204 4226 8260 4228
rect 8204 4174 8206 4226
rect 8206 4174 8258 4226
rect 8258 4174 8260 4226
rect 8204 4172 8260 4174
rect 7532 3388 7588 3444
rect 7084 2604 7140 2660
rect 7756 2492 7812 2548
rect 8092 2268 8148 2324
rect 8764 4508 8820 4564
rect 9660 4060 9716 4116
rect 8988 3948 9044 4004
rect 8764 3164 8820 3220
rect 9548 3724 9604 3780
rect 9660 3554 9716 3556
rect 9660 3502 9662 3554
rect 9662 3502 9714 3554
rect 9714 3502 9716 3554
rect 9660 3500 9716 3502
rect 10220 4338 10276 4340
rect 10220 4286 10222 4338
rect 10222 4286 10274 4338
rect 10274 4286 10276 4338
rect 10220 4284 10276 4286
rect 10220 4060 10276 4116
rect 10332 3836 10388 3892
rect 10332 3612 10388 3668
rect 9996 3276 10052 3332
rect 9884 2828 9940 2884
rect 10556 5404 10612 5460
rect 11004 5740 11060 5796
rect 11116 7420 11172 7476
rect 10780 3836 10836 3892
rect 10892 4396 10948 4452
rect 10444 3500 10500 3556
rect 11004 4226 11060 4228
rect 11004 4174 11006 4226
rect 11006 4174 11058 4226
rect 11058 4174 11060 4226
rect 11004 4172 11060 4174
rect 11228 7362 11284 7364
rect 11228 7310 11230 7362
rect 11230 7310 11282 7362
rect 11282 7310 11284 7362
rect 11228 7308 11284 7310
rect 12124 6690 12180 6692
rect 12124 6638 12126 6690
rect 12126 6638 12178 6690
rect 12178 6638 12180 6690
rect 12124 6636 12180 6638
rect 11228 5628 11284 5684
rect 11452 5292 11508 5348
rect 11452 3948 11508 4004
rect 11004 3388 11060 3444
rect 10444 3052 10500 3108
rect 10556 2380 10612 2436
rect 12012 5740 12068 5796
rect 11676 5122 11732 5124
rect 11676 5070 11678 5122
rect 11678 5070 11730 5122
rect 11730 5070 11732 5122
rect 11676 5068 11732 5070
rect 11900 4172 11956 4228
rect 12348 6860 12404 6916
rect 13132 7698 13188 7700
rect 13132 7646 13134 7698
rect 13134 7646 13186 7698
rect 13186 7646 13188 7698
rect 13132 7644 13188 7646
rect 13580 7698 13636 7700
rect 13580 7646 13582 7698
rect 13582 7646 13634 7698
rect 13634 7646 13636 7698
rect 13580 7644 13636 7646
rect 13804 7532 13860 7588
rect 12796 6636 12852 6692
rect 12684 6188 12740 6244
rect 12572 5852 12628 5908
rect 12460 5234 12516 5236
rect 12460 5182 12462 5234
rect 12462 5182 12514 5234
rect 12514 5182 12516 5234
rect 12460 5180 12516 5182
rect 12236 4396 12292 4452
rect 11676 3554 11732 3556
rect 11676 3502 11678 3554
rect 11678 3502 11730 3554
rect 11730 3502 11732 3554
rect 11676 3500 11732 3502
rect 12908 6412 12964 6468
rect 13468 7362 13524 7364
rect 13468 7310 13470 7362
rect 13470 7310 13522 7362
rect 13522 7310 13524 7362
rect 13468 7308 13524 7310
rect 13468 6860 13524 6916
rect 13580 6802 13636 6804
rect 13580 6750 13582 6802
rect 13582 6750 13634 6802
rect 13634 6750 13636 6802
rect 13580 6748 13636 6750
rect 13804 6748 13860 6804
rect 14588 11676 14644 11732
rect 14476 9938 14532 9940
rect 14476 9886 14478 9938
rect 14478 9886 14530 9938
rect 14530 9886 14532 9938
rect 14476 9884 14532 9886
rect 14364 7644 14420 7700
rect 14476 9660 14532 9716
rect 16156 23436 16212 23492
rect 15596 22482 15652 22484
rect 15596 22430 15598 22482
rect 15598 22430 15650 22482
rect 15650 22430 15652 22482
rect 15596 22428 15652 22430
rect 15484 21756 15540 21812
rect 15820 21756 15876 21812
rect 15484 21420 15540 21476
rect 14924 10780 14980 10836
rect 15372 10556 15428 10612
rect 14924 9996 14980 10052
rect 14924 9266 14980 9268
rect 14924 9214 14926 9266
rect 14926 9214 14978 9266
rect 14978 9214 14980 9266
rect 14924 9212 14980 9214
rect 15484 9884 15540 9940
rect 16044 11788 16100 11844
rect 14588 7532 14644 7588
rect 14252 6860 14308 6916
rect 14028 6524 14084 6580
rect 14252 6636 14308 6692
rect 13916 6466 13972 6468
rect 13916 6414 13918 6466
rect 13918 6414 13970 6466
rect 13970 6414 13972 6466
rect 13916 6412 13972 6414
rect 13468 6076 13524 6132
rect 13468 5516 13524 5572
rect 14140 6188 14196 6244
rect 13692 6018 13748 6020
rect 13692 5966 13694 6018
rect 13694 5966 13746 6018
rect 13746 5966 13748 6018
rect 13692 5964 13748 5966
rect 14028 5906 14084 5908
rect 14028 5854 14030 5906
rect 14030 5854 14082 5906
rect 14082 5854 14084 5906
rect 14028 5852 14084 5854
rect 13804 5628 13860 5684
rect 13020 5068 13076 5124
rect 13468 5180 13524 5236
rect 14028 5516 14084 5572
rect 13804 4844 13860 4900
rect 13916 5404 13972 5460
rect 13692 4338 13748 4340
rect 13692 4286 13694 4338
rect 13694 4286 13746 4338
rect 13746 4286 13748 4338
rect 13692 4284 13748 4286
rect 13468 3724 13524 3780
rect 13580 4060 13636 4116
rect 12572 3442 12628 3444
rect 12572 3390 12574 3442
rect 12574 3390 12626 3442
rect 12626 3390 12628 3442
rect 12572 3388 12628 3390
rect 14364 6412 14420 6468
rect 14700 6466 14756 6468
rect 14700 6414 14702 6466
rect 14702 6414 14754 6466
rect 14754 6414 14756 6466
rect 14700 6412 14756 6414
rect 14812 6300 14868 6356
rect 15148 6130 15204 6132
rect 15148 6078 15150 6130
rect 15150 6078 15202 6130
rect 15202 6078 15204 6130
rect 15148 6076 15204 6078
rect 14700 5852 14756 5908
rect 15596 8316 15652 8372
rect 15596 7586 15652 7588
rect 15596 7534 15598 7586
rect 15598 7534 15650 7586
rect 15650 7534 15652 7586
rect 15596 7532 15652 7534
rect 15820 7362 15876 7364
rect 15820 7310 15822 7362
rect 15822 7310 15874 7362
rect 15874 7310 15876 7362
rect 15820 7308 15876 7310
rect 15932 6636 15988 6692
rect 15596 5740 15652 5796
rect 14812 5292 14868 5348
rect 14588 5068 14644 5124
rect 14140 4956 14196 5012
rect 14252 4844 14308 4900
rect 14364 4732 14420 4788
rect 14140 3836 14196 3892
rect 14252 4508 14308 4564
rect 11900 2940 11956 2996
rect 12348 2604 12404 2660
rect 13020 2492 13076 2548
rect 14700 5010 14756 5012
rect 14700 4958 14702 5010
rect 14702 4958 14754 5010
rect 14754 4958 14756 5010
rect 14700 4956 14756 4958
rect 14588 4284 14644 4340
rect 14476 4226 14532 4228
rect 14476 4174 14478 4226
rect 14478 4174 14530 4226
rect 14530 4174 14532 4226
rect 14476 4172 14532 4174
rect 14924 4844 14980 4900
rect 14812 3612 14868 3668
rect 14924 4620 14980 4676
rect 15260 4898 15316 4900
rect 15260 4846 15262 4898
rect 15262 4846 15314 4898
rect 15314 4846 15316 4898
rect 15260 4844 15316 4846
rect 16828 22316 16884 22372
rect 16716 22092 16772 22148
rect 16604 13580 16660 13636
rect 16380 11676 16436 11732
rect 16268 8930 16324 8932
rect 16268 8878 16270 8930
rect 16270 8878 16322 8930
rect 16322 8878 16324 8930
rect 16268 8876 16324 8878
rect 15148 4620 15204 4676
rect 15036 4284 15092 4340
rect 15932 5122 15988 5124
rect 15932 5070 15934 5122
rect 15934 5070 15986 5122
rect 15986 5070 15988 5122
rect 15932 5068 15988 5070
rect 17052 20076 17108 20132
rect 17500 24332 17556 24388
rect 17388 23548 17444 23604
rect 17612 23378 17668 23380
rect 17612 23326 17614 23378
rect 17614 23326 17666 23378
rect 17666 23326 17668 23378
rect 17612 23324 17668 23326
rect 18060 24332 18116 24388
rect 17500 21810 17556 21812
rect 17500 21758 17502 21810
rect 17502 21758 17554 21810
rect 17554 21758 17556 21810
rect 17500 21756 17556 21758
rect 17724 21810 17780 21812
rect 17724 21758 17726 21810
rect 17726 21758 17778 21810
rect 17778 21758 17780 21810
rect 17724 21756 17780 21758
rect 17948 22204 18004 22260
rect 18172 22092 18228 22148
rect 19404 74786 19460 74788
rect 19404 74734 19406 74786
rect 19406 74734 19458 74786
rect 19458 74734 19460 74786
rect 19404 74732 19460 74734
rect 19628 75628 19684 75684
rect 21084 76690 21140 76692
rect 21084 76638 21086 76690
rect 21086 76638 21138 76690
rect 21138 76638 21140 76690
rect 21084 76636 21140 76638
rect 21980 76636 22036 76692
rect 20636 75852 20692 75908
rect 21532 75906 21588 75908
rect 21532 75854 21534 75906
rect 21534 75854 21586 75906
rect 21586 75854 21588 75906
rect 21532 75852 21588 75854
rect 20300 75682 20356 75684
rect 20300 75630 20302 75682
rect 20302 75630 20354 75682
rect 20354 75630 20356 75682
rect 20300 75628 20356 75630
rect 19836 75290 19892 75292
rect 19836 75238 19838 75290
rect 19838 75238 19890 75290
rect 19890 75238 19892 75290
rect 19836 75236 19892 75238
rect 19940 75290 19996 75292
rect 19940 75238 19942 75290
rect 19942 75238 19994 75290
rect 19994 75238 19996 75290
rect 19940 75236 19996 75238
rect 20044 75290 20100 75292
rect 20044 75238 20046 75290
rect 20046 75238 20098 75290
rect 20098 75238 20100 75290
rect 20044 75236 20100 75238
rect 23660 75740 23716 75796
rect 19836 73722 19892 73724
rect 19836 73670 19838 73722
rect 19838 73670 19890 73722
rect 19890 73670 19892 73722
rect 19836 73668 19892 73670
rect 19940 73722 19996 73724
rect 19940 73670 19942 73722
rect 19942 73670 19994 73722
rect 19994 73670 19996 73722
rect 19940 73668 19996 73670
rect 20044 73722 20100 73724
rect 20044 73670 20046 73722
rect 20046 73670 20098 73722
rect 20098 73670 20100 73722
rect 20044 73668 20100 73670
rect 19836 72154 19892 72156
rect 19836 72102 19838 72154
rect 19838 72102 19890 72154
rect 19890 72102 19892 72154
rect 19836 72100 19892 72102
rect 19940 72154 19996 72156
rect 19940 72102 19942 72154
rect 19942 72102 19994 72154
rect 19994 72102 19996 72154
rect 19940 72100 19996 72102
rect 20044 72154 20100 72156
rect 20044 72102 20046 72154
rect 20046 72102 20098 72154
rect 20098 72102 20100 72154
rect 20044 72100 20100 72102
rect 19836 70586 19892 70588
rect 19836 70534 19838 70586
rect 19838 70534 19890 70586
rect 19890 70534 19892 70586
rect 19836 70532 19892 70534
rect 19940 70586 19996 70588
rect 19940 70534 19942 70586
rect 19942 70534 19994 70586
rect 19994 70534 19996 70586
rect 19940 70532 19996 70534
rect 20044 70586 20100 70588
rect 20044 70534 20046 70586
rect 20046 70534 20098 70586
rect 20098 70534 20100 70586
rect 20044 70532 20100 70534
rect 19836 69018 19892 69020
rect 19836 68966 19838 69018
rect 19838 68966 19890 69018
rect 19890 68966 19892 69018
rect 19836 68964 19892 68966
rect 19940 69018 19996 69020
rect 19940 68966 19942 69018
rect 19942 68966 19994 69018
rect 19994 68966 19996 69018
rect 19940 68964 19996 68966
rect 20044 69018 20100 69020
rect 20044 68966 20046 69018
rect 20046 68966 20098 69018
rect 20098 68966 20100 69018
rect 20044 68964 20100 68966
rect 19836 67450 19892 67452
rect 19836 67398 19838 67450
rect 19838 67398 19890 67450
rect 19890 67398 19892 67450
rect 19836 67396 19892 67398
rect 19940 67450 19996 67452
rect 19940 67398 19942 67450
rect 19942 67398 19994 67450
rect 19994 67398 19996 67450
rect 19940 67396 19996 67398
rect 20044 67450 20100 67452
rect 20044 67398 20046 67450
rect 20046 67398 20098 67450
rect 20098 67398 20100 67450
rect 20044 67396 20100 67398
rect 19836 65882 19892 65884
rect 19836 65830 19838 65882
rect 19838 65830 19890 65882
rect 19890 65830 19892 65882
rect 19836 65828 19892 65830
rect 19940 65882 19996 65884
rect 19940 65830 19942 65882
rect 19942 65830 19994 65882
rect 19994 65830 19996 65882
rect 19940 65828 19996 65830
rect 20044 65882 20100 65884
rect 20044 65830 20046 65882
rect 20046 65830 20098 65882
rect 20098 65830 20100 65882
rect 20044 65828 20100 65830
rect 19836 64314 19892 64316
rect 19836 64262 19838 64314
rect 19838 64262 19890 64314
rect 19890 64262 19892 64314
rect 19836 64260 19892 64262
rect 19940 64314 19996 64316
rect 19940 64262 19942 64314
rect 19942 64262 19994 64314
rect 19994 64262 19996 64314
rect 19940 64260 19996 64262
rect 20044 64314 20100 64316
rect 20044 64262 20046 64314
rect 20046 64262 20098 64314
rect 20098 64262 20100 64314
rect 20044 64260 20100 64262
rect 19836 62746 19892 62748
rect 19836 62694 19838 62746
rect 19838 62694 19890 62746
rect 19890 62694 19892 62746
rect 19836 62692 19892 62694
rect 19940 62746 19996 62748
rect 19940 62694 19942 62746
rect 19942 62694 19994 62746
rect 19994 62694 19996 62746
rect 19940 62692 19996 62694
rect 20044 62746 20100 62748
rect 20044 62694 20046 62746
rect 20046 62694 20098 62746
rect 20098 62694 20100 62746
rect 20044 62692 20100 62694
rect 19836 61178 19892 61180
rect 19836 61126 19838 61178
rect 19838 61126 19890 61178
rect 19890 61126 19892 61178
rect 19836 61124 19892 61126
rect 19940 61178 19996 61180
rect 19940 61126 19942 61178
rect 19942 61126 19994 61178
rect 19994 61126 19996 61178
rect 19940 61124 19996 61126
rect 20044 61178 20100 61180
rect 20044 61126 20046 61178
rect 20046 61126 20098 61178
rect 20098 61126 20100 61178
rect 20044 61124 20100 61126
rect 19836 59610 19892 59612
rect 19836 59558 19838 59610
rect 19838 59558 19890 59610
rect 19890 59558 19892 59610
rect 19836 59556 19892 59558
rect 19940 59610 19996 59612
rect 19940 59558 19942 59610
rect 19942 59558 19994 59610
rect 19994 59558 19996 59610
rect 19940 59556 19996 59558
rect 20044 59610 20100 59612
rect 20044 59558 20046 59610
rect 20046 59558 20098 59610
rect 20098 59558 20100 59610
rect 20044 59556 20100 59558
rect 19836 58042 19892 58044
rect 19836 57990 19838 58042
rect 19838 57990 19890 58042
rect 19890 57990 19892 58042
rect 19836 57988 19892 57990
rect 19940 58042 19996 58044
rect 19940 57990 19942 58042
rect 19942 57990 19994 58042
rect 19994 57990 19996 58042
rect 19940 57988 19996 57990
rect 20044 58042 20100 58044
rect 20044 57990 20046 58042
rect 20046 57990 20098 58042
rect 20098 57990 20100 58042
rect 20044 57988 20100 57990
rect 19836 56474 19892 56476
rect 19836 56422 19838 56474
rect 19838 56422 19890 56474
rect 19890 56422 19892 56474
rect 19836 56420 19892 56422
rect 19940 56474 19996 56476
rect 19940 56422 19942 56474
rect 19942 56422 19994 56474
rect 19994 56422 19996 56474
rect 19940 56420 19996 56422
rect 20044 56474 20100 56476
rect 20044 56422 20046 56474
rect 20046 56422 20098 56474
rect 20098 56422 20100 56474
rect 20044 56420 20100 56422
rect 18396 23378 18452 23380
rect 18396 23326 18398 23378
rect 18398 23326 18450 23378
rect 18450 23326 18452 23378
rect 18396 23324 18452 23326
rect 18508 22764 18564 22820
rect 18508 21810 18564 21812
rect 18508 21758 18510 21810
rect 18510 21758 18562 21810
rect 18562 21758 18564 21810
rect 18508 21756 18564 21758
rect 18844 22316 18900 22372
rect 18620 20130 18676 20132
rect 18620 20078 18622 20130
rect 18622 20078 18674 20130
rect 18674 20078 18676 20130
rect 18620 20076 18676 20078
rect 16940 17724 16996 17780
rect 16716 6188 16772 6244
rect 16828 8540 16884 8596
rect 17948 19068 18004 19124
rect 17724 17778 17780 17780
rect 17724 17726 17726 17778
rect 17726 17726 17778 17778
rect 17778 17726 17780 17778
rect 17724 17724 17780 17726
rect 17836 17388 17892 17444
rect 16940 7698 16996 7700
rect 16940 7646 16942 7698
rect 16942 7646 16994 7698
rect 16994 7646 16996 7698
rect 16940 7644 16996 7646
rect 16828 5740 16884 5796
rect 16604 5292 16660 5348
rect 16716 5234 16772 5236
rect 16716 5182 16718 5234
rect 16718 5182 16770 5234
rect 16770 5182 16772 5234
rect 16716 5180 16772 5182
rect 16492 5068 16548 5124
rect 16044 4620 16100 4676
rect 16044 4172 16100 4228
rect 15708 3948 15764 4004
rect 16268 4060 16324 4116
rect 15372 3276 15428 3332
rect 15260 2716 15316 2772
rect 15708 3052 15764 3108
rect 17948 12066 18004 12068
rect 17948 12014 17950 12066
rect 17950 12014 18002 12066
rect 18002 12014 18004 12066
rect 17948 12012 18004 12014
rect 19836 54906 19892 54908
rect 19836 54854 19838 54906
rect 19838 54854 19890 54906
rect 19890 54854 19892 54906
rect 19836 54852 19892 54854
rect 19940 54906 19996 54908
rect 19940 54854 19942 54906
rect 19942 54854 19994 54906
rect 19994 54854 19996 54906
rect 19940 54852 19996 54854
rect 20044 54906 20100 54908
rect 20044 54854 20046 54906
rect 20046 54854 20098 54906
rect 20098 54854 20100 54906
rect 20044 54852 20100 54854
rect 19836 53338 19892 53340
rect 19836 53286 19838 53338
rect 19838 53286 19890 53338
rect 19890 53286 19892 53338
rect 19836 53284 19892 53286
rect 19940 53338 19996 53340
rect 19940 53286 19942 53338
rect 19942 53286 19994 53338
rect 19994 53286 19996 53338
rect 19940 53284 19996 53286
rect 20044 53338 20100 53340
rect 20044 53286 20046 53338
rect 20046 53286 20098 53338
rect 20098 53286 20100 53338
rect 20044 53284 20100 53286
rect 19836 51770 19892 51772
rect 19836 51718 19838 51770
rect 19838 51718 19890 51770
rect 19890 51718 19892 51770
rect 19836 51716 19892 51718
rect 19940 51770 19996 51772
rect 19940 51718 19942 51770
rect 19942 51718 19994 51770
rect 19994 51718 19996 51770
rect 19940 51716 19996 51718
rect 20044 51770 20100 51772
rect 20044 51718 20046 51770
rect 20046 51718 20098 51770
rect 20098 51718 20100 51770
rect 20044 51716 20100 51718
rect 19836 50202 19892 50204
rect 19836 50150 19838 50202
rect 19838 50150 19890 50202
rect 19890 50150 19892 50202
rect 19836 50148 19892 50150
rect 19940 50202 19996 50204
rect 19940 50150 19942 50202
rect 19942 50150 19994 50202
rect 19994 50150 19996 50202
rect 19940 50148 19996 50150
rect 20044 50202 20100 50204
rect 20044 50150 20046 50202
rect 20046 50150 20098 50202
rect 20098 50150 20100 50202
rect 20044 50148 20100 50150
rect 19836 48634 19892 48636
rect 19836 48582 19838 48634
rect 19838 48582 19890 48634
rect 19890 48582 19892 48634
rect 19836 48580 19892 48582
rect 19940 48634 19996 48636
rect 19940 48582 19942 48634
rect 19942 48582 19994 48634
rect 19994 48582 19996 48634
rect 19940 48580 19996 48582
rect 20044 48634 20100 48636
rect 20044 48582 20046 48634
rect 20046 48582 20098 48634
rect 20098 48582 20100 48634
rect 20044 48580 20100 48582
rect 19836 47066 19892 47068
rect 19836 47014 19838 47066
rect 19838 47014 19890 47066
rect 19890 47014 19892 47066
rect 19836 47012 19892 47014
rect 19940 47066 19996 47068
rect 19940 47014 19942 47066
rect 19942 47014 19994 47066
rect 19994 47014 19996 47066
rect 19940 47012 19996 47014
rect 20044 47066 20100 47068
rect 20044 47014 20046 47066
rect 20046 47014 20098 47066
rect 20098 47014 20100 47066
rect 20044 47012 20100 47014
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 20972 40460 21028 40516
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 20972 27916 21028 27972
rect 23884 75628 23940 75684
rect 31836 76300 31892 76356
rect 24780 75794 24836 75796
rect 24780 75742 24782 75794
rect 24782 75742 24834 75794
rect 24834 75742 24836 75794
rect 24780 75740 24836 75742
rect 25228 75682 25284 75684
rect 25228 75630 25230 75682
rect 25230 75630 25282 75682
rect 25282 75630 25284 75682
rect 25228 75628 25284 75630
rect 30156 75628 30212 75684
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 19292 24610 19348 24612
rect 19292 24558 19294 24610
rect 19294 24558 19346 24610
rect 19346 24558 19348 24610
rect 19292 24556 19348 24558
rect 19740 24668 19796 24724
rect 20300 24722 20356 24724
rect 20300 24670 20302 24722
rect 20302 24670 20354 24722
rect 20354 24670 20356 24722
rect 20300 24668 20356 24670
rect 21196 24668 21252 24724
rect 19740 24498 19796 24500
rect 19740 24446 19742 24498
rect 19742 24446 19794 24498
rect 19794 24446 19796 24498
rect 19740 24444 19796 24446
rect 21868 24444 21924 24500
rect 21196 23884 21252 23940
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 19292 23436 19348 23492
rect 20300 23436 20356 23492
rect 21532 23548 21588 23604
rect 19068 20076 19124 20132
rect 18956 20018 19012 20020
rect 18956 19966 18958 20018
rect 18958 19966 19010 20018
rect 19010 19966 19012 20018
rect 18956 19964 19012 19966
rect 19068 19794 19124 19796
rect 19068 19742 19070 19794
rect 19070 19742 19122 19794
rect 19122 19742 19124 19794
rect 19068 19740 19124 19742
rect 18956 19068 19012 19124
rect 18732 17724 18788 17780
rect 20076 22988 20132 23044
rect 20636 23042 20692 23044
rect 20636 22990 20638 23042
rect 20638 22990 20690 23042
rect 20690 22990 20692 23042
rect 20636 22988 20692 22990
rect 20076 22764 20132 22820
rect 20412 22652 20468 22708
rect 21420 22652 21476 22708
rect 21644 22652 21700 22708
rect 20412 22258 20468 22260
rect 20412 22206 20414 22258
rect 20414 22206 20466 22258
rect 20466 22206 20468 22258
rect 20412 22204 20468 22206
rect 19852 22092 19908 22148
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 19292 19628 19348 19684
rect 19628 20578 19684 20580
rect 19628 20526 19630 20578
rect 19630 20526 19682 20578
rect 19682 20526 19684 20578
rect 19628 20524 19684 20526
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 20524 20578 20580 20580
rect 20524 20526 20526 20578
rect 20526 20526 20578 20578
rect 20578 20526 20580 20578
rect 20524 20524 20580 20526
rect 19516 20018 19572 20020
rect 19516 19966 19518 20018
rect 19518 19966 19570 20018
rect 19570 19966 19572 20018
rect 19516 19964 19572 19966
rect 20300 20076 20356 20132
rect 19628 19852 19684 19908
rect 20748 20076 20804 20132
rect 20972 19906 21028 19908
rect 20972 19854 20974 19906
rect 20974 19854 21026 19906
rect 21026 19854 21028 19906
rect 20972 19852 21028 19854
rect 21756 20076 21812 20132
rect 19628 19068 19684 19124
rect 19516 18956 19572 19012
rect 21532 19122 21588 19124
rect 21532 19070 21534 19122
rect 21534 19070 21586 19122
rect 21586 19070 21588 19122
rect 21532 19068 21588 19070
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 21532 18732 21588 18788
rect 19404 17388 19460 17444
rect 19740 17442 19796 17444
rect 19740 17390 19742 17442
rect 19742 17390 19794 17442
rect 19794 17390 19796 17442
rect 19740 17388 19796 17390
rect 20412 17442 20468 17444
rect 20412 17390 20414 17442
rect 20414 17390 20466 17442
rect 20466 17390 20468 17442
rect 20412 17388 20468 17390
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 20412 17164 20468 17220
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 18620 13580 18676 13636
rect 18620 11116 18676 11172
rect 18284 10498 18340 10500
rect 18284 10446 18286 10498
rect 18286 10446 18338 10498
rect 18338 10446 18340 10498
rect 18284 10444 18340 10446
rect 18284 9266 18340 9268
rect 18284 9214 18286 9266
rect 18286 9214 18338 9266
rect 18338 9214 18340 9266
rect 18284 9212 18340 9214
rect 17724 8204 17780 8260
rect 18172 8930 18228 8932
rect 18172 8878 18174 8930
rect 18174 8878 18226 8930
rect 18226 8878 18228 8930
rect 18172 8876 18228 8878
rect 18172 8370 18228 8372
rect 18172 8318 18174 8370
rect 18174 8318 18226 8370
rect 18226 8318 18228 8370
rect 18172 8316 18228 8318
rect 18284 8258 18340 8260
rect 18284 8206 18286 8258
rect 18286 8206 18338 8258
rect 18338 8206 18340 8258
rect 18284 8204 18340 8206
rect 17836 7644 17892 7700
rect 17724 7474 17780 7476
rect 17724 7422 17726 7474
rect 17726 7422 17778 7474
rect 17778 7422 17780 7474
rect 17724 7420 17780 7422
rect 17724 6972 17780 7028
rect 17388 5906 17444 5908
rect 17388 5854 17390 5906
rect 17390 5854 17442 5906
rect 17442 5854 17444 5906
rect 17388 5852 17444 5854
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 21420 13692 21476 13748
rect 19628 13580 19684 13636
rect 19516 12908 19572 12964
rect 20188 12738 20244 12740
rect 20188 12686 20190 12738
rect 20190 12686 20242 12738
rect 20242 12686 20244 12738
rect 20188 12684 20244 12686
rect 19836 12570 19892 12572
rect 19516 12460 19572 12516
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19852 12236 19908 12292
rect 19292 12066 19348 12068
rect 19292 12014 19294 12066
rect 19294 12014 19346 12066
rect 19346 12014 19348 12066
rect 19292 12012 19348 12014
rect 20412 12236 20468 12292
rect 20972 12908 21028 12964
rect 19068 11340 19124 11396
rect 18732 9324 18788 9380
rect 18396 7756 18452 7812
rect 18844 8988 18900 9044
rect 18508 7532 18564 7588
rect 18508 7362 18564 7364
rect 18508 7310 18510 7362
rect 18510 7310 18562 7362
rect 18562 7310 18564 7362
rect 18508 7308 18564 7310
rect 19516 10498 19572 10500
rect 19516 10446 19518 10498
rect 19518 10446 19570 10498
rect 19570 10446 19572 10498
rect 19516 10444 19572 10446
rect 19180 9266 19236 9268
rect 19180 9214 19182 9266
rect 19182 9214 19234 9266
rect 19234 9214 19236 9266
rect 19180 9212 19236 9214
rect 19852 11452 19908 11508
rect 20300 11788 20356 11844
rect 20636 11506 20692 11508
rect 20636 11454 20638 11506
rect 20638 11454 20690 11506
rect 20690 11454 20692 11506
rect 20636 11452 20692 11454
rect 19740 11170 19796 11172
rect 19740 11118 19742 11170
rect 19742 11118 19794 11170
rect 19794 11118 19796 11170
rect 19740 11116 19796 11118
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 20188 9884 20244 9940
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 19628 9212 19684 9268
rect 19516 9042 19572 9044
rect 19516 8990 19518 9042
rect 19518 8990 19570 9042
rect 19570 8990 19572 9042
rect 19516 8988 19572 8990
rect 19180 8876 19236 8932
rect 20300 8930 20356 8932
rect 20300 8878 20302 8930
rect 20302 8878 20354 8930
rect 20354 8878 20356 8930
rect 20300 8876 20356 8878
rect 19964 8316 20020 8372
rect 20972 10220 21028 10276
rect 20748 9938 20804 9940
rect 20748 9886 20750 9938
rect 20750 9886 20802 9938
rect 20802 9886 20804 9938
rect 20748 9884 20804 9886
rect 19292 8092 19348 8148
rect 19068 6972 19124 7028
rect 19180 7756 19236 7812
rect 18844 6636 18900 6692
rect 18508 6300 18564 6356
rect 18284 6130 18340 6132
rect 18284 6078 18286 6130
rect 18286 6078 18338 6130
rect 18338 6078 18340 6130
rect 18284 6076 18340 6078
rect 18396 5964 18452 6020
rect 17388 5180 17444 5236
rect 18284 5292 18340 5348
rect 17948 4956 18004 5012
rect 17724 4396 17780 4452
rect 17052 3500 17108 3556
rect 16380 2716 16436 2772
rect 17500 4060 17556 4116
rect 17388 3164 17444 3220
rect 17276 2268 17332 2324
rect 18284 4450 18340 4452
rect 18284 4398 18286 4450
rect 18286 4398 18338 4450
rect 18338 4398 18340 4450
rect 18284 4396 18340 4398
rect 17948 4060 18004 4116
rect 17836 3948 17892 4004
rect 18396 3724 18452 3780
rect 18620 5852 18676 5908
rect 18956 6466 19012 6468
rect 18956 6414 18958 6466
rect 18958 6414 19010 6466
rect 19010 6414 19012 6466
rect 18956 6412 19012 6414
rect 18732 5180 18788 5236
rect 18956 4338 19012 4340
rect 18956 4286 18958 4338
rect 18958 4286 19010 4338
rect 19010 4286 19012 4338
rect 18956 4284 19012 4286
rect 19740 8146 19796 8148
rect 19740 8094 19742 8146
rect 19742 8094 19794 8146
rect 19794 8094 19796 8146
rect 19740 8092 19796 8094
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 19964 7644 20020 7700
rect 19628 7474 19684 7476
rect 19628 7422 19630 7474
rect 19630 7422 19682 7474
rect 19682 7422 19684 7474
rect 19628 7420 19684 7422
rect 19516 7084 19572 7140
rect 19404 6466 19460 6468
rect 19404 6414 19406 6466
rect 19406 6414 19458 6466
rect 19458 6414 19460 6466
rect 19404 6412 19460 6414
rect 19628 6636 19684 6692
rect 19852 6636 19908 6692
rect 20636 8764 20692 8820
rect 20412 7698 20468 7700
rect 20412 7646 20414 7698
rect 20414 7646 20466 7698
rect 20466 7646 20468 7698
rect 20412 7644 20468 7646
rect 19964 6412 20020 6468
rect 20188 6860 20244 6916
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 18508 3500 18564 3556
rect 18620 4060 18676 4116
rect 19404 5292 19460 5348
rect 19628 5794 19684 5796
rect 19628 5742 19630 5794
rect 19630 5742 19682 5794
rect 19682 5742 19684 5794
rect 19628 5740 19684 5742
rect 19404 5122 19460 5124
rect 19404 5070 19406 5122
rect 19406 5070 19458 5122
rect 19458 5070 19460 5122
rect 19404 5068 19460 5070
rect 20076 5068 20132 5124
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 19964 4508 20020 4564
rect 19404 4284 19460 4340
rect 19180 4060 19236 4116
rect 19068 3836 19124 3892
rect 18844 3330 18900 3332
rect 18844 3278 18846 3330
rect 18846 3278 18898 3330
rect 18898 3278 18900 3330
rect 18844 3276 18900 3278
rect 19964 4060 20020 4116
rect 19180 3554 19236 3556
rect 19180 3502 19182 3554
rect 19182 3502 19234 3554
rect 19234 3502 19236 3554
rect 19180 3500 19236 3502
rect 19404 3612 19460 3668
rect 19964 3612 20020 3668
rect 19516 3500 19572 3556
rect 20636 8428 20692 8484
rect 20412 5404 20468 5460
rect 20300 4508 20356 4564
rect 20412 4396 20468 4452
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 20748 8370 20804 8372
rect 20748 8318 20750 8370
rect 20750 8318 20802 8370
rect 20802 8318 20804 8370
rect 20748 8316 20804 8318
rect 20860 7698 20916 7700
rect 20860 7646 20862 7698
rect 20862 7646 20914 7698
rect 20914 7646 20916 7698
rect 20860 7644 20916 7646
rect 20972 6860 21028 6916
rect 20748 5346 20804 5348
rect 20748 5294 20750 5346
rect 20750 5294 20802 5346
rect 20802 5294 20804 5346
rect 20748 5292 20804 5294
rect 20636 4562 20692 4564
rect 20636 4510 20638 4562
rect 20638 4510 20690 4562
rect 20690 4510 20692 4562
rect 20636 4508 20692 4510
rect 21420 13074 21476 13076
rect 21420 13022 21422 13074
rect 21422 13022 21474 13074
rect 21474 13022 21476 13074
rect 21420 13020 21476 13022
rect 21420 12684 21476 12740
rect 21756 19234 21812 19236
rect 21756 19182 21758 19234
rect 21758 19182 21810 19234
rect 21810 19182 21812 19234
rect 21756 19180 21812 19182
rect 22092 19740 22148 19796
rect 23100 24050 23156 24052
rect 23100 23998 23102 24050
rect 23102 23998 23154 24050
rect 23154 23998 23156 24050
rect 23100 23996 23156 23998
rect 23324 23714 23380 23716
rect 23324 23662 23326 23714
rect 23326 23662 23378 23714
rect 23378 23662 23380 23714
rect 23324 23660 23380 23662
rect 22316 23548 22372 23604
rect 23772 23548 23828 23604
rect 23996 23938 24052 23940
rect 23996 23886 23998 23938
rect 23998 23886 24050 23938
rect 24050 23886 24052 23938
rect 23996 23884 24052 23886
rect 23660 23324 23716 23380
rect 23996 23324 24052 23380
rect 23548 23154 23604 23156
rect 23548 23102 23550 23154
rect 23550 23102 23602 23154
rect 23602 23102 23604 23154
rect 23548 23100 23604 23102
rect 22428 20412 22484 20468
rect 22988 20412 23044 20468
rect 23436 20524 23492 20580
rect 22764 19122 22820 19124
rect 22764 19070 22766 19122
rect 22766 19070 22818 19122
rect 22818 19070 22820 19122
rect 22764 19068 22820 19070
rect 23324 19122 23380 19124
rect 23324 19070 23326 19122
rect 23326 19070 23378 19122
rect 23378 19070 23380 19122
rect 23324 19068 23380 19070
rect 22204 18396 22260 18452
rect 21644 17724 21700 17780
rect 21644 17164 21700 17220
rect 23996 22876 24052 22932
rect 26908 40348 26964 40404
rect 26908 38892 26964 38948
rect 26908 37324 26964 37380
rect 26908 36316 26964 36372
rect 28476 33068 28532 33124
rect 28476 31612 28532 31668
rect 30156 28028 30212 28084
rect 33516 75852 33572 75908
rect 35084 76466 35140 76468
rect 35084 76414 35086 76466
rect 35086 76414 35138 76466
rect 35138 76414 35140 76466
rect 35084 76412 35140 76414
rect 35756 76412 35812 76468
rect 35196 76074 35252 76076
rect 35196 76022 35198 76074
rect 35198 76022 35250 76074
rect 35250 76022 35252 76074
rect 35196 76020 35252 76022
rect 35300 76074 35356 76076
rect 35300 76022 35302 76074
rect 35302 76022 35354 76074
rect 35354 76022 35356 76074
rect 35300 76020 35356 76022
rect 35404 76074 35460 76076
rect 35404 76022 35406 76074
rect 35406 76022 35458 76074
rect 35458 76022 35460 76074
rect 35404 76020 35460 76022
rect 33516 75682 33572 75684
rect 33516 75630 33518 75682
rect 33518 75630 33570 75682
rect 33570 75630 33572 75682
rect 33516 75628 33572 75630
rect 33964 74956 34020 75012
rect 31836 27692 31892 27748
rect 34972 75010 35028 75012
rect 34972 74958 34974 75010
rect 34974 74958 35026 75010
rect 35026 74958 35028 75010
rect 34972 74956 35028 74958
rect 35756 74786 35812 74788
rect 35756 74734 35758 74786
rect 35758 74734 35810 74786
rect 35810 74734 35812 74786
rect 35756 74732 35812 74734
rect 35196 74506 35252 74508
rect 35196 74454 35198 74506
rect 35198 74454 35250 74506
rect 35250 74454 35252 74506
rect 35196 74452 35252 74454
rect 35300 74506 35356 74508
rect 35300 74454 35302 74506
rect 35302 74454 35354 74506
rect 35354 74454 35356 74506
rect 35300 74452 35356 74454
rect 35404 74506 35460 74508
rect 35404 74454 35406 74506
rect 35406 74454 35458 74506
rect 35458 74454 35460 74506
rect 35404 74452 35460 74454
rect 35196 72938 35252 72940
rect 35196 72886 35198 72938
rect 35198 72886 35250 72938
rect 35250 72886 35252 72938
rect 35196 72884 35252 72886
rect 35300 72938 35356 72940
rect 35300 72886 35302 72938
rect 35302 72886 35354 72938
rect 35354 72886 35356 72938
rect 35300 72884 35356 72886
rect 35404 72938 35460 72940
rect 35404 72886 35406 72938
rect 35406 72886 35458 72938
rect 35458 72886 35460 72938
rect 35404 72884 35460 72886
rect 35196 71370 35252 71372
rect 35196 71318 35198 71370
rect 35198 71318 35250 71370
rect 35250 71318 35252 71370
rect 35196 71316 35252 71318
rect 35300 71370 35356 71372
rect 35300 71318 35302 71370
rect 35302 71318 35354 71370
rect 35354 71318 35356 71370
rect 35300 71316 35356 71318
rect 35404 71370 35460 71372
rect 35404 71318 35406 71370
rect 35406 71318 35458 71370
rect 35458 71318 35460 71370
rect 35404 71316 35460 71318
rect 35196 69802 35252 69804
rect 35196 69750 35198 69802
rect 35198 69750 35250 69802
rect 35250 69750 35252 69802
rect 35196 69748 35252 69750
rect 35300 69802 35356 69804
rect 35300 69750 35302 69802
rect 35302 69750 35354 69802
rect 35354 69750 35356 69802
rect 35300 69748 35356 69750
rect 35404 69802 35460 69804
rect 35404 69750 35406 69802
rect 35406 69750 35458 69802
rect 35458 69750 35460 69802
rect 35404 69748 35460 69750
rect 35196 68234 35252 68236
rect 35196 68182 35198 68234
rect 35198 68182 35250 68234
rect 35250 68182 35252 68234
rect 35196 68180 35252 68182
rect 35300 68234 35356 68236
rect 35300 68182 35302 68234
rect 35302 68182 35354 68234
rect 35354 68182 35356 68234
rect 35300 68180 35356 68182
rect 35404 68234 35460 68236
rect 35404 68182 35406 68234
rect 35406 68182 35458 68234
rect 35458 68182 35460 68234
rect 35404 68180 35460 68182
rect 35196 66666 35252 66668
rect 35196 66614 35198 66666
rect 35198 66614 35250 66666
rect 35250 66614 35252 66666
rect 35196 66612 35252 66614
rect 35300 66666 35356 66668
rect 35300 66614 35302 66666
rect 35302 66614 35354 66666
rect 35354 66614 35356 66666
rect 35300 66612 35356 66614
rect 35404 66666 35460 66668
rect 35404 66614 35406 66666
rect 35406 66614 35458 66666
rect 35458 66614 35460 66666
rect 35404 66612 35460 66614
rect 35196 65098 35252 65100
rect 35196 65046 35198 65098
rect 35198 65046 35250 65098
rect 35250 65046 35252 65098
rect 35196 65044 35252 65046
rect 35300 65098 35356 65100
rect 35300 65046 35302 65098
rect 35302 65046 35354 65098
rect 35354 65046 35356 65098
rect 35300 65044 35356 65046
rect 35404 65098 35460 65100
rect 35404 65046 35406 65098
rect 35406 65046 35458 65098
rect 35458 65046 35460 65098
rect 35404 65044 35460 65046
rect 35196 63530 35252 63532
rect 35196 63478 35198 63530
rect 35198 63478 35250 63530
rect 35250 63478 35252 63530
rect 35196 63476 35252 63478
rect 35300 63530 35356 63532
rect 35300 63478 35302 63530
rect 35302 63478 35354 63530
rect 35354 63478 35356 63530
rect 35300 63476 35356 63478
rect 35404 63530 35460 63532
rect 35404 63478 35406 63530
rect 35406 63478 35458 63530
rect 35458 63478 35460 63530
rect 35404 63476 35460 63478
rect 35196 61962 35252 61964
rect 35196 61910 35198 61962
rect 35198 61910 35250 61962
rect 35250 61910 35252 61962
rect 35196 61908 35252 61910
rect 35300 61962 35356 61964
rect 35300 61910 35302 61962
rect 35302 61910 35354 61962
rect 35354 61910 35356 61962
rect 35300 61908 35356 61910
rect 35404 61962 35460 61964
rect 35404 61910 35406 61962
rect 35406 61910 35458 61962
rect 35458 61910 35460 61962
rect 35404 61908 35460 61910
rect 35196 60394 35252 60396
rect 35196 60342 35198 60394
rect 35198 60342 35250 60394
rect 35250 60342 35252 60394
rect 35196 60340 35252 60342
rect 35300 60394 35356 60396
rect 35300 60342 35302 60394
rect 35302 60342 35354 60394
rect 35354 60342 35356 60394
rect 35300 60340 35356 60342
rect 35404 60394 35460 60396
rect 35404 60342 35406 60394
rect 35406 60342 35458 60394
rect 35458 60342 35460 60394
rect 35404 60340 35460 60342
rect 35196 58826 35252 58828
rect 35196 58774 35198 58826
rect 35198 58774 35250 58826
rect 35250 58774 35252 58826
rect 35196 58772 35252 58774
rect 35300 58826 35356 58828
rect 35300 58774 35302 58826
rect 35302 58774 35354 58826
rect 35354 58774 35356 58826
rect 35300 58772 35356 58774
rect 35404 58826 35460 58828
rect 35404 58774 35406 58826
rect 35406 58774 35458 58826
rect 35458 58774 35460 58826
rect 35404 58772 35460 58774
rect 35196 57258 35252 57260
rect 35196 57206 35198 57258
rect 35198 57206 35250 57258
rect 35250 57206 35252 57258
rect 35196 57204 35252 57206
rect 35300 57258 35356 57260
rect 35300 57206 35302 57258
rect 35302 57206 35354 57258
rect 35354 57206 35356 57258
rect 35300 57204 35356 57206
rect 35404 57258 35460 57260
rect 35404 57206 35406 57258
rect 35406 57206 35458 57258
rect 35458 57206 35460 57258
rect 35404 57204 35460 57206
rect 35196 55690 35252 55692
rect 35196 55638 35198 55690
rect 35198 55638 35250 55690
rect 35250 55638 35252 55690
rect 35196 55636 35252 55638
rect 35300 55690 35356 55692
rect 35300 55638 35302 55690
rect 35302 55638 35354 55690
rect 35354 55638 35356 55690
rect 35300 55636 35356 55638
rect 35404 55690 35460 55692
rect 35404 55638 35406 55690
rect 35406 55638 35458 55690
rect 35458 55638 35460 55690
rect 35404 55636 35460 55638
rect 33516 27580 33572 27636
rect 33852 27916 33908 27972
rect 35196 54122 35252 54124
rect 35196 54070 35198 54122
rect 35198 54070 35250 54122
rect 35250 54070 35252 54122
rect 35196 54068 35252 54070
rect 35300 54122 35356 54124
rect 35300 54070 35302 54122
rect 35302 54070 35354 54122
rect 35354 54070 35356 54122
rect 35300 54068 35356 54070
rect 35404 54122 35460 54124
rect 35404 54070 35406 54122
rect 35406 54070 35458 54122
rect 35458 54070 35460 54122
rect 35404 54068 35460 54070
rect 35196 52554 35252 52556
rect 35196 52502 35198 52554
rect 35198 52502 35250 52554
rect 35250 52502 35252 52554
rect 35196 52500 35252 52502
rect 35300 52554 35356 52556
rect 35300 52502 35302 52554
rect 35302 52502 35354 52554
rect 35354 52502 35356 52554
rect 35300 52500 35356 52502
rect 35404 52554 35460 52556
rect 35404 52502 35406 52554
rect 35406 52502 35458 52554
rect 35458 52502 35460 52554
rect 35404 52500 35460 52502
rect 35196 50986 35252 50988
rect 35196 50934 35198 50986
rect 35198 50934 35250 50986
rect 35250 50934 35252 50986
rect 35196 50932 35252 50934
rect 35300 50986 35356 50988
rect 35300 50934 35302 50986
rect 35302 50934 35354 50986
rect 35354 50934 35356 50986
rect 35300 50932 35356 50934
rect 35404 50986 35460 50988
rect 35404 50934 35406 50986
rect 35406 50934 35458 50986
rect 35458 50934 35460 50986
rect 35404 50932 35460 50934
rect 35196 49418 35252 49420
rect 35196 49366 35198 49418
rect 35198 49366 35250 49418
rect 35250 49366 35252 49418
rect 35196 49364 35252 49366
rect 35300 49418 35356 49420
rect 35300 49366 35302 49418
rect 35302 49366 35354 49418
rect 35354 49366 35356 49418
rect 35300 49364 35356 49366
rect 35404 49418 35460 49420
rect 35404 49366 35406 49418
rect 35406 49366 35458 49418
rect 35458 49366 35460 49418
rect 35404 49364 35460 49366
rect 35196 47850 35252 47852
rect 35196 47798 35198 47850
rect 35198 47798 35250 47850
rect 35250 47798 35252 47850
rect 35196 47796 35252 47798
rect 35300 47850 35356 47852
rect 35300 47798 35302 47850
rect 35302 47798 35354 47850
rect 35354 47798 35356 47850
rect 35300 47796 35356 47798
rect 35404 47850 35460 47852
rect 35404 47798 35406 47850
rect 35406 47798 35458 47850
rect 35458 47798 35460 47850
rect 35404 47796 35460 47798
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 36764 75740 36820 75796
rect 37324 75794 37380 75796
rect 37324 75742 37326 75794
rect 37326 75742 37378 75794
rect 37378 75742 37380 75794
rect 37324 75740 37380 75742
rect 37884 75794 37940 75796
rect 37884 75742 37886 75794
rect 37886 75742 37938 75794
rect 37938 75742 37940 75794
rect 37884 75740 37940 75742
rect 36092 29036 36148 29092
rect 35980 28028 36036 28084
rect 34860 27916 34916 27972
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 33740 26460 33796 26516
rect 34300 26460 34356 26516
rect 34300 26124 34356 26180
rect 25564 25676 25620 25732
rect 26572 25676 26628 25732
rect 31836 25452 31892 25508
rect 24780 24556 24836 24612
rect 25676 24610 25732 24612
rect 25676 24558 25678 24610
rect 25678 24558 25730 24610
rect 25730 24558 25732 24610
rect 25676 24556 25732 24558
rect 24332 23324 24388 23380
rect 25228 23324 25284 23380
rect 24444 23100 24500 23156
rect 26124 23378 26180 23380
rect 26124 23326 26126 23378
rect 26126 23326 26178 23378
rect 26178 23326 26180 23378
rect 26124 23324 26180 23326
rect 26572 23324 26628 23380
rect 24668 22652 24724 22708
rect 24668 21756 24724 21812
rect 25564 23154 25620 23156
rect 25564 23102 25566 23154
rect 25566 23102 25618 23154
rect 25618 23102 25620 23154
rect 25564 23100 25620 23102
rect 25340 22876 25396 22932
rect 25564 22652 25620 22708
rect 24108 20578 24164 20580
rect 24108 20526 24110 20578
rect 24110 20526 24162 20578
rect 24162 20526 24164 20578
rect 24108 20524 24164 20526
rect 23548 19010 23604 19012
rect 23548 18958 23550 19010
rect 23550 18958 23602 19010
rect 23602 18958 23604 19010
rect 23548 18956 23604 18958
rect 24668 21474 24724 21476
rect 24668 21422 24670 21474
rect 24670 21422 24722 21474
rect 24722 21422 24724 21474
rect 24668 21420 24724 21422
rect 25340 21420 25396 21476
rect 27692 24556 27748 24612
rect 30380 24610 30436 24612
rect 30380 24558 30382 24610
rect 30382 24558 30434 24610
rect 30434 24558 30436 24610
rect 30380 24556 30436 24558
rect 27580 23714 27636 23716
rect 27580 23662 27582 23714
rect 27582 23662 27634 23714
rect 27634 23662 27636 23714
rect 27580 23660 27636 23662
rect 28028 23378 28084 23380
rect 28028 23326 28030 23378
rect 28030 23326 28082 23378
rect 28082 23326 28084 23378
rect 28028 23324 28084 23326
rect 27356 23154 27412 23156
rect 27356 23102 27358 23154
rect 27358 23102 27410 23154
rect 27410 23102 27412 23154
rect 27356 23100 27412 23102
rect 27804 23154 27860 23156
rect 27804 23102 27806 23154
rect 27806 23102 27858 23154
rect 27858 23102 27860 23154
rect 27804 23100 27860 23102
rect 27916 23042 27972 23044
rect 27916 22990 27918 23042
rect 27918 22990 27970 23042
rect 27970 22990 27972 23042
rect 27916 22988 27972 22990
rect 27132 22652 27188 22708
rect 29148 23042 29204 23044
rect 29148 22990 29150 23042
rect 29150 22990 29202 23042
rect 29202 22990 29204 23042
rect 29148 22988 29204 22990
rect 31724 23154 31780 23156
rect 31724 23102 31726 23154
rect 31726 23102 31778 23154
rect 31778 23102 31780 23154
rect 31724 23100 31780 23102
rect 28364 22652 28420 22708
rect 29036 22652 29092 22708
rect 28364 22482 28420 22484
rect 28364 22430 28366 22482
rect 28366 22430 28418 22482
rect 28418 22430 28420 22482
rect 28364 22428 28420 22430
rect 29148 22482 29204 22484
rect 29148 22430 29150 22482
rect 29150 22430 29202 22482
rect 29202 22430 29204 22482
rect 29148 22428 29204 22430
rect 24220 19964 24276 20020
rect 24780 20412 24836 20468
rect 25340 20578 25396 20580
rect 25340 20526 25342 20578
rect 25342 20526 25394 20578
rect 25394 20526 25396 20578
rect 25340 20524 25396 20526
rect 25564 20578 25620 20580
rect 25564 20526 25566 20578
rect 25566 20526 25618 20578
rect 25618 20526 25620 20578
rect 25564 20524 25620 20526
rect 25228 20018 25284 20020
rect 25228 19966 25230 20018
rect 25230 19966 25282 20018
rect 25282 19966 25284 20018
rect 25228 19964 25284 19966
rect 24108 19628 24164 19684
rect 23660 18732 23716 18788
rect 23996 19068 24052 19124
rect 22316 17778 22372 17780
rect 22316 17726 22318 17778
rect 22318 17726 22370 17778
rect 22370 17726 22372 17778
rect 22316 17724 22372 17726
rect 24108 19010 24164 19012
rect 24108 18958 24110 19010
rect 24110 18958 24162 19010
rect 24162 18958 24164 19010
rect 24108 18956 24164 18958
rect 24444 19122 24500 19124
rect 24444 19070 24446 19122
rect 24446 19070 24498 19122
rect 24498 19070 24500 19122
rect 24444 19068 24500 19070
rect 24332 18732 24388 18788
rect 24668 18284 24724 18340
rect 23996 17948 24052 18004
rect 25452 19068 25508 19124
rect 25564 19180 25620 19236
rect 25340 18450 25396 18452
rect 25340 18398 25342 18450
rect 25342 18398 25394 18450
rect 25394 18398 25396 18450
rect 25340 18396 25396 18398
rect 25116 17948 25172 18004
rect 25004 17724 25060 17780
rect 23772 15820 23828 15876
rect 21756 13356 21812 13412
rect 22540 13020 22596 13076
rect 21532 11452 21588 11508
rect 22540 12012 22596 12068
rect 22092 11394 22148 11396
rect 22092 11342 22094 11394
rect 22094 11342 22146 11394
rect 22146 11342 22148 11394
rect 22092 11340 22148 11342
rect 22092 11116 22148 11172
rect 21644 8988 21700 9044
rect 21756 7084 21812 7140
rect 21532 6578 21588 6580
rect 21532 6526 21534 6578
rect 21534 6526 21586 6578
rect 21586 6526 21588 6578
rect 21532 6524 21588 6526
rect 21420 6412 21476 6468
rect 21084 5740 21140 5796
rect 20748 4060 20804 4116
rect 20524 3948 20580 4004
rect 21196 5628 21252 5684
rect 21420 5292 21476 5348
rect 21196 5180 21252 5236
rect 21308 4508 21364 4564
rect 21084 3836 21140 3892
rect 21196 4172 21252 4228
rect 21868 6748 21924 6804
rect 21868 6524 21924 6580
rect 22204 8428 22260 8484
rect 22540 10498 22596 10500
rect 22540 10446 22542 10498
rect 22542 10446 22594 10498
rect 22594 10446 22596 10498
rect 22540 10444 22596 10446
rect 23436 13746 23492 13748
rect 23436 13694 23438 13746
rect 23438 13694 23490 13746
rect 23490 13694 23492 13746
rect 23436 13692 23492 13694
rect 22988 13356 23044 13412
rect 25004 13356 25060 13412
rect 23772 13020 23828 13076
rect 25452 13244 25508 13300
rect 26124 19180 26180 19236
rect 25788 18450 25844 18452
rect 25788 18398 25790 18450
rect 25790 18398 25842 18450
rect 25842 18398 25844 18450
rect 25788 18396 25844 18398
rect 26236 19122 26292 19124
rect 26236 19070 26238 19122
rect 26238 19070 26290 19122
rect 26290 19070 26292 19122
rect 26236 19068 26292 19070
rect 26684 20076 26740 20132
rect 26572 19292 26628 19348
rect 26908 19234 26964 19236
rect 26908 19182 26910 19234
rect 26910 19182 26962 19234
rect 26962 19182 26964 19234
rect 26908 19180 26964 19182
rect 27580 19234 27636 19236
rect 27580 19182 27582 19234
rect 27582 19182 27634 19234
rect 27634 19182 27636 19234
rect 27580 19180 27636 19182
rect 26572 19010 26628 19012
rect 26572 18958 26574 19010
rect 26574 18958 26626 19010
rect 26626 18958 26628 19010
rect 26572 18956 26628 18958
rect 26012 18508 26068 18564
rect 27356 18732 27412 18788
rect 27916 18732 27972 18788
rect 26348 18396 26404 18452
rect 25900 18284 25956 18340
rect 26348 17276 26404 17332
rect 28476 18732 28532 18788
rect 28140 18396 28196 18452
rect 26796 17276 26852 17332
rect 29484 20578 29540 20580
rect 29484 20526 29486 20578
rect 29486 20526 29538 20578
rect 29538 20526 29540 20578
rect 29484 20524 29540 20526
rect 29708 20188 29764 20244
rect 29260 20076 29316 20132
rect 28700 18284 28756 18340
rect 34860 27074 34916 27076
rect 34860 27022 34862 27074
rect 34862 27022 34914 27074
rect 34914 27022 34916 27074
rect 34860 27020 34916 27022
rect 35532 27074 35588 27076
rect 35532 27022 35534 27074
rect 35534 27022 35586 27074
rect 35586 27022 35588 27074
rect 35532 27020 35588 27022
rect 34860 26348 34916 26404
rect 35532 26402 35588 26404
rect 35532 26350 35534 26402
rect 35534 26350 35586 26402
rect 35586 26350 35588 26402
rect 35532 26348 35588 26350
rect 35756 26348 35812 26404
rect 35196 26290 35252 26292
rect 35196 26238 35198 26290
rect 35198 26238 35250 26290
rect 35250 26238 35252 26290
rect 35196 26236 35252 26238
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 34748 25282 34804 25284
rect 34748 25230 34750 25282
rect 34750 25230 34802 25282
rect 34802 25230 34804 25282
rect 34748 25228 34804 25230
rect 35532 25228 35588 25284
rect 32620 24892 32676 24948
rect 30156 20076 30212 20132
rect 30156 19404 30212 19460
rect 29932 19234 29988 19236
rect 29932 19182 29934 19234
rect 29934 19182 29986 19234
rect 29986 19182 29988 19234
rect 29932 19180 29988 19182
rect 30492 19234 30548 19236
rect 30492 19182 30494 19234
rect 30494 19182 30546 19234
rect 30546 19182 30548 19234
rect 30492 19180 30548 19182
rect 29708 19122 29764 19124
rect 29708 19070 29710 19122
rect 29710 19070 29762 19122
rect 29762 19070 29764 19122
rect 29708 19068 29764 19070
rect 31276 20076 31332 20132
rect 31276 19180 31332 19236
rect 30604 19068 30660 19124
rect 29484 19010 29540 19012
rect 29484 18958 29486 19010
rect 29486 18958 29538 19010
rect 29538 18958 29540 19010
rect 29484 18956 29540 18958
rect 30716 19010 30772 19012
rect 30716 18958 30718 19010
rect 30718 18958 30770 19010
rect 30770 18958 30772 19010
rect 30716 18956 30772 18958
rect 31836 20300 31892 20356
rect 32284 20188 32340 20244
rect 31836 18844 31892 18900
rect 28700 17500 28756 17556
rect 28476 17442 28532 17444
rect 28476 17390 28478 17442
rect 28478 17390 28530 17442
rect 28530 17390 28532 17442
rect 28476 17388 28532 17390
rect 25900 16828 25956 16884
rect 26908 15820 26964 15876
rect 26796 14418 26852 14420
rect 26796 14366 26798 14418
rect 26798 14366 26850 14418
rect 26850 14366 26852 14418
rect 26796 14364 26852 14366
rect 26572 14306 26628 14308
rect 26572 14254 26574 14306
rect 26574 14254 26626 14306
rect 26626 14254 26628 14306
rect 26572 14252 26628 14254
rect 26572 13746 26628 13748
rect 26572 13694 26574 13746
rect 26574 13694 26626 13746
rect 26626 13694 26628 13746
rect 26572 13692 26628 13694
rect 26684 13522 26740 13524
rect 26684 13470 26686 13522
rect 26686 13470 26738 13522
rect 26738 13470 26740 13522
rect 26684 13468 26740 13470
rect 26124 13244 26180 13300
rect 25676 12908 25732 12964
rect 26572 13074 26628 13076
rect 26572 13022 26574 13074
rect 26574 13022 26626 13074
rect 26626 13022 26628 13074
rect 26572 13020 26628 13022
rect 24556 12236 24612 12292
rect 25452 12236 25508 12292
rect 24332 11788 24388 11844
rect 24108 11676 24164 11732
rect 25340 12066 25396 12068
rect 25340 12014 25342 12066
rect 25342 12014 25394 12066
rect 25394 12014 25396 12066
rect 25340 12012 25396 12014
rect 25228 11676 25284 11732
rect 25676 11676 25732 11732
rect 24892 11282 24948 11284
rect 24892 11230 24894 11282
rect 24894 11230 24946 11282
rect 24946 11230 24948 11282
rect 24892 11228 24948 11230
rect 24780 11170 24836 11172
rect 24780 11118 24782 11170
rect 24782 11118 24834 11170
rect 24834 11118 24836 11170
rect 24780 11116 24836 11118
rect 24220 10498 24276 10500
rect 24220 10446 24222 10498
rect 24222 10446 24274 10498
rect 24274 10446 24276 10498
rect 24220 10444 24276 10446
rect 22764 10332 22820 10388
rect 22764 9884 22820 9940
rect 23548 9714 23604 9716
rect 23548 9662 23550 9714
rect 23550 9662 23602 9714
rect 23602 9662 23604 9714
rect 23548 9660 23604 9662
rect 22540 8316 22596 8372
rect 22764 8988 22820 9044
rect 22204 7644 22260 7700
rect 21756 5906 21812 5908
rect 21756 5854 21758 5906
rect 21758 5854 21810 5906
rect 21810 5854 21812 5906
rect 21756 5852 21812 5854
rect 22540 7420 22596 7476
rect 22316 6076 22372 6132
rect 21980 5740 22036 5796
rect 21868 5404 21924 5460
rect 21868 4508 21924 4564
rect 21756 4450 21812 4452
rect 21756 4398 21758 4450
rect 21758 4398 21810 4450
rect 21810 4398 21812 4450
rect 21756 4396 21812 4398
rect 21756 4226 21812 4228
rect 21756 4174 21758 4226
rect 21758 4174 21810 4226
rect 21810 4174 21812 4226
rect 21756 4172 21812 4174
rect 21756 3948 21812 4004
rect 20860 2380 20916 2436
rect 21644 3388 21700 3444
rect 21308 1596 21364 1652
rect 22316 5292 22372 5348
rect 22540 6748 22596 6804
rect 23548 8988 23604 9044
rect 23100 8652 23156 8708
rect 23100 7698 23156 7700
rect 23100 7646 23102 7698
rect 23102 7646 23154 7698
rect 23154 7646 23156 7698
rect 23100 7644 23156 7646
rect 22652 5516 22708 5572
rect 23324 6748 23380 6804
rect 22988 6188 23044 6244
rect 23100 6412 23156 6468
rect 23772 7362 23828 7364
rect 23772 7310 23774 7362
rect 23774 7310 23826 7362
rect 23826 7310 23828 7362
rect 23772 7308 23828 7310
rect 23660 5628 23716 5684
rect 22988 5180 23044 5236
rect 22876 5122 22932 5124
rect 22876 5070 22878 5122
rect 22878 5070 22930 5122
rect 22930 5070 22932 5122
rect 22876 5068 22932 5070
rect 22428 4956 22484 5012
rect 22876 4508 22932 4564
rect 22428 3948 22484 4004
rect 22652 3442 22708 3444
rect 22652 3390 22654 3442
rect 22654 3390 22706 3442
rect 22706 3390 22708 3442
rect 22652 3388 22708 3390
rect 22316 3164 22372 3220
rect 22204 2940 22260 2996
rect 23100 4450 23156 4452
rect 23100 4398 23102 4450
rect 23102 4398 23154 4450
rect 23154 4398 23156 4450
rect 23100 4396 23156 4398
rect 22876 4284 22932 4340
rect 22988 4060 23044 4116
rect 22988 3724 23044 3780
rect 22764 1372 22820 1428
rect 23212 2828 23268 2884
rect 23548 5180 23604 5236
rect 23324 3164 23380 3220
rect 23324 2604 23380 2660
rect 23772 4620 23828 4676
rect 23996 6018 24052 6020
rect 23996 5966 23998 6018
rect 23998 5966 24050 6018
rect 24050 5966 24052 6018
rect 23996 5964 24052 5966
rect 23996 4450 24052 4452
rect 23996 4398 23998 4450
rect 23998 4398 24050 4450
rect 24050 4398 24052 4450
rect 23996 4396 24052 4398
rect 25004 10780 25060 10836
rect 24780 10610 24836 10612
rect 24780 10558 24782 10610
rect 24782 10558 24834 10610
rect 24834 10558 24836 10610
rect 24780 10556 24836 10558
rect 25228 10556 25284 10612
rect 24668 9996 24724 10052
rect 24668 9266 24724 9268
rect 24668 9214 24670 9266
rect 24670 9214 24722 9266
rect 24722 9214 24724 9266
rect 24668 9212 24724 9214
rect 25900 11452 25956 11508
rect 25788 10834 25844 10836
rect 25788 10782 25790 10834
rect 25790 10782 25842 10834
rect 25842 10782 25844 10834
rect 25788 10780 25844 10782
rect 26124 11282 26180 11284
rect 26124 11230 26126 11282
rect 26126 11230 26178 11282
rect 26178 11230 26180 11282
rect 26124 11228 26180 11230
rect 26236 10610 26292 10612
rect 26236 10558 26238 10610
rect 26238 10558 26290 10610
rect 26290 10558 26292 10610
rect 26236 10556 26292 10558
rect 26348 12124 26404 12180
rect 25340 9660 25396 9716
rect 26124 9660 26180 9716
rect 25676 9436 25732 9492
rect 25452 9212 25508 9268
rect 25004 8988 25060 9044
rect 24780 7698 24836 7700
rect 24780 7646 24782 7698
rect 24782 7646 24834 7698
rect 24834 7646 24836 7698
rect 24780 7644 24836 7646
rect 24444 6972 24500 7028
rect 24332 6860 24388 6916
rect 24332 6076 24388 6132
rect 24332 4060 24388 4116
rect 23436 2380 23492 2436
rect 24108 3052 24164 3108
rect 24668 5292 24724 5348
rect 25116 5628 25172 5684
rect 26684 11676 26740 11732
rect 27132 16828 27188 16884
rect 29596 17554 29652 17556
rect 29596 17502 29598 17554
rect 29598 17502 29650 17554
rect 29650 17502 29652 17554
rect 29596 17500 29652 17502
rect 29372 17052 29428 17108
rect 30156 16940 30212 16996
rect 27244 15820 27300 15876
rect 27356 15932 27412 15988
rect 28364 15932 28420 15988
rect 28140 15820 28196 15876
rect 27244 14306 27300 14308
rect 27244 14254 27246 14306
rect 27246 14254 27298 14306
rect 27298 14254 27300 14306
rect 27244 14252 27300 14254
rect 28252 14418 28308 14420
rect 28252 14366 28254 14418
rect 28254 14366 28306 14418
rect 28306 14366 28308 14418
rect 28252 14364 28308 14366
rect 27132 12796 27188 12852
rect 27356 13746 27412 13748
rect 27356 13694 27358 13746
rect 27358 13694 27410 13746
rect 27410 13694 27412 13746
rect 27356 13692 27412 13694
rect 27804 13746 27860 13748
rect 27804 13694 27806 13746
rect 27806 13694 27858 13746
rect 27858 13694 27860 13746
rect 27804 13692 27860 13694
rect 27916 12796 27972 12852
rect 27244 11788 27300 11844
rect 27468 11788 27524 11844
rect 26908 11116 26964 11172
rect 26908 10556 26964 10612
rect 31500 16044 31556 16100
rect 29596 15874 29652 15876
rect 29596 15822 29598 15874
rect 29598 15822 29650 15874
rect 29650 15822 29652 15874
rect 29596 15820 29652 15822
rect 29148 14418 29204 14420
rect 29148 14366 29150 14418
rect 29150 14366 29202 14418
rect 29202 14366 29204 14418
rect 29148 14364 29204 14366
rect 28588 14306 28644 14308
rect 28588 14254 28590 14306
rect 28590 14254 28642 14306
rect 28642 14254 28644 14306
rect 28588 14252 28644 14254
rect 29372 14140 29428 14196
rect 29484 14252 29540 14308
rect 29148 12850 29204 12852
rect 29148 12798 29150 12850
rect 29150 12798 29202 12850
rect 29202 12798 29204 12850
rect 29148 12796 29204 12798
rect 30156 14140 30212 14196
rect 30828 14140 30884 14196
rect 29596 13468 29652 13524
rect 31388 12684 31444 12740
rect 28252 12460 28308 12516
rect 31500 12236 31556 12292
rect 28252 11506 28308 11508
rect 28252 11454 28254 11506
rect 28254 11454 28306 11506
rect 28306 11454 28308 11506
rect 28252 11452 28308 11454
rect 28140 10668 28196 10724
rect 26572 9100 26628 9156
rect 25788 8034 25844 8036
rect 25788 7982 25790 8034
rect 25790 7982 25842 8034
rect 25842 7982 25844 8034
rect 25788 7980 25844 7982
rect 25788 7532 25844 7588
rect 25340 7474 25396 7476
rect 25340 7422 25342 7474
rect 25342 7422 25394 7474
rect 25394 7422 25396 7474
rect 25340 7420 25396 7422
rect 25340 6972 25396 7028
rect 25788 7362 25844 7364
rect 25788 7310 25790 7362
rect 25790 7310 25842 7362
rect 25842 7310 25844 7362
rect 25788 7308 25844 7310
rect 26236 7644 26292 7700
rect 26012 7532 26068 7588
rect 26348 6972 26404 7028
rect 26236 6802 26292 6804
rect 26236 6750 26238 6802
rect 26238 6750 26290 6802
rect 26290 6750 26292 6802
rect 26236 6748 26292 6750
rect 25900 6524 25956 6580
rect 25564 5852 25620 5908
rect 25788 5682 25844 5684
rect 25788 5630 25790 5682
rect 25790 5630 25842 5682
rect 25842 5630 25844 5682
rect 25788 5628 25844 5630
rect 25228 5068 25284 5124
rect 24780 3554 24836 3556
rect 24780 3502 24782 3554
rect 24782 3502 24834 3554
rect 24834 3502 24836 3554
rect 24780 3500 24836 3502
rect 25340 3500 25396 3556
rect 25788 5404 25844 5460
rect 26572 7586 26628 7588
rect 26572 7534 26574 7586
rect 26574 7534 26626 7586
rect 26626 7534 26628 7586
rect 26572 7532 26628 7534
rect 26908 8930 26964 8932
rect 26908 8878 26910 8930
rect 26910 8878 26962 8930
rect 26962 8878 26964 8930
rect 26908 8876 26964 8878
rect 26796 8428 26852 8484
rect 26908 8370 26964 8372
rect 26908 8318 26910 8370
rect 26910 8318 26962 8370
rect 26962 8318 26964 8370
rect 26908 8316 26964 8318
rect 27020 7644 27076 7700
rect 26796 6972 26852 7028
rect 26908 6748 26964 6804
rect 26348 6524 26404 6580
rect 26460 6300 26516 6356
rect 26348 6130 26404 6132
rect 26348 6078 26350 6130
rect 26350 6078 26402 6130
rect 26402 6078 26404 6130
rect 26348 6076 26404 6078
rect 26236 5628 26292 5684
rect 27020 6188 27076 6244
rect 26908 5740 26964 5796
rect 26684 5628 26740 5684
rect 26572 5404 26628 5460
rect 25452 4732 25508 4788
rect 25788 4284 25844 4340
rect 25676 3612 25732 3668
rect 24668 2716 24724 2772
rect 26012 4226 26068 4228
rect 26012 4174 26014 4226
rect 26014 4174 26066 4226
rect 26066 4174 26068 4226
rect 26012 4172 26068 4174
rect 26124 3724 26180 3780
rect 26124 3554 26180 3556
rect 26124 3502 26126 3554
rect 26126 3502 26178 3554
rect 26178 3502 26180 3554
rect 26124 3500 26180 3502
rect 26236 2828 26292 2884
rect 26348 4060 26404 4116
rect 26796 5404 26852 5460
rect 27580 8876 27636 8932
rect 27244 8652 27300 8708
rect 27356 8370 27412 8372
rect 27356 8318 27358 8370
rect 27358 8318 27410 8370
rect 27410 8318 27412 8370
rect 27356 8316 27412 8318
rect 27244 7756 27300 7812
rect 27468 7196 27524 7252
rect 27580 7084 27636 7140
rect 27804 7698 27860 7700
rect 27804 7646 27806 7698
rect 27806 7646 27858 7698
rect 27858 7646 27860 7698
rect 27804 7644 27860 7646
rect 27916 6860 27972 6916
rect 28028 10108 28084 10164
rect 27804 6748 27860 6804
rect 27132 6076 27188 6132
rect 27244 5794 27300 5796
rect 27244 5742 27246 5794
rect 27246 5742 27298 5794
rect 27298 5742 27300 5794
rect 27244 5740 27300 5742
rect 27132 5068 27188 5124
rect 27244 5404 27300 5460
rect 27132 4844 27188 4900
rect 26908 3612 26964 3668
rect 27020 3948 27076 4004
rect 27916 6690 27972 6692
rect 27916 6638 27918 6690
rect 27918 6638 27970 6690
rect 27970 6638 27972 6690
rect 27916 6636 27972 6638
rect 28252 8652 28308 8708
rect 28140 8482 28196 8484
rect 28140 8430 28142 8482
rect 28142 8430 28194 8482
rect 28194 8430 28196 8482
rect 28140 8428 28196 8430
rect 28140 7868 28196 7924
rect 31724 11900 31780 11956
rect 30044 11282 30100 11284
rect 30044 11230 30046 11282
rect 30046 11230 30098 11282
rect 30098 11230 30100 11282
rect 30044 11228 30100 11230
rect 31388 11282 31444 11284
rect 31388 11230 31390 11282
rect 31390 11230 31442 11282
rect 31442 11230 31444 11282
rect 31388 11228 31444 11230
rect 29484 10668 29540 10724
rect 28812 9772 28868 9828
rect 28476 7980 28532 8036
rect 28252 7532 28308 7588
rect 28140 7196 28196 7252
rect 28588 7420 28644 7476
rect 28700 8652 28756 8708
rect 28812 8316 28868 8372
rect 29036 9324 29092 9380
rect 29036 8930 29092 8932
rect 29036 8878 29038 8930
rect 29038 8878 29090 8930
rect 29090 8878 29092 8930
rect 29036 8876 29092 8878
rect 29036 8428 29092 8484
rect 28812 7644 28868 7700
rect 29036 7868 29092 7924
rect 28588 7196 28644 7252
rect 28140 6860 28196 6916
rect 28140 6524 28196 6580
rect 28252 6748 28308 6804
rect 28028 5516 28084 5572
rect 27804 5292 27860 5348
rect 27580 5180 27636 5236
rect 27916 5234 27972 5236
rect 27916 5182 27918 5234
rect 27918 5182 27970 5234
rect 27970 5182 27972 5234
rect 27916 5180 27972 5182
rect 28028 5068 28084 5124
rect 28588 6636 28644 6692
rect 28476 6524 28532 6580
rect 28700 6412 28756 6468
rect 28700 5180 28756 5236
rect 27692 3836 27748 3892
rect 27356 3276 27412 3332
rect 27580 2268 27636 2324
rect 28924 6972 28980 7028
rect 29260 8988 29316 9044
rect 29484 10444 29540 10500
rect 31276 11004 31332 11060
rect 30940 10780 30996 10836
rect 29820 10108 29876 10164
rect 30156 10556 30212 10612
rect 31948 18396 32004 18452
rect 32284 19010 32340 19012
rect 32284 18958 32286 19010
rect 32286 18958 32338 19010
rect 32338 18958 32340 19010
rect 32284 18956 32340 18958
rect 32508 17106 32564 17108
rect 32508 17054 32510 17106
rect 32510 17054 32562 17106
rect 32562 17054 32564 17106
rect 32508 17052 32564 17054
rect 32060 16994 32116 16996
rect 32060 16942 32062 16994
rect 32062 16942 32114 16994
rect 32114 16942 32116 16994
rect 32060 16940 32116 16942
rect 32172 16098 32228 16100
rect 32172 16046 32174 16098
rect 32174 16046 32226 16098
rect 32226 16046 32228 16098
rect 32172 16044 32228 16046
rect 34972 24722 35028 24724
rect 34972 24670 34974 24722
rect 34974 24670 35026 24722
rect 35026 24670 35028 24722
rect 34972 24668 35028 24670
rect 34076 24108 34132 24164
rect 35532 24834 35588 24836
rect 35532 24782 35534 24834
rect 35534 24782 35586 24834
rect 35586 24782 35588 24834
rect 35532 24780 35588 24782
rect 35308 24668 35364 24724
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 35756 24108 35812 24164
rect 34524 23938 34580 23940
rect 34524 23886 34526 23938
rect 34526 23886 34578 23938
rect 34578 23886 34580 23938
rect 34524 23884 34580 23886
rect 34076 23154 34132 23156
rect 34076 23102 34078 23154
rect 34078 23102 34130 23154
rect 34130 23102 34132 23154
rect 34076 23100 34132 23102
rect 33404 21532 33460 21588
rect 32956 20578 33012 20580
rect 32956 20526 32958 20578
rect 32958 20526 33010 20578
rect 33010 20526 33012 20578
rect 32956 20524 33012 20526
rect 33516 20076 33572 20132
rect 33404 19122 33460 19124
rect 33404 19070 33406 19122
rect 33406 19070 33458 19122
rect 33458 19070 33460 19122
rect 33404 19068 33460 19070
rect 34860 23548 34916 23604
rect 34860 23324 34916 23380
rect 34412 22482 34468 22484
rect 34412 22430 34414 22482
rect 34414 22430 34466 22482
rect 34466 22430 34468 22482
rect 34412 22428 34468 22430
rect 33964 22146 34020 22148
rect 33964 22094 33966 22146
rect 33966 22094 34018 22146
rect 34018 22094 34020 22146
rect 33964 22092 34020 22094
rect 33964 20860 34020 20916
rect 33740 20018 33796 20020
rect 33740 19966 33742 20018
rect 33742 19966 33794 20018
rect 33794 19966 33796 20018
rect 33740 19964 33796 19966
rect 34972 22988 35028 23044
rect 34860 22764 34916 22820
rect 35420 23714 35476 23716
rect 35420 23662 35422 23714
rect 35422 23662 35474 23714
rect 35474 23662 35476 23714
rect 35420 23660 35476 23662
rect 37100 29036 37156 29092
rect 36988 28082 37044 28084
rect 36988 28030 36990 28082
rect 36990 28030 37042 28082
rect 37042 28030 37044 28082
rect 36988 28028 37044 28030
rect 38668 76354 38724 76356
rect 38668 76302 38670 76354
rect 38670 76302 38722 76354
rect 38722 76302 38724 76354
rect 38668 76300 38724 76302
rect 38556 75852 38612 75908
rect 39004 75740 39060 75796
rect 38220 75682 38276 75684
rect 38220 75630 38222 75682
rect 38222 75630 38274 75682
rect 38274 75630 38276 75682
rect 38220 75628 38276 75630
rect 38892 75628 38948 75684
rect 41020 76690 41076 76692
rect 41020 76638 41022 76690
rect 41022 76638 41074 76690
rect 41074 76638 41076 76690
rect 41020 76636 41076 76638
rect 42028 76690 42084 76692
rect 42028 76638 42030 76690
rect 42030 76638 42082 76690
rect 42082 76638 42084 76690
rect 42028 76636 42084 76638
rect 43484 76972 43540 77028
rect 39788 74732 39844 74788
rect 40124 75628 40180 75684
rect 39788 28476 39844 28532
rect 38108 28028 38164 28084
rect 35980 25228 36036 25284
rect 35980 24780 36036 24836
rect 36316 26796 36372 26852
rect 35756 23100 35812 23156
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 35196 22316 35252 22372
rect 34972 21586 35028 21588
rect 34972 21534 34974 21586
rect 34974 21534 35026 21586
rect 35026 21534 35028 21586
rect 34972 21532 35028 21534
rect 34860 21474 34916 21476
rect 34860 21422 34862 21474
rect 34862 21422 34914 21474
rect 34914 21422 34916 21474
rect 34860 21420 34916 21422
rect 34748 21308 34804 21364
rect 35868 22258 35924 22260
rect 35868 22206 35870 22258
rect 35870 22206 35922 22258
rect 35922 22206 35924 22258
rect 35868 22204 35924 22206
rect 35756 22146 35812 22148
rect 35756 22094 35758 22146
rect 35758 22094 35810 22146
rect 35810 22094 35812 22146
rect 35756 22092 35812 22094
rect 36204 23324 36260 23380
rect 36428 26348 36484 26404
rect 38668 27580 38724 27636
rect 36988 26460 37044 26516
rect 36988 26124 37044 26180
rect 37212 26236 37268 26292
rect 36652 25452 36708 25508
rect 37212 25564 37268 25620
rect 37324 25788 37380 25844
rect 36652 25228 36708 25284
rect 36876 24946 36932 24948
rect 36876 24894 36878 24946
rect 36878 24894 36930 24946
rect 36930 24894 36932 24946
rect 36876 24892 36932 24894
rect 37212 24220 37268 24276
rect 36316 23212 36372 23268
rect 36652 23996 36708 24052
rect 36316 22988 36372 23044
rect 36316 22428 36372 22484
rect 35420 21586 35476 21588
rect 35420 21534 35422 21586
rect 35422 21534 35474 21586
rect 35474 21534 35476 21586
rect 35420 21532 35476 21534
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 34636 20690 34692 20692
rect 34636 20638 34638 20690
rect 34638 20638 34690 20690
rect 34690 20638 34692 20690
rect 34636 20636 34692 20638
rect 34860 20690 34916 20692
rect 34860 20638 34862 20690
rect 34862 20638 34914 20690
rect 34914 20638 34916 20690
rect 34860 20636 34916 20638
rect 34636 20300 34692 20356
rect 34188 19740 34244 19796
rect 34076 19628 34132 19684
rect 35084 20860 35140 20916
rect 35196 20748 35252 20804
rect 35532 20802 35588 20804
rect 35532 20750 35534 20802
rect 35534 20750 35586 20802
rect 35586 20750 35588 20802
rect 35532 20748 35588 20750
rect 35644 20636 35700 20692
rect 35756 20524 35812 20580
rect 34860 19628 34916 19684
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 35644 19404 35700 19460
rect 34972 19180 35028 19236
rect 33404 18732 33460 18788
rect 32732 18620 32788 18676
rect 33628 18450 33684 18452
rect 33628 18398 33630 18450
rect 33630 18398 33682 18450
rect 33682 18398 33684 18450
rect 33628 18396 33684 18398
rect 32956 17612 33012 17668
rect 32956 17276 33012 17332
rect 33852 18956 33908 19012
rect 34300 19068 34356 19124
rect 33852 17500 33908 17556
rect 35644 19234 35700 19236
rect 35644 19182 35646 19234
rect 35646 19182 35698 19234
rect 35698 19182 35700 19234
rect 35644 19180 35700 19182
rect 35308 19122 35364 19124
rect 35308 19070 35310 19122
rect 35310 19070 35362 19122
rect 35362 19070 35364 19122
rect 35308 19068 35364 19070
rect 35196 18284 35252 18340
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 35420 17724 35476 17780
rect 35308 17554 35364 17556
rect 35308 17502 35310 17554
rect 35310 17502 35362 17554
rect 35362 17502 35364 17554
rect 35308 17500 35364 17502
rect 35644 17724 35700 17780
rect 35980 21532 36036 21588
rect 35980 20748 36036 20804
rect 36092 20690 36148 20692
rect 36092 20638 36094 20690
rect 36094 20638 36146 20690
rect 36146 20638 36148 20690
rect 36092 20636 36148 20638
rect 36316 21308 36372 21364
rect 36540 21532 36596 21588
rect 36428 20860 36484 20916
rect 36540 20300 36596 20356
rect 37212 23884 37268 23940
rect 36988 23436 37044 23492
rect 36764 23212 36820 23268
rect 36988 22652 37044 22708
rect 36876 22204 36932 22260
rect 36652 19404 36708 19460
rect 35868 19122 35924 19124
rect 35868 19070 35870 19122
rect 35870 19070 35922 19122
rect 35922 19070 35924 19122
rect 35868 19068 35924 19070
rect 35420 17276 35476 17332
rect 34524 17052 34580 17108
rect 33516 16882 33572 16884
rect 33516 16830 33518 16882
rect 33518 16830 33570 16882
rect 33570 16830 33572 16882
rect 33516 16828 33572 16830
rect 33516 16156 33572 16212
rect 32508 15202 32564 15204
rect 32508 15150 32510 15202
rect 32510 15150 32562 15202
rect 32562 15150 32564 15202
rect 32508 15148 32564 15150
rect 31948 14476 32004 14532
rect 32060 14418 32116 14420
rect 32060 14366 32062 14418
rect 32062 14366 32114 14418
rect 32114 14366 32116 14418
rect 32060 14364 32116 14366
rect 33180 12962 33236 12964
rect 33180 12910 33182 12962
rect 33182 12910 33234 12962
rect 33234 12910 33236 12962
rect 33180 12908 33236 12910
rect 32060 12236 32116 12292
rect 31836 11452 31892 11508
rect 31500 10834 31556 10836
rect 31500 10782 31502 10834
rect 31502 10782 31554 10834
rect 31554 10782 31556 10834
rect 31500 10780 31556 10782
rect 32396 11394 32452 11396
rect 32396 11342 32398 11394
rect 32398 11342 32450 11394
rect 32450 11342 32452 11394
rect 32396 11340 32452 11342
rect 31948 11228 32004 11284
rect 30156 9884 30212 9940
rect 29484 8764 29540 8820
rect 29260 8204 29316 8260
rect 29260 7420 29316 7476
rect 29484 7644 29540 7700
rect 29596 6860 29652 6916
rect 29260 6748 29316 6804
rect 29036 6300 29092 6356
rect 29036 5964 29092 6020
rect 28924 5180 28980 5236
rect 29260 5906 29316 5908
rect 29260 5854 29262 5906
rect 29262 5854 29314 5906
rect 29314 5854 29316 5906
rect 29260 5852 29316 5854
rect 29820 8204 29876 8260
rect 32620 11282 32676 11284
rect 32620 11230 32622 11282
rect 32622 11230 32674 11282
rect 32674 11230 32676 11282
rect 32620 11228 32676 11230
rect 32172 11004 32228 11060
rect 31388 10498 31444 10500
rect 31388 10446 31390 10498
rect 31390 10446 31442 10498
rect 31442 10446 31444 10498
rect 31388 10444 31444 10446
rect 31836 9996 31892 10052
rect 30380 8428 30436 8484
rect 30044 7868 30100 7924
rect 30044 7698 30100 7700
rect 30044 7646 30046 7698
rect 30046 7646 30098 7698
rect 30098 7646 30100 7698
rect 30044 7644 30100 7646
rect 30380 7586 30436 7588
rect 30380 7534 30382 7586
rect 30382 7534 30434 7586
rect 30434 7534 30436 7586
rect 30380 7532 30436 7534
rect 30044 6860 30100 6916
rect 30156 6524 30212 6580
rect 30268 6748 30324 6804
rect 30044 6412 30100 6468
rect 30604 7084 30660 7140
rect 31724 9660 31780 9716
rect 31276 9324 31332 9380
rect 31276 8204 31332 8260
rect 30940 7308 30996 7364
rect 30828 6860 30884 6916
rect 32508 11116 32564 11172
rect 32284 9660 32340 9716
rect 32396 9212 32452 9268
rect 33068 12124 33124 12180
rect 33404 15426 33460 15428
rect 33404 15374 33406 15426
rect 33406 15374 33458 15426
rect 33458 15374 33460 15426
rect 33404 15372 33460 15374
rect 33404 14364 33460 14420
rect 33404 13970 33460 13972
rect 33404 13918 33406 13970
rect 33406 13918 33458 13970
rect 33458 13918 33460 13970
rect 33404 13916 33460 13918
rect 33628 13804 33684 13860
rect 34076 15596 34132 15652
rect 34748 16882 34804 16884
rect 34748 16830 34750 16882
rect 34750 16830 34802 16882
rect 34802 16830 34804 16882
rect 34748 16828 34804 16830
rect 34636 16716 34692 16772
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 34636 15932 34692 15988
rect 33852 15148 33908 15204
rect 34076 14476 34132 14532
rect 34412 14252 34468 14308
rect 34188 13970 34244 13972
rect 34188 13918 34190 13970
rect 34190 13918 34242 13970
rect 34242 13918 34244 13970
rect 34188 13916 34244 13918
rect 34972 15708 35028 15764
rect 34636 14028 34692 14084
rect 34860 15036 34916 15092
rect 34860 13916 34916 13972
rect 34748 13858 34804 13860
rect 34748 13806 34750 13858
rect 34750 13806 34802 13858
rect 34802 13806 34804 13858
rect 34748 13804 34804 13806
rect 34412 13692 34468 13748
rect 33292 11564 33348 11620
rect 33180 10892 33236 10948
rect 33852 12962 33908 12964
rect 33852 12910 33854 12962
rect 33854 12910 33906 12962
rect 33906 12910 33908 12962
rect 33852 12908 33908 12910
rect 34412 12962 34468 12964
rect 34412 12910 34414 12962
rect 34414 12910 34466 12962
rect 34466 12910 34468 12962
rect 34412 12908 34468 12910
rect 34748 12962 34804 12964
rect 34748 12910 34750 12962
rect 34750 12910 34802 12962
rect 34802 12910 34804 12962
rect 34748 12908 34804 12910
rect 33964 12460 34020 12516
rect 33964 12012 34020 12068
rect 33852 11788 33908 11844
rect 33740 11004 33796 11060
rect 33852 10892 33908 10948
rect 33292 10722 33348 10724
rect 33292 10670 33294 10722
rect 33294 10670 33346 10722
rect 33346 10670 33348 10722
rect 33292 10668 33348 10670
rect 33740 9714 33796 9716
rect 33740 9662 33742 9714
rect 33742 9662 33794 9714
rect 33794 9662 33796 9714
rect 33740 9660 33796 9662
rect 33292 9602 33348 9604
rect 33292 9550 33294 9602
rect 33294 9550 33346 9602
rect 33346 9550 33348 9602
rect 33292 9548 33348 9550
rect 32844 9212 32900 9268
rect 32732 8876 32788 8932
rect 32844 8092 32900 8148
rect 31836 7756 31892 7812
rect 31500 6972 31556 7028
rect 31500 6802 31556 6804
rect 31500 6750 31502 6802
rect 31502 6750 31554 6802
rect 31554 6750 31556 6802
rect 31500 6748 31556 6750
rect 30828 6690 30884 6692
rect 30828 6638 30830 6690
rect 30830 6638 30882 6690
rect 30882 6638 30884 6690
rect 30828 6636 30884 6638
rect 29260 5404 29316 5460
rect 29932 6076 29988 6132
rect 28812 4956 28868 5012
rect 28812 4450 28868 4452
rect 28812 4398 28814 4450
rect 28814 4398 28866 4450
rect 28866 4398 28868 4450
rect 28812 4396 28868 4398
rect 28588 3836 28644 3892
rect 28476 3500 28532 3556
rect 27804 2940 27860 2996
rect 28700 3388 28756 3444
rect 29596 5234 29652 5236
rect 29596 5182 29598 5234
rect 29598 5182 29650 5234
rect 29650 5182 29652 5234
rect 29596 5180 29652 5182
rect 30044 5852 30100 5908
rect 29484 5122 29540 5124
rect 29484 5070 29486 5122
rect 29486 5070 29538 5122
rect 29538 5070 29540 5122
rect 29484 5068 29540 5070
rect 28924 3052 28980 3108
rect 29932 5010 29988 5012
rect 29932 4958 29934 5010
rect 29934 4958 29986 5010
rect 29986 4958 29988 5010
rect 29932 4956 29988 4958
rect 29820 4620 29876 4676
rect 29148 2604 29204 2660
rect 29260 1820 29316 1876
rect 30604 6188 30660 6244
rect 30828 5852 30884 5908
rect 30268 5010 30324 5012
rect 30268 4958 30270 5010
rect 30270 4958 30322 5010
rect 30322 4958 30324 5010
rect 30268 4956 30324 4958
rect 30044 4396 30100 4452
rect 30268 4620 30324 4676
rect 29932 4060 29988 4116
rect 30268 4172 30324 4228
rect 30940 5740 30996 5796
rect 30604 5122 30660 5124
rect 30604 5070 30606 5122
rect 30606 5070 30658 5122
rect 30658 5070 30660 5122
rect 30604 5068 30660 5070
rect 30716 4732 30772 4788
rect 31164 6578 31220 6580
rect 31164 6526 31166 6578
rect 31166 6526 31218 6578
rect 31218 6526 31220 6578
rect 31164 6524 31220 6526
rect 31164 6300 31220 6356
rect 31388 5180 31444 5236
rect 30828 4338 30884 4340
rect 30828 4286 30830 4338
rect 30830 4286 30882 4338
rect 30882 4286 30884 4338
rect 30828 4284 30884 4286
rect 31612 5292 31668 5348
rect 32172 6860 32228 6916
rect 31836 6802 31892 6804
rect 31836 6750 31838 6802
rect 31838 6750 31890 6802
rect 31890 6750 31892 6802
rect 31836 6748 31892 6750
rect 32732 6802 32788 6804
rect 32732 6750 32734 6802
rect 32734 6750 32786 6802
rect 32786 6750 32788 6802
rect 32732 6748 32788 6750
rect 32620 6690 32676 6692
rect 32620 6638 32622 6690
rect 32622 6638 32674 6690
rect 32674 6638 32676 6690
rect 32620 6636 32676 6638
rect 34076 9212 34132 9268
rect 36428 19234 36484 19236
rect 36428 19182 36430 19234
rect 36430 19182 36482 19234
rect 36482 19182 36484 19234
rect 36428 19180 36484 19182
rect 36316 18844 36372 18900
rect 36092 17724 36148 17780
rect 36540 18172 36596 18228
rect 37660 25676 37716 25732
rect 37772 25506 37828 25508
rect 37772 25454 37774 25506
rect 37774 25454 37826 25506
rect 37826 25454 37828 25506
rect 37772 25452 37828 25454
rect 37772 25228 37828 25284
rect 37324 23154 37380 23156
rect 37324 23102 37326 23154
rect 37326 23102 37378 23154
rect 37378 23102 37380 23154
rect 37324 23100 37380 23102
rect 37212 22092 37268 22148
rect 37324 22876 37380 22932
rect 37212 21868 37268 21924
rect 38220 26348 38276 26404
rect 38332 25506 38388 25508
rect 38332 25454 38334 25506
rect 38334 25454 38386 25506
rect 38386 25454 38388 25506
rect 38332 25452 38388 25454
rect 38220 25282 38276 25284
rect 38220 25230 38222 25282
rect 38222 25230 38274 25282
rect 38274 25230 38276 25282
rect 38220 25228 38276 25230
rect 37884 24556 37940 24612
rect 37772 24444 37828 24500
rect 37660 23996 37716 24052
rect 37772 23660 37828 23716
rect 38780 26236 38836 26292
rect 38780 25452 38836 25508
rect 38668 25228 38724 25284
rect 39340 28082 39396 28084
rect 39340 28030 39342 28082
rect 39342 28030 39394 28082
rect 39394 28030 39396 28082
rect 39340 28028 39396 28030
rect 39116 26402 39172 26404
rect 39116 26350 39118 26402
rect 39118 26350 39170 26402
rect 39170 26350 39172 26402
rect 39116 26348 39172 26350
rect 37884 22876 37940 22932
rect 37436 22316 37492 22372
rect 37548 22652 37604 22708
rect 37548 21868 37604 21924
rect 37660 21756 37716 21812
rect 37436 20860 37492 20916
rect 37100 20524 37156 20580
rect 37100 19628 37156 19684
rect 37100 19292 37156 19348
rect 37436 20300 37492 20356
rect 37100 19122 37156 19124
rect 37100 19070 37102 19122
rect 37102 19070 37154 19122
rect 37154 19070 37156 19122
rect 37100 19068 37156 19070
rect 37772 20748 37828 20804
rect 38108 21980 38164 22036
rect 38108 20860 38164 20916
rect 37884 19964 37940 20020
rect 37772 19404 37828 19460
rect 37212 17724 37268 17780
rect 37660 19068 37716 19124
rect 37100 17276 37156 17332
rect 37100 16940 37156 16996
rect 37212 17164 37268 17220
rect 36988 16828 37044 16884
rect 36540 16716 36596 16772
rect 36092 16268 36148 16324
rect 36988 16268 37044 16324
rect 35644 15708 35700 15764
rect 35420 15372 35476 15428
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 37996 19628 38052 19684
rect 37884 19292 37940 19348
rect 37996 19234 38052 19236
rect 37996 19182 37998 19234
rect 37998 19182 38050 19234
rect 38050 19182 38052 19234
rect 37996 19180 38052 19182
rect 38332 22370 38388 22372
rect 38332 22318 38334 22370
rect 38334 22318 38386 22370
rect 38386 22318 38388 22370
rect 38332 22316 38388 22318
rect 38668 23212 38724 23268
rect 39228 22876 39284 22932
rect 39116 21586 39172 21588
rect 39116 21534 39118 21586
rect 39118 21534 39170 21586
rect 39170 21534 39172 21586
rect 39116 21532 39172 21534
rect 39228 21196 39284 21252
rect 38892 20860 38948 20916
rect 38332 19292 38388 19348
rect 38892 20524 38948 20580
rect 38780 20300 38836 20356
rect 38668 19068 38724 19124
rect 38220 18338 38276 18340
rect 38220 18286 38222 18338
rect 38222 18286 38274 18338
rect 38274 18286 38276 18338
rect 38220 18284 38276 18286
rect 37436 16716 37492 16772
rect 37772 16828 37828 16884
rect 38556 18396 38612 18452
rect 38108 16604 38164 16660
rect 37996 16322 38052 16324
rect 37996 16270 37998 16322
rect 37998 16270 38050 16322
rect 38050 16270 38052 16322
rect 37996 16268 38052 16270
rect 35420 14530 35476 14532
rect 35420 14478 35422 14530
rect 35422 14478 35474 14530
rect 35474 14478 35476 14530
rect 35420 14476 35476 14478
rect 35868 14530 35924 14532
rect 35868 14478 35870 14530
rect 35870 14478 35922 14530
rect 35922 14478 35924 14530
rect 35868 14476 35924 14478
rect 36092 13804 36148 13860
rect 35756 13468 35812 13524
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35084 13132 35140 13188
rect 35420 12962 35476 12964
rect 35420 12910 35422 12962
rect 35422 12910 35474 12962
rect 35474 12910 35476 12962
rect 35420 12908 35476 12910
rect 36204 12908 36260 12964
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 36988 12290 37044 12292
rect 36988 12238 36990 12290
rect 36990 12238 37042 12290
rect 37042 12238 37044 12290
rect 36988 12236 37044 12238
rect 36876 12178 36932 12180
rect 36876 12126 36878 12178
rect 36878 12126 36930 12178
rect 36930 12126 36932 12178
rect 36876 12124 36932 12126
rect 37884 15986 37940 15988
rect 37884 15934 37886 15986
rect 37886 15934 37938 15986
rect 37938 15934 37940 15986
rect 37884 15932 37940 15934
rect 37436 14476 37492 14532
rect 38668 16882 38724 16884
rect 38668 16830 38670 16882
rect 38670 16830 38722 16882
rect 38722 16830 38724 16882
rect 38668 16828 38724 16830
rect 39452 20802 39508 20804
rect 39452 20750 39454 20802
rect 39454 20750 39506 20802
rect 39506 20750 39508 20802
rect 39452 20748 39508 20750
rect 39340 20300 39396 20356
rect 39228 19516 39284 19572
rect 39228 19292 39284 19348
rect 39116 19234 39172 19236
rect 39116 19182 39118 19234
rect 39118 19182 39170 19234
rect 39170 19182 39172 19234
rect 39116 19180 39172 19182
rect 39116 19010 39172 19012
rect 39116 18958 39118 19010
rect 39118 18958 39170 19010
rect 39170 18958 39172 19010
rect 39116 18956 39172 18958
rect 38892 17164 38948 17220
rect 39116 18508 39172 18564
rect 39676 25282 39732 25284
rect 39676 25230 39678 25282
rect 39678 25230 39730 25282
rect 39730 25230 39732 25282
rect 39676 25228 39732 25230
rect 39676 24556 39732 24612
rect 39676 23266 39732 23268
rect 39676 23214 39678 23266
rect 39678 23214 39730 23266
rect 39730 23214 39732 23266
rect 39676 23212 39732 23214
rect 40012 26962 40068 26964
rect 40012 26910 40014 26962
rect 40014 26910 40066 26962
rect 40066 26910 40068 26962
rect 40012 26908 40068 26910
rect 40012 26290 40068 26292
rect 40012 26238 40014 26290
rect 40014 26238 40066 26290
rect 40066 26238 40068 26290
rect 40012 26236 40068 26238
rect 40908 75682 40964 75684
rect 40908 75630 40910 75682
rect 40910 75630 40962 75682
rect 40962 75630 40964 75682
rect 40908 75628 40964 75630
rect 41244 38946 41300 38948
rect 41244 38894 41246 38946
rect 41246 38894 41298 38946
rect 41298 38894 41300 38946
rect 41244 38892 41300 38894
rect 41580 38834 41636 38836
rect 41580 38782 41582 38834
rect 41582 38782 41634 38834
rect 41634 38782 41636 38834
rect 41580 38780 41636 38782
rect 41468 38668 41524 38724
rect 40684 28476 40740 28532
rect 40236 27916 40292 27972
rect 40348 27858 40404 27860
rect 40348 27806 40350 27858
rect 40350 27806 40402 27858
rect 40402 27806 40404 27858
rect 40348 27804 40404 27806
rect 40460 25564 40516 25620
rect 40348 24834 40404 24836
rect 40348 24782 40350 24834
rect 40350 24782 40402 24834
rect 40402 24782 40404 24834
rect 40348 24780 40404 24782
rect 40124 24332 40180 24388
rect 40012 22988 40068 23044
rect 39676 20018 39732 20020
rect 39676 19966 39678 20018
rect 39678 19966 39730 20018
rect 39730 19966 39732 20018
rect 39676 19964 39732 19966
rect 39564 19180 39620 19236
rect 39340 19068 39396 19124
rect 40348 23938 40404 23940
rect 40348 23886 40350 23938
rect 40350 23886 40402 23938
rect 40402 23886 40404 23938
rect 40348 23884 40404 23886
rect 40236 23772 40292 23828
rect 40460 23212 40516 23268
rect 40348 22652 40404 22708
rect 39900 20578 39956 20580
rect 39900 20526 39902 20578
rect 39902 20526 39954 20578
rect 39954 20526 39956 20578
rect 39900 20524 39956 20526
rect 40012 19404 40068 19460
rect 39340 18450 39396 18452
rect 39340 18398 39342 18450
rect 39342 18398 39394 18450
rect 39394 18398 39396 18450
rect 39340 18396 39396 18398
rect 40012 18844 40068 18900
rect 39900 18508 39956 18564
rect 39676 18396 39732 18452
rect 39452 18172 39508 18228
rect 39116 18060 39172 18116
rect 39116 17778 39172 17780
rect 39116 17726 39118 17778
rect 39118 17726 39170 17778
rect 39170 17726 39172 17778
rect 39116 17724 39172 17726
rect 39340 17666 39396 17668
rect 39340 17614 39342 17666
rect 39342 17614 39394 17666
rect 39394 17614 39396 17666
rect 39340 17612 39396 17614
rect 39564 17388 39620 17444
rect 42028 39058 42084 39060
rect 42028 39006 42030 39058
rect 42030 39006 42082 39058
rect 42082 39006 42084 39058
rect 42028 39004 42084 39006
rect 41692 28028 41748 28084
rect 41804 38780 41860 38836
rect 41356 27916 41412 27972
rect 41468 27858 41524 27860
rect 41468 27806 41470 27858
rect 41470 27806 41522 27858
rect 41522 27806 41524 27858
rect 41468 27804 41524 27806
rect 41692 26908 41748 26964
rect 41020 25452 41076 25508
rect 40684 20412 40740 20468
rect 40572 20076 40628 20132
rect 41356 26460 41412 26516
rect 41356 25506 41412 25508
rect 41356 25454 41358 25506
rect 41358 25454 41410 25506
rect 41410 25454 41412 25506
rect 41356 25452 41412 25454
rect 41244 24834 41300 24836
rect 41244 24782 41246 24834
rect 41246 24782 41298 24834
rect 41298 24782 41300 24834
rect 41244 24780 41300 24782
rect 41356 21586 41412 21588
rect 41356 21534 41358 21586
rect 41358 21534 41410 21586
rect 41410 21534 41412 21586
rect 41356 21532 41412 21534
rect 41356 20860 41412 20916
rect 40908 20130 40964 20132
rect 40908 20078 40910 20130
rect 40910 20078 40962 20130
rect 40962 20078 40964 20130
rect 40908 20076 40964 20078
rect 40236 19964 40292 20020
rect 41132 20018 41188 20020
rect 41132 19966 41134 20018
rect 41134 19966 41186 20018
rect 41186 19966 41188 20018
rect 41132 19964 41188 19966
rect 40572 19628 40628 19684
rect 40460 19122 40516 19124
rect 40460 19070 40462 19122
rect 40462 19070 40514 19122
rect 40514 19070 40516 19122
rect 40460 19068 40516 19070
rect 40124 17948 40180 18004
rect 40460 18844 40516 18900
rect 41132 19628 41188 19684
rect 40796 19404 40852 19460
rect 41020 19234 41076 19236
rect 41020 19182 41022 19234
rect 41022 19182 41074 19234
rect 41074 19182 41076 19234
rect 41020 19180 41076 19182
rect 40572 18284 40628 18340
rect 40012 17666 40068 17668
rect 40012 17614 40014 17666
rect 40014 17614 40066 17666
rect 40066 17614 40068 17666
rect 40012 17612 40068 17614
rect 40348 17612 40404 17668
rect 38892 16940 38948 16996
rect 39900 16994 39956 16996
rect 39900 16942 39902 16994
rect 39902 16942 39954 16994
rect 39954 16942 39956 16994
rect 39900 16940 39956 16942
rect 40124 16882 40180 16884
rect 40124 16830 40126 16882
rect 40126 16830 40178 16882
rect 40178 16830 40180 16882
rect 40124 16828 40180 16830
rect 39788 16716 39844 16772
rect 39676 16210 39732 16212
rect 39676 16158 39678 16210
rect 39678 16158 39730 16210
rect 39730 16158 39732 16210
rect 39676 16156 39732 16158
rect 40684 17666 40740 17668
rect 40684 17614 40686 17666
rect 40686 17614 40738 17666
rect 40738 17614 40740 17666
rect 40684 17612 40740 17614
rect 41020 17612 41076 17668
rect 41244 19404 41300 19460
rect 41356 19068 41412 19124
rect 41244 18450 41300 18452
rect 41244 18398 41246 18450
rect 41246 18398 41298 18450
rect 41298 18398 41300 18450
rect 41244 18396 41300 18398
rect 41244 18172 41300 18228
rect 41692 26236 41748 26292
rect 41692 24610 41748 24612
rect 41692 24558 41694 24610
rect 41694 24558 41746 24610
rect 41746 24558 41748 24610
rect 41692 24556 41748 24558
rect 41916 28028 41972 28084
rect 43932 76972 43988 77028
rect 44156 76636 44212 76692
rect 44492 76972 44548 77028
rect 42140 27132 42196 27188
rect 43820 75628 43876 75684
rect 43596 41804 43652 41860
rect 43148 40572 43204 40628
rect 42588 40348 42644 40404
rect 43036 38946 43092 38948
rect 43036 38894 43038 38946
rect 43038 38894 43090 38946
rect 43090 38894 43092 38946
rect 43036 38892 43092 38894
rect 42924 38834 42980 38836
rect 42924 38782 42926 38834
rect 42926 38782 42978 38834
rect 42978 38782 42980 38834
rect 42924 38780 42980 38782
rect 42588 28476 42644 28532
rect 42476 28082 42532 28084
rect 42476 28030 42478 28082
rect 42478 28030 42530 28082
rect 42530 28030 42532 28082
rect 42476 28028 42532 28030
rect 42028 26236 42084 26292
rect 42476 27580 42532 27636
rect 41916 25676 41972 25732
rect 42028 25564 42084 25620
rect 42364 26514 42420 26516
rect 42364 26462 42366 26514
rect 42366 26462 42418 26514
rect 42418 26462 42420 26514
rect 42364 26460 42420 26462
rect 42252 25228 42308 25284
rect 43036 27186 43092 27188
rect 43036 27134 43038 27186
rect 43038 27134 43090 27186
rect 43090 27134 43092 27186
rect 43036 27132 43092 27134
rect 42924 26290 42980 26292
rect 42924 26238 42926 26290
rect 42926 26238 42978 26290
rect 42978 26238 42980 26290
rect 42924 26236 42980 26238
rect 43036 25676 43092 25732
rect 42812 25228 42868 25284
rect 42140 21362 42196 21364
rect 42140 21310 42142 21362
rect 42142 21310 42194 21362
rect 42194 21310 42196 21362
rect 42140 21308 42196 21310
rect 42700 24332 42756 24388
rect 42476 22370 42532 22372
rect 42476 22318 42478 22370
rect 42478 22318 42530 22370
rect 42530 22318 42532 22370
rect 42476 22316 42532 22318
rect 42476 21586 42532 21588
rect 42476 21534 42478 21586
rect 42478 21534 42530 21586
rect 42530 21534 42532 21586
rect 42476 21532 42532 21534
rect 42364 21084 42420 21140
rect 41580 19404 41636 19460
rect 41580 18844 41636 18900
rect 41356 17388 41412 17444
rect 41804 18956 41860 19012
rect 41916 18396 41972 18452
rect 42140 19068 42196 19124
rect 41916 18226 41972 18228
rect 41916 18174 41918 18226
rect 41918 18174 41970 18226
rect 41970 18174 41972 18226
rect 41916 18172 41972 18174
rect 41468 16828 41524 16884
rect 41916 16828 41972 16884
rect 38892 15484 38948 15540
rect 39452 15538 39508 15540
rect 39452 15486 39454 15538
rect 39454 15486 39506 15538
rect 39506 15486 39508 15538
rect 39452 15484 39508 15486
rect 38556 14812 38612 14868
rect 39228 15148 39284 15204
rect 37212 14364 37268 14420
rect 38444 14252 38500 14308
rect 37660 13916 37716 13972
rect 37436 13132 37492 13188
rect 36988 12012 37044 12068
rect 35980 11340 36036 11396
rect 37212 11676 37268 11732
rect 37324 12124 37380 12180
rect 36428 11170 36484 11172
rect 36428 11118 36430 11170
rect 36430 11118 36482 11170
rect 36482 11118 36484 11170
rect 36428 11116 36484 11118
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 34860 9938 34916 9940
rect 34860 9886 34862 9938
rect 34862 9886 34914 9938
rect 34914 9886 34916 9938
rect 34860 9884 34916 9886
rect 36876 9772 36932 9828
rect 34524 9100 34580 9156
rect 33516 8930 33572 8932
rect 33516 8878 33518 8930
rect 33518 8878 33570 8930
rect 33570 8878 33572 8930
rect 33516 8876 33572 8878
rect 34300 8764 34356 8820
rect 33292 7980 33348 8036
rect 32172 5852 32228 5908
rect 31724 5180 31780 5236
rect 31836 5292 31892 5348
rect 30604 3164 30660 3220
rect 30604 2156 30660 2212
rect 30940 3330 30996 3332
rect 30940 3278 30942 3330
rect 30942 3278 30994 3330
rect 30994 3278 30996 3330
rect 30940 3276 30996 3278
rect 31836 3724 31892 3780
rect 31500 1708 31556 1764
rect 31612 1484 31668 1540
rect 32284 5122 32340 5124
rect 32284 5070 32286 5122
rect 32286 5070 32338 5122
rect 32338 5070 32340 5122
rect 32284 5068 32340 5070
rect 33068 7308 33124 7364
rect 33068 7084 33124 7140
rect 32620 5628 32676 5684
rect 33292 6748 33348 6804
rect 33964 7698 34020 7700
rect 33964 7646 33966 7698
rect 33966 7646 34018 7698
rect 34018 7646 34020 7698
rect 33964 7644 34020 7646
rect 33852 7586 33908 7588
rect 33852 7534 33854 7586
rect 33854 7534 33906 7586
rect 33906 7534 33908 7586
rect 33852 7532 33908 7534
rect 33740 7420 33796 7476
rect 34748 8930 34804 8932
rect 34748 8878 34750 8930
rect 34750 8878 34802 8930
rect 34802 8878 34804 8930
rect 34748 8876 34804 8878
rect 37884 13692 37940 13748
rect 38444 13522 38500 13524
rect 38444 13470 38446 13522
rect 38446 13470 38498 13522
rect 38498 13470 38500 13522
rect 38444 13468 38500 13470
rect 37996 12460 38052 12516
rect 37436 11900 37492 11956
rect 38220 11340 38276 11396
rect 39004 13746 39060 13748
rect 39004 13694 39006 13746
rect 39006 13694 39058 13746
rect 39058 13694 39060 13746
rect 39004 13692 39060 13694
rect 39340 14028 39396 14084
rect 39676 13916 39732 13972
rect 39228 13132 39284 13188
rect 40124 15820 40180 15876
rect 40236 13970 40292 13972
rect 40236 13918 40238 13970
rect 40238 13918 40290 13970
rect 40290 13918 40292 13970
rect 40236 13916 40292 13918
rect 40012 13858 40068 13860
rect 40012 13806 40014 13858
rect 40014 13806 40066 13858
rect 40066 13806 40068 13858
rect 40012 13804 40068 13806
rect 39788 13468 39844 13524
rect 40796 13468 40852 13524
rect 39564 12460 39620 12516
rect 39228 12012 39284 12068
rect 40684 12124 40740 12180
rect 40908 12460 40964 12516
rect 41468 16210 41524 16212
rect 41468 16158 41470 16210
rect 41470 16158 41522 16210
rect 41522 16158 41524 16210
rect 41468 16156 41524 16158
rect 41244 16044 41300 16100
rect 43596 40348 43652 40404
rect 43260 39340 43316 39396
rect 45388 76690 45444 76692
rect 45388 76638 45390 76690
rect 45390 76638 45442 76690
rect 45442 76638 45444 76690
rect 45388 76636 45444 76638
rect 45836 76636 45892 76692
rect 46172 76636 46228 76692
rect 47404 76690 47460 76692
rect 47404 76638 47406 76690
rect 47406 76638 47458 76690
rect 47458 76638 47460 76690
rect 47404 76636 47460 76638
rect 47852 76636 47908 76692
rect 46844 75852 46900 75908
rect 47852 76354 47908 76356
rect 47852 76302 47854 76354
rect 47854 76302 47906 76354
rect 47906 76302 47908 76354
rect 47852 76300 47908 76302
rect 48188 76636 48244 76692
rect 48412 75852 48468 75908
rect 43820 27356 43876 27412
rect 43484 25676 43540 25732
rect 43708 25564 43764 25620
rect 43372 25506 43428 25508
rect 43372 25454 43374 25506
rect 43374 25454 43426 25506
rect 43426 25454 43428 25506
rect 43372 25452 43428 25454
rect 43036 21532 43092 21588
rect 42812 21420 42868 21476
rect 42924 21308 42980 21364
rect 43260 21698 43316 21700
rect 43260 21646 43262 21698
rect 43262 21646 43314 21698
rect 43314 21646 43316 21698
rect 43260 21644 43316 21646
rect 43260 21084 43316 21140
rect 43148 20412 43204 20468
rect 42588 18396 42644 18452
rect 42364 16492 42420 16548
rect 42700 16940 42756 16996
rect 44044 38834 44100 38836
rect 44044 38782 44046 38834
rect 44046 38782 44098 38834
rect 44098 38782 44100 38834
rect 44044 38780 44100 38782
rect 44828 36370 44884 36372
rect 44828 36318 44830 36370
rect 44830 36318 44882 36370
rect 44882 36318 44884 36370
rect 44828 36316 44884 36318
rect 44268 36204 44324 36260
rect 44940 36258 44996 36260
rect 44940 36206 44942 36258
rect 44942 36206 44994 36258
rect 44994 36206 44996 36258
rect 44940 36204 44996 36206
rect 44716 35698 44772 35700
rect 44716 35646 44718 35698
rect 44718 35646 44770 35698
rect 44770 35646 44772 35698
rect 44716 35644 44772 35646
rect 46508 38892 46564 38948
rect 45388 36370 45444 36372
rect 45388 36318 45390 36370
rect 45390 36318 45442 36370
rect 45442 36318 45444 36370
rect 45388 36316 45444 36318
rect 45388 35698 45444 35700
rect 45388 35646 45390 35698
rect 45390 35646 45442 35698
rect 45442 35646 45444 35698
rect 45388 35644 45444 35646
rect 45612 35586 45668 35588
rect 45612 35534 45614 35586
rect 45614 35534 45666 35586
rect 45666 35534 45668 35586
rect 45612 35532 45668 35534
rect 44380 34690 44436 34692
rect 44380 34638 44382 34690
rect 44382 34638 44434 34690
rect 44434 34638 44436 34690
rect 44380 34636 44436 34638
rect 44156 34242 44212 34244
rect 44156 34190 44158 34242
rect 44158 34190 44210 34242
rect 44210 34190 44212 34242
rect 44156 34188 44212 34190
rect 44492 33292 44548 33348
rect 44380 31666 44436 31668
rect 44380 31614 44382 31666
rect 44382 31614 44434 31666
rect 44434 31614 44436 31666
rect 44380 31612 44436 31614
rect 44156 31106 44212 31108
rect 44156 31054 44158 31106
rect 44158 31054 44210 31106
rect 44210 31054 44212 31106
rect 44156 31052 44212 31054
rect 45612 34914 45668 34916
rect 45612 34862 45614 34914
rect 45614 34862 45666 34914
rect 45666 34862 45668 34914
rect 45612 34860 45668 34862
rect 44828 34636 44884 34692
rect 45836 35810 45892 35812
rect 45836 35758 45838 35810
rect 45838 35758 45890 35810
rect 45890 35758 45892 35810
rect 45836 35756 45892 35758
rect 45388 33346 45444 33348
rect 45388 33294 45390 33346
rect 45390 33294 45442 33346
rect 45442 33294 45444 33346
rect 45388 33292 45444 33294
rect 45500 32732 45556 32788
rect 45724 34076 45780 34132
rect 45836 33346 45892 33348
rect 45836 33294 45838 33346
rect 45838 33294 45890 33346
rect 45890 33294 45892 33346
rect 45836 33292 45892 33294
rect 46396 33292 46452 33348
rect 45276 31890 45332 31892
rect 45276 31838 45278 31890
rect 45278 31838 45330 31890
rect 45330 31838 45332 31890
rect 45276 31836 45332 31838
rect 44940 31778 44996 31780
rect 44940 31726 44942 31778
rect 44942 31726 44994 31778
rect 44994 31726 44996 31778
rect 44940 31724 44996 31726
rect 45724 31778 45780 31780
rect 45724 31726 45726 31778
rect 45726 31726 45778 31778
rect 45778 31726 45780 31778
rect 45724 31724 45780 31726
rect 44828 31666 44884 31668
rect 44828 31614 44830 31666
rect 44830 31614 44882 31666
rect 44882 31614 44884 31666
rect 44828 31612 44884 31614
rect 45500 31106 45556 31108
rect 45500 31054 45502 31106
rect 45502 31054 45554 31106
rect 45554 31054 45556 31106
rect 45500 31052 45556 31054
rect 45276 30994 45332 30996
rect 45276 30942 45278 30994
rect 45278 30942 45330 30994
rect 45330 30942 45332 30994
rect 45276 30940 45332 30942
rect 45612 30940 45668 30996
rect 45500 30716 45556 30772
rect 44492 30156 44548 30212
rect 44940 30044 44996 30100
rect 44604 29538 44660 29540
rect 44604 29486 44606 29538
rect 44606 29486 44658 29538
rect 44658 29486 44660 29538
rect 44604 29484 44660 29486
rect 44716 28476 44772 28532
rect 45052 28476 45108 28532
rect 44828 27244 44884 27300
rect 44044 27132 44100 27188
rect 45388 27244 45444 27300
rect 44940 26962 44996 26964
rect 44940 26910 44942 26962
rect 44942 26910 44994 26962
rect 44994 26910 44996 26962
rect 44940 26908 44996 26910
rect 46620 35810 46676 35812
rect 46620 35758 46622 35810
rect 46622 35758 46674 35810
rect 46674 35758 46676 35810
rect 46620 35756 46676 35758
rect 46956 36204 47012 36260
rect 46844 35586 46900 35588
rect 46844 35534 46846 35586
rect 46846 35534 46898 35586
rect 46898 35534 46900 35586
rect 46844 35532 46900 35534
rect 46508 32732 46564 32788
rect 45948 31778 46004 31780
rect 45948 31726 45950 31778
rect 45950 31726 46002 31778
rect 46002 31726 46004 31778
rect 45948 31724 46004 31726
rect 45948 30882 46004 30884
rect 45948 30830 45950 30882
rect 45950 30830 46002 30882
rect 46002 30830 46004 30882
rect 45948 30828 46004 30830
rect 44268 25452 44324 25508
rect 43596 23996 43652 24052
rect 43708 23324 43764 23380
rect 44268 23324 44324 23380
rect 43820 22764 43876 22820
rect 43708 22258 43764 22260
rect 43708 22206 43710 22258
rect 43710 22206 43762 22258
rect 43762 22206 43764 22258
rect 43708 22204 43764 22206
rect 45052 26290 45108 26292
rect 45052 26238 45054 26290
rect 45054 26238 45106 26290
rect 45106 26238 45108 26290
rect 45052 26236 45108 26238
rect 44940 26012 44996 26068
rect 44940 25506 44996 25508
rect 44940 25454 44942 25506
rect 44942 25454 44994 25506
rect 44994 25454 44996 25506
rect 44940 25452 44996 25454
rect 44604 25228 44660 25284
rect 44828 24780 44884 24836
rect 44604 24556 44660 24612
rect 45164 24834 45220 24836
rect 45164 24782 45166 24834
rect 45166 24782 45218 24834
rect 45218 24782 45220 24834
rect 45164 24780 45220 24782
rect 44940 24050 44996 24052
rect 44940 23998 44942 24050
rect 44942 23998 44994 24050
rect 44994 23998 44996 24050
rect 44940 23996 44996 23998
rect 44828 23884 44884 23940
rect 45164 23884 45220 23940
rect 45052 23660 45108 23716
rect 43484 20076 43540 20132
rect 43932 21980 43988 22036
rect 43036 19292 43092 19348
rect 43148 18338 43204 18340
rect 43148 18286 43150 18338
rect 43150 18286 43202 18338
rect 43202 18286 43204 18338
rect 43148 18284 43204 18286
rect 43036 17724 43092 17780
rect 43148 17666 43204 17668
rect 43148 17614 43150 17666
rect 43150 17614 43202 17666
rect 43202 17614 43204 17666
rect 43148 17612 43204 17614
rect 42588 16380 42644 16436
rect 38556 11004 38612 11060
rect 39676 11340 39732 11396
rect 38668 11116 38724 11172
rect 39564 10892 39620 10948
rect 37996 9996 38052 10052
rect 37548 9884 37604 9940
rect 37324 9714 37380 9716
rect 37324 9662 37326 9714
rect 37326 9662 37378 9714
rect 37378 9662 37380 9714
rect 37324 9660 37380 9662
rect 38780 9996 38836 10052
rect 40348 11340 40404 11396
rect 40348 10892 40404 10948
rect 39788 9772 39844 9828
rect 37660 9660 37716 9716
rect 39004 9660 39060 9716
rect 36876 8764 36932 8820
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 34412 7474 34468 7476
rect 34412 7422 34414 7474
rect 34414 7422 34466 7474
rect 34466 7422 34468 7474
rect 34412 7420 34468 7422
rect 34188 6636 34244 6692
rect 34412 6860 34468 6916
rect 34972 7644 35028 7700
rect 37324 8204 37380 8260
rect 35308 7756 35364 7812
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 34636 6748 34692 6804
rect 35644 6076 35700 6132
rect 34300 5964 34356 6020
rect 33516 5852 33572 5908
rect 33852 5906 33908 5908
rect 33852 5854 33854 5906
rect 33854 5854 33906 5906
rect 33906 5854 33908 5906
rect 33852 5852 33908 5854
rect 33292 5516 33348 5572
rect 33180 5068 33236 5124
rect 32396 4562 32452 4564
rect 32396 4510 32398 4562
rect 32398 4510 32450 4562
rect 32450 4510 32452 4562
rect 32396 4508 32452 4510
rect 32732 4396 32788 4452
rect 32508 3612 32564 3668
rect 32396 3554 32452 3556
rect 32396 3502 32398 3554
rect 32398 3502 32450 3554
rect 32450 3502 32452 3554
rect 32396 3500 32452 3502
rect 32956 4338 33012 4340
rect 32956 4286 32958 4338
rect 32958 4286 33010 4338
rect 33010 4286 33012 4338
rect 32956 4284 33012 4286
rect 33292 4844 33348 4900
rect 33404 4620 33460 4676
rect 33516 5068 33572 5124
rect 33180 4284 33236 4340
rect 33404 4284 33460 4340
rect 33068 2828 33124 2884
rect 33180 4060 33236 4116
rect 33516 2716 33572 2772
rect 34300 5794 34356 5796
rect 34300 5742 34302 5794
rect 34302 5742 34354 5794
rect 34354 5742 34356 5794
rect 34300 5740 34356 5742
rect 33852 5682 33908 5684
rect 33852 5630 33854 5682
rect 33854 5630 33906 5682
rect 33906 5630 33908 5682
rect 33852 5628 33908 5630
rect 33740 5516 33796 5572
rect 33740 3612 33796 3668
rect 33852 5180 33908 5236
rect 33628 1372 33684 1428
rect 34076 5180 34132 5236
rect 34524 4620 34580 4676
rect 34188 4508 34244 4564
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 35308 5010 35364 5012
rect 35308 4958 35310 5010
rect 35310 4958 35362 5010
rect 35362 4958 35364 5010
rect 35308 4956 35364 4958
rect 34972 4172 35028 4228
rect 34524 3554 34580 3556
rect 34524 3502 34526 3554
rect 34526 3502 34578 3554
rect 34578 3502 34580 3554
rect 34524 3500 34580 3502
rect 34748 4060 34804 4116
rect 34860 3836 34916 3892
rect 34972 3724 35028 3780
rect 35532 4172 35588 4228
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 34524 2268 34580 2324
rect 37100 8034 37156 8036
rect 37100 7982 37102 8034
rect 37102 7982 37154 8034
rect 37154 7982 37156 8034
rect 37100 7980 37156 7982
rect 37324 7532 37380 7588
rect 36428 7420 36484 7476
rect 36428 6860 36484 6916
rect 36540 6636 36596 6692
rect 37660 7868 37716 7924
rect 37996 9602 38052 9604
rect 37996 9550 37998 9602
rect 37998 9550 38050 9602
rect 38050 9550 38052 9602
rect 37996 9548 38052 9550
rect 37772 7420 37828 7476
rect 38556 9436 38612 9492
rect 38332 8204 38388 8260
rect 38668 9100 38724 9156
rect 38892 8204 38948 8260
rect 39452 9714 39508 9716
rect 39452 9662 39454 9714
rect 39454 9662 39506 9714
rect 39506 9662 39508 9714
rect 39452 9660 39508 9662
rect 39788 9100 39844 9156
rect 40908 9660 40964 9716
rect 41692 15148 41748 15204
rect 42028 15148 42084 15204
rect 41468 14028 41524 14084
rect 41580 13804 41636 13860
rect 42252 15874 42308 15876
rect 42252 15822 42254 15874
rect 42254 15822 42306 15874
rect 42306 15822 42308 15874
rect 42252 15820 42308 15822
rect 42588 15820 42644 15876
rect 42924 16156 42980 16212
rect 43036 16098 43092 16100
rect 43036 16046 43038 16098
rect 43038 16046 43090 16098
rect 43090 16046 43092 16098
rect 43036 16044 43092 16046
rect 42700 15596 42756 15652
rect 44268 21698 44324 21700
rect 44268 21646 44270 21698
rect 44270 21646 44322 21698
rect 44322 21646 44324 21698
rect 44268 21644 44324 21646
rect 44044 21532 44100 21588
rect 44156 20188 44212 20244
rect 43372 18060 43428 18116
rect 43372 16604 43428 16660
rect 43932 17948 43988 18004
rect 43708 16604 43764 16660
rect 43820 17724 43876 17780
rect 43820 17164 43876 17220
rect 43596 16268 43652 16324
rect 43484 16156 43540 16212
rect 43260 15596 43316 15652
rect 42700 14700 42756 14756
rect 42924 14418 42980 14420
rect 42924 14366 42926 14418
rect 42926 14366 42978 14418
rect 42978 14366 42980 14418
rect 42924 14364 42980 14366
rect 42476 13916 42532 13972
rect 42364 12962 42420 12964
rect 42364 12910 42366 12962
rect 42366 12910 42418 12962
rect 42418 12910 42420 12962
rect 42364 12908 42420 12910
rect 42028 12796 42084 12852
rect 41580 12178 41636 12180
rect 41580 12126 41582 12178
rect 41582 12126 41634 12178
rect 41634 12126 41636 12178
rect 41580 12124 41636 12126
rect 41468 12012 41524 12068
rect 41692 11340 41748 11396
rect 38892 7756 38948 7812
rect 38668 7586 38724 7588
rect 38668 7534 38670 7586
rect 38670 7534 38722 7586
rect 38722 7534 38724 7586
rect 38668 7532 38724 7534
rect 38444 6748 38500 6804
rect 36540 5292 36596 5348
rect 36764 5628 36820 5684
rect 36092 4508 36148 4564
rect 36428 4732 36484 4788
rect 35868 3724 35924 3780
rect 36316 3836 36372 3892
rect 36652 4450 36708 4452
rect 36652 4398 36654 4450
rect 36654 4398 36706 4450
rect 36706 4398 36708 4450
rect 36652 4396 36708 4398
rect 36540 4338 36596 4340
rect 36540 4286 36542 4338
rect 36542 4286 36594 4338
rect 36594 4286 36596 4338
rect 36540 4284 36596 4286
rect 35084 3164 35140 3220
rect 35980 2380 36036 2436
rect 35868 1820 35924 1876
rect 36876 3836 36932 3892
rect 37548 5852 37604 5908
rect 37324 5122 37380 5124
rect 37324 5070 37326 5122
rect 37326 5070 37378 5122
rect 37378 5070 37380 5122
rect 37324 5068 37380 5070
rect 38108 5740 38164 5796
rect 37884 5068 37940 5124
rect 38332 5292 38388 5348
rect 39116 7644 39172 7700
rect 39228 6972 39284 7028
rect 39788 8204 39844 8260
rect 39676 7698 39732 7700
rect 39676 7646 39678 7698
rect 39678 7646 39730 7698
rect 39730 7646 39732 7698
rect 39676 7644 39732 7646
rect 39564 6636 39620 6692
rect 39788 6188 39844 6244
rect 39452 5292 39508 5348
rect 40124 6972 40180 7028
rect 40908 8146 40964 8148
rect 40908 8094 40910 8146
rect 40910 8094 40962 8146
rect 40962 8094 40964 8146
rect 40908 8092 40964 8094
rect 41020 7756 41076 7812
rect 40908 7644 40964 7700
rect 40684 6466 40740 6468
rect 40684 6414 40686 6466
rect 40686 6414 40738 6466
rect 40738 6414 40740 6466
rect 40684 6412 40740 6414
rect 40012 5740 40068 5796
rect 39676 5068 39732 5124
rect 40012 5122 40068 5124
rect 40012 5070 40014 5122
rect 40014 5070 40066 5122
rect 40066 5070 40068 5122
rect 40012 5068 40068 5070
rect 39788 4844 39844 4900
rect 40460 5122 40516 5124
rect 40460 5070 40462 5122
rect 40462 5070 40514 5122
rect 40514 5070 40516 5122
rect 40460 5068 40516 5070
rect 40236 4956 40292 5012
rect 38556 3388 38612 3444
rect 37436 3052 37492 3108
rect 36988 2940 37044 2996
rect 37212 2156 37268 2212
rect 37884 1708 37940 1764
rect 38668 3276 38724 3332
rect 39340 3948 39396 4004
rect 39900 3612 39956 3668
rect 38892 1596 38948 1652
rect 39004 1484 39060 1540
rect 39228 2828 39284 2884
rect 40572 4060 40628 4116
rect 41580 9884 41636 9940
rect 41804 9938 41860 9940
rect 41804 9886 41806 9938
rect 41806 9886 41858 9938
rect 41858 9886 41860 9938
rect 41804 9884 41860 9886
rect 41244 7756 41300 7812
rect 42364 12402 42420 12404
rect 42364 12350 42366 12402
rect 42366 12350 42418 12402
rect 42418 12350 42420 12402
rect 42364 12348 42420 12350
rect 42364 10220 42420 10276
rect 42364 9884 42420 9940
rect 42700 13692 42756 13748
rect 43148 12796 43204 12852
rect 42588 9996 42644 10052
rect 42588 9826 42644 9828
rect 42588 9774 42590 9826
rect 42590 9774 42642 9826
rect 42642 9774 42644 9826
rect 42588 9772 42644 9774
rect 42140 9602 42196 9604
rect 42140 9550 42142 9602
rect 42142 9550 42194 9602
rect 42194 9550 42196 9602
rect 42140 9548 42196 9550
rect 43148 9602 43204 9604
rect 43148 9550 43150 9602
rect 43150 9550 43202 9602
rect 43202 9550 43204 9602
rect 43148 9548 43204 9550
rect 42364 8146 42420 8148
rect 42364 8094 42366 8146
rect 42366 8094 42418 8146
rect 42418 8094 42420 8146
rect 42364 8092 42420 8094
rect 43036 8258 43092 8260
rect 43036 8206 43038 8258
rect 43038 8206 43090 8258
rect 43090 8206 43092 8258
rect 43036 8204 43092 8206
rect 43372 9996 43428 10052
rect 43372 9436 43428 9492
rect 43596 8092 43652 8148
rect 42476 7756 42532 7812
rect 41356 7420 41412 7476
rect 41468 7532 41524 7588
rect 43036 7420 43092 7476
rect 43036 6748 43092 6804
rect 44044 17836 44100 17892
rect 44044 15874 44100 15876
rect 44044 15822 44046 15874
rect 44046 15822 44098 15874
rect 44098 15822 44100 15874
rect 44044 15820 44100 15822
rect 43932 9602 43988 9604
rect 43932 9550 43934 9602
rect 43934 9550 43986 9602
rect 43986 9550 43988 9602
rect 43932 9548 43988 9550
rect 43932 8876 43988 8932
rect 44492 20130 44548 20132
rect 44492 20078 44494 20130
rect 44494 20078 44546 20130
rect 44546 20078 44548 20130
rect 44492 20076 44548 20078
rect 45500 26012 45556 26068
rect 45500 25676 45556 25732
rect 45724 30210 45780 30212
rect 45724 30158 45726 30210
rect 45726 30158 45778 30210
rect 45778 30158 45780 30210
rect 45724 30156 45780 30158
rect 45612 25452 45668 25508
rect 46060 30380 46116 30436
rect 46172 30210 46228 30212
rect 46172 30158 46174 30210
rect 46174 30158 46226 30210
rect 46226 30158 46228 30210
rect 46172 30156 46228 30158
rect 46284 31052 46340 31108
rect 46508 30716 46564 30772
rect 46284 30268 46340 30324
rect 46732 30268 46788 30324
rect 45388 24556 45444 24612
rect 45836 28476 45892 28532
rect 46956 30210 47012 30212
rect 46956 30158 46958 30210
rect 46958 30158 47010 30210
rect 47010 30158 47012 30210
rect 46956 30156 47012 30158
rect 47180 30210 47236 30212
rect 47180 30158 47182 30210
rect 47182 30158 47234 30210
rect 47234 30158 47236 30210
rect 47180 30156 47236 30158
rect 47292 30098 47348 30100
rect 47292 30046 47294 30098
rect 47294 30046 47346 30098
rect 47346 30046 47348 30098
rect 47292 30044 47348 30046
rect 45836 27186 45892 27188
rect 45836 27134 45838 27186
rect 45838 27134 45890 27186
rect 45890 27134 45892 27186
rect 45836 27132 45892 27134
rect 46060 26460 46116 26516
rect 46172 26402 46228 26404
rect 46172 26350 46174 26402
rect 46174 26350 46226 26402
rect 46226 26350 46228 26402
rect 46172 26348 46228 26350
rect 46396 26290 46452 26292
rect 46396 26238 46398 26290
rect 46398 26238 46450 26290
rect 46450 26238 46452 26290
rect 46396 26236 46452 26238
rect 45836 25564 45892 25620
rect 45836 25228 45892 25284
rect 45388 23714 45444 23716
rect 45388 23662 45390 23714
rect 45390 23662 45442 23714
rect 45442 23662 45444 23714
rect 45388 23660 45444 23662
rect 45388 21756 45444 21812
rect 45724 23938 45780 23940
rect 45724 23886 45726 23938
rect 45726 23886 45778 23938
rect 45778 23886 45780 23938
rect 45724 23884 45780 23886
rect 46620 27244 46676 27300
rect 46732 26460 46788 26516
rect 46844 26402 46900 26404
rect 46844 26350 46846 26402
rect 46846 26350 46898 26402
rect 46898 26350 46900 26402
rect 46844 26348 46900 26350
rect 47516 27074 47572 27076
rect 47516 27022 47518 27074
rect 47518 27022 47570 27074
rect 47570 27022 47572 27074
rect 47516 27020 47572 27022
rect 47292 26908 47348 26964
rect 46620 26290 46676 26292
rect 46620 26238 46622 26290
rect 46622 26238 46674 26290
rect 46674 26238 46676 26290
rect 46620 26236 46676 26238
rect 47740 26402 47796 26404
rect 47740 26350 47742 26402
rect 47742 26350 47794 26402
rect 47794 26350 47796 26402
rect 47740 26348 47796 26350
rect 46508 25564 46564 25620
rect 46060 25452 46116 25508
rect 46956 26124 47012 26180
rect 47852 26124 47908 26180
rect 47516 26012 47572 26068
rect 46956 25394 47012 25396
rect 46956 25342 46958 25394
rect 46958 25342 47010 25394
rect 47010 25342 47012 25394
rect 46956 25340 47012 25342
rect 47516 25394 47572 25396
rect 47516 25342 47518 25394
rect 47518 25342 47570 25394
rect 47570 25342 47572 25394
rect 47516 25340 47572 25342
rect 46060 23714 46116 23716
rect 46060 23662 46062 23714
rect 46062 23662 46114 23714
rect 46114 23662 46116 23714
rect 46060 23660 46116 23662
rect 46396 23548 46452 23604
rect 45836 23212 45892 23268
rect 46844 23378 46900 23380
rect 46844 23326 46846 23378
rect 46846 23326 46898 23378
rect 46898 23326 46900 23378
rect 46844 23324 46900 23326
rect 45948 22370 46004 22372
rect 45948 22318 45950 22370
rect 45950 22318 46002 22370
rect 46002 22318 46004 22370
rect 45948 22316 46004 22318
rect 46284 23100 46340 23156
rect 46844 22930 46900 22932
rect 46844 22878 46846 22930
rect 46846 22878 46898 22930
rect 46898 22878 46900 22930
rect 46844 22876 46900 22878
rect 47964 24332 48020 24388
rect 48076 29148 48132 29204
rect 47292 23884 47348 23940
rect 46956 22540 47012 22596
rect 45612 21586 45668 21588
rect 45612 21534 45614 21586
rect 45614 21534 45666 21586
rect 45666 21534 45668 21586
rect 45612 21532 45668 21534
rect 45500 21308 45556 21364
rect 45052 20188 45108 20244
rect 44716 18172 44772 18228
rect 45052 18732 45108 18788
rect 44940 17724 44996 17780
rect 44940 17164 44996 17220
rect 44268 16156 44324 16212
rect 45612 18450 45668 18452
rect 45612 18398 45614 18450
rect 45614 18398 45666 18450
rect 45666 18398 45668 18450
rect 45612 18396 45668 18398
rect 45500 18338 45556 18340
rect 45500 18286 45502 18338
rect 45502 18286 45554 18338
rect 45554 18286 45556 18338
rect 45500 18284 45556 18286
rect 45388 17836 45444 17892
rect 45052 17612 45108 17668
rect 45612 16994 45668 16996
rect 45612 16942 45614 16994
rect 45614 16942 45666 16994
rect 45666 16942 45668 16994
rect 45612 16940 45668 16942
rect 47068 23548 47124 23604
rect 47404 23660 47460 23716
rect 47964 23266 48020 23268
rect 47964 23214 47966 23266
rect 47966 23214 48018 23266
rect 48018 23214 48020 23266
rect 47964 23212 48020 23214
rect 47292 23154 47348 23156
rect 47292 23102 47294 23154
rect 47294 23102 47346 23154
rect 47346 23102 47348 23154
rect 47292 23100 47348 23102
rect 47068 22316 47124 22372
rect 46396 22092 46452 22148
rect 46172 21644 46228 21700
rect 46396 21756 46452 21812
rect 46284 21532 46340 21588
rect 46172 21084 46228 21140
rect 45948 19516 46004 19572
rect 45388 16268 45444 16324
rect 45500 16492 45556 16548
rect 45164 14754 45220 14756
rect 45164 14702 45166 14754
rect 45166 14702 45218 14754
rect 45218 14702 45220 14754
rect 45164 14700 45220 14702
rect 45500 14252 45556 14308
rect 45388 13746 45444 13748
rect 45388 13694 45390 13746
rect 45390 13694 45442 13746
rect 45442 13694 45444 13746
rect 45388 13692 45444 13694
rect 45276 13468 45332 13524
rect 45164 11116 45220 11172
rect 45164 10220 45220 10276
rect 46060 16492 46116 16548
rect 45836 16268 45892 16324
rect 45724 15708 45780 15764
rect 45836 15820 45892 15876
rect 45612 11788 45668 11844
rect 45836 9772 45892 9828
rect 45276 8930 45332 8932
rect 45276 8878 45278 8930
rect 45278 8878 45330 8930
rect 45330 8878 45332 8930
rect 45276 8876 45332 8878
rect 44716 8258 44772 8260
rect 44716 8206 44718 8258
rect 44718 8206 44770 8258
rect 44770 8206 44772 8258
rect 44716 8204 44772 8206
rect 43932 7980 43988 8036
rect 44044 7532 44100 7588
rect 44380 8092 44436 8148
rect 45052 8146 45108 8148
rect 45052 8094 45054 8146
rect 45054 8094 45106 8146
rect 45106 8094 45108 8146
rect 45052 8092 45108 8094
rect 44940 7644 44996 7700
rect 44492 7586 44548 7588
rect 44492 7534 44494 7586
rect 44494 7534 44546 7586
rect 44546 7534 44548 7586
rect 44492 7532 44548 7534
rect 44268 6972 44324 7028
rect 44380 6188 44436 6244
rect 42252 6018 42308 6020
rect 42252 5966 42254 6018
rect 42254 5966 42306 6018
rect 42306 5966 42308 6018
rect 42252 5964 42308 5966
rect 41804 5906 41860 5908
rect 41804 5854 41806 5906
rect 41806 5854 41858 5906
rect 41858 5854 41860 5906
rect 41804 5852 41860 5854
rect 42476 5852 42532 5908
rect 41580 4844 41636 4900
rect 41804 5068 41860 5124
rect 42140 5180 42196 5236
rect 40796 4060 40852 4116
rect 41244 4060 41300 4116
rect 40236 3612 40292 3668
rect 41132 3836 41188 3892
rect 40572 3500 40628 3556
rect 41916 3836 41972 3892
rect 42252 3500 42308 3556
rect 42476 4956 42532 5012
rect 42700 4284 42756 4340
rect 42588 3724 42644 3780
rect 42476 3164 42532 3220
rect 44268 5906 44324 5908
rect 44268 5854 44270 5906
rect 44270 5854 44322 5906
rect 44322 5854 44324 5906
rect 44268 5852 44324 5854
rect 43260 5180 43316 5236
rect 43148 4172 43204 4228
rect 43036 3948 43092 4004
rect 43036 3388 43092 3444
rect 43708 4508 43764 4564
rect 43932 3948 43988 4004
rect 45164 6018 45220 6020
rect 45164 5966 45166 6018
rect 45166 5966 45218 6018
rect 45218 5966 45220 6018
rect 45164 5964 45220 5966
rect 44828 5852 44884 5908
rect 45164 5516 45220 5572
rect 44604 3612 44660 3668
rect 45724 6748 45780 6804
rect 45500 5180 45556 5236
rect 45612 5964 45668 6020
rect 45388 4844 45444 4900
rect 45612 4508 45668 4564
rect 47180 21532 47236 21588
rect 47068 20802 47124 20804
rect 47068 20750 47070 20802
rect 47070 20750 47122 20802
rect 47122 20750 47124 20802
rect 47068 20748 47124 20750
rect 46396 20188 46452 20244
rect 46732 19292 46788 19348
rect 46284 19180 46340 19236
rect 46620 19234 46676 19236
rect 46620 19182 46622 19234
rect 46622 19182 46674 19234
rect 46674 19182 46676 19234
rect 46620 19180 46676 19182
rect 46620 19010 46676 19012
rect 46620 18958 46622 19010
rect 46622 18958 46674 19010
rect 46674 18958 46676 19010
rect 46620 18956 46676 18958
rect 46620 18620 46676 18676
rect 46284 18508 46340 18564
rect 46284 15932 46340 15988
rect 46732 17724 46788 17780
rect 46396 15874 46452 15876
rect 46396 15822 46398 15874
rect 46398 15822 46450 15874
rect 46450 15822 46452 15874
rect 46396 15820 46452 15822
rect 46396 15596 46452 15652
rect 47068 19740 47124 19796
rect 46956 19180 47012 19236
rect 46956 17666 47012 17668
rect 46956 17614 46958 17666
rect 46958 17614 47010 17666
rect 47010 17614 47012 17666
rect 46956 17612 47012 17614
rect 47180 18844 47236 18900
rect 47068 16882 47124 16884
rect 47068 16830 47070 16882
rect 47070 16830 47122 16882
rect 47122 16830 47124 16882
rect 47068 16828 47124 16830
rect 47180 16716 47236 16772
rect 47628 22876 47684 22932
rect 47964 22652 48020 22708
rect 47628 22540 47684 22596
rect 47404 21698 47460 21700
rect 47404 21646 47406 21698
rect 47406 21646 47458 21698
rect 47458 21646 47460 21698
rect 47404 21644 47460 21646
rect 47404 20188 47460 20244
rect 47404 19852 47460 19908
rect 47292 15372 47348 15428
rect 47068 14588 47124 14644
rect 47628 21698 47684 21700
rect 47628 21646 47630 21698
rect 47630 21646 47682 21698
rect 47682 21646 47684 21698
rect 47628 21644 47684 21646
rect 47628 20802 47684 20804
rect 47628 20750 47630 20802
rect 47630 20750 47682 20802
rect 47682 20750 47684 20802
rect 47628 20748 47684 20750
rect 48076 22092 48132 22148
rect 48188 21756 48244 21812
rect 47852 20748 47908 20804
rect 48188 20972 48244 21028
rect 48188 20524 48244 20580
rect 48076 19964 48132 20020
rect 47740 17948 47796 18004
rect 47740 16716 47796 16772
rect 48076 16828 48132 16884
rect 49196 76690 49252 76692
rect 49196 76638 49198 76690
rect 49198 76638 49250 76690
rect 49250 76638 49252 76690
rect 49196 76636 49252 76638
rect 50556 76858 50612 76860
rect 50556 76806 50558 76858
rect 50558 76806 50610 76858
rect 50610 76806 50612 76858
rect 50556 76804 50612 76806
rect 50660 76858 50716 76860
rect 50660 76806 50662 76858
rect 50662 76806 50714 76858
rect 50714 76806 50716 76858
rect 50660 76804 50716 76806
rect 50764 76858 50820 76860
rect 50764 76806 50766 76858
rect 50766 76806 50818 76858
rect 50818 76806 50820 76858
rect 50764 76804 50820 76806
rect 50204 76636 50260 76692
rect 51212 76690 51268 76692
rect 51212 76638 51214 76690
rect 51214 76638 51266 76690
rect 51266 76638 51268 76690
rect 51212 76636 51268 76638
rect 50092 75740 50148 75796
rect 50764 75794 50820 75796
rect 50764 75742 50766 75794
rect 50766 75742 50818 75794
rect 50818 75742 50820 75794
rect 50764 75740 50820 75742
rect 50540 75628 50596 75684
rect 50556 75290 50612 75292
rect 50556 75238 50558 75290
rect 50558 75238 50610 75290
rect 50610 75238 50612 75290
rect 50556 75236 50612 75238
rect 50660 75290 50716 75292
rect 50660 75238 50662 75290
rect 50662 75238 50714 75290
rect 50714 75238 50716 75290
rect 50660 75236 50716 75238
rect 50764 75290 50820 75292
rect 50764 75238 50766 75290
rect 50766 75238 50818 75290
rect 50818 75238 50820 75290
rect 50764 75236 50820 75238
rect 50556 73722 50612 73724
rect 50556 73670 50558 73722
rect 50558 73670 50610 73722
rect 50610 73670 50612 73722
rect 50556 73668 50612 73670
rect 50660 73722 50716 73724
rect 50660 73670 50662 73722
rect 50662 73670 50714 73722
rect 50714 73670 50716 73722
rect 50660 73668 50716 73670
rect 50764 73722 50820 73724
rect 50764 73670 50766 73722
rect 50766 73670 50818 73722
rect 50818 73670 50820 73722
rect 50764 73668 50820 73670
rect 50556 72154 50612 72156
rect 50556 72102 50558 72154
rect 50558 72102 50610 72154
rect 50610 72102 50612 72154
rect 50556 72100 50612 72102
rect 50660 72154 50716 72156
rect 50660 72102 50662 72154
rect 50662 72102 50714 72154
rect 50714 72102 50716 72154
rect 50660 72100 50716 72102
rect 50764 72154 50820 72156
rect 50764 72102 50766 72154
rect 50766 72102 50818 72154
rect 50818 72102 50820 72154
rect 50764 72100 50820 72102
rect 50556 70586 50612 70588
rect 50556 70534 50558 70586
rect 50558 70534 50610 70586
rect 50610 70534 50612 70586
rect 50556 70532 50612 70534
rect 50660 70586 50716 70588
rect 50660 70534 50662 70586
rect 50662 70534 50714 70586
rect 50714 70534 50716 70586
rect 50660 70532 50716 70534
rect 50764 70586 50820 70588
rect 50764 70534 50766 70586
rect 50766 70534 50818 70586
rect 50818 70534 50820 70586
rect 50764 70532 50820 70534
rect 50556 69018 50612 69020
rect 50556 68966 50558 69018
rect 50558 68966 50610 69018
rect 50610 68966 50612 69018
rect 50556 68964 50612 68966
rect 50660 69018 50716 69020
rect 50660 68966 50662 69018
rect 50662 68966 50714 69018
rect 50714 68966 50716 69018
rect 50660 68964 50716 68966
rect 50764 69018 50820 69020
rect 50764 68966 50766 69018
rect 50766 68966 50818 69018
rect 50818 68966 50820 69018
rect 50764 68964 50820 68966
rect 50556 67450 50612 67452
rect 50556 67398 50558 67450
rect 50558 67398 50610 67450
rect 50610 67398 50612 67450
rect 50556 67396 50612 67398
rect 50660 67450 50716 67452
rect 50660 67398 50662 67450
rect 50662 67398 50714 67450
rect 50714 67398 50716 67450
rect 50660 67396 50716 67398
rect 50764 67450 50820 67452
rect 50764 67398 50766 67450
rect 50766 67398 50818 67450
rect 50818 67398 50820 67450
rect 50764 67396 50820 67398
rect 50556 65882 50612 65884
rect 50556 65830 50558 65882
rect 50558 65830 50610 65882
rect 50610 65830 50612 65882
rect 50556 65828 50612 65830
rect 50660 65882 50716 65884
rect 50660 65830 50662 65882
rect 50662 65830 50714 65882
rect 50714 65830 50716 65882
rect 50660 65828 50716 65830
rect 50764 65882 50820 65884
rect 50764 65830 50766 65882
rect 50766 65830 50818 65882
rect 50818 65830 50820 65882
rect 50764 65828 50820 65830
rect 50556 64314 50612 64316
rect 50556 64262 50558 64314
rect 50558 64262 50610 64314
rect 50610 64262 50612 64314
rect 50556 64260 50612 64262
rect 50660 64314 50716 64316
rect 50660 64262 50662 64314
rect 50662 64262 50714 64314
rect 50714 64262 50716 64314
rect 50660 64260 50716 64262
rect 50764 64314 50820 64316
rect 50764 64262 50766 64314
rect 50766 64262 50818 64314
rect 50818 64262 50820 64314
rect 50764 64260 50820 64262
rect 50556 62746 50612 62748
rect 50556 62694 50558 62746
rect 50558 62694 50610 62746
rect 50610 62694 50612 62746
rect 50556 62692 50612 62694
rect 50660 62746 50716 62748
rect 50660 62694 50662 62746
rect 50662 62694 50714 62746
rect 50714 62694 50716 62746
rect 50660 62692 50716 62694
rect 50764 62746 50820 62748
rect 50764 62694 50766 62746
rect 50766 62694 50818 62746
rect 50818 62694 50820 62746
rect 50764 62692 50820 62694
rect 50556 61178 50612 61180
rect 50556 61126 50558 61178
rect 50558 61126 50610 61178
rect 50610 61126 50612 61178
rect 50556 61124 50612 61126
rect 50660 61178 50716 61180
rect 50660 61126 50662 61178
rect 50662 61126 50714 61178
rect 50714 61126 50716 61178
rect 50660 61124 50716 61126
rect 50764 61178 50820 61180
rect 50764 61126 50766 61178
rect 50766 61126 50818 61178
rect 50818 61126 50820 61178
rect 50764 61124 50820 61126
rect 50556 59610 50612 59612
rect 50556 59558 50558 59610
rect 50558 59558 50610 59610
rect 50610 59558 50612 59610
rect 50556 59556 50612 59558
rect 50660 59610 50716 59612
rect 50660 59558 50662 59610
rect 50662 59558 50714 59610
rect 50714 59558 50716 59610
rect 50660 59556 50716 59558
rect 50764 59610 50820 59612
rect 50764 59558 50766 59610
rect 50766 59558 50818 59610
rect 50818 59558 50820 59610
rect 50764 59556 50820 59558
rect 50556 58042 50612 58044
rect 50556 57990 50558 58042
rect 50558 57990 50610 58042
rect 50610 57990 50612 58042
rect 50556 57988 50612 57990
rect 50660 58042 50716 58044
rect 50660 57990 50662 58042
rect 50662 57990 50714 58042
rect 50714 57990 50716 58042
rect 50660 57988 50716 57990
rect 50764 58042 50820 58044
rect 50764 57990 50766 58042
rect 50766 57990 50818 58042
rect 50818 57990 50820 58042
rect 50764 57988 50820 57990
rect 50556 56474 50612 56476
rect 50556 56422 50558 56474
rect 50558 56422 50610 56474
rect 50610 56422 50612 56474
rect 50556 56420 50612 56422
rect 50660 56474 50716 56476
rect 50660 56422 50662 56474
rect 50662 56422 50714 56474
rect 50714 56422 50716 56474
rect 50660 56420 50716 56422
rect 50764 56474 50820 56476
rect 50764 56422 50766 56474
rect 50766 56422 50818 56474
rect 50818 56422 50820 56474
rect 50764 56420 50820 56422
rect 52892 76636 52948 76692
rect 52780 75122 52836 75124
rect 52780 75070 52782 75122
rect 52782 75070 52834 75122
rect 52834 75070 52836 75122
rect 52780 75068 52836 75070
rect 53900 76690 53956 76692
rect 53900 76638 53902 76690
rect 53902 76638 53954 76690
rect 53954 76638 53956 76690
rect 53900 76636 53956 76638
rect 53004 75068 53060 75124
rect 52892 73836 52948 73892
rect 53340 73836 53396 73892
rect 50556 54906 50612 54908
rect 50556 54854 50558 54906
rect 50558 54854 50610 54906
rect 50610 54854 50612 54906
rect 50556 54852 50612 54854
rect 50660 54906 50716 54908
rect 50660 54854 50662 54906
rect 50662 54854 50714 54906
rect 50714 54854 50716 54906
rect 50660 54852 50716 54854
rect 50764 54906 50820 54908
rect 50764 54854 50766 54906
rect 50766 54854 50818 54906
rect 50818 54854 50820 54906
rect 50764 54852 50820 54854
rect 50556 53338 50612 53340
rect 50556 53286 50558 53338
rect 50558 53286 50610 53338
rect 50610 53286 50612 53338
rect 50556 53284 50612 53286
rect 50660 53338 50716 53340
rect 50660 53286 50662 53338
rect 50662 53286 50714 53338
rect 50714 53286 50716 53338
rect 50660 53284 50716 53286
rect 50764 53338 50820 53340
rect 50764 53286 50766 53338
rect 50766 53286 50818 53338
rect 50818 53286 50820 53338
rect 50764 53284 50820 53286
rect 50556 51770 50612 51772
rect 50556 51718 50558 51770
rect 50558 51718 50610 51770
rect 50610 51718 50612 51770
rect 50556 51716 50612 51718
rect 50660 51770 50716 51772
rect 50660 51718 50662 51770
rect 50662 51718 50714 51770
rect 50714 51718 50716 51770
rect 50660 51716 50716 51718
rect 50764 51770 50820 51772
rect 50764 51718 50766 51770
rect 50766 51718 50818 51770
rect 50818 51718 50820 51770
rect 50764 51716 50820 51718
rect 50556 50202 50612 50204
rect 50556 50150 50558 50202
rect 50558 50150 50610 50202
rect 50610 50150 50612 50202
rect 50556 50148 50612 50150
rect 50660 50202 50716 50204
rect 50660 50150 50662 50202
rect 50662 50150 50714 50202
rect 50714 50150 50716 50202
rect 50660 50148 50716 50150
rect 50764 50202 50820 50204
rect 50764 50150 50766 50202
rect 50766 50150 50818 50202
rect 50818 50150 50820 50202
rect 50764 50148 50820 50150
rect 50556 48634 50612 48636
rect 50556 48582 50558 48634
rect 50558 48582 50610 48634
rect 50610 48582 50612 48634
rect 50556 48580 50612 48582
rect 50660 48634 50716 48636
rect 50660 48582 50662 48634
rect 50662 48582 50714 48634
rect 50714 48582 50716 48634
rect 50660 48580 50716 48582
rect 50764 48634 50820 48636
rect 50764 48582 50766 48634
rect 50766 48582 50818 48634
rect 50818 48582 50820 48634
rect 50764 48580 50820 48582
rect 50556 47066 50612 47068
rect 50556 47014 50558 47066
rect 50558 47014 50610 47066
rect 50610 47014 50612 47066
rect 50556 47012 50612 47014
rect 50660 47066 50716 47068
rect 50660 47014 50662 47066
rect 50662 47014 50714 47066
rect 50714 47014 50716 47066
rect 50660 47012 50716 47014
rect 50764 47066 50820 47068
rect 50764 47014 50766 47066
rect 50766 47014 50818 47066
rect 50818 47014 50820 47066
rect 50764 47012 50820 47014
rect 50556 45498 50612 45500
rect 50556 45446 50558 45498
rect 50558 45446 50610 45498
rect 50610 45446 50612 45498
rect 50556 45444 50612 45446
rect 50660 45498 50716 45500
rect 50660 45446 50662 45498
rect 50662 45446 50714 45498
rect 50714 45446 50716 45498
rect 50660 45444 50716 45446
rect 50764 45498 50820 45500
rect 50764 45446 50766 45498
rect 50766 45446 50818 45498
rect 50818 45446 50820 45498
rect 50764 45444 50820 45446
rect 50556 43930 50612 43932
rect 50556 43878 50558 43930
rect 50558 43878 50610 43930
rect 50610 43878 50612 43930
rect 50556 43876 50612 43878
rect 50660 43930 50716 43932
rect 50660 43878 50662 43930
rect 50662 43878 50714 43930
rect 50714 43878 50716 43930
rect 50660 43876 50716 43878
rect 50764 43930 50820 43932
rect 50764 43878 50766 43930
rect 50766 43878 50818 43930
rect 50818 43878 50820 43930
rect 50764 43876 50820 43878
rect 49756 29372 49812 29428
rect 50092 30492 50148 30548
rect 49196 28588 49252 28644
rect 48972 27244 49028 27300
rect 49084 27132 49140 27188
rect 48860 26514 48916 26516
rect 48860 26462 48862 26514
rect 48862 26462 48914 26514
rect 48914 26462 48916 26514
rect 48860 26460 48916 26462
rect 48748 26290 48804 26292
rect 48748 26238 48750 26290
rect 48750 26238 48802 26290
rect 48802 26238 48804 26290
rect 48748 26236 48804 26238
rect 48524 23938 48580 23940
rect 48524 23886 48526 23938
rect 48526 23886 48578 23938
rect 48578 23886 48580 23938
rect 48524 23884 48580 23886
rect 48636 22370 48692 22372
rect 48636 22318 48638 22370
rect 48638 22318 48690 22370
rect 48690 22318 48692 22370
rect 48636 22316 48692 22318
rect 48412 20972 48468 21028
rect 48972 24332 49028 24388
rect 48972 23714 49028 23716
rect 48972 23662 48974 23714
rect 48974 23662 49026 23714
rect 49026 23662 49028 23714
rect 48972 23660 49028 23662
rect 49532 27074 49588 27076
rect 49532 27022 49534 27074
rect 49534 27022 49586 27074
rect 49586 27022 49588 27074
rect 49532 27020 49588 27022
rect 49644 26962 49700 26964
rect 49644 26910 49646 26962
rect 49646 26910 49698 26962
rect 49698 26910 49700 26962
rect 49644 26908 49700 26910
rect 48972 23378 49028 23380
rect 48972 23326 48974 23378
rect 48974 23326 49026 23378
rect 49026 23326 49028 23378
rect 48972 23324 49028 23326
rect 48860 22540 48916 22596
rect 48860 21084 48916 21140
rect 48972 22370 49028 22372
rect 48972 22318 48974 22370
rect 48974 22318 49026 22370
rect 49026 22318 49028 22370
rect 48972 22316 49028 22318
rect 48972 20802 49028 20804
rect 48972 20750 48974 20802
rect 48974 20750 49026 20802
rect 49026 20750 49028 20802
rect 48972 20748 49028 20750
rect 48524 20076 48580 20132
rect 48524 19852 48580 19908
rect 48972 20300 49028 20356
rect 48524 19346 48580 19348
rect 48524 19294 48526 19346
rect 48526 19294 48578 19346
rect 48578 19294 48580 19346
rect 48524 19292 48580 19294
rect 48300 18732 48356 18788
rect 48524 18844 48580 18900
rect 48748 20018 48804 20020
rect 48748 19966 48750 20018
rect 48750 19966 48802 20018
rect 48802 19966 48804 20018
rect 48748 19964 48804 19966
rect 49420 26402 49476 26404
rect 49420 26350 49422 26402
rect 49422 26350 49474 26402
rect 49474 26350 49476 26402
rect 49420 26348 49476 26350
rect 49308 26012 49364 26068
rect 50204 27186 50260 27188
rect 50204 27134 50206 27186
rect 50206 27134 50258 27186
rect 50258 27134 50260 27186
rect 50204 27132 50260 27134
rect 50092 26514 50148 26516
rect 50092 26462 50094 26514
rect 50094 26462 50146 26514
rect 50146 26462 50148 26514
rect 50092 26460 50148 26462
rect 49644 26290 49700 26292
rect 49644 26238 49646 26290
rect 49646 26238 49698 26290
rect 49698 26238 49700 26290
rect 49644 26236 49700 26238
rect 49980 26236 50036 26292
rect 49756 26124 49812 26180
rect 49420 23266 49476 23268
rect 49420 23214 49422 23266
rect 49422 23214 49474 23266
rect 49474 23214 49476 23266
rect 49420 23212 49476 23214
rect 49420 22876 49476 22932
rect 49756 23324 49812 23380
rect 49420 22316 49476 22372
rect 49532 21586 49588 21588
rect 49532 21534 49534 21586
rect 49534 21534 49586 21586
rect 49586 21534 49588 21586
rect 49532 21532 49588 21534
rect 49532 21084 49588 21140
rect 49420 20130 49476 20132
rect 49420 20078 49422 20130
rect 49422 20078 49474 20130
rect 49474 20078 49476 20130
rect 49420 20076 49476 20078
rect 49308 20018 49364 20020
rect 49308 19966 49310 20018
rect 49310 19966 49362 20018
rect 49362 19966 49364 20018
rect 49308 19964 49364 19966
rect 48972 19180 49028 19236
rect 48972 18732 49028 18788
rect 48748 18284 48804 18340
rect 48748 16828 48804 16884
rect 47852 15708 47908 15764
rect 47740 15596 47796 15652
rect 46956 13468 47012 13524
rect 46508 11228 46564 11284
rect 46172 8204 46228 8260
rect 45948 8034 46004 8036
rect 45948 7982 45950 8034
rect 45950 7982 46002 8034
rect 46002 7982 46004 8034
rect 45948 7980 46004 7982
rect 47292 10892 47348 10948
rect 46732 7756 46788 7812
rect 46508 7308 46564 7364
rect 46060 6076 46116 6132
rect 45948 5292 46004 5348
rect 45276 3554 45332 3556
rect 45276 3502 45278 3554
rect 45278 3502 45330 3554
rect 45330 3502 45332 3554
rect 45276 3500 45332 3502
rect 45388 3442 45444 3444
rect 45388 3390 45390 3442
rect 45390 3390 45442 3442
rect 45442 3390 45444 3442
rect 45388 3388 45444 3390
rect 46396 5068 46452 5124
rect 47068 7362 47124 7364
rect 47068 7310 47070 7362
rect 47070 7310 47122 7362
rect 47122 7310 47124 7362
rect 47068 7308 47124 7310
rect 46844 5122 46900 5124
rect 46844 5070 46846 5122
rect 46846 5070 46898 5122
rect 46898 5070 46900 5122
rect 46844 5068 46900 5070
rect 46620 4844 46676 4900
rect 46620 4508 46676 4564
rect 48076 15820 48132 15876
rect 48188 15596 48244 15652
rect 49084 18284 49140 18340
rect 49308 19180 49364 19236
rect 49308 17388 49364 17444
rect 48972 15314 49028 15316
rect 48972 15262 48974 15314
rect 48974 15262 49026 15314
rect 49026 15262 49028 15314
rect 48972 15260 49028 15262
rect 50556 42362 50612 42364
rect 50556 42310 50558 42362
rect 50558 42310 50610 42362
rect 50610 42310 50612 42362
rect 50556 42308 50612 42310
rect 50660 42362 50716 42364
rect 50660 42310 50662 42362
rect 50662 42310 50714 42362
rect 50714 42310 50716 42362
rect 50660 42308 50716 42310
rect 50764 42362 50820 42364
rect 50764 42310 50766 42362
rect 50766 42310 50818 42362
rect 50818 42310 50820 42362
rect 50764 42308 50820 42310
rect 50556 40794 50612 40796
rect 50556 40742 50558 40794
rect 50558 40742 50610 40794
rect 50610 40742 50612 40794
rect 50556 40740 50612 40742
rect 50660 40794 50716 40796
rect 50660 40742 50662 40794
rect 50662 40742 50714 40794
rect 50714 40742 50716 40794
rect 50660 40740 50716 40742
rect 50764 40794 50820 40796
rect 50764 40742 50766 40794
rect 50766 40742 50818 40794
rect 50818 40742 50820 40794
rect 50764 40740 50820 40742
rect 50556 39226 50612 39228
rect 50556 39174 50558 39226
rect 50558 39174 50610 39226
rect 50610 39174 50612 39226
rect 50556 39172 50612 39174
rect 50660 39226 50716 39228
rect 50660 39174 50662 39226
rect 50662 39174 50714 39226
rect 50714 39174 50716 39226
rect 50660 39172 50716 39174
rect 50764 39226 50820 39228
rect 50764 39174 50766 39226
rect 50766 39174 50818 39226
rect 50818 39174 50820 39226
rect 50764 39172 50820 39174
rect 50556 37658 50612 37660
rect 50556 37606 50558 37658
rect 50558 37606 50610 37658
rect 50610 37606 50612 37658
rect 50556 37604 50612 37606
rect 50660 37658 50716 37660
rect 50660 37606 50662 37658
rect 50662 37606 50714 37658
rect 50714 37606 50716 37658
rect 50660 37604 50716 37606
rect 50764 37658 50820 37660
rect 50764 37606 50766 37658
rect 50766 37606 50818 37658
rect 50818 37606 50820 37658
rect 50764 37604 50820 37606
rect 50556 36090 50612 36092
rect 50556 36038 50558 36090
rect 50558 36038 50610 36090
rect 50610 36038 50612 36090
rect 50556 36036 50612 36038
rect 50660 36090 50716 36092
rect 50660 36038 50662 36090
rect 50662 36038 50714 36090
rect 50714 36038 50716 36090
rect 50660 36036 50716 36038
rect 50764 36090 50820 36092
rect 50764 36038 50766 36090
rect 50766 36038 50818 36090
rect 50818 36038 50820 36090
rect 50764 36036 50820 36038
rect 50556 34522 50612 34524
rect 50556 34470 50558 34522
rect 50558 34470 50610 34522
rect 50610 34470 50612 34522
rect 50556 34468 50612 34470
rect 50660 34522 50716 34524
rect 50660 34470 50662 34522
rect 50662 34470 50714 34522
rect 50714 34470 50716 34522
rect 50660 34468 50716 34470
rect 50764 34522 50820 34524
rect 50764 34470 50766 34522
rect 50766 34470 50818 34522
rect 50818 34470 50820 34522
rect 50764 34468 50820 34470
rect 50556 32954 50612 32956
rect 50556 32902 50558 32954
rect 50558 32902 50610 32954
rect 50610 32902 50612 32954
rect 50556 32900 50612 32902
rect 50660 32954 50716 32956
rect 50660 32902 50662 32954
rect 50662 32902 50714 32954
rect 50714 32902 50716 32954
rect 50660 32900 50716 32902
rect 50764 32954 50820 32956
rect 50764 32902 50766 32954
rect 50766 32902 50818 32954
rect 50818 32902 50820 32954
rect 50764 32900 50820 32902
rect 50556 31386 50612 31388
rect 50556 31334 50558 31386
rect 50558 31334 50610 31386
rect 50610 31334 50612 31386
rect 50556 31332 50612 31334
rect 50660 31386 50716 31388
rect 50660 31334 50662 31386
rect 50662 31334 50714 31386
rect 50714 31334 50716 31386
rect 50660 31332 50716 31334
rect 50764 31386 50820 31388
rect 50764 31334 50766 31386
rect 50766 31334 50818 31386
rect 50818 31334 50820 31386
rect 50764 31332 50820 31334
rect 50540 30716 50596 30772
rect 50876 30210 50932 30212
rect 50876 30158 50878 30210
rect 50878 30158 50930 30210
rect 50930 30158 50932 30210
rect 50876 30156 50932 30158
rect 50556 29818 50612 29820
rect 50556 29766 50558 29818
rect 50558 29766 50610 29818
rect 50610 29766 50612 29818
rect 50556 29764 50612 29766
rect 50660 29818 50716 29820
rect 50660 29766 50662 29818
rect 50662 29766 50714 29818
rect 50714 29766 50716 29818
rect 50660 29764 50716 29766
rect 50764 29818 50820 29820
rect 50764 29766 50766 29818
rect 50766 29766 50818 29818
rect 50818 29766 50820 29818
rect 50764 29764 50820 29766
rect 50556 28250 50612 28252
rect 50556 28198 50558 28250
rect 50558 28198 50610 28250
rect 50610 28198 50612 28250
rect 50556 28196 50612 28198
rect 50660 28250 50716 28252
rect 50660 28198 50662 28250
rect 50662 28198 50714 28250
rect 50714 28198 50716 28250
rect 50660 28196 50716 28198
rect 50764 28250 50820 28252
rect 50764 28198 50766 28250
rect 50766 28198 50818 28250
rect 50818 28198 50820 28250
rect 50764 28196 50820 28198
rect 50876 27356 50932 27412
rect 50652 26962 50708 26964
rect 50652 26910 50654 26962
rect 50654 26910 50706 26962
rect 50706 26910 50708 26962
rect 50652 26908 50708 26910
rect 50556 26682 50612 26684
rect 50556 26630 50558 26682
rect 50558 26630 50610 26682
rect 50610 26630 50612 26682
rect 50556 26628 50612 26630
rect 50660 26682 50716 26684
rect 50660 26630 50662 26682
rect 50662 26630 50714 26682
rect 50714 26630 50716 26682
rect 50660 26628 50716 26630
rect 50764 26682 50820 26684
rect 50764 26630 50766 26682
rect 50766 26630 50818 26682
rect 50818 26630 50820 26682
rect 50764 26628 50820 26630
rect 50428 26460 50484 26516
rect 50556 25114 50612 25116
rect 50556 25062 50558 25114
rect 50558 25062 50610 25114
rect 50610 25062 50612 25114
rect 50556 25060 50612 25062
rect 50660 25114 50716 25116
rect 50660 25062 50662 25114
rect 50662 25062 50714 25114
rect 50714 25062 50716 25114
rect 50660 25060 50716 25062
rect 50764 25114 50820 25116
rect 50764 25062 50766 25114
rect 50766 25062 50818 25114
rect 50818 25062 50820 25114
rect 50764 25060 50820 25062
rect 50556 23546 50612 23548
rect 50556 23494 50558 23546
rect 50558 23494 50610 23546
rect 50610 23494 50612 23546
rect 50556 23492 50612 23494
rect 50660 23546 50716 23548
rect 50660 23494 50662 23546
rect 50662 23494 50714 23546
rect 50714 23494 50716 23546
rect 50660 23492 50716 23494
rect 50764 23546 50820 23548
rect 50764 23494 50766 23546
rect 50766 23494 50818 23546
rect 50818 23494 50820 23546
rect 50764 23492 50820 23494
rect 50988 23436 51044 23492
rect 50764 23378 50820 23380
rect 50764 23326 50766 23378
rect 50766 23326 50818 23378
rect 50818 23326 50820 23378
rect 50764 23324 50820 23326
rect 50556 21978 50612 21980
rect 50556 21926 50558 21978
rect 50558 21926 50610 21978
rect 50610 21926 50612 21978
rect 50556 21924 50612 21926
rect 50660 21978 50716 21980
rect 50660 21926 50662 21978
rect 50662 21926 50714 21978
rect 50714 21926 50716 21978
rect 50660 21924 50716 21926
rect 50764 21978 50820 21980
rect 50764 21926 50766 21978
rect 50766 21926 50818 21978
rect 50818 21926 50820 21978
rect 50764 21924 50820 21926
rect 49980 20690 50036 20692
rect 49980 20638 49982 20690
rect 49982 20638 50034 20690
rect 50034 20638 50036 20690
rect 49980 20636 50036 20638
rect 48300 15036 48356 15092
rect 48748 14530 48804 14532
rect 48748 14478 48750 14530
rect 48750 14478 48802 14530
rect 48802 14478 48804 14530
rect 48748 14476 48804 14478
rect 47964 9548 48020 9604
rect 49420 14812 49476 14868
rect 49420 14140 49476 14196
rect 48412 9100 48468 9156
rect 48860 11788 48916 11844
rect 47292 6412 47348 6468
rect 47516 5852 47572 5908
rect 47180 4508 47236 4564
rect 47404 4620 47460 4676
rect 46620 4172 46676 4228
rect 47964 6130 48020 6132
rect 47964 6078 47966 6130
rect 47966 6078 48018 6130
rect 48018 6078 48020 6130
rect 47964 6076 48020 6078
rect 48636 6076 48692 6132
rect 47628 5516 47684 5572
rect 48076 5404 48132 5460
rect 47964 5180 48020 5236
rect 49532 7980 49588 8036
rect 48860 5964 48916 6020
rect 48748 5180 48804 5236
rect 48188 5068 48244 5124
rect 48972 5068 49028 5124
rect 49196 5292 49252 5348
rect 48748 4562 48804 4564
rect 48748 4510 48750 4562
rect 48750 4510 48802 4562
rect 48802 4510 48804 4562
rect 48748 4508 48804 4510
rect 48524 4284 48580 4340
rect 48972 4172 49028 4228
rect 49084 4338 49140 4340
rect 49084 4286 49086 4338
rect 49086 4286 49138 4338
rect 49138 4286 49140 4338
rect 49084 4284 49140 4286
rect 48860 4060 48916 4116
rect 48748 3836 48804 3892
rect 50204 21756 50260 21812
rect 50204 21308 50260 21364
rect 50316 20802 50372 20804
rect 50316 20750 50318 20802
rect 50318 20750 50370 20802
rect 50370 20750 50372 20802
rect 50316 20748 50372 20750
rect 50764 21308 50820 21364
rect 51660 38780 51716 38836
rect 51324 38668 51380 38724
rect 51212 30098 51268 30100
rect 51212 30046 51214 30098
rect 51214 30046 51266 30098
rect 51266 30046 51268 30098
rect 51212 30044 51268 30046
rect 51436 31778 51492 31780
rect 51436 31726 51438 31778
rect 51438 31726 51490 31778
rect 51490 31726 51492 31778
rect 51436 31724 51492 31726
rect 51548 31666 51604 31668
rect 51548 31614 51550 31666
rect 51550 31614 51602 31666
rect 51602 31614 51604 31666
rect 51548 31612 51604 31614
rect 51436 30828 51492 30884
rect 50652 20636 50708 20692
rect 50204 19516 50260 19572
rect 50556 20410 50612 20412
rect 50556 20358 50558 20410
rect 50558 20358 50610 20410
rect 50610 20358 50612 20410
rect 50556 20356 50612 20358
rect 50660 20410 50716 20412
rect 50660 20358 50662 20410
rect 50662 20358 50714 20410
rect 50714 20358 50716 20410
rect 50660 20356 50716 20358
rect 50764 20410 50820 20412
rect 50764 20358 50766 20410
rect 50766 20358 50818 20410
rect 50818 20358 50820 20410
rect 50764 20356 50820 20358
rect 50988 20690 51044 20692
rect 50988 20638 50990 20690
rect 50990 20638 51042 20690
rect 51042 20638 51044 20690
rect 50988 20636 51044 20638
rect 51100 20130 51156 20132
rect 51100 20078 51102 20130
rect 51102 20078 51154 20130
rect 51154 20078 51156 20130
rect 51100 20076 51156 20078
rect 50876 19852 50932 19908
rect 50428 19180 50484 19236
rect 50556 18842 50612 18844
rect 50556 18790 50558 18842
rect 50558 18790 50610 18842
rect 50610 18790 50612 18842
rect 50556 18788 50612 18790
rect 50660 18842 50716 18844
rect 50660 18790 50662 18842
rect 50662 18790 50714 18842
rect 50714 18790 50716 18842
rect 50660 18788 50716 18790
rect 50764 18842 50820 18844
rect 50764 18790 50766 18842
rect 50766 18790 50818 18842
rect 50818 18790 50820 18842
rect 50764 18788 50820 18790
rect 50988 18508 51044 18564
rect 50876 17388 50932 17444
rect 50556 17274 50612 17276
rect 50556 17222 50558 17274
rect 50558 17222 50610 17274
rect 50610 17222 50612 17274
rect 50556 17220 50612 17222
rect 50660 17274 50716 17276
rect 50660 17222 50662 17274
rect 50662 17222 50714 17274
rect 50714 17222 50716 17274
rect 50660 17220 50716 17222
rect 50764 17274 50820 17276
rect 50764 17222 50766 17274
rect 50766 17222 50818 17274
rect 50818 17222 50820 17274
rect 50764 17220 50820 17222
rect 49868 13356 49924 13412
rect 49756 7980 49812 8036
rect 50988 17052 51044 17108
rect 50316 15708 50372 15764
rect 50092 14642 50148 14644
rect 50092 14590 50094 14642
rect 50094 14590 50146 14642
rect 50146 14590 50148 14642
rect 50092 14588 50148 14590
rect 50316 14588 50372 14644
rect 50556 15706 50612 15708
rect 50556 15654 50558 15706
rect 50558 15654 50610 15706
rect 50610 15654 50612 15706
rect 50556 15652 50612 15654
rect 50660 15706 50716 15708
rect 50660 15654 50662 15706
rect 50662 15654 50714 15706
rect 50714 15654 50716 15706
rect 50660 15652 50716 15654
rect 50764 15706 50820 15708
rect 50764 15654 50766 15706
rect 50766 15654 50818 15706
rect 50818 15654 50820 15706
rect 50764 15652 50820 15654
rect 50652 15426 50708 15428
rect 50652 15374 50654 15426
rect 50654 15374 50706 15426
rect 50706 15374 50708 15426
rect 50652 15372 50708 15374
rect 50876 15036 50932 15092
rect 51436 22652 51492 22708
rect 51548 23436 51604 23492
rect 51548 21756 51604 21812
rect 51324 20076 51380 20132
rect 52332 34524 52388 34580
rect 51772 30268 51828 30324
rect 51772 22540 51828 22596
rect 52556 31948 52612 32004
rect 52444 30380 52500 30436
rect 51996 30098 52052 30100
rect 51996 30046 51998 30098
rect 51998 30046 52050 30098
rect 52050 30046 52052 30098
rect 51996 30044 52052 30046
rect 51884 21586 51940 21588
rect 51884 21534 51886 21586
rect 51886 21534 51938 21586
rect 51938 21534 51940 21586
rect 51884 21532 51940 21534
rect 51884 20972 51940 21028
rect 51436 16044 51492 16100
rect 51772 20018 51828 20020
rect 51772 19966 51774 20018
rect 51774 19966 51826 20018
rect 51826 19966 51828 20018
rect 51772 19964 51828 19966
rect 51436 15874 51492 15876
rect 51436 15822 51438 15874
rect 51438 15822 51490 15874
rect 51490 15822 51492 15874
rect 51436 15820 51492 15822
rect 51324 14812 51380 14868
rect 50428 14476 50484 14532
rect 51324 14530 51380 14532
rect 51324 14478 51326 14530
rect 51326 14478 51378 14530
rect 51378 14478 51380 14530
rect 51324 14476 51380 14478
rect 50316 14028 50372 14084
rect 50556 14138 50612 14140
rect 50556 14086 50558 14138
rect 50558 14086 50610 14138
rect 50610 14086 50612 14138
rect 50556 14084 50612 14086
rect 50660 14138 50716 14140
rect 50660 14086 50662 14138
rect 50662 14086 50714 14138
rect 50714 14086 50716 14138
rect 50660 14084 50716 14086
rect 50764 14138 50820 14140
rect 50764 14086 50766 14138
rect 50766 14086 50818 14138
rect 50818 14086 50820 14138
rect 50764 14084 50820 14086
rect 50556 12570 50612 12572
rect 50556 12518 50558 12570
rect 50558 12518 50610 12570
rect 50610 12518 50612 12570
rect 50556 12516 50612 12518
rect 50660 12570 50716 12572
rect 50660 12518 50662 12570
rect 50662 12518 50714 12570
rect 50714 12518 50716 12570
rect 50660 12516 50716 12518
rect 50764 12570 50820 12572
rect 50764 12518 50766 12570
rect 50766 12518 50818 12570
rect 50818 12518 50820 12570
rect 50764 12516 50820 12518
rect 50556 11002 50612 11004
rect 50556 10950 50558 11002
rect 50558 10950 50610 11002
rect 50610 10950 50612 11002
rect 50556 10948 50612 10950
rect 50660 11002 50716 11004
rect 50660 10950 50662 11002
rect 50662 10950 50714 11002
rect 50714 10950 50716 11002
rect 50660 10948 50716 10950
rect 50764 11002 50820 11004
rect 50764 10950 50766 11002
rect 50766 10950 50818 11002
rect 50818 10950 50820 11002
rect 50764 10948 50820 10950
rect 50556 9434 50612 9436
rect 50556 9382 50558 9434
rect 50558 9382 50610 9434
rect 50610 9382 50612 9434
rect 50556 9380 50612 9382
rect 50660 9434 50716 9436
rect 50660 9382 50662 9434
rect 50662 9382 50714 9434
rect 50714 9382 50716 9434
rect 50660 9380 50716 9382
rect 50764 9434 50820 9436
rect 50764 9382 50766 9434
rect 50766 9382 50818 9434
rect 50818 9382 50820 9434
rect 50764 9380 50820 9382
rect 50988 8428 51044 8484
rect 50556 7866 50612 7868
rect 50556 7814 50558 7866
rect 50558 7814 50610 7866
rect 50610 7814 50612 7866
rect 50556 7812 50612 7814
rect 50660 7866 50716 7868
rect 50660 7814 50662 7866
rect 50662 7814 50714 7866
rect 50714 7814 50716 7866
rect 50660 7812 50716 7814
rect 50764 7866 50820 7868
rect 50764 7814 50766 7866
rect 50766 7814 50818 7866
rect 50818 7814 50820 7866
rect 50764 7812 50820 7814
rect 49980 7532 50036 7588
rect 49980 6690 50036 6692
rect 49980 6638 49982 6690
rect 49982 6638 50034 6690
rect 50034 6638 50036 6690
rect 49980 6636 50036 6638
rect 49644 6130 49700 6132
rect 49644 6078 49646 6130
rect 49646 6078 49698 6130
rect 49698 6078 49700 6130
rect 49644 6076 49700 6078
rect 51324 13746 51380 13748
rect 51324 13694 51326 13746
rect 51326 13694 51378 13746
rect 51378 13694 51380 13746
rect 51324 13692 51380 13694
rect 51772 19180 51828 19236
rect 51772 17388 51828 17444
rect 52332 30268 52388 30324
rect 52780 35980 52836 36036
rect 53004 34130 53060 34132
rect 53004 34078 53006 34130
rect 53006 34078 53058 34130
rect 53058 34078 53060 34130
rect 53004 34076 53060 34078
rect 52780 31612 52836 31668
rect 53004 33740 53060 33796
rect 52892 30882 52948 30884
rect 52892 30830 52894 30882
rect 52894 30830 52946 30882
rect 52946 30830 52948 30882
rect 52892 30828 52948 30830
rect 52892 30322 52948 30324
rect 52892 30270 52894 30322
rect 52894 30270 52946 30322
rect 52946 30270 52948 30322
rect 52892 30268 52948 30270
rect 52780 23436 52836 23492
rect 52556 22652 52612 22708
rect 52108 20018 52164 20020
rect 52108 19966 52110 20018
rect 52110 19966 52162 20018
rect 52162 19966 52164 20018
rect 52108 19964 52164 19966
rect 52108 19740 52164 19796
rect 51884 16828 51940 16884
rect 51996 19180 52052 19236
rect 51996 15260 52052 15316
rect 51660 15202 51716 15204
rect 51660 15150 51662 15202
rect 51662 15150 51714 15202
rect 51714 15150 51716 15202
rect 51660 15148 51716 15150
rect 52444 19964 52500 20020
rect 52444 19740 52500 19796
rect 52668 21532 52724 21588
rect 52780 21308 52836 21364
rect 52780 20578 52836 20580
rect 52780 20526 52782 20578
rect 52782 20526 52834 20578
rect 52834 20526 52836 20578
rect 52780 20524 52836 20526
rect 52892 20018 52948 20020
rect 52892 19966 52894 20018
rect 52894 19966 52946 20018
rect 52946 19966 52948 20018
rect 52892 19964 52948 19966
rect 52668 19234 52724 19236
rect 52668 19182 52670 19234
rect 52670 19182 52722 19234
rect 52722 19182 52724 19234
rect 52668 19180 52724 19182
rect 52556 18172 52612 18228
rect 52780 17388 52836 17444
rect 52668 16882 52724 16884
rect 52668 16830 52670 16882
rect 52670 16830 52722 16882
rect 52722 16830 52724 16882
rect 52668 16828 52724 16830
rect 52668 16098 52724 16100
rect 52668 16046 52670 16098
rect 52670 16046 52722 16098
rect 52722 16046 52724 16098
rect 52668 16044 52724 16046
rect 52668 14530 52724 14532
rect 52668 14478 52670 14530
rect 52670 14478 52722 14530
rect 52722 14478 52724 14530
rect 52668 14476 52724 14478
rect 53340 34242 53396 34244
rect 53340 34190 53342 34242
rect 53342 34190 53394 34242
rect 53394 34190 53396 34242
rect 53340 34188 53396 34190
rect 53788 40796 53844 40852
rect 53788 38668 53844 38724
rect 53788 36092 53844 36148
rect 53564 34914 53620 34916
rect 53564 34862 53566 34914
rect 53566 34862 53618 34914
rect 53618 34862 53620 34914
rect 53564 34860 53620 34862
rect 53788 34188 53844 34244
rect 53564 33740 53620 33796
rect 53676 32732 53732 32788
rect 53676 31948 53732 32004
rect 53340 30828 53396 30884
rect 53340 21586 53396 21588
rect 53340 21534 53342 21586
rect 53342 21534 53394 21586
rect 53394 21534 53396 21586
rect 53340 21532 53396 21534
rect 53228 20130 53284 20132
rect 53228 20078 53230 20130
rect 53230 20078 53282 20130
rect 53282 20078 53284 20130
rect 53228 20076 53284 20078
rect 53564 20300 53620 20356
rect 53228 18562 53284 18564
rect 53228 18510 53230 18562
rect 53230 18510 53282 18562
rect 53282 18510 53284 18562
rect 53228 18508 53284 18510
rect 53452 20076 53508 20132
rect 53788 23436 53844 23492
rect 53788 21810 53844 21812
rect 53788 21758 53790 21810
rect 53790 21758 53842 21810
rect 53842 21758 53844 21810
rect 53788 21756 53844 21758
rect 55132 76690 55188 76692
rect 55132 76638 55134 76690
rect 55134 76638 55186 76690
rect 55186 76638 55188 76690
rect 55132 76636 55188 76638
rect 54012 34188 54068 34244
rect 55692 76300 55748 76356
rect 56924 76636 56980 76692
rect 57484 76412 57540 76468
rect 54348 39004 54404 39060
rect 54908 41858 54964 41860
rect 54908 41806 54910 41858
rect 54910 41806 54962 41858
rect 54962 41806 54964 41858
rect 54908 41804 54964 41806
rect 55020 40796 55076 40852
rect 55356 41356 55412 41412
rect 55356 40796 55412 40852
rect 55132 40684 55188 40740
rect 55580 41410 55636 41412
rect 55580 41358 55582 41410
rect 55582 41358 55634 41410
rect 55634 41358 55636 41410
rect 55580 41356 55636 41358
rect 54460 35532 54516 35588
rect 54236 35308 54292 35364
rect 54796 34860 54852 34916
rect 54572 34300 54628 34356
rect 54012 20802 54068 20804
rect 54012 20750 54014 20802
rect 54014 20750 54066 20802
rect 54066 20750 54068 20802
rect 54012 20748 54068 20750
rect 53340 18284 53396 18340
rect 53452 17612 53508 17668
rect 53452 17276 53508 17332
rect 52780 14364 52836 14420
rect 51884 9548 51940 9604
rect 50540 6578 50596 6580
rect 50540 6526 50542 6578
rect 50542 6526 50594 6578
rect 50594 6526 50596 6578
rect 50540 6524 50596 6526
rect 51772 9212 51828 9268
rect 51436 6690 51492 6692
rect 51436 6638 51438 6690
rect 51438 6638 51490 6690
rect 51490 6638 51492 6690
rect 51436 6636 51492 6638
rect 51324 6524 51380 6580
rect 50556 6298 50612 6300
rect 50556 6246 50558 6298
rect 50558 6246 50610 6298
rect 50610 6246 50612 6298
rect 50556 6244 50612 6246
rect 50660 6298 50716 6300
rect 50660 6246 50662 6298
rect 50662 6246 50714 6298
rect 50714 6246 50716 6298
rect 50660 6244 50716 6246
rect 50764 6298 50820 6300
rect 50764 6246 50766 6298
rect 50766 6246 50818 6298
rect 50818 6246 50820 6298
rect 50764 6244 50820 6246
rect 49980 6076 50036 6132
rect 50764 6130 50820 6132
rect 50764 6078 50766 6130
rect 50766 6078 50818 6130
rect 50818 6078 50820 6130
rect 50764 6076 50820 6078
rect 49868 5906 49924 5908
rect 49868 5854 49870 5906
rect 49870 5854 49922 5906
rect 49922 5854 49924 5906
rect 49868 5852 49924 5854
rect 50092 5740 50148 5796
rect 49756 5292 49812 5348
rect 50540 5292 50596 5348
rect 51212 5292 51268 5348
rect 48972 3948 49028 4004
rect 49308 4060 49364 4116
rect 49420 3724 49476 3780
rect 49532 3500 49588 3556
rect 49868 4844 49924 4900
rect 50556 4730 50612 4732
rect 50556 4678 50558 4730
rect 50558 4678 50610 4730
rect 50610 4678 50612 4730
rect 50556 4676 50612 4678
rect 50660 4730 50716 4732
rect 50660 4678 50662 4730
rect 50662 4678 50714 4730
rect 50714 4678 50716 4730
rect 50660 4676 50716 4678
rect 50764 4730 50820 4732
rect 50764 4678 50766 4730
rect 50766 4678 50818 4730
rect 50818 4678 50820 4730
rect 50764 4676 50820 4678
rect 50540 4114 50596 4116
rect 50540 4062 50542 4114
rect 50542 4062 50594 4114
rect 50594 4062 50596 4114
rect 50540 4060 50596 4062
rect 50092 3948 50148 4004
rect 51100 3836 51156 3892
rect 51548 3724 51604 3780
rect 50092 3612 50148 3668
rect 50652 3666 50708 3668
rect 50652 3614 50654 3666
rect 50654 3614 50706 3666
rect 50706 3614 50708 3666
rect 50652 3612 50708 3614
rect 51324 3612 51380 3668
rect 50876 3500 50932 3556
rect 49980 3388 50036 3444
rect 50556 3162 50612 3164
rect 50556 3110 50558 3162
rect 50558 3110 50610 3162
rect 50610 3110 50612 3162
rect 50556 3108 50612 3110
rect 50660 3162 50716 3164
rect 50660 3110 50662 3162
rect 50662 3110 50714 3162
rect 50714 3110 50716 3162
rect 50660 3108 50716 3110
rect 50764 3162 50820 3164
rect 50764 3110 50766 3162
rect 50766 3110 50818 3162
rect 50818 3110 50820 3162
rect 50764 3108 50820 3110
rect 51212 3442 51268 3444
rect 51212 3390 51214 3442
rect 51214 3390 51266 3442
rect 51266 3390 51268 3442
rect 51212 3388 51268 3390
rect 51884 8428 51940 8484
rect 51660 3388 51716 3444
rect 51884 3388 51940 3444
rect 51996 3724 52052 3780
rect 54236 20076 54292 20132
rect 54348 21532 54404 21588
rect 54348 20690 54404 20692
rect 54348 20638 54350 20690
rect 54350 20638 54402 20690
rect 54402 20638 54404 20690
rect 54348 20636 54404 20638
rect 55580 35026 55636 35028
rect 55580 34974 55582 35026
rect 55582 34974 55634 35026
rect 55634 34974 55636 35026
rect 55580 34972 55636 34974
rect 55468 34354 55524 34356
rect 55468 34302 55470 34354
rect 55470 34302 55522 34354
rect 55522 34302 55524 34354
rect 55468 34300 55524 34302
rect 54908 21756 54964 21812
rect 55132 20860 55188 20916
rect 55020 20690 55076 20692
rect 55020 20638 55022 20690
rect 55022 20638 55074 20690
rect 55074 20638 55076 20690
rect 55020 20636 55076 20638
rect 54124 18508 54180 18564
rect 54012 17612 54068 17668
rect 53676 15148 53732 15204
rect 52556 10780 52612 10836
rect 52332 6076 52388 6132
rect 52220 4172 52276 4228
rect 52332 3554 52388 3556
rect 52332 3502 52334 3554
rect 52334 3502 52386 3554
rect 52386 3502 52388 3554
rect 52332 3500 52388 3502
rect 53676 9324 53732 9380
rect 53452 7308 53508 7364
rect 52556 4338 52612 4340
rect 52556 4286 52558 4338
rect 52558 4286 52610 4338
rect 52610 4286 52612 4338
rect 52556 4284 52612 4286
rect 52668 4060 52724 4116
rect 53228 3724 53284 3780
rect 53004 3612 53060 3668
rect 53340 3612 53396 3668
rect 52780 3442 52836 3444
rect 52780 3390 52782 3442
rect 52782 3390 52834 3442
rect 52834 3390 52836 3442
rect 52780 3388 52836 3390
rect 53900 11564 53956 11620
rect 54572 16380 54628 16436
rect 54908 18450 54964 18452
rect 54908 18398 54910 18450
rect 54910 18398 54962 18450
rect 54962 18398 54964 18450
rect 54908 18396 54964 18398
rect 54684 15820 54740 15876
rect 54236 15314 54292 15316
rect 54236 15262 54238 15314
rect 54238 15262 54290 15314
rect 54290 15262 54292 15314
rect 54236 15260 54292 15262
rect 54460 14700 54516 14756
rect 54796 13804 54852 13860
rect 55132 18562 55188 18564
rect 55132 18510 55134 18562
rect 55134 18510 55186 18562
rect 55186 18510 55188 18562
rect 55132 18508 55188 18510
rect 56924 73164 56980 73220
rect 56028 45276 56084 45332
rect 58716 76748 58772 76804
rect 58156 75516 58212 75572
rect 57036 43426 57092 43428
rect 57036 43374 57038 43426
rect 57038 43374 57090 43426
rect 57090 43374 57092 43426
rect 57036 43372 57092 43374
rect 58492 45276 58548 45332
rect 58156 42866 58212 42868
rect 58156 42814 58158 42866
rect 58158 42814 58210 42866
rect 58210 42814 58212 42866
rect 58156 42812 58212 42814
rect 56364 41692 56420 41748
rect 56924 41356 56980 41412
rect 56364 38780 56420 38836
rect 57148 41692 57204 41748
rect 57820 41356 57876 41412
rect 57148 40962 57204 40964
rect 57148 40910 57150 40962
rect 57150 40910 57202 40962
rect 57202 40910 57204 40962
rect 57148 40908 57204 40910
rect 58492 41186 58548 41188
rect 58492 41134 58494 41186
rect 58494 41134 58546 41186
rect 58546 41134 58548 41186
rect 58492 41132 58548 41134
rect 58268 40908 58324 40964
rect 57148 40572 57204 40628
rect 58828 76466 58884 76468
rect 58828 76414 58830 76466
rect 58830 76414 58882 76466
rect 58882 76414 58884 76466
rect 58828 76412 58884 76414
rect 59836 76690 59892 76692
rect 59836 76638 59838 76690
rect 59838 76638 59890 76690
rect 59890 76638 59892 76690
rect 59836 76636 59892 76638
rect 59612 76412 59668 76468
rect 58940 75404 58996 75460
rect 59388 75570 59444 75572
rect 59388 75518 59390 75570
rect 59390 75518 59442 75570
rect 59442 75518 59444 75570
rect 59388 75516 59444 75518
rect 61628 76972 61684 77028
rect 60284 75516 60340 75572
rect 61180 75570 61236 75572
rect 61180 75518 61182 75570
rect 61182 75518 61234 75570
rect 61234 75518 61236 75570
rect 61180 75516 61236 75518
rect 59612 70532 59668 70588
rect 60508 75458 60564 75460
rect 60508 75406 60510 75458
rect 60510 75406 60562 75458
rect 60562 75406 60564 75458
rect 60508 75404 60564 75406
rect 61292 75404 61348 75460
rect 59836 70588 59892 70644
rect 60844 74620 60900 74676
rect 59500 43372 59556 43428
rect 60396 55020 60452 55076
rect 59948 42812 60004 42868
rect 59164 41916 59220 41972
rect 58716 37660 58772 37716
rect 57036 37548 57092 37604
rect 57036 36540 57092 36596
rect 59388 41186 59444 41188
rect 59388 41134 59390 41186
rect 59390 41134 59442 41186
rect 59442 41134 59444 41186
rect 59388 41132 59444 41134
rect 57036 34300 57092 34356
rect 59612 40124 59668 40180
rect 58604 26124 58660 26180
rect 56812 23772 56868 23828
rect 55804 21756 55860 21812
rect 55468 20300 55524 20356
rect 55356 19516 55412 19572
rect 56476 20802 56532 20804
rect 56476 20750 56478 20802
rect 56478 20750 56530 20802
rect 56530 20750 56532 20802
rect 56476 20748 56532 20750
rect 56924 20914 56980 20916
rect 56924 20862 56926 20914
rect 56926 20862 56978 20914
rect 56978 20862 56980 20914
rect 56924 20860 56980 20862
rect 56700 20018 56756 20020
rect 56700 19966 56702 20018
rect 56702 19966 56754 20018
rect 56754 19966 56756 20018
rect 56700 19964 56756 19966
rect 56028 19906 56084 19908
rect 56028 19854 56030 19906
rect 56030 19854 56082 19906
rect 56082 19854 56084 19906
rect 56028 19852 56084 19854
rect 56588 19516 56644 19572
rect 56364 18844 56420 18900
rect 56140 18508 56196 18564
rect 55916 18172 55972 18228
rect 55244 17612 55300 17668
rect 55132 17276 55188 17332
rect 56700 18450 56756 18452
rect 56700 18398 56702 18450
rect 56702 18398 56754 18450
rect 56754 18398 56756 18450
rect 56700 18396 56756 18398
rect 56812 17666 56868 17668
rect 56812 17614 56814 17666
rect 56814 17614 56866 17666
rect 56866 17614 56868 17666
rect 56812 17612 56868 17614
rect 55244 15202 55300 15204
rect 55244 15150 55246 15202
rect 55246 15150 55298 15202
rect 55298 15150 55300 15202
rect 55244 15148 55300 15150
rect 54908 11116 54964 11172
rect 55020 11452 55076 11508
rect 53788 4508 53844 4564
rect 54012 5180 54068 5236
rect 53900 4114 53956 4116
rect 53900 4062 53902 4114
rect 53902 4062 53954 4114
rect 53954 4062 53956 4114
rect 53900 4060 53956 4062
rect 53564 3948 53620 4004
rect 53676 3724 53732 3780
rect 54348 5740 54404 5796
rect 55244 7756 55300 7812
rect 55468 14588 55524 14644
rect 56588 11676 56644 11732
rect 56028 6412 56084 6468
rect 55356 5852 55412 5908
rect 55244 5234 55300 5236
rect 55244 5182 55246 5234
rect 55246 5182 55298 5234
rect 55298 5182 55300 5234
rect 55244 5180 55300 5182
rect 56140 5180 56196 5236
rect 55020 4956 55076 5012
rect 54236 3554 54292 3556
rect 54236 3502 54238 3554
rect 54238 3502 54290 3554
rect 54290 3502 54292 3554
rect 54236 3500 54292 3502
rect 55916 4956 55972 5012
rect 56028 3666 56084 3668
rect 56028 3614 56030 3666
rect 56030 3614 56082 3666
rect 56082 3614 56084 3666
rect 56028 3612 56084 3614
rect 55356 3500 55412 3556
rect 54684 3388 54740 3444
rect 57260 20412 57316 20468
rect 57596 20130 57652 20132
rect 57596 20078 57598 20130
rect 57598 20078 57650 20130
rect 57650 20078 57652 20130
rect 57596 20076 57652 20078
rect 57260 19628 57316 19684
rect 58828 18396 58884 18452
rect 57148 18338 57204 18340
rect 57148 18286 57150 18338
rect 57150 18286 57202 18338
rect 57202 18286 57204 18338
rect 57148 18284 57204 18286
rect 57036 9660 57092 9716
rect 57148 17612 57204 17668
rect 58716 17666 58772 17668
rect 58716 17614 58718 17666
rect 58718 17614 58770 17666
rect 58770 17614 58772 17666
rect 58716 17612 58772 17614
rect 57148 8876 57204 8932
rect 57708 7644 57764 7700
rect 58156 13356 58212 13412
rect 56588 4338 56644 4340
rect 56588 4286 56590 4338
rect 56590 4286 56642 4338
rect 56642 4286 56644 4338
rect 56588 4284 56644 4286
rect 56700 5628 56756 5684
rect 56924 6412 56980 6468
rect 59500 12796 59556 12852
rect 60172 41132 60228 41188
rect 60060 40402 60116 40404
rect 60060 40350 60062 40402
rect 60062 40350 60114 40402
rect 60114 40350 60116 40402
rect 60060 40348 60116 40350
rect 60620 41804 60676 41860
rect 60508 41186 60564 41188
rect 60508 41134 60510 41186
rect 60510 41134 60562 41186
rect 60562 41134 60564 41186
rect 60508 41132 60564 41134
rect 62972 77084 63028 77140
rect 62636 76972 62692 77028
rect 63644 76972 63700 77028
rect 63980 77084 64036 77140
rect 62076 76466 62132 76468
rect 62076 76414 62078 76466
rect 62078 76414 62130 76466
rect 62130 76414 62132 76466
rect 62076 76412 62132 76414
rect 61740 75516 61796 75572
rect 61628 74620 61684 74676
rect 64652 76972 64708 77028
rect 64316 76188 64372 76244
rect 63756 74956 63812 75012
rect 61068 41970 61124 41972
rect 61068 41918 61070 41970
rect 61070 41918 61122 41970
rect 61122 41918 61124 41970
rect 61068 41916 61124 41918
rect 61628 41970 61684 41972
rect 61628 41918 61630 41970
rect 61630 41918 61682 41970
rect 61682 41918 61684 41970
rect 61628 41916 61684 41918
rect 61628 41186 61684 41188
rect 61628 41134 61630 41186
rect 61630 41134 61682 41186
rect 61682 41134 61684 41186
rect 61628 41132 61684 41134
rect 61628 40348 61684 40404
rect 62300 40236 62356 40292
rect 62524 41020 62580 41076
rect 62860 41186 62916 41188
rect 62860 41134 62862 41186
rect 62862 41134 62914 41186
rect 62914 41134 62916 41186
rect 62860 41132 62916 41134
rect 62860 40908 62916 40964
rect 67004 76972 67060 77028
rect 65324 75740 65380 75796
rect 65548 75458 65604 75460
rect 65548 75406 65550 75458
rect 65550 75406 65602 75458
rect 65602 75406 65604 75458
rect 65548 75404 65604 75406
rect 63756 43484 63812 43540
rect 64540 55916 64596 55972
rect 64428 41970 64484 41972
rect 64428 41918 64430 41970
rect 64430 41918 64482 41970
rect 64482 41918 64484 41970
rect 64428 41916 64484 41918
rect 64428 41356 64484 41412
rect 63532 41244 63588 41300
rect 63308 41132 63364 41188
rect 63420 41020 63476 41076
rect 64316 41186 64372 41188
rect 64316 41134 64318 41186
rect 64318 41134 64370 41186
rect 64370 41134 64372 41186
rect 64316 41132 64372 41134
rect 62412 39788 62468 39844
rect 61852 38946 61908 38948
rect 61852 38894 61854 38946
rect 61854 38894 61906 38946
rect 61906 38894 61908 38946
rect 61852 38892 61908 38894
rect 62524 38834 62580 38836
rect 62524 38782 62526 38834
rect 62526 38782 62578 38834
rect 62578 38782 62580 38834
rect 62524 38780 62580 38782
rect 60620 36316 60676 36372
rect 61740 36204 61796 36260
rect 60284 28700 60340 28756
rect 60396 31052 60452 31108
rect 60396 27020 60452 27076
rect 60172 23996 60228 24052
rect 61628 21196 61684 21252
rect 60172 9996 60228 10052
rect 59612 9548 59668 9604
rect 60060 9884 60116 9940
rect 58156 6188 58212 6244
rect 60060 6412 60116 6468
rect 57932 5682 57988 5684
rect 57932 5630 57934 5682
rect 57934 5630 57986 5682
rect 57986 5630 57988 5682
rect 57932 5628 57988 5630
rect 59388 5628 59444 5684
rect 58156 5234 58212 5236
rect 58156 5182 58158 5234
rect 58158 5182 58210 5234
rect 58210 5182 58212 5234
rect 58156 5180 58212 5182
rect 58716 4844 58772 4900
rect 58044 4284 58100 4340
rect 57372 4060 57428 4116
rect 57596 3388 57652 3444
rect 58044 3388 58100 3444
rect 59052 3666 59108 3668
rect 59052 3614 59054 3666
rect 59054 3614 59106 3666
rect 59106 3614 59108 3666
rect 59052 3612 59108 3614
rect 59724 4114 59780 4116
rect 59724 4062 59726 4114
rect 59726 4062 59778 4114
rect 59778 4062 59780 4114
rect 59724 4060 59780 4062
rect 61516 6466 61572 6468
rect 61516 6414 61518 6466
rect 61518 6414 61570 6466
rect 61570 6414 61572 6466
rect 61516 6412 61572 6414
rect 60844 5682 60900 5684
rect 60844 5630 60846 5682
rect 60846 5630 60898 5682
rect 60898 5630 60900 5682
rect 60844 5628 60900 5630
rect 60732 5180 60788 5236
rect 61516 4898 61572 4900
rect 61516 4846 61518 4898
rect 61518 4846 61570 4898
rect 61570 4846 61572 4898
rect 61516 4844 61572 4846
rect 62076 33180 62132 33236
rect 62076 30044 62132 30100
rect 62860 39788 62916 39844
rect 63196 40402 63252 40404
rect 63196 40350 63198 40402
rect 63198 40350 63250 40402
rect 63250 40350 63252 40402
rect 63196 40348 63252 40350
rect 64204 40572 64260 40628
rect 63532 40348 63588 40404
rect 63756 40236 63812 40292
rect 63868 39004 63924 39060
rect 64204 26460 64260 26516
rect 64652 40626 64708 40628
rect 64652 40574 64654 40626
rect 64654 40574 64706 40626
rect 64706 40574 64708 40626
rect 64652 40572 64708 40574
rect 64652 39004 64708 39060
rect 65100 41916 65156 41972
rect 64988 41468 65044 41524
rect 64988 41298 65044 41300
rect 64988 41246 64990 41298
rect 64990 41246 65042 41298
rect 65042 41246 65044 41298
rect 64988 41244 65044 41246
rect 65916 76074 65972 76076
rect 65916 76022 65918 76074
rect 65918 76022 65970 76074
rect 65970 76022 65972 76074
rect 65916 76020 65972 76022
rect 66020 76074 66076 76076
rect 66020 76022 66022 76074
rect 66022 76022 66074 76074
rect 66074 76022 66076 76074
rect 66020 76020 66076 76022
rect 66124 76074 66180 76076
rect 66124 76022 66126 76074
rect 66126 76022 66178 76074
rect 66178 76022 66180 76074
rect 66124 76020 66180 76022
rect 65996 75794 66052 75796
rect 65996 75742 65998 75794
rect 65998 75742 66050 75794
rect 66050 75742 66052 75794
rect 65996 75740 66052 75742
rect 66108 75404 66164 75460
rect 65916 74506 65972 74508
rect 65916 74454 65918 74506
rect 65918 74454 65970 74506
rect 65970 74454 65972 74506
rect 65916 74452 65972 74454
rect 66020 74506 66076 74508
rect 66020 74454 66022 74506
rect 66022 74454 66074 74506
rect 66074 74454 66076 74506
rect 66020 74452 66076 74454
rect 66124 74506 66180 74508
rect 66124 74454 66126 74506
rect 66126 74454 66178 74506
rect 66178 74454 66180 74506
rect 66124 74452 66180 74454
rect 65916 72938 65972 72940
rect 65916 72886 65918 72938
rect 65918 72886 65970 72938
rect 65970 72886 65972 72938
rect 65916 72884 65972 72886
rect 66020 72938 66076 72940
rect 66020 72886 66022 72938
rect 66022 72886 66074 72938
rect 66074 72886 66076 72938
rect 66020 72884 66076 72886
rect 66124 72938 66180 72940
rect 66124 72886 66126 72938
rect 66126 72886 66178 72938
rect 66178 72886 66180 72938
rect 66124 72884 66180 72886
rect 65916 71370 65972 71372
rect 65916 71318 65918 71370
rect 65918 71318 65970 71370
rect 65970 71318 65972 71370
rect 65916 71316 65972 71318
rect 66020 71370 66076 71372
rect 66020 71318 66022 71370
rect 66022 71318 66074 71370
rect 66074 71318 66076 71370
rect 66020 71316 66076 71318
rect 66124 71370 66180 71372
rect 66124 71318 66126 71370
rect 66126 71318 66178 71370
rect 66178 71318 66180 71370
rect 66124 71316 66180 71318
rect 65916 69802 65972 69804
rect 65916 69750 65918 69802
rect 65918 69750 65970 69802
rect 65970 69750 65972 69802
rect 65916 69748 65972 69750
rect 66020 69802 66076 69804
rect 66020 69750 66022 69802
rect 66022 69750 66074 69802
rect 66074 69750 66076 69802
rect 66020 69748 66076 69750
rect 66124 69802 66180 69804
rect 66124 69750 66126 69802
rect 66126 69750 66178 69802
rect 66178 69750 66180 69802
rect 66124 69748 66180 69750
rect 65916 68234 65972 68236
rect 65916 68182 65918 68234
rect 65918 68182 65970 68234
rect 65970 68182 65972 68234
rect 65916 68180 65972 68182
rect 66020 68234 66076 68236
rect 66020 68182 66022 68234
rect 66022 68182 66074 68234
rect 66074 68182 66076 68234
rect 66020 68180 66076 68182
rect 66124 68234 66180 68236
rect 66124 68182 66126 68234
rect 66126 68182 66178 68234
rect 66178 68182 66180 68234
rect 66124 68180 66180 68182
rect 65916 66666 65972 66668
rect 65916 66614 65918 66666
rect 65918 66614 65970 66666
rect 65970 66614 65972 66666
rect 65916 66612 65972 66614
rect 66020 66666 66076 66668
rect 66020 66614 66022 66666
rect 66022 66614 66074 66666
rect 66074 66614 66076 66666
rect 66020 66612 66076 66614
rect 66124 66666 66180 66668
rect 66124 66614 66126 66666
rect 66126 66614 66178 66666
rect 66178 66614 66180 66666
rect 66124 66612 66180 66614
rect 65916 65098 65972 65100
rect 65916 65046 65918 65098
rect 65918 65046 65970 65098
rect 65970 65046 65972 65098
rect 65916 65044 65972 65046
rect 66020 65098 66076 65100
rect 66020 65046 66022 65098
rect 66022 65046 66074 65098
rect 66074 65046 66076 65098
rect 66020 65044 66076 65046
rect 66124 65098 66180 65100
rect 66124 65046 66126 65098
rect 66126 65046 66178 65098
rect 66178 65046 66180 65098
rect 66124 65044 66180 65046
rect 65916 63530 65972 63532
rect 65916 63478 65918 63530
rect 65918 63478 65970 63530
rect 65970 63478 65972 63530
rect 65916 63476 65972 63478
rect 66020 63530 66076 63532
rect 66020 63478 66022 63530
rect 66022 63478 66074 63530
rect 66074 63478 66076 63530
rect 66020 63476 66076 63478
rect 66124 63530 66180 63532
rect 66124 63478 66126 63530
rect 66126 63478 66178 63530
rect 66178 63478 66180 63530
rect 66124 63476 66180 63478
rect 65916 61962 65972 61964
rect 65916 61910 65918 61962
rect 65918 61910 65970 61962
rect 65970 61910 65972 61962
rect 65916 61908 65972 61910
rect 66020 61962 66076 61964
rect 66020 61910 66022 61962
rect 66022 61910 66074 61962
rect 66074 61910 66076 61962
rect 66020 61908 66076 61910
rect 66124 61962 66180 61964
rect 66124 61910 66126 61962
rect 66126 61910 66178 61962
rect 66178 61910 66180 61962
rect 66124 61908 66180 61910
rect 65916 60394 65972 60396
rect 65916 60342 65918 60394
rect 65918 60342 65970 60394
rect 65970 60342 65972 60394
rect 65916 60340 65972 60342
rect 66020 60394 66076 60396
rect 66020 60342 66022 60394
rect 66022 60342 66074 60394
rect 66074 60342 66076 60394
rect 66020 60340 66076 60342
rect 66124 60394 66180 60396
rect 66124 60342 66126 60394
rect 66126 60342 66178 60394
rect 66178 60342 66180 60394
rect 66124 60340 66180 60342
rect 65916 58826 65972 58828
rect 65916 58774 65918 58826
rect 65918 58774 65970 58826
rect 65970 58774 65972 58826
rect 65916 58772 65972 58774
rect 66020 58826 66076 58828
rect 66020 58774 66022 58826
rect 66022 58774 66074 58826
rect 66074 58774 66076 58826
rect 66020 58772 66076 58774
rect 66124 58826 66180 58828
rect 66124 58774 66126 58826
rect 66126 58774 66178 58826
rect 66178 58774 66180 58826
rect 66124 58772 66180 58774
rect 65916 57258 65972 57260
rect 65916 57206 65918 57258
rect 65918 57206 65970 57258
rect 65970 57206 65972 57258
rect 65916 57204 65972 57206
rect 66020 57258 66076 57260
rect 66020 57206 66022 57258
rect 66022 57206 66074 57258
rect 66074 57206 66076 57258
rect 66020 57204 66076 57206
rect 66124 57258 66180 57260
rect 66124 57206 66126 57258
rect 66126 57206 66178 57258
rect 66178 57206 66180 57258
rect 66124 57204 66180 57206
rect 65916 55690 65972 55692
rect 65916 55638 65918 55690
rect 65918 55638 65970 55690
rect 65970 55638 65972 55690
rect 65916 55636 65972 55638
rect 66020 55690 66076 55692
rect 66020 55638 66022 55690
rect 66022 55638 66074 55690
rect 66074 55638 66076 55690
rect 66020 55636 66076 55638
rect 66124 55690 66180 55692
rect 66124 55638 66126 55690
rect 66126 55638 66178 55690
rect 66178 55638 66180 55690
rect 66124 55636 66180 55638
rect 65916 54122 65972 54124
rect 65916 54070 65918 54122
rect 65918 54070 65970 54122
rect 65970 54070 65972 54122
rect 65916 54068 65972 54070
rect 66020 54122 66076 54124
rect 66020 54070 66022 54122
rect 66022 54070 66074 54122
rect 66074 54070 66076 54122
rect 66020 54068 66076 54070
rect 66124 54122 66180 54124
rect 66124 54070 66126 54122
rect 66126 54070 66178 54122
rect 66178 54070 66180 54122
rect 66124 54068 66180 54070
rect 65916 52554 65972 52556
rect 65916 52502 65918 52554
rect 65918 52502 65970 52554
rect 65970 52502 65972 52554
rect 65916 52500 65972 52502
rect 66020 52554 66076 52556
rect 66020 52502 66022 52554
rect 66022 52502 66074 52554
rect 66074 52502 66076 52554
rect 66020 52500 66076 52502
rect 66124 52554 66180 52556
rect 66124 52502 66126 52554
rect 66126 52502 66178 52554
rect 66178 52502 66180 52554
rect 66124 52500 66180 52502
rect 65916 50986 65972 50988
rect 65916 50934 65918 50986
rect 65918 50934 65970 50986
rect 65970 50934 65972 50986
rect 65916 50932 65972 50934
rect 66020 50986 66076 50988
rect 66020 50934 66022 50986
rect 66022 50934 66074 50986
rect 66074 50934 66076 50986
rect 66020 50932 66076 50934
rect 66124 50986 66180 50988
rect 66124 50934 66126 50986
rect 66126 50934 66178 50986
rect 66178 50934 66180 50986
rect 66124 50932 66180 50934
rect 65916 49418 65972 49420
rect 65916 49366 65918 49418
rect 65918 49366 65970 49418
rect 65970 49366 65972 49418
rect 65916 49364 65972 49366
rect 66020 49418 66076 49420
rect 66020 49366 66022 49418
rect 66022 49366 66074 49418
rect 66074 49366 66076 49418
rect 66020 49364 66076 49366
rect 66124 49418 66180 49420
rect 66124 49366 66126 49418
rect 66126 49366 66178 49418
rect 66178 49366 66180 49418
rect 66124 49364 66180 49366
rect 65916 47850 65972 47852
rect 65916 47798 65918 47850
rect 65918 47798 65970 47850
rect 65970 47798 65972 47850
rect 65916 47796 65972 47798
rect 66020 47850 66076 47852
rect 66020 47798 66022 47850
rect 66022 47798 66074 47850
rect 66074 47798 66076 47850
rect 66020 47796 66076 47798
rect 66124 47850 66180 47852
rect 66124 47798 66126 47850
rect 66126 47798 66178 47850
rect 66178 47798 66180 47850
rect 66124 47796 66180 47798
rect 65916 46282 65972 46284
rect 65916 46230 65918 46282
rect 65918 46230 65970 46282
rect 65970 46230 65972 46282
rect 65916 46228 65972 46230
rect 66020 46282 66076 46284
rect 66020 46230 66022 46282
rect 66022 46230 66074 46282
rect 66074 46230 66076 46282
rect 66020 46228 66076 46230
rect 66124 46282 66180 46284
rect 66124 46230 66126 46282
rect 66126 46230 66178 46282
rect 66178 46230 66180 46282
rect 66124 46228 66180 46230
rect 65916 44714 65972 44716
rect 65916 44662 65918 44714
rect 65918 44662 65970 44714
rect 65970 44662 65972 44714
rect 65916 44660 65972 44662
rect 66020 44714 66076 44716
rect 66020 44662 66022 44714
rect 66022 44662 66074 44714
rect 66074 44662 66076 44714
rect 66020 44660 66076 44662
rect 66124 44714 66180 44716
rect 66124 44662 66126 44714
rect 66126 44662 66178 44714
rect 66178 44662 66180 44714
rect 66124 44660 66180 44662
rect 65916 43146 65972 43148
rect 65916 43094 65918 43146
rect 65918 43094 65970 43146
rect 65970 43094 65972 43146
rect 65916 43092 65972 43094
rect 66020 43146 66076 43148
rect 66020 43094 66022 43146
rect 66022 43094 66074 43146
rect 66074 43094 66076 43146
rect 66020 43092 66076 43094
rect 66124 43146 66180 43148
rect 66124 43094 66126 43146
rect 66126 43094 66178 43146
rect 66178 43094 66180 43146
rect 66124 43092 66180 43094
rect 65772 42140 65828 42196
rect 65660 41468 65716 41524
rect 65884 41970 65940 41972
rect 65884 41918 65886 41970
rect 65886 41918 65938 41970
rect 65938 41918 65940 41970
rect 65884 41916 65940 41918
rect 65916 41578 65972 41580
rect 65916 41526 65918 41578
rect 65918 41526 65970 41578
rect 65970 41526 65972 41578
rect 65916 41524 65972 41526
rect 66020 41578 66076 41580
rect 66020 41526 66022 41578
rect 66022 41526 66074 41578
rect 66074 41526 66076 41578
rect 66020 41524 66076 41526
rect 66124 41578 66180 41580
rect 66124 41526 66126 41578
rect 66126 41526 66178 41578
rect 66178 41526 66180 41578
rect 66124 41524 66180 41526
rect 67788 76972 67844 77028
rect 68348 76636 68404 76692
rect 68012 76524 68068 76580
rect 66332 40572 66388 40628
rect 65212 39618 65268 39620
rect 65212 39566 65214 39618
rect 65214 39566 65266 39618
rect 65266 39566 65268 39618
rect 65212 39564 65268 39566
rect 65916 40010 65972 40012
rect 65916 39958 65918 40010
rect 65918 39958 65970 40010
rect 65970 39958 65972 40010
rect 65916 39956 65972 39958
rect 66020 40010 66076 40012
rect 66020 39958 66022 40010
rect 66022 39958 66074 40010
rect 66074 39958 66076 40010
rect 66020 39956 66076 39958
rect 66124 40010 66180 40012
rect 66124 39958 66126 40010
rect 66126 39958 66178 40010
rect 66178 39958 66180 40010
rect 66124 39956 66180 39958
rect 65772 39676 65828 39732
rect 65772 39506 65828 39508
rect 65772 39454 65774 39506
rect 65774 39454 65826 39506
rect 65826 39454 65828 39506
rect 65772 39452 65828 39454
rect 66332 39564 66388 39620
rect 65884 39116 65940 39172
rect 65324 39058 65380 39060
rect 65324 39006 65326 39058
rect 65326 39006 65378 39058
rect 65378 39006 65380 39058
rect 65324 39004 65380 39006
rect 65916 38442 65972 38444
rect 65916 38390 65918 38442
rect 65918 38390 65970 38442
rect 65970 38390 65972 38442
rect 65916 38388 65972 38390
rect 66020 38442 66076 38444
rect 66020 38390 66022 38442
rect 66022 38390 66074 38442
rect 66074 38390 66076 38442
rect 66020 38388 66076 38390
rect 66124 38442 66180 38444
rect 66124 38390 66126 38442
rect 66126 38390 66178 38442
rect 66178 38390 66180 38442
rect 66124 38388 66180 38390
rect 64764 37996 64820 38052
rect 65916 36874 65972 36876
rect 65916 36822 65918 36874
rect 65918 36822 65970 36874
rect 65970 36822 65972 36874
rect 65916 36820 65972 36822
rect 66020 36874 66076 36876
rect 66020 36822 66022 36874
rect 66022 36822 66074 36874
rect 66074 36822 66076 36874
rect 66020 36820 66076 36822
rect 66124 36874 66180 36876
rect 66124 36822 66126 36874
rect 66126 36822 66178 36874
rect 66178 36822 66180 36874
rect 66124 36820 66180 36822
rect 65916 35306 65972 35308
rect 65916 35254 65918 35306
rect 65918 35254 65970 35306
rect 65970 35254 65972 35306
rect 65916 35252 65972 35254
rect 66020 35306 66076 35308
rect 66020 35254 66022 35306
rect 66022 35254 66074 35306
rect 66074 35254 66076 35306
rect 66020 35252 66076 35254
rect 66124 35306 66180 35308
rect 66124 35254 66126 35306
rect 66126 35254 66178 35306
rect 66178 35254 66180 35306
rect 66124 35252 66180 35254
rect 64540 28364 64596 28420
rect 64652 33852 64708 33908
rect 64428 25452 64484 25508
rect 63196 25116 63252 25172
rect 63308 25004 63364 25060
rect 65916 33738 65972 33740
rect 65916 33686 65918 33738
rect 65918 33686 65970 33738
rect 65970 33686 65972 33738
rect 65916 33684 65972 33686
rect 66020 33738 66076 33740
rect 66020 33686 66022 33738
rect 66022 33686 66074 33738
rect 66074 33686 66076 33738
rect 66020 33684 66076 33686
rect 66124 33738 66180 33740
rect 66124 33686 66126 33738
rect 66126 33686 66178 33738
rect 66178 33686 66180 33738
rect 66124 33684 66180 33686
rect 65916 32170 65972 32172
rect 65916 32118 65918 32170
rect 65918 32118 65970 32170
rect 65970 32118 65972 32170
rect 65916 32116 65972 32118
rect 66020 32170 66076 32172
rect 66020 32118 66022 32170
rect 66022 32118 66074 32170
rect 66074 32118 66076 32170
rect 66020 32116 66076 32118
rect 66124 32170 66180 32172
rect 66124 32118 66126 32170
rect 66126 32118 66178 32170
rect 66178 32118 66180 32170
rect 66124 32116 66180 32118
rect 64652 25004 64708 25060
rect 64764 31724 64820 31780
rect 63420 24610 63476 24612
rect 63420 24558 63422 24610
rect 63422 24558 63474 24610
rect 63474 24558 63476 24610
rect 63420 24556 63476 24558
rect 63532 24220 63588 24276
rect 63420 23996 63476 24052
rect 61740 17724 61796 17780
rect 61852 23100 61908 23156
rect 61628 4396 61684 4452
rect 61404 3836 61460 3892
rect 64092 24050 64148 24052
rect 64092 23998 64094 24050
rect 64094 23998 64146 24050
rect 64146 23998 64148 24050
rect 64092 23996 64148 23998
rect 63756 22988 63812 23044
rect 63644 21756 63700 21812
rect 62636 21420 62692 21476
rect 62188 7980 62244 8036
rect 62188 6300 62244 6356
rect 62524 4450 62580 4452
rect 62524 4398 62526 4450
rect 62526 4398 62578 4450
rect 62578 4398 62580 4450
rect 62524 4396 62580 4398
rect 63532 20188 63588 20244
rect 62076 3724 62132 3780
rect 62748 6412 62804 6468
rect 63196 6018 63252 6020
rect 63196 5966 63198 6018
rect 63198 5966 63250 6018
rect 63250 5966 63252 6018
rect 63196 5964 63252 5966
rect 64652 18956 64708 19012
rect 64540 17948 64596 18004
rect 63868 9100 63924 9156
rect 64428 6466 64484 6468
rect 64428 6414 64430 6466
rect 64430 6414 64482 6466
rect 64482 6414 64484 6466
rect 64428 6412 64484 6414
rect 64428 5234 64484 5236
rect 64428 5182 64430 5234
rect 64430 5182 64482 5234
rect 64482 5182 64484 5234
rect 64428 5180 64484 5182
rect 63756 5068 63812 5124
rect 65916 30602 65972 30604
rect 65916 30550 65918 30602
rect 65918 30550 65970 30602
rect 65970 30550 65972 30602
rect 65916 30548 65972 30550
rect 66020 30602 66076 30604
rect 66020 30550 66022 30602
rect 66022 30550 66074 30602
rect 66074 30550 66076 30602
rect 66020 30548 66076 30550
rect 66124 30602 66180 30604
rect 66124 30550 66126 30602
rect 66126 30550 66178 30602
rect 66178 30550 66180 30602
rect 66124 30548 66180 30550
rect 65916 29034 65972 29036
rect 65916 28982 65918 29034
rect 65918 28982 65970 29034
rect 65970 28982 65972 29034
rect 65916 28980 65972 28982
rect 66020 29034 66076 29036
rect 66020 28982 66022 29034
rect 66022 28982 66074 29034
rect 66074 28982 66076 29034
rect 66020 28980 66076 28982
rect 66124 29034 66180 29036
rect 66124 28982 66126 29034
rect 66126 28982 66178 29034
rect 66178 28982 66180 29034
rect 66124 28980 66180 28982
rect 65916 27466 65972 27468
rect 65916 27414 65918 27466
rect 65918 27414 65970 27466
rect 65970 27414 65972 27466
rect 65916 27412 65972 27414
rect 66020 27466 66076 27468
rect 66020 27414 66022 27466
rect 66022 27414 66074 27466
rect 66074 27414 66076 27466
rect 66020 27412 66076 27414
rect 66124 27466 66180 27468
rect 66124 27414 66126 27466
rect 66126 27414 66178 27466
rect 66178 27414 66180 27466
rect 66124 27412 66180 27414
rect 65916 25898 65972 25900
rect 65916 25846 65918 25898
rect 65918 25846 65970 25898
rect 65970 25846 65972 25898
rect 65916 25844 65972 25846
rect 66020 25898 66076 25900
rect 66020 25846 66022 25898
rect 66022 25846 66074 25898
rect 66074 25846 66076 25898
rect 66020 25844 66076 25846
rect 66124 25898 66180 25900
rect 66124 25846 66126 25898
rect 66126 25846 66178 25898
rect 66178 25846 66180 25898
rect 66124 25844 66180 25846
rect 65916 24330 65972 24332
rect 65916 24278 65918 24330
rect 65918 24278 65970 24330
rect 65970 24278 65972 24330
rect 65916 24276 65972 24278
rect 66020 24330 66076 24332
rect 66020 24278 66022 24330
rect 66022 24278 66074 24330
rect 66074 24278 66076 24330
rect 66020 24276 66076 24278
rect 66124 24330 66180 24332
rect 66124 24278 66126 24330
rect 66126 24278 66178 24330
rect 66178 24278 66180 24330
rect 66124 24276 66180 24278
rect 65916 22762 65972 22764
rect 65916 22710 65918 22762
rect 65918 22710 65970 22762
rect 65970 22710 65972 22762
rect 65916 22708 65972 22710
rect 66020 22762 66076 22764
rect 66020 22710 66022 22762
rect 66022 22710 66074 22762
rect 66074 22710 66076 22762
rect 66020 22708 66076 22710
rect 66124 22762 66180 22764
rect 66124 22710 66126 22762
rect 66126 22710 66178 22762
rect 66178 22710 66180 22762
rect 66124 22708 66180 22710
rect 66444 21644 66500 21700
rect 65916 21194 65972 21196
rect 65916 21142 65918 21194
rect 65918 21142 65970 21194
rect 65970 21142 65972 21194
rect 65916 21140 65972 21142
rect 66020 21194 66076 21196
rect 66020 21142 66022 21194
rect 66022 21142 66074 21194
rect 66074 21142 66076 21194
rect 66020 21140 66076 21142
rect 66124 21194 66180 21196
rect 66124 21142 66126 21194
rect 66126 21142 66178 21194
rect 66178 21142 66180 21194
rect 66124 21140 66180 21142
rect 66668 39618 66724 39620
rect 66668 39566 66670 39618
rect 66670 39566 66722 39618
rect 66722 39566 66724 39618
rect 66668 39564 66724 39566
rect 67452 40626 67508 40628
rect 67452 40574 67454 40626
rect 67454 40574 67506 40626
rect 67506 40574 67508 40626
rect 67452 40572 67508 40574
rect 67564 40348 67620 40404
rect 67116 39730 67172 39732
rect 67116 39678 67118 39730
rect 67118 39678 67170 39730
rect 67170 39678 67172 39730
rect 67116 39676 67172 39678
rect 67116 38946 67172 38948
rect 67116 38894 67118 38946
rect 67118 38894 67170 38946
rect 67170 38894 67172 38946
rect 67116 38892 67172 38894
rect 67900 41356 67956 41412
rect 67900 41020 67956 41076
rect 67676 39452 67732 39508
rect 67340 38668 67396 38724
rect 68012 39004 68068 39060
rect 67788 37826 67844 37828
rect 67788 37774 67790 37826
rect 67790 37774 67842 37826
rect 67842 37774 67844 37826
rect 67788 37772 67844 37774
rect 67564 36204 67620 36260
rect 67004 32844 67060 32900
rect 66668 28924 66724 28980
rect 68236 40402 68292 40404
rect 68236 40350 68238 40402
rect 68238 40350 68290 40402
rect 68290 40350 68292 40402
rect 68236 40348 68292 40350
rect 68460 39788 68516 39844
rect 68460 39506 68516 39508
rect 68460 39454 68462 39506
rect 68462 39454 68514 39506
rect 68514 39454 68516 39506
rect 68460 39452 68516 39454
rect 68572 39116 68628 39172
rect 69132 76690 69188 76692
rect 69132 76638 69134 76690
rect 69134 76638 69186 76690
rect 69186 76638 69188 76690
rect 69132 76636 69188 76638
rect 68796 76578 68852 76580
rect 68796 76526 68798 76578
rect 68798 76526 68850 76578
rect 68850 76526 68852 76578
rect 68796 76524 68852 76526
rect 68684 39004 68740 39060
rect 68908 58156 68964 58212
rect 68236 38668 68292 38724
rect 68684 37772 68740 37828
rect 68012 32844 68068 32900
rect 67788 23324 67844 23380
rect 66556 20860 66612 20916
rect 67116 22204 67172 22260
rect 65916 19626 65972 19628
rect 65916 19574 65918 19626
rect 65918 19574 65970 19626
rect 65970 19574 65972 19626
rect 65916 19572 65972 19574
rect 66020 19626 66076 19628
rect 66020 19574 66022 19626
rect 66022 19574 66074 19626
rect 66074 19574 66076 19626
rect 66020 19572 66076 19574
rect 66124 19626 66180 19628
rect 66124 19574 66126 19626
rect 66126 19574 66178 19626
rect 66178 19574 66180 19626
rect 66124 19572 66180 19574
rect 70364 76972 70420 77028
rect 69692 76524 69748 76580
rect 69356 75964 69412 76020
rect 70924 76578 70980 76580
rect 70924 76526 70926 76578
rect 70926 76526 70978 76578
rect 70978 76526 70980 76578
rect 70924 76524 70980 76526
rect 70476 76076 70532 76132
rect 70028 66220 70084 66276
rect 69580 41356 69636 41412
rect 69356 40572 69412 40628
rect 69020 40348 69076 40404
rect 69356 39394 69412 39396
rect 69356 39342 69358 39394
rect 69358 39342 69410 39394
rect 69410 39342 69412 39394
rect 69356 39340 69412 39342
rect 69020 39116 69076 39172
rect 69020 38780 69076 38836
rect 69244 39058 69300 39060
rect 69244 39006 69246 39058
rect 69246 39006 69298 39058
rect 69298 39006 69300 39058
rect 69244 39004 69300 39006
rect 69020 36258 69076 36260
rect 69020 36206 69022 36258
rect 69022 36206 69074 36258
rect 69074 36206 69076 36258
rect 69020 36204 69076 36206
rect 68908 28140 68964 28196
rect 68908 23548 68964 23604
rect 68908 22428 68964 22484
rect 69356 36204 69412 36260
rect 69244 22428 69300 22484
rect 69692 39452 69748 39508
rect 69692 38946 69748 38948
rect 69692 38894 69694 38946
rect 69694 38894 69746 38946
rect 69746 38894 69748 38946
rect 69692 38892 69748 38894
rect 69580 38332 69636 38388
rect 69804 38668 69860 38724
rect 69804 38108 69860 38164
rect 69692 37772 69748 37828
rect 70476 42252 70532 42308
rect 70812 53004 70868 53060
rect 70252 40796 70308 40852
rect 70476 41580 70532 41636
rect 70700 41244 70756 41300
rect 70700 40684 70756 40740
rect 70476 40460 70532 40516
rect 70700 40460 70756 40516
rect 70140 40124 70196 40180
rect 70700 39676 70756 39732
rect 70364 39618 70420 39620
rect 70364 39566 70366 39618
rect 70366 39566 70418 39618
rect 70418 39566 70420 39618
rect 70364 39564 70420 39566
rect 70028 39506 70084 39508
rect 70028 39454 70030 39506
rect 70030 39454 70082 39506
rect 70082 39454 70084 39506
rect 70028 39452 70084 39454
rect 70028 38780 70084 38836
rect 70140 38220 70196 38276
rect 69916 32844 69972 32900
rect 70476 39340 70532 39396
rect 70364 38834 70420 38836
rect 70364 38782 70366 38834
rect 70366 38782 70418 38834
rect 70418 38782 70420 38834
rect 70364 38780 70420 38782
rect 70700 38834 70756 38836
rect 70700 38782 70702 38834
rect 70702 38782 70754 38834
rect 70754 38782 70756 38834
rect 70700 38780 70756 38782
rect 70588 38162 70644 38164
rect 70588 38110 70590 38162
rect 70590 38110 70642 38162
rect 70642 38110 70644 38162
rect 70588 38108 70644 38110
rect 70588 37772 70644 37828
rect 70588 37378 70644 37380
rect 70588 37326 70590 37378
rect 70590 37326 70642 37378
rect 70642 37326 70644 37378
rect 70588 37324 70644 37326
rect 70588 35532 70644 35588
rect 70588 31948 70644 32004
rect 71148 41692 71204 41748
rect 70924 40796 70980 40852
rect 71372 41298 71428 41300
rect 71372 41246 71374 41298
rect 71374 41246 71426 41298
rect 71426 41246 71428 41298
rect 71372 41244 71428 41246
rect 71372 40626 71428 40628
rect 71372 40574 71374 40626
rect 71374 40574 71426 40626
rect 71426 40574 71428 40626
rect 71372 40572 71428 40574
rect 71260 40236 71316 40292
rect 70924 39676 70980 39732
rect 70924 39506 70980 39508
rect 70924 39454 70926 39506
rect 70926 39454 70978 39506
rect 70978 39454 70980 39506
rect 70924 39452 70980 39454
rect 71708 76524 71764 76580
rect 71820 76972 71876 77028
rect 72268 76188 72324 76244
rect 73052 76636 73108 76692
rect 72156 68796 72212 68852
rect 71596 41692 71652 41748
rect 71708 41468 71764 41524
rect 71484 39564 71540 39620
rect 70924 37884 70980 37940
rect 71260 39340 71316 39396
rect 72044 45836 72100 45892
rect 71932 39788 71988 39844
rect 71260 38780 71316 38836
rect 71260 38050 71316 38052
rect 71260 37998 71262 38050
rect 71262 37998 71314 38050
rect 71314 37998 71316 38050
rect 71260 37996 71316 37998
rect 71260 37378 71316 37380
rect 71260 37326 71262 37378
rect 71262 37326 71314 37378
rect 71314 37326 71316 37378
rect 71260 37324 71316 37326
rect 71932 38108 71988 38164
rect 71820 37996 71876 38052
rect 71596 37938 71652 37940
rect 71596 37886 71598 37938
rect 71598 37886 71650 37938
rect 71650 37886 71652 37938
rect 71596 37884 71652 37886
rect 71708 35586 71764 35588
rect 71708 35534 71710 35586
rect 71710 35534 71762 35586
rect 71762 35534 71764 35586
rect 71708 35532 71764 35534
rect 73164 76524 73220 76580
rect 73724 76524 73780 76580
rect 74060 76690 74116 76692
rect 74060 76638 74062 76690
rect 74062 76638 74114 76690
rect 74114 76638 74116 76690
rect 74060 76636 74116 76638
rect 73836 75628 73892 75684
rect 73724 73948 73780 74004
rect 72156 41804 72212 41860
rect 72604 48524 72660 48580
rect 72268 40460 72324 40516
rect 72380 40236 72436 40292
rect 72380 39340 72436 39396
rect 72492 38834 72548 38836
rect 72492 38782 72494 38834
rect 72494 38782 72546 38834
rect 72546 38782 72548 38834
rect 72492 38780 72548 38782
rect 72268 38220 72324 38276
rect 72492 38556 72548 38612
rect 72268 37884 72324 37940
rect 72268 37378 72324 37380
rect 72268 37326 72270 37378
rect 72270 37326 72322 37378
rect 72322 37326 72324 37378
rect 72268 37324 72324 37326
rect 73164 45612 73220 45668
rect 72940 40684 72996 40740
rect 72828 39564 72884 39620
rect 73276 41074 73332 41076
rect 73276 41022 73278 41074
rect 73278 41022 73330 41074
rect 73330 41022 73332 41074
rect 73276 41020 73332 41022
rect 73388 40402 73444 40404
rect 73388 40350 73390 40402
rect 73390 40350 73442 40402
rect 73442 40350 73444 40402
rect 73388 40348 73444 40350
rect 73276 39676 73332 39732
rect 72940 39116 72996 39172
rect 72604 38108 72660 38164
rect 72940 38162 72996 38164
rect 72940 38110 72942 38162
rect 72942 38110 72994 38162
rect 72994 38110 72996 38162
rect 72940 38108 72996 38110
rect 72828 37938 72884 37940
rect 72828 37886 72830 37938
rect 72830 37886 72882 37938
rect 72882 37886 72884 37938
rect 72828 37884 72884 37886
rect 73612 41916 73668 41972
rect 73612 40514 73668 40516
rect 73612 40462 73614 40514
rect 73614 40462 73666 40514
rect 73666 40462 73668 40514
rect 73612 40460 73668 40462
rect 74060 75404 74116 75460
rect 73836 45276 73892 45332
rect 74172 74732 74228 74788
rect 74060 41970 74116 41972
rect 74060 41918 74062 41970
rect 74062 41918 74114 41970
rect 74114 41918 74116 41970
rect 74060 41916 74116 41918
rect 74508 76524 74564 76580
rect 74508 75516 74564 75572
rect 74620 74060 74676 74116
rect 74396 41468 74452 41524
rect 73836 41074 73892 41076
rect 73836 41022 73838 41074
rect 73838 41022 73890 41074
rect 73890 41022 73892 41074
rect 73836 41020 73892 41022
rect 73724 38834 73780 38836
rect 73724 38782 73726 38834
rect 73726 38782 73778 38834
rect 73778 38782 73780 38834
rect 73724 38780 73780 38782
rect 73388 38556 73444 38612
rect 73948 40348 74004 40404
rect 74172 41298 74228 41300
rect 74172 41246 74174 41298
rect 74174 41246 74226 41298
rect 74226 41246 74228 41298
rect 74172 41244 74228 41246
rect 74060 40124 74116 40180
rect 74284 40514 74340 40516
rect 74284 40462 74286 40514
rect 74286 40462 74338 40514
rect 74338 40462 74340 40514
rect 74284 40460 74340 40462
rect 74172 39564 74228 39620
rect 74172 38892 74228 38948
rect 73164 38108 73220 38164
rect 72716 37772 72772 37828
rect 71484 35196 71540 35252
rect 71260 34972 71316 35028
rect 70924 34802 70980 34804
rect 70924 34750 70926 34802
rect 70926 34750 70978 34802
rect 70978 34750 70980 34802
rect 70924 34748 70980 34750
rect 70812 34300 70868 34356
rect 70700 30492 70756 30548
rect 70700 30268 70756 30324
rect 70140 27356 70196 27412
rect 70924 29036 70980 29092
rect 70812 28588 70868 28644
rect 70700 27858 70756 27860
rect 70700 27806 70702 27858
rect 70702 27806 70754 27858
rect 70754 27806 70756 27858
rect 70700 27804 70756 27806
rect 70700 27468 70756 27524
rect 70252 25004 70308 25060
rect 70476 25394 70532 25396
rect 70476 25342 70478 25394
rect 70478 25342 70530 25394
rect 70530 25342 70532 25394
rect 70476 25340 70532 25342
rect 70476 24332 70532 24388
rect 71932 34972 71988 35028
rect 71596 34914 71652 34916
rect 71596 34862 71598 34914
rect 71598 34862 71650 34914
rect 71650 34862 71652 34914
rect 71596 34860 71652 34862
rect 71820 34914 71876 34916
rect 71820 34862 71822 34914
rect 71822 34862 71874 34914
rect 71874 34862 71876 34914
rect 71820 34860 71876 34862
rect 71932 34690 71988 34692
rect 71932 34638 71934 34690
rect 71934 34638 71986 34690
rect 71986 34638 71988 34690
rect 71932 34636 71988 34638
rect 71260 34300 71316 34356
rect 71372 34242 71428 34244
rect 71372 34190 71374 34242
rect 71374 34190 71426 34242
rect 71426 34190 71428 34242
rect 71372 34188 71428 34190
rect 71260 32562 71316 32564
rect 71260 32510 71262 32562
rect 71262 32510 71314 32562
rect 71314 32510 71316 32562
rect 71260 32508 71316 32510
rect 71372 31836 71428 31892
rect 71372 30940 71428 30996
rect 72156 34972 72212 35028
rect 73164 37772 73220 37828
rect 73612 37772 73668 37828
rect 72604 37100 72660 37156
rect 72492 36482 72548 36484
rect 72492 36430 72494 36482
rect 72494 36430 72546 36482
rect 72546 36430 72548 36482
rect 72492 36428 72548 36430
rect 73052 37324 73108 37380
rect 73388 37324 73444 37380
rect 73276 37154 73332 37156
rect 73276 37102 73278 37154
rect 73278 37102 73330 37154
rect 73330 37102 73332 37154
rect 73276 37100 73332 37102
rect 72268 34636 72324 34692
rect 72380 34802 72436 34804
rect 72380 34750 72382 34802
rect 72382 34750 72434 34802
rect 72434 34750 72436 34802
rect 72380 34748 72436 34750
rect 72604 35532 72660 35588
rect 72044 33404 72100 33460
rect 71596 32450 71652 32452
rect 71596 32398 71598 32450
rect 71598 32398 71650 32450
rect 71650 32398 71652 32450
rect 71596 32396 71652 32398
rect 71708 30940 71764 30996
rect 71372 30156 71428 30212
rect 71148 29986 71204 29988
rect 71148 29934 71150 29986
rect 71150 29934 71202 29986
rect 71202 29934 71204 29986
rect 71148 29932 71204 29934
rect 71484 28476 71540 28532
rect 70924 26236 70980 26292
rect 70588 23772 70644 23828
rect 70924 25506 70980 25508
rect 70924 25454 70926 25506
rect 70926 25454 70978 25506
rect 70978 25454 70980 25506
rect 70924 25452 70980 25454
rect 71036 25004 71092 25060
rect 71036 23660 71092 23716
rect 70700 22876 70756 22932
rect 71036 22876 71092 22932
rect 69468 22316 69524 22372
rect 68012 21532 68068 21588
rect 70252 22204 70308 22260
rect 67116 18956 67172 19012
rect 68572 18844 68628 18900
rect 65916 18058 65972 18060
rect 65916 18006 65918 18058
rect 65918 18006 65970 18058
rect 65970 18006 65972 18058
rect 65916 18004 65972 18006
rect 66020 18058 66076 18060
rect 66020 18006 66022 18058
rect 66022 18006 66074 18058
rect 66074 18006 66076 18058
rect 66020 18004 66076 18006
rect 66124 18058 66180 18060
rect 66124 18006 66126 18058
rect 66126 18006 66178 18058
rect 66178 18006 66180 18058
rect 66124 18004 66180 18006
rect 65916 16490 65972 16492
rect 65916 16438 65918 16490
rect 65918 16438 65970 16490
rect 65970 16438 65972 16490
rect 65916 16436 65972 16438
rect 66020 16490 66076 16492
rect 66020 16438 66022 16490
rect 66022 16438 66074 16490
rect 66074 16438 66076 16490
rect 66020 16436 66076 16438
rect 66124 16490 66180 16492
rect 66124 16438 66126 16490
rect 66126 16438 66178 16490
rect 66178 16438 66180 16490
rect 66124 16436 66180 16438
rect 65916 14922 65972 14924
rect 65916 14870 65918 14922
rect 65918 14870 65970 14922
rect 65970 14870 65972 14922
rect 65916 14868 65972 14870
rect 66020 14922 66076 14924
rect 66020 14870 66022 14922
rect 66022 14870 66074 14922
rect 66074 14870 66076 14922
rect 66020 14868 66076 14870
rect 66124 14922 66180 14924
rect 66124 14870 66126 14922
rect 66126 14870 66178 14922
rect 66178 14870 66180 14922
rect 66124 14868 66180 14870
rect 65916 13354 65972 13356
rect 65916 13302 65918 13354
rect 65918 13302 65970 13354
rect 65970 13302 65972 13354
rect 65916 13300 65972 13302
rect 66020 13354 66076 13356
rect 66020 13302 66022 13354
rect 66022 13302 66074 13354
rect 66074 13302 66076 13354
rect 66020 13300 66076 13302
rect 66124 13354 66180 13356
rect 66124 13302 66126 13354
rect 66126 13302 66178 13354
rect 66178 13302 66180 13354
rect 66124 13300 66180 13302
rect 65916 11786 65972 11788
rect 65916 11734 65918 11786
rect 65918 11734 65970 11786
rect 65970 11734 65972 11786
rect 65916 11732 65972 11734
rect 66020 11786 66076 11788
rect 66020 11734 66022 11786
rect 66022 11734 66074 11786
rect 66074 11734 66076 11786
rect 66020 11732 66076 11734
rect 66124 11786 66180 11788
rect 66124 11734 66126 11786
rect 66126 11734 66178 11786
rect 66178 11734 66180 11786
rect 66124 11732 66180 11734
rect 67452 11228 67508 11284
rect 65916 10218 65972 10220
rect 65916 10166 65918 10218
rect 65918 10166 65970 10218
rect 65970 10166 65972 10218
rect 65916 10164 65972 10166
rect 66020 10218 66076 10220
rect 66020 10166 66022 10218
rect 66022 10166 66074 10218
rect 66074 10166 66076 10218
rect 66020 10164 66076 10166
rect 66124 10218 66180 10220
rect 66124 10166 66126 10218
rect 66126 10166 66178 10218
rect 66178 10166 66180 10218
rect 66124 10164 66180 10166
rect 64764 9772 64820 9828
rect 67116 9212 67172 9268
rect 65916 8650 65972 8652
rect 65916 8598 65918 8650
rect 65918 8598 65970 8650
rect 65970 8598 65972 8650
rect 65916 8596 65972 8598
rect 66020 8650 66076 8652
rect 66020 8598 66022 8650
rect 66022 8598 66074 8650
rect 66074 8598 66076 8650
rect 66020 8596 66076 8598
rect 66124 8650 66180 8652
rect 66124 8598 66126 8650
rect 66126 8598 66178 8650
rect 66178 8598 66180 8650
rect 66124 8596 66180 8598
rect 66668 7586 66724 7588
rect 66668 7534 66670 7586
rect 66670 7534 66722 7586
rect 66722 7534 66724 7586
rect 66668 7532 66724 7534
rect 65916 7082 65972 7084
rect 65916 7030 65918 7082
rect 65918 7030 65970 7082
rect 65970 7030 65972 7082
rect 65916 7028 65972 7030
rect 66020 7082 66076 7084
rect 66020 7030 66022 7082
rect 66022 7030 66074 7082
rect 66074 7030 66076 7082
rect 66020 7028 66076 7030
rect 66124 7082 66180 7084
rect 66124 7030 66126 7082
rect 66126 7030 66178 7082
rect 66178 7030 66180 7082
rect 66124 7028 66180 7030
rect 67340 6188 67396 6244
rect 64652 5180 64708 5236
rect 65916 5514 65972 5516
rect 65916 5462 65918 5514
rect 65918 5462 65970 5514
rect 65970 5462 65972 5514
rect 65916 5460 65972 5462
rect 66020 5514 66076 5516
rect 66020 5462 66022 5514
rect 66022 5462 66074 5514
rect 66074 5462 66076 5514
rect 66020 5460 66076 5462
rect 66124 5514 66180 5516
rect 66124 5462 66126 5514
rect 66126 5462 66178 5514
rect 66178 5462 66180 5514
rect 66124 5460 66180 5462
rect 65548 5068 65604 5124
rect 66332 5292 66388 5348
rect 64540 4338 64596 4340
rect 64540 4286 64542 4338
rect 64542 4286 64594 4338
rect 64594 4286 64596 4338
rect 64540 4284 64596 4286
rect 65660 4284 65716 4340
rect 64092 4060 64148 4116
rect 63868 3388 63924 3444
rect 65548 3836 65604 3892
rect 65916 3946 65972 3948
rect 65916 3894 65918 3946
rect 65918 3894 65970 3946
rect 65970 3894 65972 3946
rect 65916 3892 65972 3894
rect 66020 3946 66076 3948
rect 66020 3894 66022 3946
rect 66022 3894 66074 3946
rect 66074 3894 66076 3946
rect 66020 3892 66076 3894
rect 66124 3946 66180 3948
rect 66124 3894 66126 3946
rect 66126 3894 66178 3946
rect 66178 3894 66180 3946
rect 66124 3892 66180 3894
rect 65436 3500 65492 3556
rect 64764 3388 64820 3444
rect 66444 5234 66500 5236
rect 66444 5182 66446 5234
rect 66446 5182 66498 5234
rect 66498 5182 66500 5234
rect 66444 5180 66500 5182
rect 66780 5068 66836 5124
rect 67564 6412 67620 6468
rect 67452 3778 67508 3780
rect 67452 3726 67454 3778
rect 67454 3726 67506 3778
rect 67506 3726 67508 3778
rect 67452 3724 67508 3726
rect 67900 6300 67956 6356
rect 68460 6188 68516 6244
rect 67788 5068 67844 5124
rect 68124 5180 68180 5236
rect 70476 20636 70532 20692
rect 70476 19404 70532 19460
rect 70588 17836 70644 17892
rect 71372 25788 71428 25844
rect 71260 25730 71316 25732
rect 71260 25678 71262 25730
rect 71262 25678 71314 25730
rect 71314 25678 71316 25730
rect 71260 25676 71316 25678
rect 73724 37212 73780 37268
rect 72940 36764 72996 36820
rect 72940 35084 72996 35140
rect 73724 35308 73780 35364
rect 72828 34748 72884 34804
rect 73276 34914 73332 34916
rect 73276 34862 73278 34914
rect 73278 34862 73330 34914
rect 73330 34862 73332 34914
rect 73276 34860 73332 34862
rect 73500 34914 73556 34916
rect 73500 34862 73502 34914
rect 73502 34862 73554 34914
rect 73554 34862 73556 34914
rect 73500 34860 73556 34862
rect 72940 34412 72996 34468
rect 73276 34300 73332 34356
rect 73388 34636 73444 34692
rect 74284 38050 74340 38052
rect 74284 37998 74286 38050
rect 74286 37998 74338 38050
rect 74338 37998 74340 38050
rect 74284 37996 74340 37998
rect 73948 37436 74004 37492
rect 73948 36370 74004 36372
rect 73948 36318 73950 36370
rect 73950 36318 74002 36370
rect 74002 36318 74004 36370
rect 73948 36316 74004 36318
rect 73948 35756 74004 35812
rect 74284 36988 74340 37044
rect 74284 36764 74340 36820
rect 74956 76524 75012 76580
rect 74732 73948 74788 74004
rect 74844 75740 74900 75796
rect 75404 76748 75460 76804
rect 75404 75852 75460 75908
rect 75628 75628 75684 75684
rect 75404 75180 75460 75236
rect 74956 75122 75012 75124
rect 74956 75070 74958 75122
rect 74958 75070 75010 75122
rect 75010 75070 75012 75122
rect 74956 75068 75012 75070
rect 75292 74226 75348 74228
rect 75292 74174 75294 74226
rect 75294 74174 75346 74226
rect 75346 74174 75348 74226
rect 75292 74172 75348 74174
rect 76076 76578 76132 76580
rect 76076 76526 76078 76578
rect 76078 76526 76130 76578
rect 76130 76526 76132 76578
rect 76076 76524 76132 76526
rect 76076 75292 76132 75348
rect 75964 75180 76020 75236
rect 76188 75068 76244 75124
rect 76412 75852 76468 75908
rect 76300 74786 76356 74788
rect 76300 74734 76302 74786
rect 76302 74734 76354 74786
rect 76354 74734 76356 74786
rect 76300 74732 76356 74734
rect 76524 75740 76580 75796
rect 76524 74732 76580 74788
rect 76748 76354 76804 76356
rect 76748 76302 76750 76354
rect 76750 76302 76802 76354
rect 76802 76302 76804 76354
rect 76748 76300 76804 76302
rect 76860 75516 76916 75572
rect 76972 76860 77028 76916
rect 77196 78988 77252 79044
rect 77980 77980 78036 78036
rect 77084 75292 77140 75348
rect 76972 74114 77028 74116
rect 76972 74062 76974 74114
rect 76974 74062 77026 74114
rect 77026 74062 77028 74114
rect 76972 74060 77028 74062
rect 76412 72492 76468 72548
rect 74956 42140 75012 42196
rect 74732 41580 74788 41636
rect 75852 59052 75908 59108
rect 75740 45276 75796 45332
rect 75740 42588 75796 42644
rect 75068 41916 75124 41972
rect 75292 42476 75348 42532
rect 75068 41580 75124 41636
rect 74620 40626 74676 40628
rect 74620 40574 74622 40626
rect 74622 40574 74674 40626
rect 74674 40574 74676 40626
rect 74620 40572 74676 40574
rect 75068 40684 75124 40740
rect 75292 41298 75348 41300
rect 75292 41246 75294 41298
rect 75294 41246 75346 41298
rect 75346 41246 75348 41298
rect 75292 41244 75348 41246
rect 74620 39730 74676 39732
rect 74620 39678 74622 39730
rect 74622 39678 74674 39730
rect 74674 39678 74676 39730
rect 74620 39676 74676 39678
rect 75068 39618 75124 39620
rect 75068 39566 75070 39618
rect 75070 39566 75122 39618
rect 75122 39566 75124 39618
rect 75068 39564 75124 39566
rect 74508 39004 74564 39060
rect 75068 39340 75124 39396
rect 74844 38668 74900 38724
rect 74620 38050 74676 38052
rect 74620 37998 74622 38050
rect 74622 37998 74674 38050
rect 74674 37998 74676 38050
rect 74620 37996 74676 37998
rect 74620 36876 74676 36932
rect 74396 36370 74452 36372
rect 74396 36318 74398 36370
rect 74398 36318 74450 36370
rect 74450 36318 74452 36370
rect 74396 36316 74452 36318
rect 75292 40348 75348 40404
rect 75292 40178 75348 40180
rect 75292 40126 75294 40178
rect 75294 40126 75346 40178
rect 75346 40126 75348 40178
rect 75292 40124 75348 40126
rect 75292 39564 75348 39620
rect 77868 75964 77924 76020
rect 77756 75292 77812 75348
rect 77532 75010 77588 75012
rect 77532 74958 77534 75010
rect 77534 74958 77586 75010
rect 77586 74958 77588 75010
rect 77532 74956 77588 74958
rect 77308 74732 77364 74788
rect 77420 73554 77476 73556
rect 77420 73502 77422 73554
rect 77422 73502 77474 73554
rect 77474 73502 77476 73554
rect 77420 73500 77476 73502
rect 77644 73218 77700 73220
rect 77644 73166 77646 73218
rect 77646 73166 77698 73218
rect 77698 73166 77700 73218
rect 77644 73164 77700 73166
rect 78204 76076 78260 76132
rect 78092 75682 78148 75684
rect 78092 75630 78094 75682
rect 78094 75630 78146 75682
rect 78146 75630 78148 75682
rect 78092 75628 78148 75630
rect 78428 75516 78484 75572
rect 78092 75404 78148 75460
rect 79100 75180 79156 75236
rect 78092 74620 78148 74676
rect 78092 74172 78148 74228
rect 78204 73554 78260 73556
rect 78204 73502 78206 73554
rect 78206 73502 78258 73554
rect 78258 73502 78260 73554
rect 78204 73500 78260 73502
rect 77868 72492 77924 72548
rect 77644 72434 77700 72436
rect 77644 72382 77646 72434
rect 77646 72382 77698 72434
rect 77698 72382 77700 72434
rect 77644 72380 77700 72382
rect 78204 72434 78260 72436
rect 78204 72382 78206 72434
rect 78206 72382 78258 72434
rect 78258 72382 78260 72434
rect 78204 72380 78260 72382
rect 77868 71874 77924 71876
rect 77868 71822 77870 71874
rect 77870 71822 77922 71874
rect 77922 71822 77924 71874
rect 77868 71820 77924 71822
rect 77644 71762 77700 71764
rect 77644 71710 77646 71762
rect 77646 71710 77698 71762
rect 77698 71710 77700 71762
rect 77644 71708 77700 71710
rect 77756 71090 77812 71092
rect 77756 71038 77758 71090
rect 77758 71038 77810 71090
rect 77810 71038 77812 71090
rect 77756 71036 77812 71038
rect 77420 70754 77476 70756
rect 77420 70702 77422 70754
rect 77422 70702 77474 70754
rect 77474 70702 77476 70754
rect 77420 70700 77476 70702
rect 77644 69020 77700 69076
rect 77084 68796 77140 68852
rect 77420 68514 77476 68516
rect 77420 68462 77422 68514
rect 77422 68462 77474 68514
rect 77474 68462 77476 68514
rect 77420 68460 77476 68462
rect 77644 67788 77700 67844
rect 77644 66780 77700 66836
rect 77644 66274 77700 66276
rect 77644 66222 77646 66274
rect 77646 66222 77698 66274
rect 77698 66222 77700 66274
rect 77644 66220 77700 66222
rect 77420 65660 77476 65716
rect 77644 64706 77700 64708
rect 77644 64654 77646 64706
rect 77646 64654 77698 64706
rect 77698 64654 77700 64706
rect 77644 64652 77700 64654
rect 77420 64594 77476 64596
rect 77420 64542 77422 64594
rect 77422 64542 77474 64594
rect 77474 64542 77476 64594
rect 77420 64540 77476 64542
rect 77644 63922 77700 63924
rect 77644 63870 77646 63922
rect 77646 63870 77698 63922
rect 77698 63870 77700 63922
rect 77644 63868 77700 63870
rect 77420 62914 77476 62916
rect 77420 62862 77422 62914
rect 77422 62862 77474 62914
rect 77474 62862 77476 62914
rect 77420 62860 77476 62862
rect 77644 61180 77700 61236
rect 77644 60786 77700 60788
rect 77644 60734 77646 60786
rect 77646 60734 77698 60786
rect 77698 60734 77700 60786
rect 77644 60732 77700 60734
rect 77644 59106 77700 59108
rect 77644 59054 77646 59106
rect 77646 59054 77698 59106
rect 77698 59054 77700 59106
rect 77644 59052 77700 59054
rect 77420 58940 77476 58996
rect 77644 57820 77700 57876
rect 77644 56754 77700 56756
rect 77644 56702 77646 56754
rect 77646 56702 77698 56754
rect 77698 56702 77700 56754
rect 77644 56700 77700 56702
rect 77644 55970 77700 55972
rect 77644 55918 77646 55970
rect 77646 55918 77698 55970
rect 77698 55918 77700 55970
rect 77644 55916 77700 55918
rect 77420 55580 77476 55636
rect 78540 71820 78596 71876
rect 78204 71762 78260 71764
rect 78204 71710 78206 71762
rect 78206 71710 78258 71762
rect 78258 71710 78260 71762
rect 78204 71708 78260 71710
rect 78204 71260 78260 71316
rect 78204 70754 78260 70756
rect 78204 70702 78206 70754
rect 78206 70702 78258 70754
rect 78258 70702 78260 70754
rect 78204 70700 78260 70702
rect 78204 70140 78260 70196
rect 78204 69020 78260 69076
rect 78204 68460 78260 68516
rect 78204 67900 78260 67956
rect 77868 67170 77924 67172
rect 77868 67118 77870 67170
rect 77870 67118 77922 67170
rect 77922 67118 77924 67170
rect 77868 67116 77924 67118
rect 78204 66780 78260 66836
rect 78204 65660 78260 65716
rect 78204 64594 78260 64596
rect 78204 64542 78206 64594
rect 78206 64542 78258 64594
rect 78258 64542 78260 64594
rect 78204 64540 78260 64542
rect 78204 63922 78260 63924
rect 78204 63870 78206 63922
rect 78206 63870 78258 63922
rect 78258 63870 78260 63922
rect 78204 63868 78260 63870
rect 78204 63420 78260 63476
rect 78204 62914 78260 62916
rect 78204 62862 78206 62914
rect 78206 62862 78258 62914
rect 78258 62862 78260 62914
rect 78204 62860 78260 62862
rect 78204 62300 78260 62356
rect 77868 62188 77924 62244
rect 77868 61346 77924 61348
rect 77868 61294 77870 61346
rect 77870 61294 77922 61346
rect 77922 61294 77924 61346
rect 77868 61292 77924 61294
rect 78204 61180 78260 61236
rect 78204 60786 78260 60788
rect 78204 60734 78206 60786
rect 78206 60734 78258 60786
rect 78258 60734 78260 60786
rect 78204 60732 78260 60734
rect 78204 60060 78260 60116
rect 78204 58940 78260 58996
rect 77868 58210 77924 58212
rect 77868 58158 77870 58210
rect 77870 58158 77922 58210
rect 77922 58158 77924 58210
rect 77868 58156 77924 58158
rect 78204 57820 78260 57876
rect 78204 56754 78260 56756
rect 78204 56702 78206 56754
rect 78206 56702 78258 56754
rect 78258 56702 78260 56754
rect 78204 56700 78260 56702
rect 77868 56642 77924 56644
rect 77868 56590 77870 56642
rect 77870 56590 77922 56642
rect 77922 56590 77924 56642
rect 77868 56588 77924 56590
rect 78204 55580 78260 55636
rect 77644 55186 77700 55188
rect 77644 55134 77646 55186
rect 77646 55134 77698 55186
rect 77698 55134 77700 55186
rect 77644 55132 77700 55134
rect 78204 55186 78260 55188
rect 78204 55134 78206 55186
rect 78206 55134 78258 55186
rect 78258 55134 78260 55186
rect 78204 55132 78260 55134
rect 77868 55074 77924 55076
rect 77868 55022 77870 55074
rect 77870 55022 77922 55074
rect 77922 55022 77924 55074
rect 77868 55020 77924 55022
rect 78204 54460 78260 54516
rect 77644 53340 77700 53396
rect 78204 53340 78260 53396
rect 77868 53058 77924 53060
rect 77868 53006 77870 53058
rect 77870 53006 77922 53058
rect 77922 53006 77924 53058
rect 77868 53004 77924 53006
rect 76076 41356 76132 41412
rect 75628 40124 75684 40180
rect 76300 42530 76356 42532
rect 76300 42478 76302 42530
rect 76302 42478 76354 42530
rect 76354 42478 76356 42530
rect 76300 42476 76356 42478
rect 76188 40796 76244 40852
rect 75180 38668 75236 38724
rect 74956 37938 75012 37940
rect 74956 37886 74958 37938
rect 74958 37886 75010 37938
rect 75010 37886 75012 37938
rect 74956 37884 75012 37886
rect 75068 37772 75124 37828
rect 74956 36876 75012 36932
rect 74844 36652 74900 36708
rect 74060 35308 74116 35364
rect 74172 35196 74228 35252
rect 73388 34076 73444 34132
rect 72716 33458 72772 33460
rect 72716 33406 72718 33458
rect 72718 33406 72770 33458
rect 72770 33406 72772 33458
rect 72716 33404 72772 33406
rect 72604 33292 72660 33348
rect 72380 32620 72436 32676
rect 72380 32450 72436 32452
rect 72380 32398 72382 32450
rect 72382 32398 72434 32450
rect 72434 32398 72436 32450
rect 72380 32396 72436 32398
rect 71932 31836 71988 31892
rect 72268 30994 72324 30996
rect 72268 30942 72270 30994
rect 72270 30942 72322 30994
rect 72322 30942 72324 30994
rect 72268 30940 72324 30942
rect 72044 30828 72100 30884
rect 71932 30716 71988 30772
rect 71820 29708 71876 29764
rect 71820 28530 71876 28532
rect 71820 28478 71822 28530
rect 71822 28478 71874 28530
rect 71874 28478 71876 28530
rect 71820 28476 71876 28478
rect 71820 28252 71876 28308
rect 72156 29932 72212 29988
rect 71932 27804 71988 27860
rect 72268 27186 72324 27188
rect 72268 27134 72270 27186
rect 72270 27134 72322 27186
rect 72322 27134 72324 27186
rect 72268 27132 72324 27134
rect 72828 32562 72884 32564
rect 72828 32510 72830 32562
rect 72830 32510 72882 32562
rect 72882 32510 72884 32562
rect 72828 32508 72884 32510
rect 72716 31666 72772 31668
rect 72716 31614 72718 31666
rect 72718 31614 72770 31666
rect 72770 31614 72772 31666
rect 72716 31612 72772 31614
rect 72604 31388 72660 31444
rect 72828 30434 72884 30436
rect 72828 30382 72830 30434
rect 72830 30382 72882 30434
rect 72882 30382 72884 30434
rect 72828 30380 72884 30382
rect 73500 33740 73556 33796
rect 73276 33292 73332 33348
rect 73164 32508 73220 32564
rect 73836 34354 73892 34356
rect 73836 34302 73838 34354
rect 73838 34302 73890 34354
rect 73890 34302 73892 34354
rect 73836 34300 73892 34302
rect 73724 32284 73780 32340
rect 73836 33740 73892 33796
rect 74172 34300 74228 34356
rect 74396 34748 74452 34804
rect 74396 34076 74452 34132
rect 74396 33180 74452 33236
rect 73388 31388 73444 31444
rect 74732 34748 74788 34804
rect 74956 34860 75012 34916
rect 74732 34130 74788 34132
rect 74732 34078 74734 34130
rect 74734 34078 74786 34130
rect 74786 34078 74788 34130
rect 74732 34076 74788 34078
rect 74508 32956 74564 33012
rect 75180 37266 75236 37268
rect 75180 37214 75182 37266
rect 75182 37214 75234 37266
rect 75234 37214 75236 37266
rect 75180 37212 75236 37214
rect 75404 38668 75460 38724
rect 75516 39004 75572 39060
rect 75628 38834 75684 38836
rect 75628 38782 75630 38834
rect 75630 38782 75682 38834
rect 75682 38782 75684 38834
rect 75628 38780 75684 38782
rect 75516 38108 75572 38164
rect 75404 37772 75460 37828
rect 75516 37660 75572 37716
rect 75404 36482 75460 36484
rect 75404 36430 75406 36482
rect 75406 36430 75458 36482
rect 75458 36430 75460 36482
rect 75404 36428 75460 36430
rect 75292 35756 75348 35812
rect 75404 35420 75460 35476
rect 75964 38668 76020 38724
rect 76524 41804 76580 41860
rect 76524 41244 76580 41300
rect 76636 41020 76692 41076
rect 76748 40572 76804 40628
rect 76412 39900 76468 39956
rect 76524 39618 76580 39620
rect 76524 39566 76526 39618
rect 76526 39566 76578 39618
rect 76578 39566 76580 39618
rect 76524 39564 76580 39566
rect 75852 38444 75908 38500
rect 75852 36540 75908 36596
rect 76412 38556 76468 38612
rect 76524 38444 76580 38500
rect 76188 38220 76244 38276
rect 76188 38050 76244 38052
rect 76188 37998 76190 38050
rect 76190 37998 76242 38050
rect 76242 37998 76244 38050
rect 76188 37996 76244 37998
rect 76636 38220 76692 38276
rect 78204 52220 78260 52276
rect 77420 48524 77476 48580
rect 77644 51100 77700 51156
rect 78204 51100 78260 51156
rect 77644 50482 77700 50484
rect 77644 50430 77646 50482
rect 77646 50430 77698 50482
rect 77698 50430 77700 50482
rect 77644 50428 77700 50430
rect 78204 50482 78260 50484
rect 78204 50430 78206 50482
rect 78206 50430 78258 50482
rect 78258 50430 78260 50482
rect 78204 50428 78260 50430
rect 77868 50370 77924 50372
rect 77868 50318 77870 50370
rect 77870 50318 77922 50370
rect 77922 50318 77924 50370
rect 77868 50316 77924 50318
rect 78204 49980 78260 50036
rect 77644 48914 77700 48916
rect 77644 48862 77646 48914
rect 77646 48862 77698 48914
rect 77698 48862 77700 48914
rect 77644 48860 77700 48862
rect 78204 48914 78260 48916
rect 78204 48862 78206 48914
rect 78206 48862 78258 48914
rect 78258 48862 78260 48914
rect 78204 48860 78260 48862
rect 77868 48802 77924 48804
rect 77868 48750 77870 48802
rect 77870 48750 77922 48802
rect 77922 48750 77924 48802
rect 77868 48748 77924 48750
rect 77644 48242 77700 48244
rect 77644 48190 77646 48242
rect 77646 48190 77698 48242
rect 77698 48190 77700 48242
rect 77644 48188 77700 48190
rect 77644 47234 77700 47236
rect 77644 47182 77646 47234
rect 77646 47182 77698 47234
rect 77698 47182 77700 47234
rect 77644 47180 77700 47182
rect 77644 45500 77700 45556
rect 77420 45276 77476 45332
rect 77644 44994 77700 44996
rect 77644 44942 77646 44994
rect 77646 44942 77698 44994
rect 77698 44942 77700 44994
rect 77644 44940 77700 44942
rect 77420 43538 77476 43540
rect 77420 43486 77422 43538
rect 77422 43486 77474 43538
rect 77474 43486 77476 43538
rect 77420 43484 77476 43486
rect 76972 41356 77028 41412
rect 76748 38108 76804 38164
rect 76188 37266 76244 37268
rect 76188 37214 76190 37266
rect 76190 37214 76242 37266
rect 76242 37214 76244 37266
rect 76188 37212 76244 37214
rect 76636 37772 76692 37828
rect 76636 37324 76692 37380
rect 75740 35698 75796 35700
rect 75740 35646 75742 35698
rect 75742 35646 75794 35698
rect 75794 35646 75796 35698
rect 75740 35644 75796 35646
rect 75628 34860 75684 34916
rect 74956 33852 75012 33908
rect 74732 32732 74788 32788
rect 74956 32674 75012 32676
rect 74956 32622 74958 32674
rect 74958 32622 75010 32674
rect 75010 32622 75012 32674
rect 74956 32620 75012 32622
rect 74060 32060 74116 32116
rect 74508 32284 74564 32340
rect 73948 31948 74004 32004
rect 73724 31554 73780 31556
rect 73724 31502 73726 31554
rect 73726 31502 73778 31554
rect 73778 31502 73780 31554
rect 73724 31500 73780 31502
rect 72492 28812 72548 28868
rect 72828 28700 72884 28756
rect 72604 28588 72660 28644
rect 72492 28364 72548 28420
rect 72716 28476 72772 28532
rect 73500 29426 73556 29428
rect 73500 29374 73502 29426
rect 73502 29374 73554 29426
rect 73554 29374 73556 29426
rect 73500 29372 73556 29374
rect 72828 28028 72884 28084
rect 73500 28754 73556 28756
rect 73500 28702 73502 28754
rect 73502 28702 73554 28754
rect 73554 28702 73556 28754
rect 73500 28700 73556 28702
rect 72716 27580 72772 27636
rect 72716 27020 72772 27076
rect 72492 26514 72548 26516
rect 72492 26462 72494 26514
rect 72494 26462 72546 26514
rect 72546 26462 72548 26514
rect 72492 26460 72548 26462
rect 72604 25900 72660 25956
rect 72604 25676 72660 25732
rect 71932 25452 71988 25508
rect 71596 25228 71652 25284
rect 71708 25116 71764 25172
rect 71820 25004 71876 25060
rect 71372 24610 71428 24612
rect 71372 24558 71374 24610
rect 71374 24558 71426 24610
rect 71426 24558 71428 24610
rect 71372 24556 71428 24558
rect 71820 23884 71876 23940
rect 71708 23378 71764 23380
rect 71708 23326 71710 23378
rect 71710 23326 71762 23378
rect 71762 23326 71764 23378
rect 71708 23324 71764 23326
rect 71820 23212 71876 23268
rect 72156 25116 72212 25172
rect 72268 25004 72324 25060
rect 72156 23938 72212 23940
rect 72156 23886 72158 23938
rect 72158 23886 72210 23938
rect 72210 23886 72212 23938
rect 72156 23884 72212 23886
rect 72044 23100 72100 23156
rect 72156 23324 72212 23380
rect 72380 23548 72436 23604
rect 72492 23772 72548 23828
rect 71932 22482 71988 22484
rect 71932 22430 71934 22482
rect 71934 22430 71986 22482
rect 71986 22430 71988 22482
rect 71932 22428 71988 22430
rect 72268 22204 72324 22260
rect 71708 21698 71764 21700
rect 71708 21646 71710 21698
rect 71710 21646 71762 21698
rect 71762 21646 71764 21698
rect 71708 21644 71764 21646
rect 72156 21644 72212 21700
rect 71260 20914 71316 20916
rect 71260 20862 71262 20914
rect 71262 20862 71314 20914
rect 71314 20862 71316 20914
rect 71260 20860 71316 20862
rect 72268 20690 72324 20692
rect 72268 20638 72270 20690
rect 72270 20638 72322 20690
rect 72322 20638 72324 20690
rect 72268 20636 72324 20638
rect 72716 24668 72772 24724
rect 73164 27858 73220 27860
rect 73164 27806 73166 27858
rect 73166 27806 73218 27858
rect 73218 27806 73220 27858
rect 73164 27804 73220 27806
rect 73164 27074 73220 27076
rect 73164 27022 73166 27074
rect 73166 27022 73218 27074
rect 73218 27022 73220 27074
rect 73164 27020 73220 27022
rect 73724 29372 73780 29428
rect 73724 28642 73780 28644
rect 73724 28590 73726 28642
rect 73726 28590 73778 28642
rect 73778 28590 73780 28642
rect 73724 28588 73780 28590
rect 74060 31218 74116 31220
rect 74060 31166 74062 31218
rect 74062 31166 74114 31218
rect 74114 31166 74116 31218
rect 74060 31164 74116 31166
rect 74172 31106 74228 31108
rect 74172 31054 74174 31106
rect 74174 31054 74226 31106
rect 74226 31054 74228 31106
rect 74172 31052 74228 31054
rect 73948 30492 74004 30548
rect 74284 30380 74340 30436
rect 74396 29932 74452 29988
rect 74060 29202 74116 29204
rect 74060 29150 74062 29202
rect 74062 29150 74114 29202
rect 74114 29150 74116 29202
rect 74060 29148 74116 29150
rect 74396 28812 74452 28868
rect 73836 28476 73892 28532
rect 73948 28140 74004 28196
rect 73724 28028 73780 28084
rect 73724 27692 73780 27748
rect 73500 27074 73556 27076
rect 73500 27022 73502 27074
rect 73502 27022 73554 27074
rect 73554 27022 73556 27074
rect 73500 27020 73556 27022
rect 74060 27074 74116 27076
rect 74060 27022 74062 27074
rect 74062 27022 74114 27074
rect 74114 27022 74116 27074
rect 74060 27020 74116 27022
rect 72940 26684 72996 26740
rect 73276 26460 73332 26516
rect 73164 26178 73220 26180
rect 73164 26126 73166 26178
rect 73166 26126 73218 26178
rect 73218 26126 73220 26178
rect 73164 26124 73220 26126
rect 72940 25618 72996 25620
rect 72940 25566 72942 25618
rect 72942 25566 72994 25618
rect 72994 25566 72996 25618
rect 72940 25564 72996 25566
rect 72940 25228 72996 25284
rect 72716 23938 72772 23940
rect 72716 23886 72718 23938
rect 72718 23886 72770 23938
rect 72770 23886 72772 23938
rect 72716 23884 72772 23886
rect 73500 25900 73556 25956
rect 74060 26796 74116 26852
rect 73836 26460 73892 26516
rect 74396 28140 74452 28196
rect 74284 27692 74340 27748
rect 74284 26684 74340 26740
rect 73724 24780 73780 24836
rect 74060 24892 74116 24948
rect 73612 24668 73668 24724
rect 73500 24556 73556 24612
rect 73164 24050 73220 24052
rect 73164 23998 73166 24050
rect 73166 23998 73218 24050
rect 73218 23998 73220 24050
rect 73164 23996 73220 23998
rect 73276 23938 73332 23940
rect 73276 23886 73278 23938
rect 73278 23886 73330 23938
rect 73330 23886 73332 23938
rect 73276 23884 73332 23886
rect 73388 21868 73444 21924
rect 74060 24162 74116 24164
rect 74060 24110 74062 24162
rect 74062 24110 74114 24162
rect 74114 24110 74116 24162
rect 74060 24108 74116 24110
rect 73836 23996 73892 24052
rect 73948 23212 74004 23268
rect 74060 22930 74116 22932
rect 74060 22878 74062 22930
rect 74062 22878 74114 22930
rect 74114 22878 74116 22930
rect 74060 22876 74116 22878
rect 74060 22370 74116 22372
rect 74060 22318 74062 22370
rect 74062 22318 74114 22370
rect 74114 22318 74116 22370
rect 74060 22316 74116 22318
rect 75292 33964 75348 34020
rect 75740 34636 75796 34692
rect 75740 34300 75796 34356
rect 75628 33516 75684 33572
rect 75180 33180 75236 33236
rect 76412 35980 76468 36036
rect 77308 42642 77364 42644
rect 77308 42590 77310 42642
rect 77310 42590 77362 42642
rect 77362 42590 77364 42642
rect 77308 42588 77364 42590
rect 77308 42252 77364 42308
rect 77196 39788 77252 39844
rect 77532 41186 77588 41188
rect 77532 41134 77534 41186
rect 77534 41134 77586 41186
rect 77586 41134 77588 41186
rect 77532 41132 77588 41134
rect 77420 40572 77476 40628
rect 78204 48242 78260 48244
rect 78204 48190 78206 48242
rect 78206 48190 78258 48242
rect 78258 48190 78260 48242
rect 78204 48188 78260 48190
rect 78204 47740 78260 47796
rect 78204 47180 78260 47236
rect 78204 46620 78260 46676
rect 77868 45836 77924 45892
rect 77868 45666 77924 45668
rect 77868 45614 77870 45666
rect 77870 45614 77922 45666
rect 77922 45614 77924 45666
rect 77868 45612 77924 45614
rect 78204 45500 78260 45556
rect 78204 44940 78260 44996
rect 78204 44380 78260 44436
rect 78204 43426 78260 43428
rect 78204 43374 78206 43426
rect 78206 43374 78258 43426
rect 78258 43374 78260 43426
rect 78204 43372 78260 43374
rect 78092 43260 78148 43316
rect 77980 42140 78036 42196
rect 78092 41298 78148 41300
rect 78092 41246 78094 41298
rect 78094 41246 78146 41298
rect 78146 41246 78148 41298
rect 78092 41244 78148 41246
rect 77868 40684 77924 40740
rect 77980 40572 78036 40628
rect 77196 38668 77252 38724
rect 77196 38444 77252 38500
rect 77308 38332 77364 38388
rect 77308 37436 77364 37492
rect 77644 39788 77700 39844
rect 78092 40124 78148 40180
rect 77644 38946 77700 38948
rect 77644 38894 77646 38946
rect 77646 38894 77698 38946
rect 77698 38894 77700 38946
rect 77644 38892 77700 38894
rect 77756 38780 77812 38836
rect 77644 38220 77700 38276
rect 77644 37324 77700 37380
rect 77308 36652 77364 36708
rect 77420 36092 77476 36148
rect 76860 35810 76916 35812
rect 76860 35758 76862 35810
rect 76862 35758 76914 35810
rect 76914 35758 76916 35810
rect 76860 35756 76916 35758
rect 76748 35420 76804 35476
rect 76524 34524 76580 34580
rect 76636 34412 76692 34468
rect 75964 34354 76020 34356
rect 75964 34302 75966 34354
rect 75966 34302 76018 34354
rect 76018 34302 76020 34354
rect 75964 34300 76020 34302
rect 75852 33068 75908 33124
rect 76300 34242 76356 34244
rect 76300 34190 76302 34242
rect 76302 34190 76354 34242
rect 76354 34190 76356 34242
rect 76300 34188 76356 34190
rect 76412 34130 76468 34132
rect 76412 34078 76414 34130
rect 76414 34078 76466 34130
rect 76466 34078 76468 34130
rect 76412 34076 76468 34078
rect 76972 34076 77028 34132
rect 76860 33852 76916 33908
rect 76524 33458 76580 33460
rect 76524 33406 76526 33458
rect 76526 33406 76578 33458
rect 76578 33406 76580 33458
rect 76524 33404 76580 33406
rect 75180 32620 75236 32676
rect 75740 32620 75796 32676
rect 75068 32172 75124 32228
rect 75292 32396 75348 32452
rect 74844 32060 74900 32116
rect 74732 31890 74788 31892
rect 74732 31838 74734 31890
rect 74734 31838 74786 31890
rect 74786 31838 74788 31890
rect 74732 31836 74788 31838
rect 75180 31948 75236 32004
rect 75068 31778 75124 31780
rect 75068 31726 75070 31778
rect 75070 31726 75122 31778
rect 75122 31726 75124 31778
rect 75068 31724 75124 31726
rect 75292 31836 75348 31892
rect 75180 30940 75236 30996
rect 74620 30716 74676 30772
rect 75404 31276 75460 31332
rect 75740 31276 75796 31332
rect 75404 30940 75460 30996
rect 75628 30882 75684 30884
rect 75628 30830 75630 30882
rect 75630 30830 75682 30882
rect 75682 30830 75684 30882
rect 75628 30828 75684 30830
rect 75516 30044 75572 30100
rect 74732 28924 74788 28980
rect 74732 28588 74788 28644
rect 75068 28812 75124 28868
rect 75180 28364 75236 28420
rect 74956 27916 75012 27972
rect 74732 27692 74788 27748
rect 74620 27132 74676 27188
rect 74732 26908 74788 26964
rect 74956 27020 75012 27076
rect 74620 26572 74676 26628
rect 74620 26402 74676 26404
rect 74620 26350 74622 26402
rect 74622 26350 74674 26402
rect 74674 26350 74676 26402
rect 74620 26348 74676 26350
rect 74732 26124 74788 26180
rect 74508 24050 74564 24052
rect 74508 23998 74510 24050
rect 74510 23998 74562 24050
rect 74562 23998 74564 24050
rect 74508 23996 74564 23998
rect 74396 23938 74452 23940
rect 74396 23886 74398 23938
rect 74398 23886 74450 23938
rect 74450 23886 74452 23938
rect 74396 23884 74452 23886
rect 74956 23548 75012 23604
rect 74284 22594 74340 22596
rect 74284 22542 74286 22594
rect 74286 22542 74338 22594
rect 74338 22542 74340 22594
rect 74284 22540 74340 22542
rect 73500 21420 73556 21476
rect 73276 20972 73332 21028
rect 72716 20076 72772 20132
rect 74060 20690 74116 20692
rect 74060 20638 74062 20690
rect 74062 20638 74114 20690
rect 74114 20638 74116 20690
rect 74060 20636 74116 20638
rect 73836 19292 73892 19348
rect 74284 18844 74340 18900
rect 75628 29596 75684 29652
rect 75628 29426 75684 29428
rect 75628 29374 75630 29426
rect 75630 29374 75682 29426
rect 75682 29374 75684 29426
rect 75628 29372 75684 29374
rect 75516 28924 75572 28980
rect 75404 28418 75460 28420
rect 75404 28366 75406 28418
rect 75406 28366 75458 28418
rect 75458 28366 75460 28418
rect 75404 28364 75460 28366
rect 75292 27074 75348 27076
rect 75292 27022 75294 27074
rect 75294 27022 75346 27074
rect 75346 27022 75348 27074
rect 75292 27020 75348 27022
rect 75628 28476 75684 28532
rect 76076 32450 76132 32452
rect 76076 32398 76078 32450
rect 76078 32398 76130 32450
rect 76130 32398 76132 32450
rect 76076 32396 76132 32398
rect 76412 31778 76468 31780
rect 76412 31726 76414 31778
rect 76414 31726 76466 31778
rect 76466 31726 76468 31778
rect 76412 31724 76468 31726
rect 76300 31554 76356 31556
rect 76300 31502 76302 31554
rect 76302 31502 76354 31554
rect 76354 31502 76356 31554
rect 76300 31500 76356 31502
rect 76860 32674 76916 32676
rect 76860 32622 76862 32674
rect 76862 32622 76914 32674
rect 76914 32622 76916 32674
rect 76860 32620 76916 32622
rect 77084 34188 77140 34244
rect 77084 33234 77140 33236
rect 77084 33182 77086 33234
rect 77086 33182 77138 33234
rect 77138 33182 77140 33234
rect 77084 33180 77140 33182
rect 77644 36988 77700 37044
rect 77644 36540 77700 36596
rect 77980 38108 78036 38164
rect 77868 36876 77924 36932
rect 77868 35868 77924 35924
rect 77980 35756 78036 35812
rect 77308 34972 77364 35028
rect 77308 34018 77364 34020
rect 77308 33966 77310 34018
rect 77310 33966 77362 34018
rect 77362 33966 77364 34018
rect 77308 33964 77364 33966
rect 76748 31164 76804 31220
rect 76860 31276 76916 31332
rect 77868 35138 77924 35140
rect 77868 35086 77870 35138
rect 77870 35086 77922 35138
rect 77922 35086 77924 35138
rect 77868 35084 77924 35086
rect 77532 34972 77588 35028
rect 77532 34524 77588 34580
rect 77644 34130 77700 34132
rect 77644 34078 77646 34130
rect 77646 34078 77698 34130
rect 77698 34078 77700 34130
rect 77644 34076 77700 34078
rect 77868 33516 77924 33572
rect 78316 36764 78372 36820
rect 78316 35420 78372 35476
rect 78204 34914 78260 34916
rect 78204 34862 78206 34914
rect 78206 34862 78258 34914
rect 78258 34862 78260 34914
rect 78204 34860 78260 34862
rect 78092 34412 78148 34468
rect 77532 32002 77588 32004
rect 77532 31950 77534 32002
rect 77534 31950 77586 32002
rect 77586 31950 77588 32002
rect 77532 31948 77588 31950
rect 77532 31724 77588 31780
rect 77868 32172 77924 32228
rect 77308 31218 77364 31220
rect 77308 31166 77310 31218
rect 77310 31166 77362 31218
rect 77362 31166 77364 31218
rect 77308 31164 77364 31166
rect 76412 30268 76468 30324
rect 76076 30044 76132 30100
rect 76300 29986 76356 29988
rect 76300 29934 76302 29986
rect 76302 29934 76354 29986
rect 76354 29934 76356 29986
rect 76300 29932 76356 29934
rect 76076 29538 76132 29540
rect 76076 29486 76078 29538
rect 76078 29486 76130 29538
rect 76130 29486 76132 29538
rect 76076 29484 76132 29486
rect 75964 29372 76020 29428
rect 76076 28642 76132 28644
rect 76076 28590 76078 28642
rect 76078 28590 76130 28642
rect 76130 28590 76132 28642
rect 76076 28588 76132 28590
rect 75852 27970 75908 27972
rect 75852 27918 75854 27970
rect 75854 27918 75906 27970
rect 75906 27918 75908 27970
rect 75852 27916 75908 27918
rect 76524 30098 76580 30100
rect 76524 30046 76526 30098
rect 76526 30046 76578 30098
rect 76578 30046 76580 30098
rect 76524 30044 76580 30046
rect 77308 30044 77364 30100
rect 76972 29708 77028 29764
rect 76524 29484 76580 29540
rect 76524 28642 76580 28644
rect 76524 28590 76526 28642
rect 76526 28590 76578 28642
rect 76578 28590 76580 28642
rect 76524 28588 76580 28590
rect 77084 28588 77140 28644
rect 76636 28364 76692 28420
rect 76748 27804 76804 27860
rect 76860 27580 76916 27636
rect 76524 27468 76580 27524
rect 76860 27298 76916 27300
rect 76860 27246 76862 27298
rect 76862 27246 76914 27298
rect 76914 27246 76916 27298
rect 76860 27244 76916 27246
rect 76188 26962 76244 26964
rect 76188 26910 76190 26962
rect 76190 26910 76242 26962
rect 76242 26910 76244 26962
rect 76188 26908 76244 26910
rect 75404 25340 75460 25396
rect 75180 24722 75236 24724
rect 75180 24670 75182 24722
rect 75182 24670 75234 24722
rect 75234 24670 75236 24722
rect 75180 24668 75236 24670
rect 75292 24050 75348 24052
rect 75292 23998 75294 24050
rect 75294 23998 75346 24050
rect 75346 23998 75348 24050
rect 75292 23996 75348 23998
rect 74956 21586 75012 21588
rect 74956 21534 74958 21586
rect 74958 21534 75010 21586
rect 75010 21534 75012 21586
rect 74956 21532 75012 21534
rect 74732 20188 74788 20244
rect 75068 20130 75124 20132
rect 75068 20078 75070 20130
rect 75070 20078 75122 20130
rect 75122 20078 75124 20130
rect 75068 20076 75124 20078
rect 74844 19740 74900 19796
rect 74620 18060 74676 18116
rect 72156 16940 72212 16996
rect 75292 21420 75348 21476
rect 75404 20972 75460 21028
rect 75404 19906 75460 19908
rect 75404 19854 75406 19906
rect 75406 19854 75458 19906
rect 75458 19854 75460 19906
rect 75404 19852 75460 19854
rect 75404 19010 75460 19012
rect 75404 18958 75406 19010
rect 75406 18958 75458 19010
rect 75458 18958 75460 19010
rect 75404 18956 75460 18958
rect 75292 17388 75348 17444
rect 71036 16268 71092 16324
rect 70252 16156 70308 16212
rect 69692 15148 69748 15204
rect 71372 14364 71428 14420
rect 69692 6636 69748 6692
rect 69804 9324 69860 9380
rect 69244 6524 69300 6580
rect 69356 6466 69412 6468
rect 69356 6414 69358 6466
rect 69358 6414 69410 6466
rect 69410 6414 69412 6466
rect 69356 6412 69412 6414
rect 69244 6300 69300 6356
rect 68572 6076 68628 6132
rect 68348 4114 68404 4116
rect 68348 4062 68350 4114
rect 68350 4062 68402 4114
rect 68402 4062 68404 4114
rect 68348 4060 68404 4062
rect 68796 3836 68852 3892
rect 69356 5346 69412 5348
rect 69356 5294 69358 5346
rect 69358 5294 69410 5346
rect 69410 5294 69412 5346
rect 69356 5292 69412 5294
rect 68908 3500 68964 3556
rect 69468 3724 69524 3780
rect 71260 6690 71316 6692
rect 71260 6638 71262 6690
rect 71262 6638 71314 6690
rect 71314 6638 71316 6690
rect 71260 6636 71316 6638
rect 70476 6412 70532 6468
rect 70476 5794 70532 5796
rect 70476 5742 70478 5794
rect 70478 5742 70530 5794
rect 70530 5742 70532 5794
rect 70476 5740 70532 5742
rect 70476 5292 70532 5348
rect 70812 5628 70868 5684
rect 70476 3948 70532 4004
rect 73052 12684 73108 12740
rect 71708 7756 71764 7812
rect 72380 7756 72436 7812
rect 72268 6466 72324 6468
rect 72268 6414 72270 6466
rect 72270 6414 72322 6466
rect 72322 6414 72324 6466
rect 72268 6412 72324 6414
rect 71708 5906 71764 5908
rect 71708 5854 71710 5906
rect 71710 5854 71762 5906
rect 71762 5854 71764 5906
rect 71708 5852 71764 5854
rect 72268 5906 72324 5908
rect 72268 5854 72270 5906
rect 72270 5854 72322 5906
rect 72322 5854 72324 5906
rect 72268 5852 72324 5854
rect 72828 5740 72884 5796
rect 72268 5234 72324 5236
rect 72268 5182 72270 5234
rect 72270 5182 72322 5234
rect 72322 5182 72324 5234
rect 72268 5180 72324 5182
rect 72156 5068 72212 5124
rect 71708 4562 71764 4564
rect 71708 4510 71710 4562
rect 71710 4510 71762 4562
rect 71762 4510 71764 4562
rect 71708 4508 71764 4510
rect 71484 4060 71540 4116
rect 71260 3666 71316 3668
rect 71260 3614 71262 3666
rect 71262 3614 71314 3666
rect 71314 3614 71316 3666
rect 71260 3612 71316 3614
rect 72268 4508 72324 4564
rect 73612 8316 73668 8372
rect 73612 6188 73668 6244
rect 73276 5682 73332 5684
rect 73276 5630 73278 5682
rect 73278 5630 73330 5682
rect 73330 5630 73332 5682
rect 73276 5628 73332 5630
rect 73052 4172 73108 4228
rect 73500 5180 73556 5236
rect 73276 3836 73332 3892
rect 76188 26514 76244 26516
rect 76188 26462 76190 26514
rect 76190 26462 76242 26514
rect 76242 26462 76244 26514
rect 76188 26460 76244 26462
rect 75740 25116 75796 25172
rect 75852 26124 75908 26180
rect 75628 24892 75684 24948
rect 76972 25788 77028 25844
rect 77196 27298 77252 27300
rect 77196 27246 77198 27298
rect 77198 27246 77250 27298
rect 77250 27246 77252 27298
rect 77196 27244 77252 27246
rect 77532 30492 77588 30548
rect 77644 30380 77700 30436
rect 78204 34354 78260 34356
rect 78204 34302 78206 34354
rect 78206 34302 78258 34354
rect 78258 34302 78260 34354
rect 78204 34300 78260 34302
rect 78204 33458 78260 33460
rect 78204 33406 78206 33458
rect 78206 33406 78258 33458
rect 78258 33406 78260 33458
rect 78204 33404 78260 33406
rect 78092 31164 78148 31220
rect 78540 38332 78596 38388
rect 78540 37436 78596 37492
rect 78652 35756 78708 35812
rect 78876 71036 78932 71092
rect 78764 34412 78820 34468
rect 78876 64652 78932 64708
rect 78540 33404 78596 33460
rect 77868 29820 77924 29876
rect 77756 29650 77812 29652
rect 77756 29598 77758 29650
rect 77758 29598 77810 29650
rect 77810 29598 77812 29650
rect 77756 29596 77812 29598
rect 77420 28924 77476 28980
rect 77420 28252 77476 28308
rect 77644 28642 77700 28644
rect 77644 28590 77646 28642
rect 77646 28590 77698 28642
rect 77698 28590 77700 28642
rect 77644 28588 77700 28590
rect 77868 28476 77924 28532
rect 77756 27970 77812 27972
rect 77756 27918 77758 27970
rect 77758 27918 77810 27970
rect 77810 27918 77812 27970
rect 77756 27916 77812 27918
rect 77532 27244 77588 27300
rect 77420 27020 77476 27076
rect 76524 25452 76580 25508
rect 78092 30716 78148 30772
rect 78428 32620 78484 32676
rect 78204 30210 78260 30212
rect 78204 30158 78206 30210
rect 78206 30158 78258 30210
rect 78258 30158 78260 30210
rect 78204 30156 78260 30158
rect 78204 29036 78260 29092
rect 78540 33180 78596 33236
rect 78540 30156 78596 30212
rect 78988 50316 79044 50372
rect 78988 48748 79044 48804
rect 78988 35196 79044 35252
rect 79324 34972 79380 35028
rect 79436 38332 79492 38388
rect 79100 33516 79156 33572
rect 78876 30044 78932 30100
rect 79100 28924 79156 28980
rect 77868 27074 77924 27076
rect 77868 27022 77870 27074
rect 77870 27022 77922 27074
rect 77922 27022 77924 27074
rect 77868 27020 77924 27022
rect 78204 27580 78260 27636
rect 77756 26684 77812 26740
rect 77644 26290 77700 26292
rect 77644 26238 77646 26290
rect 77646 26238 77698 26290
rect 77698 26238 77700 26290
rect 77644 26236 77700 26238
rect 77420 25506 77476 25508
rect 77420 25454 77422 25506
rect 77422 25454 77474 25506
rect 77474 25454 77476 25506
rect 77420 25452 77476 25454
rect 76188 25228 76244 25284
rect 75628 24668 75684 24724
rect 75740 24444 75796 24500
rect 75740 24220 75796 24276
rect 76524 25004 76580 25060
rect 76524 24668 76580 24724
rect 76412 24444 76468 24500
rect 76188 23826 76244 23828
rect 76188 23774 76190 23826
rect 76190 23774 76242 23826
rect 76242 23774 76244 23826
rect 76188 23772 76244 23774
rect 76188 23436 76244 23492
rect 75740 21980 75796 22036
rect 76300 21980 76356 22036
rect 76076 21698 76132 21700
rect 76076 21646 76078 21698
rect 76078 21646 76130 21698
rect 76130 21646 76132 21698
rect 76076 21644 76132 21646
rect 75740 21586 75796 21588
rect 75740 21534 75742 21586
rect 75742 21534 75794 21586
rect 75794 21534 75796 21586
rect 75740 21532 75796 21534
rect 75740 19964 75796 20020
rect 75964 19852 76020 19908
rect 75964 19068 76020 19124
rect 76076 19292 76132 19348
rect 75628 16940 75684 16996
rect 74620 14700 74676 14756
rect 76300 21644 76356 21700
rect 76860 24498 76916 24500
rect 76860 24446 76862 24498
rect 76862 24446 76914 24498
rect 76914 24446 76916 24498
rect 76860 24444 76916 24446
rect 77644 26012 77700 26068
rect 77084 25116 77140 25172
rect 77868 25788 77924 25844
rect 78204 25676 78260 25732
rect 77756 24892 77812 24948
rect 76748 23772 76804 23828
rect 77644 24668 77700 24724
rect 77196 23548 77252 23604
rect 77644 23714 77700 23716
rect 77644 23662 77646 23714
rect 77646 23662 77698 23714
rect 77698 23662 77700 23714
rect 77644 23660 77700 23662
rect 76860 22988 76916 23044
rect 76636 21698 76692 21700
rect 76636 21646 76638 21698
rect 76638 21646 76690 21698
rect 76690 21646 76692 21698
rect 76636 21644 76692 21646
rect 76524 21026 76580 21028
rect 76524 20974 76526 21026
rect 76526 20974 76578 21026
rect 76578 20974 76580 21026
rect 76524 20972 76580 20974
rect 76412 20412 76468 20468
rect 77644 23100 77700 23156
rect 77868 22092 77924 22148
rect 77868 21756 77924 21812
rect 77756 21698 77812 21700
rect 77756 21646 77758 21698
rect 77758 21646 77810 21698
rect 77810 21646 77812 21698
rect 77756 21644 77812 21646
rect 78540 24220 78596 24276
rect 78316 23436 78372 23492
rect 76412 19964 76468 20020
rect 76524 19292 76580 19348
rect 78204 23100 78260 23156
rect 77308 20914 77364 20916
rect 77308 20862 77310 20914
rect 77310 20862 77362 20914
rect 77362 20862 77364 20914
rect 77308 20860 77364 20862
rect 76860 19964 76916 20020
rect 77532 20802 77588 20804
rect 77532 20750 77534 20802
rect 77534 20750 77586 20802
rect 77586 20750 77588 20802
rect 77532 20748 77588 20750
rect 77980 20860 78036 20916
rect 76972 20188 77028 20244
rect 76524 19122 76580 19124
rect 76524 19070 76526 19122
rect 76526 19070 76578 19122
rect 76578 19070 76580 19122
rect 76524 19068 76580 19070
rect 76748 18956 76804 19012
rect 76636 18844 76692 18900
rect 76748 18674 76804 18676
rect 76748 18622 76750 18674
rect 76750 18622 76802 18674
rect 76802 18622 76804 18674
rect 76748 18620 76804 18622
rect 76524 18508 76580 18564
rect 76972 17554 77028 17556
rect 76972 17502 76974 17554
rect 76974 17502 77026 17554
rect 77026 17502 77028 17554
rect 76972 17500 77028 17502
rect 77196 18844 77252 18900
rect 77644 20130 77700 20132
rect 77644 20078 77646 20130
rect 77646 20078 77698 20130
rect 77698 20078 77700 20130
rect 77644 20076 77700 20078
rect 77420 20018 77476 20020
rect 77420 19966 77422 20018
rect 77422 19966 77474 20018
rect 77474 19966 77476 20018
rect 77420 19964 77476 19966
rect 77644 19906 77700 19908
rect 77644 19854 77646 19906
rect 77646 19854 77698 19906
rect 77698 19854 77700 19906
rect 77644 19852 77700 19854
rect 77532 19122 77588 19124
rect 77532 19070 77534 19122
rect 77534 19070 77586 19122
rect 77586 19070 77588 19122
rect 77532 19068 77588 19070
rect 77980 19068 78036 19124
rect 78092 20748 78148 20804
rect 77868 19010 77924 19012
rect 77868 18958 77870 19010
rect 77870 18958 77922 19010
rect 77922 18958 77924 19010
rect 77868 18956 77924 18958
rect 78428 21980 78484 22036
rect 78204 19234 78260 19236
rect 78204 19182 78206 19234
rect 78206 19182 78258 19234
rect 78258 19182 78260 19234
rect 78204 19180 78260 19182
rect 78204 18844 78260 18900
rect 77532 18620 77588 18676
rect 78204 18620 78260 18676
rect 77420 18562 77476 18564
rect 77420 18510 77422 18562
rect 77422 18510 77474 18562
rect 77474 18510 77476 18562
rect 77420 18508 77476 18510
rect 77756 18450 77812 18452
rect 77756 18398 77758 18450
rect 77758 18398 77810 18450
rect 77810 18398 77812 18450
rect 77756 18396 77812 18398
rect 77756 18226 77812 18228
rect 77756 18174 77758 18226
rect 77758 18174 77810 18226
rect 77810 18174 77812 18226
rect 77756 18172 77812 18174
rect 77644 17612 77700 17668
rect 77532 17554 77588 17556
rect 77532 17502 77534 17554
rect 77534 17502 77586 17554
rect 77586 17502 77588 17554
rect 77532 17500 77588 17502
rect 77308 17276 77364 17332
rect 77532 17164 77588 17220
rect 77308 16940 77364 16996
rect 77196 16882 77252 16884
rect 77196 16830 77198 16882
rect 77198 16830 77250 16882
rect 77250 16830 77252 16882
rect 77196 16828 77252 16830
rect 77308 14364 77364 14420
rect 77420 16716 77476 16772
rect 76300 13916 76356 13972
rect 76076 13468 76132 13524
rect 75180 12348 75236 12404
rect 75964 12402 76020 12404
rect 75964 12350 75966 12402
rect 75966 12350 76018 12402
rect 76018 12350 76020 12402
rect 75964 12348 76020 12350
rect 75516 11340 75572 11396
rect 75292 9602 75348 9604
rect 75292 9550 75294 9602
rect 75294 9550 75346 9602
rect 75346 9550 75348 9602
rect 75292 9548 75348 9550
rect 75292 9324 75348 9380
rect 74060 8092 74116 8148
rect 73948 5068 74004 5124
rect 73612 3442 73668 3444
rect 73612 3390 73614 3442
rect 73614 3390 73666 3442
rect 73666 3390 73668 3442
rect 73612 3388 73668 3390
rect 74172 4172 74228 4228
rect 74060 3948 74116 4004
rect 74060 2940 74116 2996
rect 74732 7644 74788 7700
rect 74956 6524 75012 6580
rect 75628 8204 75684 8260
rect 75292 7644 75348 7700
rect 75180 6860 75236 6916
rect 76188 9324 76244 9380
rect 76412 11394 76468 11396
rect 76412 11342 76414 11394
rect 76414 11342 76466 11394
rect 76466 11342 76468 11394
rect 76412 11340 76468 11342
rect 75292 6748 75348 6804
rect 75068 5404 75124 5460
rect 75180 5292 75236 5348
rect 74620 924 74676 980
rect 75068 3778 75124 3780
rect 75068 3726 75070 3778
rect 75070 3726 75122 3778
rect 75122 3726 75124 3778
rect 75068 3724 75124 3726
rect 74844 3388 74900 3444
rect 75516 6466 75572 6468
rect 75516 6414 75518 6466
rect 75518 6414 75570 6466
rect 75570 6414 75572 6466
rect 75516 6412 75572 6414
rect 75516 6188 75572 6244
rect 76188 8204 76244 8260
rect 77084 13916 77140 13972
rect 76524 8204 76580 8260
rect 76860 8316 76916 8372
rect 76412 8092 76468 8148
rect 75628 5794 75684 5796
rect 75628 5742 75630 5794
rect 75630 5742 75682 5794
rect 75682 5742 75684 5794
rect 75628 5740 75684 5742
rect 76412 6802 76468 6804
rect 76412 6750 76414 6802
rect 76414 6750 76466 6802
rect 76466 6750 76468 6802
rect 76412 6748 76468 6750
rect 77980 18396 78036 18452
rect 77868 17276 77924 17332
rect 77644 15874 77700 15876
rect 77644 15822 77646 15874
rect 77646 15822 77698 15874
rect 77698 15822 77700 15874
rect 77644 15820 77700 15822
rect 77644 14140 77700 14196
rect 78428 19180 78484 19236
rect 78204 17666 78260 17668
rect 78204 17614 78206 17666
rect 78206 17614 78258 17666
rect 78258 17614 78260 17666
rect 78204 17612 78260 17614
rect 78204 17388 78260 17444
rect 78092 16882 78148 16884
rect 78092 16830 78094 16882
rect 78094 16830 78146 16882
rect 78146 16830 78148 16882
rect 78092 16828 78148 16830
rect 78204 15820 78260 15876
rect 78204 15260 78260 15316
rect 78652 22092 78708 22148
rect 78652 17276 78708 17332
rect 77868 14418 77924 14420
rect 77868 14366 77870 14418
rect 77870 14366 77922 14418
rect 77922 14366 77924 14418
rect 77868 14364 77924 14366
rect 78204 14140 78260 14196
rect 78092 13468 78148 13524
rect 77756 13132 77812 13188
rect 77644 11900 77700 11956
rect 77644 10780 77700 10836
rect 77196 8316 77252 8372
rect 77644 9714 77700 9716
rect 77644 9662 77646 9714
rect 77646 9662 77698 9714
rect 77698 9662 77700 9714
rect 77644 9660 77700 9662
rect 77868 8930 77924 8932
rect 77868 8878 77870 8930
rect 77870 8878 77922 8930
rect 77922 8878 77924 8930
rect 77868 8876 77924 8878
rect 77868 8204 77924 8260
rect 77532 7420 77588 7476
rect 77196 6860 77252 6916
rect 76860 6524 76916 6580
rect 76300 5180 76356 5236
rect 76860 6300 76916 6356
rect 76972 5068 77028 5124
rect 77532 6748 77588 6804
rect 77420 6412 77476 6468
rect 77308 6076 77364 6132
rect 76188 4114 76244 4116
rect 76188 4062 76190 4114
rect 76190 4062 76242 4114
rect 76242 4062 76244 4114
rect 76188 4060 76244 4062
rect 78204 11900 78260 11956
rect 78204 10780 78260 10836
rect 78204 9714 78260 9716
rect 78204 9662 78206 9714
rect 78206 9662 78258 9714
rect 78258 9662 78260 9714
rect 78204 9660 78260 9662
rect 78092 9548 78148 9604
rect 78092 8540 78148 8596
rect 78092 6802 78148 6804
rect 78092 6750 78094 6802
rect 78094 6750 78146 6802
rect 78146 6750 78148 6802
rect 78092 6748 78148 6750
rect 78204 6130 78260 6132
rect 78204 6078 78206 6130
rect 78206 6078 78258 6130
rect 78258 6078 78260 6130
rect 78204 6076 78260 6078
rect 78428 8876 78484 8932
rect 78092 5180 78148 5236
rect 78316 5068 78372 5124
rect 78428 4060 78484 4116
rect 75516 1820 75572 1876
<< metal3 >>
rect 79200 79156 80000 79184
rect 77196 79100 80000 79156
rect 77196 79044 77252 79100
rect 79200 79072 80000 79100
rect 77186 78988 77196 79044
rect 77252 78988 77262 79044
rect 79200 78036 80000 78064
rect 77970 77980 77980 78036
rect 78036 77980 80000 78036
rect 79200 77952 80000 77980
rect 0 77364 800 77392
rect 0 77308 2156 77364
rect 2212 77308 2222 77364
rect 0 77280 800 77308
rect 62962 77084 62972 77140
rect 63028 77084 63980 77140
rect 64036 77084 64046 77140
rect 43474 76972 43484 77028
rect 43540 76972 43932 77028
rect 43988 76972 44492 77028
rect 44548 76972 44558 77028
rect 61618 76972 61628 77028
rect 61684 76972 62636 77028
rect 62692 76972 62702 77028
rect 63634 76972 63644 77028
rect 63700 76972 64652 77028
rect 64708 76972 64718 77028
rect 66994 76972 67004 77028
rect 67060 76972 67788 77028
rect 67844 76972 67854 77028
rect 70354 76972 70364 77028
rect 70420 76972 71820 77028
rect 71876 76972 71886 77028
rect 79200 76916 80000 76944
rect 76962 76860 76972 76916
rect 77028 76860 80000 76916
rect 19826 76804 19836 76860
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 20100 76804 20110 76860
rect 50546 76804 50556 76860
rect 50612 76804 50660 76860
rect 50716 76804 50764 76860
rect 50820 76804 50830 76860
rect 79200 76832 80000 76860
rect 58706 76748 58716 76804
rect 58772 76748 75404 76804
rect 75460 76748 75470 76804
rect 15362 76636 15372 76692
rect 15428 76636 16604 76692
rect 16660 76636 16670 76692
rect 21074 76636 21084 76692
rect 21140 76636 21980 76692
rect 22036 76636 22046 76692
rect 41010 76636 41020 76692
rect 41076 76636 42028 76692
rect 42084 76636 42094 76692
rect 44146 76636 44156 76692
rect 44212 76636 45388 76692
rect 45444 76636 45836 76692
rect 45892 76636 45902 76692
rect 46162 76636 46172 76692
rect 46228 76636 47404 76692
rect 47460 76636 47852 76692
rect 47908 76636 47918 76692
rect 48178 76636 48188 76692
rect 48244 76636 49196 76692
rect 49252 76636 49262 76692
rect 50194 76636 50204 76692
rect 50260 76636 51212 76692
rect 51268 76636 51278 76692
rect 52882 76636 52892 76692
rect 52948 76636 53900 76692
rect 53956 76636 55132 76692
rect 55188 76636 55198 76692
rect 56914 76636 56924 76692
rect 56980 76636 59836 76692
rect 59892 76636 59902 76692
rect 68338 76636 68348 76692
rect 68404 76636 69132 76692
rect 69188 76636 69198 76692
rect 73042 76636 73052 76692
rect 73108 76636 74060 76692
rect 74116 76636 74126 76692
rect 68002 76524 68012 76580
rect 68068 76524 68796 76580
rect 68852 76524 68862 76580
rect 69682 76524 69692 76580
rect 69748 76524 70924 76580
rect 70980 76524 70990 76580
rect 71698 76524 71708 76580
rect 71764 76524 73164 76580
rect 73220 76524 73230 76580
rect 73714 76524 73724 76580
rect 73780 76524 74508 76580
rect 74564 76524 74956 76580
rect 75012 76524 75022 76580
rect 76038 76524 76076 76580
rect 76132 76524 76142 76580
rect 35074 76412 35084 76468
rect 35140 76412 35756 76468
rect 35812 76412 35822 76468
rect 57474 76412 57484 76468
rect 57540 76412 58828 76468
rect 58884 76412 58894 76468
rect 59602 76412 59612 76468
rect 59668 76412 62076 76468
rect 62132 76412 62142 76468
rect 8306 76300 8316 76356
rect 8372 76300 12124 76356
rect 12180 76300 13356 76356
rect 13412 76300 13422 76356
rect 16370 76300 16380 76356
rect 16436 76300 17164 76356
rect 17220 76300 17230 76356
rect 31826 76300 31836 76356
rect 31892 76300 38668 76356
rect 38724 76300 38734 76356
rect 47058 76300 47068 76356
rect 47124 76300 47852 76356
rect 47908 76300 47918 76356
rect 55682 76300 55692 76356
rect 55748 76300 76748 76356
rect 76804 76300 76814 76356
rect 0 76244 800 76272
rect 0 76188 1932 76244
rect 1988 76188 1998 76244
rect 64306 76188 64316 76244
rect 64372 76188 72268 76244
rect 72324 76188 72334 76244
rect 0 76160 800 76188
rect 70466 76076 70476 76132
rect 70532 76076 78204 76132
rect 78260 76076 78270 76132
rect 4466 76020 4476 76076
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4740 76020 4750 76076
rect 35186 76020 35196 76076
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35460 76020 35470 76076
rect 65906 76020 65916 76076
rect 65972 76020 66020 76076
rect 66076 76020 66124 76076
rect 66180 76020 66190 76076
rect 69346 75964 69356 76020
rect 69412 75964 77868 76020
rect 77924 75964 77934 76020
rect 11890 75852 11900 75908
rect 11956 75852 12572 75908
rect 12628 75852 12638 75908
rect 20626 75852 20636 75908
rect 20692 75852 21532 75908
rect 21588 75852 21598 75908
rect 33506 75852 33516 75908
rect 33572 75852 38556 75908
rect 38612 75852 38622 75908
rect 46834 75852 46844 75908
rect 46900 75852 48412 75908
rect 48468 75852 48478 75908
rect 75394 75852 75404 75908
rect 75460 75852 76412 75908
rect 76468 75852 77140 75908
rect 23650 75740 23660 75796
rect 23716 75740 24780 75796
rect 24836 75740 24846 75796
rect 36754 75740 36764 75796
rect 36820 75740 37324 75796
rect 37380 75740 37390 75796
rect 37874 75740 37884 75796
rect 37940 75740 39004 75796
rect 39060 75740 39070 75796
rect 50082 75740 50092 75796
rect 50148 75740 50764 75796
rect 50820 75740 50830 75796
rect 65314 75740 65324 75796
rect 65380 75740 65996 75796
rect 66052 75740 66062 75796
rect 74834 75740 74844 75796
rect 74900 75740 76524 75796
rect 76580 75740 76590 75796
rect 12674 75628 12684 75684
rect 12740 75628 13580 75684
rect 13636 75628 13646 75684
rect 19618 75628 19628 75684
rect 19684 75628 20300 75684
rect 20356 75628 20366 75684
rect 23874 75628 23884 75684
rect 23940 75628 25228 75684
rect 25284 75628 25294 75684
rect 30146 75628 30156 75684
rect 30212 75628 33516 75684
rect 33572 75628 33582 75684
rect 38210 75628 38220 75684
rect 38276 75628 38892 75684
rect 38948 75628 38958 75684
rect 40114 75628 40124 75684
rect 40180 75628 40908 75684
rect 40964 75628 40974 75684
rect 43810 75628 43820 75684
rect 43876 75628 50540 75684
rect 50596 75628 50606 75684
rect 73826 75628 73836 75684
rect 73892 75628 75628 75684
rect 75684 75628 75694 75684
rect 77084 75572 77140 75852
rect 79200 75796 80000 75824
rect 78092 75740 80000 75796
rect 78092 75684 78148 75740
rect 79200 75712 80000 75740
rect 78082 75628 78092 75684
rect 78148 75628 78158 75684
rect 11554 75516 11564 75572
rect 11620 75516 13916 75572
rect 13972 75516 13982 75572
rect 17938 75516 17948 75572
rect 18004 75516 19180 75572
rect 19236 75516 19246 75572
rect 58146 75516 58156 75572
rect 58212 75516 59388 75572
rect 59444 75516 59454 75572
rect 60274 75516 60284 75572
rect 60340 75516 61180 75572
rect 61236 75516 61740 75572
rect 61796 75516 61806 75572
rect 74498 75516 74508 75572
rect 74564 75516 76860 75572
rect 76916 75516 76926 75572
rect 77084 75516 78428 75572
rect 78484 75516 78494 75572
rect 58930 75404 58940 75460
rect 58996 75404 60508 75460
rect 60564 75404 61292 75460
rect 61348 75404 61358 75460
rect 65538 75404 65548 75460
rect 65604 75404 66108 75460
rect 66164 75404 66174 75460
rect 74050 75404 74060 75460
rect 74116 75404 78092 75460
rect 78148 75404 78158 75460
rect 1922 75292 1932 75348
rect 1988 75292 1998 75348
rect 76066 75292 76076 75348
rect 76132 75292 77084 75348
rect 77140 75292 77756 75348
rect 77812 75292 77822 75348
rect 0 75124 800 75152
rect 1932 75124 1988 75292
rect 19826 75236 19836 75292
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 20100 75236 20110 75292
rect 50546 75236 50556 75292
rect 50612 75236 50660 75292
rect 50716 75236 50764 75292
rect 50820 75236 50830 75292
rect 75394 75180 75404 75236
rect 75460 75180 75964 75236
rect 76020 75180 79100 75236
rect 79156 75180 79166 75236
rect 0 75068 1988 75124
rect 52770 75068 52780 75124
rect 52836 75068 53004 75124
rect 53060 75068 53070 75124
rect 74946 75068 74956 75124
rect 75012 75068 76188 75124
rect 76244 75068 76254 75124
rect 0 75040 800 75068
rect 33954 74956 33964 75012
rect 34020 74956 34972 75012
rect 35028 74956 35038 75012
rect 63746 74956 63756 75012
rect 63812 74956 77532 75012
rect 77588 74956 77598 75012
rect 9986 74844 9996 74900
rect 10052 74844 13468 74900
rect 13524 74844 14252 74900
rect 14308 74844 14318 74900
rect 11666 74732 11676 74788
rect 11732 74732 19404 74788
rect 19460 74732 19470 74788
rect 35746 74732 35756 74788
rect 35812 74732 39788 74788
rect 39844 74732 39854 74788
rect 74162 74732 74172 74788
rect 74228 74732 76300 74788
rect 76356 74732 76366 74788
rect 76514 74732 76524 74788
rect 76580 74732 77308 74788
rect 77364 74732 77374 74788
rect 79200 74676 80000 74704
rect 60834 74620 60844 74676
rect 60900 74620 61628 74676
rect 61684 74620 61694 74676
rect 78082 74620 78092 74676
rect 78148 74620 80000 74676
rect 79200 74592 80000 74620
rect 4466 74452 4476 74508
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4740 74452 4750 74508
rect 35186 74452 35196 74508
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35460 74452 35470 74508
rect 65906 74452 65916 74508
rect 65972 74452 66020 74508
rect 66076 74452 66124 74508
rect 66180 74452 66190 74508
rect 1922 74172 1932 74228
rect 1988 74172 1998 74228
rect 75282 74172 75292 74228
rect 75348 74172 78092 74228
rect 78148 74172 78158 74228
rect 0 74004 800 74032
rect 1932 74004 1988 74172
rect 14018 74060 14028 74116
rect 14084 74060 16380 74116
rect 16436 74060 16446 74116
rect 74610 74060 74620 74116
rect 74676 74060 76972 74116
rect 77028 74060 77038 74116
rect 0 73948 1988 74004
rect 12898 73948 12908 74004
rect 12964 73948 14364 74004
rect 14420 73948 14430 74004
rect 73714 73948 73724 74004
rect 73780 73948 74732 74004
rect 74788 73948 74798 74004
rect 0 73920 800 73948
rect 52882 73836 52892 73892
rect 52948 73836 53340 73892
rect 53396 73836 53406 73892
rect 19826 73668 19836 73724
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 20100 73668 20110 73724
rect 50546 73668 50556 73724
rect 50612 73668 50660 73724
rect 50716 73668 50764 73724
rect 50820 73668 50830 73724
rect 79200 73556 80000 73584
rect 77410 73500 77420 73556
rect 77476 73500 78204 73556
rect 78260 73500 80000 73556
rect 79200 73472 80000 73500
rect 56914 73164 56924 73220
rect 56980 73164 77644 73220
rect 77700 73164 77710 73220
rect 1922 73052 1932 73108
rect 1988 73052 1998 73108
rect 0 72884 800 72912
rect 1932 72884 1988 73052
rect 4466 72884 4476 72940
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4740 72884 4750 72940
rect 35186 72884 35196 72940
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35460 72884 35470 72940
rect 65906 72884 65916 72940
rect 65972 72884 66020 72940
rect 66076 72884 66124 72940
rect 66180 72884 66190 72940
rect 0 72828 1988 72884
rect 0 72800 800 72828
rect 2930 72492 2940 72548
rect 2996 72492 4956 72548
rect 5012 72492 5740 72548
rect 5796 72492 5806 72548
rect 76402 72492 76412 72548
rect 76468 72492 77868 72548
rect 77924 72492 77934 72548
rect 79200 72436 80000 72464
rect 77634 72380 77644 72436
rect 77700 72380 78204 72436
rect 78260 72380 80000 72436
rect 79200 72352 80000 72380
rect 19826 72100 19836 72156
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 20100 72100 20110 72156
rect 50546 72100 50556 72156
rect 50612 72100 50660 72156
rect 50716 72100 50764 72156
rect 50820 72100 50830 72156
rect 1922 71932 1932 71988
rect 1988 71932 1998 71988
rect 3154 71932 3164 71988
rect 3220 71932 3948 71988
rect 4004 71932 4014 71988
rect 0 71764 800 71792
rect 1932 71764 1988 71932
rect 77858 71820 77868 71876
rect 77924 71820 78540 71876
rect 78596 71820 78606 71876
rect 0 71708 1988 71764
rect 77634 71708 77644 71764
rect 77700 71708 78204 71764
rect 78260 71708 78270 71764
rect 0 71680 800 71708
rect 4466 71316 4476 71372
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4740 71316 4750 71372
rect 35186 71316 35196 71372
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35460 71316 35470 71372
rect 65906 71316 65916 71372
rect 65972 71316 66020 71372
rect 66076 71316 66124 71372
rect 66180 71316 66190 71372
rect 79200 71316 80000 71344
rect 78194 71260 78204 71316
rect 78260 71260 80000 71316
rect 79200 71232 80000 71260
rect 77746 71036 77756 71092
rect 77812 71036 78876 71092
rect 78932 71036 78942 71092
rect 77410 70700 77420 70756
rect 77476 70700 78204 70756
rect 78260 70700 78270 70756
rect 0 70644 800 70672
rect 0 70588 1932 70644
rect 1988 70588 1998 70644
rect 59612 70588 59836 70644
rect 59892 70588 59902 70644
rect 0 70560 800 70588
rect 19826 70532 19836 70588
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 20100 70532 20110 70588
rect 50546 70532 50556 70588
rect 50612 70532 50660 70588
rect 50716 70532 50764 70588
rect 50820 70532 50830 70588
rect 59602 70532 59612 70588
rect 59668 70532 59678 70588
rect 79200 70196 80000 70224
rect 2706 70140 2716 70196
rect 2772 70140 3836 70196
rect 3892 70140 3902 70196
rect 78194 70140 78204 70196
rect 78260 70140 80000 70196
rect 79200 70112 80000 70140
rect 4466 69748 4476 69804
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4740 69748 4750 69804
rect 35186 69748 35196 69804
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35460 69748 35470 69804
rect 65906 69748 65916 69804
rect 65972 69748 66020 69804
rect 66076 69748 66124 69804
rect 66180 69748 66190 69804
rect 0 69524 800 69552
rect 0 69468 1932 69524
rect 1988 69468 1998 69524
rect 0 69440 800 69468
rect 79200 69076 80000 69104
rect 77634 69020 77644 69076
rect 77700 69020 78204 69076
rect 78260 69020 80000 69076
rect 19826 68964 19836 69020
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 20100 68964 20110 69020
rect 50546 68964 50556 69020
rect 50612 68964 50660 69020
rect 50716 68964 50764 69020
rect 50820 68964 50830 69020
rect 79200 68992 80000 69020
rect 72146 68796 72156 68852
rect 72212 68796 77084 68852
rect 77140 68796 77150 68852
rect 77410 68460 77420 68516
rect 77476 68460 78204 68516
rect 78260 68460 78270 68516
rect 0 68404 800 68432
rect 0 68348 2716 68404
rect 2772 68348 2782 68404
rect 0 68320 800 68348
rect 4466 68180 4476 68236
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4740 68180 4750 68236
rect 35186 68180 35196 68236
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35460 68180 35470 68236
rect 65906 68180 65916 68236
rect 65972 68180 66020 68236
rect 66076 68180 66124 68236
rect 66180 68180 66190 68236
rect 79200 67956 80000 67984
rect 78194 67900 78204 67956
rect 78260 67900 80000 67956
rect 79200 67872 80000 67900
rect 76290 67788 76300 67844
rect 76356 67788 77644 67844
rect 77700 67788 77710 67844
rect 19826 67396 19836 67452
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 20100 67396 20110 67452
rect 50546 67396 50556 67452
rect 50612 67396 50660 67452
rect 50716 67396 50764 67452
rect 50820 67396 50830 67452
rect 0 67284 800 67312
rect 0 67228 1932 67284
rect 1988 67228 1998 67284
rect 0 67200 800 67228
rect 2706 67116 2716 67172
rect 2772 67116 3724 67172
rect 3780 67116 4284 67172
rect 4340 67116 4350 67172
rect 75842 67116 75852 67172
rect 75908 67116 77868 67172
rect 77924 67116 77934 67172
rect 2258 67004 2268 67060
rect 2324 67004 3388 67060
rect 3444 67004 3454 67060
rect 79200 66836 80000 66864
rect 77634 66780 77644 66836
rect 77700 66780 78204 66836
rect 78260 66780 80000 66836
rect 79200 66752 80000 66780
rect 4466 66612 4476 66668
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4740 66612 4750 66668
rect 35186 66612 35196 66668
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35460 66612 35470 66668
rect 65906 66612 65916 66668
rect 65972 66612 66020 66668
rect 66076 66612 66124 66668
rect 66180 66612 66190 66668
rect 1922 66332 1932 66388
rect 1988 66332 1998 66388
rect 0 66164 800 66192
rect 1932 66164 1988 66332
rect 3042 66220 3052 66276
rect 3108 66220 3836 66276
rect 3892 66220 3902 66276
rect 70018 66220 70028 66276
rect 70084 66220 77644 66276
rect 77700 66220 77710 66276
rect 0 66108 1988 66164
rect 0 66080 800 66108
rect 19826 65828 19836 65884
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 20100 65828 20110 65884
rect 50546 65828 50556 65884
rect 50612 65828 50660 65884
rect 50716 65828 50764 65884
rect 50820 65828 50830 65884
rect 79200 65716 80000 65744
rect 77410 65660 77420 65716
rect 77476 65660 78204 65716
rect 78260 65660 80000 65716
rect 79200 65632 80000 65660
rect 2706 65212 2716 65268
rect 2772 65212 2782 65268
rect 0 65044 800 65072
rect 2716 65044 2772 65212
rect 4466 65044 4476 65100
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4740 65044 4750 65100
rect 35186 65044 35196 65100
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35460 65044 35470 65100
rect 65906 65044 65916 65100
rect 65972 65044 66020 65100
rect 66076 65044 66124 65100
rect 66180 65044 66190 65100
rect 0 64988 2772 65044
rect 0 64960 800 64988
rect 77634 64652 77644 64708
rect 77700 64652 78876 64708
rect 78932 64652 78942 64708
rect 79200 64596 80000 64624
rect 77410 64540 77420 64596
rect 77476 64540 78204 64596
rect 78260 64540 80000 64596
rect 79200 64512 80000 64540
rect 19826 64260 19836 64316
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 20100 64260 20110 64316
rect 50546 64260 50556 64316
rect 50612 64260 50660 64316
rect 50716 64260 50764 64316
rect 50820 64260 50830 64316
rect 2818 63980 2828 64036
rect 2884 63980 3724 64036
rect 3780 63980 3790 64036
rect 0 63924 800 63952
rect 0 63868 1932 63924
rect 1988 63868 1998 63924
rect 77634 63868 77644 63924
rect 77700 63868 78204 63924
rect 78260 63868 78270 63924
rect 0 63840 800 63868
rect 4466 63476 4476 63532
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4740 63476 4750 63532
rect 35186 63476 35196 63532
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35460 63476 35470 63532
rect 65906 63476 65916 63532
rect 65972 63476 66020 63532
rect 66076 63476 66124 63532
rect 66180 63476 66190 63532
rect 79200 63476 80000 63504
rect 78194 63420 78204 63476
rect 78260 63420 80000 63476
rect 79200 63392 80000 63420
rect 77410 62860 77420 62916
rect 77476 62860 78204 62916
rect 78260 62860 78270 62916
rect 0 62804 800 62832
rect 0 62748 1932 62804
rect 1988 62748 1998 62804
rect 0 62720 800 62748
rect 19826 62692 19836 62748
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 20100 62692 20110 62748
rect 50546 62692 50556 62748
rect 50612 62692 50660 62748
rect 50716 62692 50764 62748
rect 50820 62692 50830 62748
rect 79200 62356 80000 62384
rect 78194 62300 78204 62356
rect 78260 62300 80000 62356
rect 79200 62272 80000 62300
rect 76402 62188 76412 62244
rect 76468 62188 77868 62244
rect 77924 62188 77934 62244
rect 2818 62076 2828 62132
rect 2884 62076 3612 62132
rect 3668 62076 3678 62132
rect 4466 61908 4476 61964
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4740 61908 4750 61964
rect 35186 61908 35196 61964
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35460 61908 35470 61964
rect 65906 61908 65916 61964
rect 65972 61908 66020 61964
rect 66076 61908 66124 61964
rect 66180 61908 66190 61964
rect 0 61684 800 61712
rect 0 61628 1932 61684
rect 1988 61628 1998 61684
rect 0 61600 800 61628
rect 2818 61292 2828 61348
rect 2884 61292 4172 61348
rect 4228 61292 4238 61348
rect 76962 61292 76972 61348
rect 77028 61292 77868 61348
rect 77924 61292 77934 61348
rect 79200 61236 80000 61264
rect 77634 61180 77644 61236
rect 77700 61180 78204 61236
rect 78260 61180 80000 61236
rect 19826 61124 19836 61180
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 20100 61124 20110 61180
rect 50546 61124 50556 61180
rect 50612 61124 50660 61180
rect 50716 61124 50764 61180
rect 50820 61124 50830 61180
rect 79200 61152 80000 61180
rect 77634 60732 77644 60788
rect 77700 60732 78204 60788
rect 78260 60732 78270 60788
rect 0 60564 800 60592
rect 0 60508 2716 60564
rect 2772 60508 2782 60564
rect 0 60480 800 60508
rect 4466 60340 4476 60396
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4740 60340 4750 60396
rect 35186 60340 35196 60396
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35460 60340 35470 60396
rect 65906 60340 65916 60396
rect 65972 60340 66020 60396
rect 66076 60340 66124 60396
rect 66180 60340 66190 60396
rect 79200 60116 80000 60144
rect 78194 60060 78204 60116
rect 78260 60060 80000 60116
rect 79200 60032 80000 60060
rect 2706 59948 2716 60004
rect 2772 59948 3836 60004
rect 3892 59948 3902 60004
rect 19826 59556 19836 59612
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 20100 59556 20110 59612
rect 50546 59556 50556 59612
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50820 59556 50830 59612
rect 0 59444 800 59472
rect 0 59388 1932 59444
rect 1988 59388 1998 59444
rect 0 59360 800 59388
rect 2146 59164 2156 59220
rect 2212 59164 2940 59220
rect 2996 59164 3500 59220
rect 3556 59164 3566 59220
rect 75842 59052 75852 59108
rect 75908 59052 77644 59108
rect 77700 59052 77710 59108
rect 79200 58996 80000 59024
rect 77410 58940 77420 58996
rect 77476 58940 78204 58996
rect 78260 58940 80000 58996
rect 79200 58912 80000 58940
rect 4466 58772 4476 58828
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4740 58772 4750 58828
rect 35186 58772 35196 58828
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35460 58772 35470 58828
rect 65906 58772 65916 58828
rect 65972 58772 66020 58828
rect 66076 58772 66124 58828
rect 66180 58772 66190 58828
rect 0 58324 800 58352
rect 0 58268 2772 58324
rect 0 58240 800 58268
rect 2716 58212 2772 58268
rect 2706 58156 2716 58212
rect 2772 58156 2782 58212
rect 68898 58156 68908 58212
rect 68964 58156 77868 58212
rect 77924 58156 77934 58212
rect 19826 57988 19836 58044
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 20100 57988 20110 58044
rect 50546 57988 50556 58044
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50820 57988 50830 58044
rect 79200 57876 80000 57904
rect 77634 57820 77644 57876
rect 77700 57820 78204 57876
rect 78260 57820 80000 57876
rect 79200 57792 80000 57820
rect 1922 57372 1932 57428
rect 1988 57372 1998 57428
rect 0 57204 800 57232
rect 1932 57204 1988 57372
rect 4466 57204 4476 57260
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4740 57204 4750 57260
rect 35186 57204 35196 57260
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35460 57204 35470 57260
rect 65906 57204 65916 57260
rect 65972 57204 66020 57260
rect 66076 57204 66124 57260
rect 66180 57204 66190 57260
rect 0 57148 1988 57204
rect 0 57120 800 57148
rect 79200 56756 80000 56784
rect 77634 56700 77644 56756
rect 77700 56700 78204 56756
rect 78260 56700 80000 56756
rect 79200 56672 80000 56700
rect 74050 56588 74060 56644
rect 74116 56588 77868 56644
rect 77924 56588 77934 56644
rect 19826 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20110 56476
rect 50546 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50830 56476
rect 2706 56140 2716 56196
rect 2772 56140 3388 56196
rect 3444 56140 4844 56196
rect 4900 56140 4910 56196
rect 0 56084 800 56112
rect 0 56028 1932 56084
rect 1988 56028 1998 56084
rect 0 56000 800 56028
rect 64530 55916 64540 55972
rect 64596 55916 77644 55972
rect 77700 55916 77710 55972
rect 4466 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4750 55692
rect 35186 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35470 55692
rect 65906 55636 65916 55692
rect 65972 55636 66020 55692
rect 66076 55636 66124 55692
rect 66180 55636 66190 55692
rect 79200 55636 80000 55664
rect 77410 55580 77420 55636
rect 77476 55580 78204 55636
rect 78260 55580 80000 55636
rect 79200 55552 80000 55580
rect 77634 55132 77644 55188
rect 77700 55132 78204 55188
rect 78260 55132 78270 55188
rect 2706 55020 2716 55076
rect 2772 55020 2782 55076
rect 60386 55020 60396 55076
rect 60452 55020 77868 55076
rect 77924 55020 77934 55076
rect 0 54964 800 54992
rect 2716 54964 2772 55020
rect 0 54908 2772 54964
rect 0 54880 800 54908
rect 19826 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20110 54908
rect 50546 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50830 54908
rect 79200 54516 80000 54544
rect 78194 54460 78204 54516
rect 78260 54460 80000 54516
rect 79200 54432 80000 54460
rect 4466 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4750 54124
rect 35186 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35470 54124
rect 65906 54068 65916 54124
rect 65972 54068 66020 54124
rect 66076 54068 66124 54124
rect 66180 54068 66190 54124
rect 0 53844 800 53872
rect 0 53788 1932 53844
rect 1988 53788 1998 53844
rect 0 53760 800 53788
rect 3154 53564 3164 53620
rect 3220 53564 3948 53620
rect 4004 53564 4014 53620
rect 2482 53452 2492 53508
rect 2548 53452 2940 53508
rect 2996 53452 3836 53508
rect 3892 53452 3902 53508
rect 79200 53396 80000 53424
rect 77634 53340 77644 53396
rect 77700 53340 78204 53396
rect 78260 53340 80000 53396
rect 19826 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20110 53340
rect 50546 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50830 53340
rect 79200 53312 80000 53340
rect 70802 53004 70812 53060
rect 70868 53004 77868 53060
rect 77924 53004 77934 53060
rect 0 52724 800 52752
rect 0 52668 1932 52724
rect 1988 52668 1998 52724
rect 0 52640 800 52668
rect 4466 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4750 52556
rect 35186 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35470 52556
rect 65906 52500 65916 52556
rect 65972 52500 66020 52556
rect 66076 52500 66124 52556
rect 66180 52500 66190 52556
rect 79200 52276 80000 52304
rect 78194 52220 78204 52276
rect 78260 52220 80000 52276
rect 79200 52192 80000 52220
rect 19826 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20110 51772
rect 50546 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50830 51772
rect 0 51604 800 51632
rect 0 51548 1932 51604
rect 1988 51548 1998 51604
rect 0 51520 800 51548
rect 79200 51156 80000 51184
rect 77634 51100 77644 51156
rect 77700 51100 78204 51156
rect 78260 51100 80000 51156
rect 79200 51072 80000 51100
rect 4466 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4750 50988
rect 35186 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35470 50988
rect 65906 50932 65916 50988
rect 65972 50932 66020 50988
rect 66076 50932 66124 50988
rect 66180 50932 66190 50988
rect 1922 50652 1932 50708
rect 1988 50652 1998 50708
rect 0 50484 800 50512
rect 1932 50484 1988 50652
rect 2818 50540 2828 50596
rect 2884 50540 3836 50596
rect 3892 50540 3902 50596
rect 0 50428 1988 50484
rect 77634 50428 77644 50484
rect 77700 50428 78204 50484
rect 78260 50428 78270 50484
rect 0 50400 800 50428
rect 77858 50316 77868 50372
rect 77924 50316 78988 50372
rect 79044 50316 79054 50372
rect 19826 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20110 50204
rect 50546 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50830 50204
rect 79200 50036 80000 50064
rect 78194 49980 78204 50036
rect 78260 49980 80000 50036
rect 79200 49952 80000 49980
rect 1922 49532 1932 49588
rect 1988 49532 1998 49588
rect 3154 49532 3164 49588
rect 3220 49532 3612 49588
rect 3668 49532 3678 49588
rect 0 49364 800 49392
rect 1932 49364 1988 49532
rect 4466 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4750 49420
rect 35186 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35470 49420
rect 65906 49364 65916 49420
rect 65972 49364 66020 49420
rect 66076 49364 66124 49420
rect 66180 49364 66190 49420
rect 0 49308 1988 49364
rect 0 49280 800 49308
rect 2706 48972 2716 49028
rect 2772 48972 3836 49028
rect 3892 48972 3902 49028
rect 79200 48916 80000 48944
rect 77634 48860 77644 48916
rect 77700 48860 78204 48916
rect 78260 48860 80000 48916
rect 79200 48832 80000 48860
rect 77858 48748 77868 48804
rect 77924 48748 78988 48804
rect 79044 48748 79054 48804
rect 19826 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20110 48636
rect 50546 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50830 48636
rect 72594 48524 72604 48580
rect 72660 48524 77420 48580
rect 77476 48524 77486 48580
rect 0 48244 800 48272
rect 0 48188 1932 48244
rect 1988 48188 1998 48244
rect 2370 48188 2380 48244
rect 2436 48188 2940 48244
rect 2996 48188 3006 48244
rect 77634 48188 77644 48244
rect 77700 48188 78204 48244
rect 78260 48188 78270 48244
rect 0 48160 800 48188
rect 4466 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4750 47852
rect 35186 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35470 47852
rect 65906 47796 65916 47852
rect 65972 47796 66020 47852
rect 66076 47796 66124 47852
rect 66180 47796 66190 47852
rect 79200 47796 80000 47824
rect 78194 47740 78204 47796
rect 78260 47740 80000 47796
rect 79200 47712 80000 47740
rect 2706 47180 2716 47236
rect 2772 47180 2782 47236
rect 77634 47180 77644 47236
rect 77700 47180 78204 47236
rect 78260 47180 78270 47236
rect 0 47124 800 47152
rect 2716 47124 2772 47180
rect 0 47068 2772 47124
rect 0 47040 800 47068
rect 19826 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20110 47068
rect 50546 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50830 47068
rect 79200 46676 80000 46704
rect 78194 46620 78204 46676
rect 78260 46620 80000 46676
rect 79200 46592 80000 46620
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 65906 46228 65916 46284
rect 65972 46228 66020 46284
rect 66076 46228 66124 46284
rect 66180 46228 66190 46284
rect 0 46004 800 46032
rect 0 45948 1932 46004
rect 1988 45948 1998 46004
rect 0 45920 800 45948
rect 2706 45836 2716 45892
rect 2772 45836 3276 45892
rect 3332 45836 4284 45892
rect 4340 45836 4350 45892
rect 72034 45836 72044 45892
rect 72100 45836 77868 45892
rect 77924 45836 77934 45892
rect 2370 45724 2380 45780
rect 2436 45724 3052 45780
rect 3108 45724 3612 45780
rect 3668 45724 3678 45780
rect 73154 45612 73164 45668
rect 73220 45612 77868 45668
rect 77924 45612 77934 45668
rect 79200 45556 80000 45584
rect 77634 45500 77644 45556
rect 77700 45500 78204 45556
rect 78260 45500 80000 45556
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 50546 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50830 45500
rect 79200 45472 80000 45500
rect 56018 45276 56028 45332
rect 56084 45276 58492 45332
rect 58548 45276 58558 45332
rect 73826 45276 73836 45332
rect 73892 45276 75740 45332
rect 75796 45276 75806 45332
rect 77410 45276 77420 45332
rect 77476 45276 77486 45332
rect 77420 45108 77476 45276
rect 72594 45052 72604 45108
rect 72660 45052 77476 45108
rect 77634 44940 77644 44996
rect 77700 44940 78204 44996
rect 78260 44940 78270 44996
rect 0 44884 800 44912
rect 0 44828 2716 44884
rect 2772 44828 2782 44884
rect 0 44800 800 44828
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 65906 44660 65916 44716
rect 65972 44660 66020 44716
rect 66076 44660 66124 44716
rect 66180 44660 66190 44716
rect 79200 44436 80000 44464
rect 78194 44380 78204 44436
rect 78260 44380 80000 44436
rect 79200 44352 80000 44380
rect 2706 44044 2716 44100
rect 2772 44044 2782 44100
rect 0 43764 800 43792
rect 2716 43764 2772 44044
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 50546 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50830 43932
rect 0 43708 2772 43764
rect 0 43680 800 43708
rect 2258 43484 2268 43540
rect 2324 43484 2828 43540
rect 2884 43484 2894 43540
rect 63746 43484 63756 43540
rect 63812 43484 77420 43540
rect 77476 43484 77486 43540
rect 77420 43428 77476 43484
rect 57026 43372 57036 43428
rect 57092 43372 59500 43428
rect 59556 43372 59566 43428
rect 77420 43372 78204 43428
rect 78260 43372 78270 43428
rect 79200 43316 80000 43344
rect 78082 43260 78092 43316
rect 78148 43260 80000 43316
rect 79200 43232 80000 43260
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 65906 43092 65916 43148
rect 65972 43092 66020 43148
rect 66076 43092 66124 43148
rect 66180 43092 66190 43148
rect 1922 42812 1932 42868
rect 1988 42812 1998 42868
rect 58146 42812 58156 42868
rect 58212 42812 59948 42868
rect 60004 42812 60014 42868
rect 0 42644 800 42672
rect 1932 42644 1988 42812
rect 2706 42700 2716 42756
rect 2772 42700 3836 42756
rect 3892 42700 3902 42756
rect 0 42588 1988 42644
rect 75730 42588 75740 42644
rect 75796 42588 77308 42644
rect 77364 42588 77374 42644
rect 0 42560 800 42588
rect 75282 42476 75292 42532
rect 75348 42476 76300 42532
rect 76356 42476 76366 42532
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 50546 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50830 42364
rect 70466 42252 70476 42308
rect 70532 42252 77308 42308
rect 77364 42252 77374 42308
rect 79200 42196 80000 42224
rect 65734 42140 65772 42196
rect 65828 42140 65838 42196
rect 74946 42140 74956 42196
rect 75012 42140 75348 42196
rect 77970 42140 77980 42196
rect 78036 42140 80000 42196
rect 75292 41972 75348 42140
rect 79200 42112 80000 42140
rect 1698 41916 1708 41972
rect 1764 41916 3836 41972
rect 3892 41916 4732 41972
rect 4788 41916 4798 41972
rect 59154 41916 59164 41972
rect 59220 41916 61068 41972
rect 61124 41916 61134 41972
rect 61618 41916 61628 41972
rect 61684 41916 64428 41972
rect 64484 41916 64494 41972
rect 65090 41916 65100 41972
rect 65156 41916 65884 41972
rect 65940 41916 65950 41972
rect 73602 41916 73612 41972
rect 73668 41916 74060 41972
rect 74116 41916 75068 41972
rect 75124 41916 75134 41972
rect 75292 41916 76188 41972
rect 76244 41916 76254 41972
rect 61628 41860 61684 41916
rect 43586 41804 43596 41860
rect 43652 41804 54908 41860
rect 54964 41804 54974 41860
rect 60610 41804 60620 41860
rect 60676 41804 61684 41860
rect 72146 41804 72156 41860
rect 72212 41804 76524 41860
rect 76580 41804 76590 41860
rect 1922 41692 1932 41748
rect 1988 41692 1998 41748
rect 56354 41692 56364 41748
rect 56420 41692 57148 41748
rect 57204 41692 71148 41748
rect 71204 41692 71596 41748
rect 71652 41692 71662 41748
rect 0 41524 800 41552
rect 1932 41524 1988 41692
rect 70466 41580 70476 41636
rect 70532 41580 74620 41636
rect 74676 41580 74732 41636
rect 74788 41580 75068 41636
rect 75124 41580 75134 41636
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 65906 41524 65916 41580
rect 65972 41524 66020 41580
rect 66076 41524 66124 41580
rect 66180 41524 66190 41580
rect 0 41468 1988 41524
rect 64978 41468 64988 41524
rect 65044 41468 65660 41524
rect 65716 41468 65726 41524
rect 71698 41468 71708 41524
rect 71764 41468 74396 41524
rect 74452 41468 74462 41524
rect 0 41440 800 41468
rect 55346 41356 55356 41412
rect 55412 41356 55580 41412
rect 55636 41356 56924 41412
rect 56980 41356 57820 41412
rect 57876 41356 57886 41412
rect 64418 41356 64428 41412
rect 64484 41356 67900 41412
rect 67956 41356 67966 41412
rect 69570 41356 69580 41412
rect 69636 41356 76076 41412
rect 76132 41356 76972 41412
rect 77028 41356 77038 41412
rect 63522 41244 63532 41300
rect 63588 41244 64988 41300
rect 65044 41244 65054 41300
rect 70690 41244 70700 41300
rect 70756 41244 71372 41300
rect 71428 41244 71438 41300
rect 74162 41244 74172 41300
rect 74228 41244 75292 41300
rect 75348 41244 75358 41300
rect 76514 41244 76524 41300
rect 76580 41244 78092 41300
rect 78148 41244 78158 41300
rect 58482 41132 58492 41188
rect 58548 41132 59388 41188
rect 59444 41132 60172 41188
rect 60228 41132 60508 41188
rect 60564 41132 60574 41188
rect 61618 41132 61628 41188
rect 61684 41132 62860 41188
rect 62916 41132 62926 41188
rect 63298 41132 63308 41188
rect 63364 41132 64316 41188
rect 64372 41132 64382 41188
rect 76188 41132 77532 41188
rect 77588 41132 77598 41188
rect 76188 41076 76244 41132
rect 79200 41076 80000 41104
rect 62514 41020 62524 41076
rect 62580 41020 63420 41076
rect 63476 41020 63486 41076
rect 67890 41020 67900 41076
rect 67956 41020 73276 41076
rect 73332 41020 73342 41076
rect 73826 41020 73836 41076
rect 73892 41020 76244 41076
rect 76626 41020 76636 41076
rect 76692 41020 80000 41076
rect 62860 40964 62916 41020
rect 79200 40992 80000 41020
rect 57138 40908 57148 40964
rect 57204 40908 58268 40964
rect 58324 40908 62692 40964
rect 62850 40908 62860 40964
rect 62916 40908 62926 40964
rect 62636 40852 62692 40908
rect 53778 40796 53788 40852
rect 53844 40796 55020 40852
rect 55076 40796 55356 40852
rect 55412 40796 62580 40852
rect 62636 40796 70252 40852
rect 70308 40796 70924 40852
rect 70980 40796 70990 40852
rect 73892 40796 76188 40852
rect 76244 40796 76254 40852
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 50546 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50830 40796
rect 62524 40740 62580 40796
rect 73892 40740 73948 40796
rect 55122 40684 55132 40740
rect 55188 40684 62188 40740
rect 62524 40684 70700 40740
rect 70756 40684 70766 40740
rect 72930 40684 72940 40740
rect 72996 40684 73948 40740
rect 75058 40684 75068 40740
rect 75124 40684 77868 40740
rect 77924 40684 77934 40740
rect 2258 40572 2268 40628
rect 2324 40572 5404 40628
rect 5460 40572 8428 40628
rect 43138 40572 43148 40628
rect 43204 40572 57148 40628
rect 57204 40572 57214 40628
rect 8372 40516 8428 40572
rect 62132 40516 62188 40684
rect 64194 40572 64204 40628
rect 64260 40572 64652 40628
rect 64708 40572 64718 40628
rect 66322 40572 66332 40628
rect 66388 40572 67452 40628
rect 67508 40572 67518 40628
rect 69346 40572 69356 40628
rect 69412 40572 71372 40628
rect 71428 40572 71438 40628
rect 74610 40572 74620 40628
rect 74676 40572 75068 40628
rect 75124 40572 76748 40628
rect 76804 40572 76814 40628
rect 77410 40572 77420 40628
rect 77476 40572 77980 40628
rect 78036 40572 78046 40628
rect 4050 40460 4060 40516
rect 4116 40460 4508 40516
rect 4564 40460 5180 40516
rect 5236 40460 5246 40516
rect 8372 40460 20972 40516
rect 21028 40460 21038 40516
rect 62132 40460 70476 40516
rect 70532 40460 70542 40516
rect 70690 40460 70700 40516
rect 70756 40460 72268 40516
rect 72324 40460 73612 40516
rect 73668 40460 74284 40516
rect 74340 40460 74350 40516
rect 0 40404 800 40432
rect 0 40348 1932 40404
rect 1988 40348 1998 40404
rect 3154 40348 3164 40404
rect 3220 40348 4956 40404
rect 5012 40348 26908 40404
rect 26964 40348 26974 40404
rect 42578 40348 42588 40404
rect 42644 40348 43596 40404
rect 43652 40348 43662 40404
rect 60050 40348 60060 40404
rect 60116 40348 61628 40404
rect 61684 40348 61694 40404
rect 63186 40348 63196 40404
rect 63252 40348 63532 40404
rect 63588 40348 63598 40404
rect 67554 40348 67564 40404
rect 67620 40348 68236 40404
rect 68292 40348 69020 40404
rect 69076 40348 69086 40404
rect 73378 40348 73388 40404
rect 73444 40348 73948 40404
rect 74004 40348 75292 40404
rect 75348 40348 75358 40404
rect 0 40320 800 40348
rect 62290 40236 62300 40292
rect 62356 40236 63756 40292
rect 63812 40236 63822 40292
rect 71250 40236 71260 40292
rect 71316 40236 72380 40292
rect 72436 40236 72446 40292
rect 59602 40124 59612 40180
rect 59668 40124 70140 40180
rect 70196 40124 70206 40180
rect 74050 40124 74060 40180
rect 74116 40124 75292 40180
rect 75348 40124 75358 40180
rect 75618 40124 75628 40180
rect 75684 40124 78092 40180
rect 78148 40124 78158 40180
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 65906 39956 65916 40012
rect 65972 39956 66020 40012
rect 66076 39956 66124 40012
rect 66180 39956 66190 40012
rect 79200 39956 80000 39984
rect 76402 39900 76412 39956
rect 76468 39900 80000 39956
rect 79200 39872 80000 39900
rect 62402 39788 62412 39844
rect 62468 39788 62860 39844
rect 62916 39788 62926 39844
rect 68450 39788 68460 39844
rect 68516 39788 71932 39844
rect 71988 39788 71998 39844
rect 77186 39788 77196 39844
rect 77252 39788 77644 39844
rect 77700 39788 77710 39844
rect 65762 39676 65772 39732
rect 65828 39676 67116 39732
rect 67172 39676 67182 39732
rect 70690 39676 70700 39732
rect 70756 39676 70924 39732
rect 70980 39676 70990 39732
rect 73266 39676 73276 39732
rect 73332 39676 74620 39732
rect 74676 39676 74686 39732
rect 2594 39564 2604 39620
rect 2660 39564 3836 39620
rect 3892 39564 4732 39620
rect 4788 39564 4798 39620
rect 65202 39564 65212 39620
rect 65268 39564 66332 39620
rect 66388 39564 66668 39620
rect 66724 39564 66734 39620
rect 70354 39564 70364 39620
rect 70420 39564 71484 39620
rect 71540 39564 71550 39620
rect 72790 39564 72828 39620
rect 72884 39564 72894 39620
rect 74162 39564 74172 39620
rect 74228 39564 75068 39620
rect 75124 39564 75134 39620
rect 75282 39564 75292 39620
rect 75348 39564 76524 39620
rect 76580 39564 76590 39620
rect 65734 39452 65772 39508
rect 65828 39452 65838 39508
rect 67666 39452 67676 39508
rect 67732 39452 68460 39508
rect 68516 39452 68526 39508
rect 69682 39452 69692 39508
rect 69748 39452 70028 39508
rect 70084 39452 70924 39508
rect 70980 39452 70990 39508
rect 5170 39340 5180 39396
rect 5236 39340 43260 39396
rect 43316 39340 43326 39396
rect 69346 39340 69356 39396
rect 69412 39340 70476 39396
rect 70532 39340 70542 39396
rect 71250 39340 71260 39396
rect 71316 39340 72380 39396
rect 72436 39340 72446 39396
rect 75030 39340 75068 39396
rect 75124 39340 75134 39396
rect 0 39284 800 39312
rect 0 39228 1932 39284
rect 1988 39228 1998 39284
rect 62132 39228 77700 39284
rect 0 39200 800 39228
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 50546 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50830 39228
rect 62132 39060 62188 39228
rect 65874 39116 65884 39172
rect 65940 39116 68572 39172
rect 68628 39116 69020 39172
rect 69076 39116 69086 39172
rect 72706 39116 72716 39172
rect 72772 39116 72940 39172
rect 72996 39116 73006 39172
rect 2930 39004 2940 39060
rect 2996 39004 3276 39060
rect 3332 39004 42028 39060
rect 42084 39004 42094 39060
rect 54338 39004 54348 39060
rect 54404 39004 62188 39060
rect 63858 39004 63868 39060
rect 63924 39004 64652 39060
rect 64708 39004 65324 39060
rect 65380 39004 65390 39060
rect 68002 39004 68012 39060
rect 68068 39004 68684 39060
rect 68740 39004 69244 39060
rect 69300 39004 69310 39060
rect 74498 39004 74508 39060
rect 74564 39004 75516 39060
rect 75572 39004 75582 39060
rect 77644 38948 77700 39228
rect 26898 38892 26908 38948
rect 26964 38892 41244 38948
rect 41300 38892 41310 38948
rect 43026 38892 43036 38948
rect 43092 38892 43708 38948
rect 46498 38892 46508 38948
rect 46564 38892 61852 38948
rect 61908 38892 62188 38948
rect 67106 38892 67116 38948
rect 67172 38892 69692 38948
rect 69748 38892 69758 38948
rect 73724 38892 74172 38948
rect 74228 38892 74238 38948
rect 77634 38892 77644 38948
rect 77700 38892 77710 38948
rect 43652 38836 43708 38892
rect 62132 38836 62188 38892
rect 73724 38836 73780 38892
rect 79200 38836 80000 38864
rect 41570 38780 41580 38836
rect 41636 38780 41804 38836
rect 41860 38780 42924 38836
rect 42980 38780 42990 38836
rect 43652 38780 44044 38836
rect 44100 38780 51660 38836
rect 51716 38780 56364 38836
rect 56420 38780 56430 38836
rect 62132 38780 62524 38836
rect 62580 38780 68516 38836
rect 69010 38780 69020 38836
rect 69076 38780 70028 38836
rect 70084 38780 70364 38836
rect 70420 38780 70430 38836
rect 70690 38780 70700 38836
rect 70756 38780 71260 38836
rect 71316 38780 71326 38836
rect 72482 38780 72492 38836
rect 72548 38780 73108 38836
rect 73686 38780 73724 38836
rect 73780 38780 73790 38836
rect 73892 38780 75068 38836
rect 75124 38780 75628 38836
rect 75684 38780 75694 38836
rect 77746 38780 77756 38836
rect 77812 38780 80000 38836
rect 68460 38724 68516 38780
rect 73052 38724 73108 38780
rect 73892 38724 73948 38780
rect 74844 38724 74900 38780
rect 79200 38752 80000 38780
rect 41458 38668 41468 38724
rect 41524 38668 51324 38724
rect 51380 38668 53788 38724
rect 53844 38668 53854 38724
rect 67330 38668 67340 38724
rect 67396 38668 68236 38724
rect 68292 38668 68302 38724
rect 68460 38668 69804 38724
rect 69860 38668 69870 38724
rect 73052 38668 73948 38724
rect 74834 38668 74844 38724
rect 74900 38668 74910 38724
rect 75170 38668 75180 38724
rect 75236 38668 75404 38724
rect 75460 38668 75964 38724
rect 76020 38668 77196 38724
rect 77252 38668 77262 38724
rect 72482 38556 72492 38612
rect 72548 38556 72828 38612
rect 72884 38556 72894 38612
rect 73350 38556 73388 38612
rect 73444 38556 73454 38612
rect 76402 38556 76412 38612
rect 76468 38556 77252 38612
rect 77196 38500 77252 38556
rect 75842 38444 75852 38500
rect 75908 38444 76524 38500
rect 76580 38444 76590 38500
rect 77186 38444 77196 38500
rect 77252 38444 77262 38500
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 65906 38388 65916 38444
rect 65972 38388 66020 38444
rect 66076 38388 66124 38444
rect 66180 38388 66190 38444
rect 69570 38332 69580 38388
rect 69636 38332 77308 38388
rect 77364 38332 77374 38388
rect 78530 38332 78540 38388
rect 78596 38332 79436 38388
rect 79492 38332 79502 38388
rect 70130 38220 70140 38276
rect 70196 38220 72268 38276
rect 72324 38220 72334 38276
rect 76150 38220 76188 38276
rect 76244 38220 76254 38276
rect 76626 38220 76636 38276
rect 76692 38220 77644 38276
rect 77700 38220 77710 38276
rect 0 38164 800 38192
rect 0 38108 3388 38164
rect 3444 38108 3454 38164
rect 69794 38108 69804 38164
rect 69860 38108 70588 38164
rect 70644 38108 70654 38164
rect 71260 38108 71932 38164
rect 71988 38108 71998 38164
rect 72566 38108 72604 38164
rect 72660 38108 72670 38164
rect 72902 38108 72940 38164
rect 72996 38108 73006 38164
rect 73154 38108 73164 38164
rect 73220 38108 75516 38164
rect 75572 38108 75582 38164
rect 76738 38108 76748 38164
rect 76804 38108 77980 38164
rect 78036 38108 78046 38164
rect 0 38080 800 38108
rect 71260 38052 71316 38108
rect 64754 37996 64764 38052
rect 64820 37996 71260 38052
rect 71316 37996 71326 38052
rect 71810 37996 71820 38052
rect 71876 37996 74284 38052
rect 74340 37996 74620 38052
rect 74676 37996 76188 38052
rect 76244 37996 76254 38052
rect 70914 37884 70924 37940
rect 70980 37884 71596 37940
rect 71652 37884 72268 37940
rect 72324 37884 72828 37940
rect 72884 37884 72894 37940
rect 73892 37884 74956 37940
rect 75012 37884 75022 37940
rect 67778 37772 67788 37828
rect 67844 37772 68684 37828
rect 68740 37772 69692 37828
rect 69748 37772 70588 37828
rect 70644 37772 70654 37828
rect 72706 37772 72716 37828
rect 72772 37772 73164 37828
rect 73220 37772 73612 37828
rect 73668 37772 73678 37828
rect 73892 37716 73948 37884
rect 75058 37772 75068 37828
rect 75124 37772 75404 37828
rect 75460 37772 76636 37828
rect 76692 37772 76702 37828
rect 79200 37716 80000 37744
rect 58706 37660 58716 37716
rect 58772 37660 73948 37716
rect 74004 37660 74014 37716
rect 75506 37660 75516 37716
rect 75572 37660 80000 37716
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 50546 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50830 37660
rect 79200 37632 80000 37660
rect 57026 37548 57036 37604
rect 57092 37548 76244 37604
rect 73938 37436 73948 37492
rect 74004 37436 74396 37492
rect 74452 37436 74462 37492
rect 2034 37324 2044 37380
rect 2100 37324 26908 37380
rect 26964 37324 26974 37380
rect 70578 37324 70588 37380
rect 70644 37324 71260 37380
rect 71316 37324 71326 37380
rect 72258 37324 72268 37380
rect 72324 37324 73052 37380
rect 73108 37324 73118 37380
rect 73350 37324 73388 37380
rect 73444 37324 73454 37380
rect 76188 37268 76244 37548
rect 77298 37436 77308 37492
rect 77364 37436 78540 37492
rect 78596 37436 78606 37492
rect 76626 37324 76636 37380
rect 76692 37324 77644 37380
rect 77700 37324 77710 37380
rect 73686 37212 73724 37268
rect 73780 37212 73790 37268
rect 75170 37212 75180 37268
rect 75236 37212 75964 37268
rect 76020 37212 76030 37268
rect 76178 37212 76188 37268
rect 76244 37212 76636 37268
rect 76692 37212 76702 37268
rect 72594 37100 72604 37156
rect 72660 37100 73276 37156
rect 73332 37100 73342 37156
rect 0 37044 800 37072
rect 0 36988 1708 37044
rect 1764 36988 2492 37044
rect 2548 36988 2558 37044
rect 74274 36988 74284 37044
rect 74340 36988 77644 37044
rect 77700 36988 77710 37044
rect 0 36960 800 36988
rect 74610 36876 74620 36932
rect 74676 36876 74956 36932
rect 75012 36876 77868 36932
rect 77924 36876 77934 36932
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 65906 36820 65916 36876
rect 65972 36820 66020 36876
rect 66076 36820 66124 36876
rect 66180 36820 66190 36876
rect 72902 36764 72940 36820
rect 72996 36764 73006 36820
rect 74274 36764 74284 36820
rect 74340 36764 78316 36820
rect 78372 36764 78382 36820
rect 74834 36652 74844 36708
rect 74900 36652 77308 36708
rect 77364 36652 77374 36708
rect 79200 36596 80000 36624
rect 57026 36540 57036 36596
rect 57092 36540 75852 36596
rect 75908 36540 75918 36596
rect 77634 36540 77644 36596
rect 77700 36540 80000 36596
rect 79200 36512 80000 36540
rect 72482 36428 72492 36484
rect 72548 36428 75404 36484
rect 75460 36428 75470 36484
rect 26898 36316 26908 36372
rect 26964 36316 44828 36372
rect 44884 36316 45388 36372
rect 45444 36316 45454 36372
rect 60610 36316 60620 36372
rect 60676 36316 73276 36372
rect 73332 36316 73342 36372
rect 73938 36316 73948 36372
rect 74004 36316 74042 36372
rect 74358 36316 74396 36372
rect 74452 36316 74462 36372
rect 2034 36204 2044 36260
rect 2100 36204 44268 36260
rect 44324 36204 44334 36260
rect 44930 36204 44940 36260
rect 44996 36204 46956 36260
rect 47012 36204 47022 36260
rect 61730 36204 61740 36260
rect 61796 36204 67564 36260
rect 67620 36204 69020 36260
rect 69076 36204 69356 36260
rect 69412 36204 69422 36260
rect 53778 36092 53788 36148
rect 53844 36092 77420 36148
rect 77476 36092 77486 36148
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 50546 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50830 36092
rect 52770 35980 52780 36036
rect 52836 35980 76412 36036
rect 76468 35980 76478 36036
rect 0 35924 800 35952
rect 0 35868 1708 35924
rect 1764 35868 2492 35924
rect 2548 35868 2558 35924
rect 77830 35868 77868 35924
rect 77924 35868 77934 35924
rect 0 35840 800 35868
rect 45826 35756 45836 35812
rect 45892 35756 46620 35812
rect 46676 35756 46686 35812
rect 73938 35756 73948 35812
rect 74004 35756 75292 35812
rect 75348 35756 75358 35812
rect 76850 35756 76860 35812
rect 76916 35756 77980 35812
rect 78036 35756 78652 35812
rect 78708 35756 78718 35812
rect 44706 35644 44716 35700
rect 44772 35644 45388 35700
rect 45444 35644 45454 35700
rect 73892 35644 75740 35700
rect 75796 35644 75806 35700
rect 73892 35588 73948 35644
rect 45602 35532 45612 35588
rect 45668 35532 45678 35588
rect 46834 35532 46844 35588
rect 46900 35532 54460 35588
rect 54516 35532 54526 35588
rect 70578 35532 70588 35588
rect 70644 35532 71708 35588
rect 71764 35532 72604 35588
rect 72660 35532 73948 35588
rect 45612 35364 45668 35532
rect 79200 35476 80000 35504
rect 75394 35420 75404 35476
rect 75460 35420 76748 35476
rect 76804 35420 76814 35476
rect 78306 35420 78316 35476
rect 78372 35420 80000 35476
rect 79200 35392 80000 35420
rect 45612 35308 54236 35364
rect 54292 35308 54302 35364
rect 73714 35308 73724 35364
rect 73780 35308 74060 35364
rect 74116 35308 74126 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 65906 35252 65916 35308
rect 65972 35252 66020 35308
rect 66076 35252 66124 35308
rect 66180 35252 66190 35308
rect 71474 35196 71484 35252
rect 71540 35196 72268 35252
rect 72324 35196 72334 35252
rect 72706 35196 72716 35252
rect 72772 35196 72782 35252
rect 74162 35196 74172 35252
rect 74228 35196 78988 35252
rect 79044 35196 79054 35252
rect 72716 35140 72772 35196
rect 62132 35084 72772 35140
rect 72902 35084 72940 35140
rect 72996 35084 73006 35140
rect 77830 35084 77868 35140
rect 77924 35084 77934 35140
rect 62132 35028 62188 35084
rect 55412 34972 55580 35028
rect 55636 34972 62188 35028
rect 71250 34972 71260 35028
rect 71316 34972 71932 35028
rect 71988 34972 71998 35028
rect 72146 34972 72156 35028
rect 72212 34972 77308 35028
rect 77364 34972 77374 35028
rect 77522 34972 77532 35028
rect 77588 34972 79324 35028
rect 79380 34972 79390 35028
rect 55412 34916 55468 34972
rect 45602 34860 45612 34916
rect 45668 34860 53564 34916
rect 53620 34860 53630 34916
rect 54786 34860 54796 34916
rect 54852 34860 55468 34916
rect 71586 34860 71596 34916
rect 71652 34860 71820 34916
rect 71876 34860 73276 34916
rect 73332 34860 73500 34916
rect 73556 34860 73566 34916
rect 0 34804 800 34832
rect 0 34748 1708 34804
rect 1764 34748 2492 34804
rect 2548 34748 2558 34804
rect 70914 34748 70924 34804
rect 70980 34748 72380 34804
rect 72436 34748 72828 34804
rect 72884 34748 72894 34804
rect 0 34720 800 34748
rect 73892 34692 73948 34972
rect 74918 34860 74956 34916
rect 75012 34860 75022 34916
rect 75618 34860 75628 34916
rect 75684 34860 78204 34916
rect 78260 34860 78270 34916
rect 74386 34748 74396 34804
rect 74452 34748 74732 34804
rect 74788 34748 79044 34804
rect 2034 34636 2044 34692
rect 2100 34636 44380 34692
rect 44436 34636 44828 34692
rect 44884 34636 44894 34692
rect 70802 34636 70812 34692
rect 70868 34636 71932 34692
rect 71988 34636 71998 34692
rect 72258 34636 72268 34692
rect 72324 34636 72380 34692
rect 72436 34636 72446 34692
rect 73378 34636 73388 34692
rect 73444 34636 73948 34692
rect 75730 34636 75740 34692
rect 75796 34636 77588 34692
rect 77532 34580 77588 34636
rect 52322 34524 52332 34580
rect 52388 34524 76524 34580
rect 76580 34524 76590 34580
rect 77522 34524 77532 34580
rect 77588 34524 77598 34580
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 50546 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50830 34524
rect 70532 34412 72940 34468
rect 72996 34412 73006 34468
rect 76626 34412 76636 34468
rect 76692 34412 78092 34468
rect 78148 34412 78764 34468
rect 78820 34412 78830 34468
rect 54562 34300 54572 34356
rect 54628 34300 55468 34356
rect 55524 34300 57036 34356
rect 57092 34300 57102 34356
rect 2034 34188 2044 34244
rect 2100 34188 44156 34244
rect 44212 34188 44222 34244
rect 53330 34188 53340 34244
rect 53396 34188 53788 34244
rect 53844 34188 54012 34244
rect 54068 34188 54078 34244
rect 45714 34076 45724 34132
rect 45780 34076 53004 34132
rect 53060 34076 53070 34132
rect 70532 33908 70588 34412
rect 78988 34356 79044 34748
rect 79200 34356 80000 34384
rect 70802 34300 70812 34356
rect 70868 34300 71260 34356
rect 71316 34300 71326 34356
rect 73266 34300 73276 34356
rect 73332 34300 73836 34356
rect 73892 34300 74172 34356
rect 74228 34300 74238 34356
rect 75730 34300 75740 34356
rect 75796 34300 75806 34356
rect 75926 34300 75964 34356
rect 76020 34300 76030 34356
rect 76178 34300 76188 34356
rect 76244 34300 78204 34356
rect 78260 34300 78270 34356
rect 78988 34300 80000 34356
rect 75740 34244 75796 34300
rect 79200 34272 80000 34300
rect 71362 34188 71372 34244
rect 71428 34188 75796 34244
rect 76290 34188 76300 34244
rect 76356 34188 77084 34244
rect 77140 34188 77150 34244
rect 73378 34076 73388 34132
rect 73444 34076 74396 34132
rect 74452 34076 74462 34132
rect 74722 34076 74732 34132
rect 74788 34076 76412 34132
rect 76468 34076 76478 34132
rect 76962 34076 76972 34132
rect 77028 34076 77644 34132
rect 77700 34076 77710 34132
rect 75282 33964 75292 34020
rect 75348 33964 77308 34020
rect 77364 33964 77374 34020
rect 64642 33852 64652 33908
rect 64708 33852 70588 33908
rect 74946 33852 74956 33908
rect 75012 33852 76860 33908
rect 76916 33852 76926 33908
rect 52994 33740 53004 33796
rect 53060 33740 53564 33796
rect 53620 33740 53630 33796
rect 73490 33740 73500 33796
rect 73556 33740 73836 33796
rect 73892 33740 73902 33796
rect 0 33684 800 33712
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 65906 33684 65916 33740
rect 65972 33684 66020 33740
rect 66076 33684 66124 33740
rect 66180 33684 66190 33740
rect 0 33628 1708 33684
rect 1764 33628 2492 33684
rect 2548 33628 2558 33684
rect 0 33600 800 33628
rect 75618 33516 75628 33572
rect 75684 33516 77868 33572
rect 77924 33516 77934 33572
rect 78764 33516 79100 33572
rect 79156 33516 79166 33572
rect 72034 33404 72044 33460
rect 72100 33404 72716 33460
rect 72772 33404 73948 33460
rect 76514 33404 76524 33460
rect 76580 33404 76636 33460
rect 76692 33404 76702 33460
rect 78194 33404 78204 33460
rect 78260 33404 78540 33460
rect 78596 33404 78606 33460
rect 73892 33348 73948 33404
rect 78764 33348 78820 33516
rect 44482 33292 44492 33348
rect 44548 33292 45388 33348
rect 45444 33292 45454 33348
rect 45826 33292 45836 33348
rect 45892 33292 46396 33348
rect 46452 33292 46462 33348
rect 72566 33292 72604 33348
rect 72660 33292 72670 33348
rect 72930 33292 72940 33348
rect 72996 33292 73276 33348
rect 73332 33292 73342 33348
rect 73892 33292 78820 33348
rect 79200 33236 80000 33264
rect 62066 33180 62076 33236
rect 62132 33180 74396 33236
rect 74452 33180 74462 33236
rect 75170 33180 75180 33236
rect 75236 33180 77084 33236
rect 77140 33180 77150 33236
rect 78530 33180 78540 33236
rect 78596 33180 80000 33236
rect 79200 33152 80000 33180
rect 2034 33068 2044 33124
rect 2100 33068 28476 33124
rect 28532 33068 28542 33124
rect 75618 33068 75628 33124
rect 75684 33068 75852 33124
rect 75908 33068 75918 33124
rect 74470 32956 74508 33012
rect 74564 32956 74574 33012
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 50546 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50830 32956
rect 66994 32844 67004 32900
rect 67060 32844 68012 32900
rect 68068 32844 68078 32900
rect 69906 32844 69916 32900
rect 69972 32844 75796 32900
rect 45490 32732 45500 32788
rect 45556 32732 46508 32788
rect 46564 32732 46574 32788
rect 53666 32732 53676 32788
rect 53732 32732 74732 32788
rect 74788 32732 74798 32788
rect 75740 32676 75796 32844
rect 72342 32620 72380 32676
rect 72436 32620 72446 32676
rect 74946 32620 74956 32676
rect 75012 32620 75180 32676
rect 75236 32620 75246 32676
rect 75730 32620 75740 32676
rect 75796 32620 75806 32676
rect 76850 32620 76860 32676
rect 76916 32620 78428 32676
rect 78484 32620 78494 32676
rect 0 32564 800 32592
rect 0 32508 1708 32564
rect 1764 32508 2492 32564
rect 2548 32508 2558 32564
rect 71250 32508 71260 32564
rect 71316 32508 72828 32564
rect 72884 32508 73164 32564
rect 73220 32508 73230 32564
rect 0 32480 800 32508
rect 71558 32396 71596 32452
rect 71652 32396 71662 32452
rect 72370 32396 72380 32452
rect 72436 32396 72604 32452
rect 72660 32396 72670 32452
rect 75282 32396 75292 32452
rect 75348 32396 76076 32452
rect 76132 32396 76142 32452
rect 73714 32284 73724 32340
rect 73780 32284 74508 32340
rect 74564 32284 74574 32340
rect 75058 32172 75068 32228
rect 75124 32172 77868 32228
rect 77924 32172 77934 32228
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 65906 32116 65916 32172
rect 65972 32116 66020 32172
rect 66076 32116 66124 32172
rect 66180 32116 66190 32172
rect 79200 32116 80000 32144
rect 74050 32060 74060 32116
rect 74116 32060 74844 32116
rect 74900 32060 80000 32116
rect 79200 32032 80000 32060
rect 52546 31948 52556 32004
rect 52612 31948 53676 32004
rect 53732 31948 53742 32004
rect 70578 31948 70588 32004
rect 70644 31948 72436 32004
rect 73938 31948 73948 32004
rect 74004 31948 75180 32004
rect 75236 31948 75246 32004
rect 77074 31948 77084 32004
rect 77140 31948 77532 32004
rect 77588 31948 77598 32004
rect 72380 31892 72436 31948
rect 31892 31836 45276 31892
rect 45332 31836 45342 31892
rect 71362 31836 71372 31892
rect 71428 31836 71932 31892
rect 71988 31836 71998 31892
rect 72370 31836 72380 31892
rect 72436 31836 74732 31892
rect 74788 31836 75292 31892
rect 75348 31836 75358 31892
rect 31892 31780 31948 31836
rect 77532 31780 77588 31948
rect 2034 31724 2044 31780
rect 2100 31724 31948 31780
rect 44930 31724 44940 31780
rect 44996 31724 45724 31780
rect 45780 31724 45790 31780
rect 45938 31724 45948 31780
rect 46004 31724 51436 31780
rect 51492 31724 51502 31780
rect 64754 31724 64764 31780
rect 64820 31724 75068 31780
rect 75124 31724 75134 31780
rect 76290 31724 76300 31780
rect 76356 31724 76412 31780
rect 76468 31724 76478 31780
rect 77522 31724 77532 31780
rect 77588 31724 77598 31780
rect 76300 31668 76356 31724
rect 28466 31612 28476 31668
rect 28532 31612 44380 31668
rect 44436 31612 44828 31668
rect 44884 31612 44894 31668
rect 51538 31612 51548 31668
rect 51604 31612 52780 31668
rect 52836 31612 52846 31668
rect 72706 31612 72716 31668
rect 72772 31612 76356 31668
rect 73714 31500 73724 31556
rect 73780 31500 73948 31556
rect 0 31444 800 31472
rect 0 31388 1708 31444
rect 1764 31388 2492 31444
rect 2548 31388 2558 31444
rect 72482 31388 72492 31444
rect 72548 31388 72604 31444
rect 72660 31388 73388 31444
rect 73444 31388 73454 31444
rect 0 31360 800 31388
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 50546 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50830 31388
rect 73892 31332 73948 31500
rect 74284 31500 76300 31556
rect 76356 31500 76366 31556
rect 74284 31332 74340 31500
rect 73892 31276 74340 31332
rect 75394 31276 75404 31332
rect 75460 31276 75740 31332
rect 75796 31276 76860 31332
rect 76916 31276 76926 31332
rect 74050 31164 74060 31220
rect 74116 31164 76748 31220
rect 76804 31164 76814 31220
rect 77298 31164 77308 31220
rect 77364 31164 78092 31220
rect 78148 31164 78158 31220
rect 2034 31052 2044 31108
rect 2100 31052 44156 31108
rect 44212 31052 44222 31108
rect 45490 31052 45500 31108
rect 45556 31052 46284 31108
rect 46340 31052 46350 31108
rect 60386 31052 60396 31108
rect 60452 31052 74172 31108
rect 74228 31052 74238 31108
rect 79200 30996 80000 31024
rect 45266 30940 45276 30996
rect 45332 30940 45612 30996
rect 45668 30940 45678 30996
rect 71362 30940 71372 30996
rect 71428 30940 71708 30996
rect 71764 30940 72268 30996
rect 72324 30940 72334 30996
rect 75170 30940 75180 30996
rect 75236 30940 75404 30996
rect 75460 30940 80000 30996
rect 79200 30912 80000 30940
rect 1698 30828 1708 30884
rect 1764 30828 2492 30884
rect 2548 30828 2558 30884
rect 45938 30828 45948 30884
rect 46004 30828 51436 30884
rect 51492 30828 51502 30884
rect 52882 30828 52892 30884
rect 52948 30828 53340 30884
rect 53396 30828 53406 30884
rect 72034 30828 72044 30884
rect 72100 30828 75628 30884
rect 75684 30828 75694 30884
rect 45490 30716 45500 30772
rect 45556 30716 46508 30772
rect 46564 30716 46574 30772
rect 50530 30716 50540 30772
rect 50596 30716 71932 30772
rect 71988 30716 71998 30772
rect 74610 30716 74620 30772
rect 74676 30716 78092 30772
rect 78148 30716 78158 30772
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 65906 30548 65916 30604
rect 65972 30548 66020 30604
rect 66076 30548 66124 30604
rect 66180 30548 66190 30604
rect 50082 30492 50092 30548
rect 50148 30492 58828 30548
rect 70690 30492 70700 30548
rect 70756 30492 71820 30548
rect 71876 30492 71886 30548
rect 73938 30492 73948 30548
rect 74004 30492 77532 30548
rect 77588 30492 77598 30548
rect 58772 30436 58828 30492
rect 46050 30380 46060 30436
rect 46116 30380 52444 30436
rect 52500 30380 52510 30436
rect 58772 30380 72828 30436
rect 72884 30380 72894 30436
rect 74274 30380 74284 30436
rect 74340 30380 77644 30436
rect 77700 30380 77710 30436
rect 0 30324 800 30352
rect 0 30268 1708 30324
rect 1764 30268 1774 30324
rect 46274 30268 46284 30324
rect 46340 30268 46732 30324
rect 46788 30268 46798 30324
rect 51762 30268 51772 30324
rect 51828 30268 52332 30324
rect 52388 30268 52892 30324
rect 52948 30268 52958 30324
rect 70690 30268 70700 30324
rect 70756 30268 76412 30324
rect 76468 30268 76478 30324
rect 0 30240 800 30268
rect 44482 30156 44492 30212
rect 44548 30156 45724 30212
rect 45780 30156 45790 30212
rect 46162 30156 46172 30212
rect 46228 30156 46956 30212
rect 47012 30156 47022 30212
rect 47170 30156 47180 30212
rect 47236 30156 50876 30212
rect 50932 30156 50942 30212
rect 71362 30156 71372 30212
rect 71428 30156 76860 30212
rect 76916 30156 76926 30212
rect 78194 30156 78204 30212
rect 78260 30156 78540 30212
rect 78596 30156 78606 30212
rect 44930 30044 44940 30100
rect 44996 30044 47292 30100
rect 47348 30044 47358 30100
rect 51202 30044 51212 30100
rect 51268 30044 51996 30100
rect 52052 30044 62076 30100
rect 62132 30044 62142 30100
rect 75506 30044 75516 30100
rect 75572 30044 76076 30100
rect 76132 30044 76142 30100
rect 76514 30044 76524 30100
rect 76580 30044 77308 30100
rect 77364 30044 78876 30100
rect 78932 30044 78942 30100
rect 71138 29932 71148 29988
rect 71204 29932 72156 29988
rect 72212 29932 72222 29988
rect 74386 29932 74396 29988
rect 74452 29932 76300 29988
rect 76356 29932 76366 29988
rect 79200 29876 80000 29904
rect 77858 29820 77868 29876
rect 77924 29820 80000 29876
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 50546 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50830 29820
rect 79200 29792 80000 29820
rect 71810 29708 71820 29764
rect 71876 29708 76972 29764
rect 77028 29708 77038 29764
rect 75618 29596 75628 29652
rect 75684 29596 77756 29652
rect 77812 29596 77822 29652
rect 2034 29484 2044 29540
rect 2100 29484 44604 29540
rect 44660 29484 44670 29540
rect 76066 29484 76076 29540
rect 76132 29484 76524 29540
rect 76580 29484 76590 29540
rect 49718 29372 49756 29428
rect 49812 29372 49822 29428
rect 72258 29372 72268 29428
rect 72324 29372 73500 29428
rect 73556 29372 73566 29428
rect 73714 29372 73724 29428
rect 73780 29372 75628 29428
rect 75684 29372 75694 29428
rect 75842 29372 75852 29428
rect 75908 29372 75964 29428
rect 76020 29372 76030 29428
rect 0 29204 800 29232
rect 0 29148 1708 29204
rect 1764 29148 2492 29204
rect 2548 29148 2558 29204
rect 48066 29148 48076 29204
rect 48132 29148 74060 29204
rect 74116 29148 74126 29204
rect 0 29120 800 29148
rect 36082 29036 36092 29092
rect 36148 29036 37100 29092
rect 37156 29036 37166 29092
rect 70914 29036 70924 29092
rect 70980 29036 78204 29092
rect 78260 29036 78270 29092
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 65906 28980 65916 29036
rect 65972 28980 66020 29036
rect 66076 28980 66124 29036
rect 66180 28980 66190 29036
rect 66658 28924 66668 28980
rect 66724 28924 72716 28980
rect 72772 28924 72782 28980
rect 74722 28924 74732 28980
rect 74788 28924 75516 28980
rect 75572 28924 75582 28980
rect 77410 28924 77420 28980
rect 77476 28924 79100 28980
rect 79156 28924 79166 28980
rect 72482 28812 72492 28868
rect 72548 28812 74396 28868
rect 74452 28812 75068 28868
rect 75124 28812 75134 28868
rect 79200 28756 80000 28784
rect 2034 28700 2044 28756
rect 2100 28700 38668 28756
rect 60274 28700 60284 28756
rect 60340 28700 72828 28756
rect 72884 28700 73500 28756
rect 73556 28700 73566 28756
rect 73892 28700 80000 28756
rect 38612 28644 38668 28700
rect 73892 28644 73948 28700
rect 79200 28672 80000 28700
rect 38612 28588 43708 28644
rect 49186 28588 49196 28644
rect 49252 28588 70812 28644
rect 70868 28588 70878 28644
rect 72594 28588 72604 28644
rect 72660 28588 73724 28644
rect 73780 28588 73948 28644
rect 74722 28588 74732 28644
rect 74788 28588 76076 28644
rect 76132 28588 76142 28644
rect 76514 28588 76524 28644
rect 76580 28588 76860 28644
rect 76916 28588 76926 28644
rect 77074 28588 77084 28644
rect 77140 28588 77644 28644
rect 77700 28588 77710 28644
rect 43652 28532 43708 28588
rect 39778 28476 39788 28532
rect 39844 28476 40684 28532
rect 40740 28476 42588 28532
rect 42644 28476 42654 28532
rect 43652 28476 44716 28532
rect 44772 28476 44782 28532
rect 45042 28476 45052 28532
rect 45108 28476 45836 28532
rect 45892 28476 45902 28532
rect 71474 28476 71484 28532
rect 71540 28476 71820 28532
rect 71876 28476 72380 28532
rect 72436 28476 72446 28532
rect 72706 28476 72716 28532
rect 72772 28476 73836 28532
rect 73892 28476 73902 28532
rect 75618 28476 75628 28532
rect 75684 28476 76524 28532
rect 76580 28476 77868 28532
rect 77924 28476 77934 28532
rect 64530 28364 64540 28420
rect 64596 28364 72492 28420
rect 72548 28364 72558 28420
rect 75170 28364 75180 28420
rect 75236 28364 75404 28420
rect 75460 28364 76636 28420
rect 76692 28364 76702 28420
rect 71810 28252 71820 28308
rect 71876 28252 74676 28308
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 50546 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50830 28252
rect 68898 28140 68908 28196
rect 68964 28140 73948 28196
rect 74004 28140 74396 28196
rect 74452 28140 74462 28196
rect 0 28084 800 28112
rect 74620 28084 74676 28252
rect 77196 28252 77420 28308
rect 77476 28252 77486 28308
rect 77196 28196 77252 28252
rect 75628 28140 77252 28196
rect 75628 28084 75684 28140
rect 0 28028 1708 28084
rect 1764 28028 2492 28084
rect 2548 28028 2558 28084
rect 30146 28028 30156 28084
rect 30212 28028 35812 28084
rect 35970 28028 35980 28084
rect 36036 28028 36988 28084
rect 37044 28028 37054 28084
rect 38098 28028 38108 28084
rect 38164 28028 39340 28084
rect 39396 28028 39406 28084
rect 41682 28028 41692 28084
rect 41748 28028 41916 28084
rect 41972 28028 42476 28084
rect 42532 28028 42542 28084
rect 50372 28028 68068 28084
rect 72818 28028 72828 28084
rect 72884 28028 73724 28084
rect 73780 28028 73790 28084
rect 74620 28028 75684 28084
rect 0 28000 800 28028
rect 35756 27972 35812 28028
rect 50372 27972 50428 28028
rect 20962 27916 20972 27972
rect 21028 27916 31948 27972
rect 33842 27916 33852 27972
rect 33908 27916 34860 27972
rect 34916 27916 34926 27972
rect 35756 27916 40236 27972
rect 40292 27916 40302 27972
rect 41346 27916 41356 27972
rect 41412 27916 50428 27972
rect 31892 27860 31948 27916
rect 31892 27804 40124 27860
rect 40180 27804 40190 27860
rect 40338 27804 40348 27860
rect 40404 27804 41468 27860
rect 41524 27804 41534 27860
rect 40348 27748 40404 27804
rect 31826 27692 31836 27748
rect 31892 27692 40404 27748
rect 68012 27748 68068 28028
rect 70700 27916 73948 27972
rect 74946 27916 74956 27972
rect 75012 27916 75628 27972
rect 75684 27916 75694 27972
rect 75842 27916 75852 27972
rect 75908 27916 77756 27972
rect 77812 27916 77822 27972
rect 70700 27860 70756 27916
rect 73892 27860 73948 27916
rect 70690 27804 70700 27860
rect 70756 27804 70766 27860
rect 71894 27804 71932 27860
rect 71988 27804 71998 27860
rect 73154 27804 73164 27860
rect 73220 27804 73230 27860
rect 73892 27804 76748 27860
rect 76804 27804 76814 27860
rect 68012 27692 72268 27748
rect 72324 27692 72334 27748
rect 73164 27636 73220 27804
rect 73686 27692 73724 27748
rect 73780 27692 73790 27748
rect 74274 27692 74284 27748
rect 74340 27692 74732 27748
rect 74788 27692 74798 27748
rect 79200 27636 80000 27664
rect 33506 27580 33516 27636
rect 33572 27580 38668 27636
rect 38724 27580 38734 27636
rect 40114 27580 40124 27636
rect 40180 27580 42476 27636
rect 42532 27580 42542 27636
rect 68124 27580 72716 27636
rect 72772 27580 72782 27636
rect 73164 27580 74060 27636
rect 74116 27580 74126 27636
rect 76850 27580 76860 27636
rect 76916 27580 76972 27636
rect 77028 27580 77038 27636
rect 78194 27580 78204 27636
rect 78260 27580 80000 27636
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 65906 27412 65916 27468
rect 65972 27412 66020 27468
rect 66076 27412 66124 27468
rect 66180 27412 66190 27468
rect 43810 27356 43820 27412
rect 43876 27356 50876 27412
rect 50932 27356 50942 27412
rect 2034 27244 2044 27300
rect 2100 27244 44828 27300
rect 44884 27244 45388 27300
rect 45444 27244 45454 27300
rect 46610 27244 46620 27300
rect 46676 27244 48972 27300
rect 49028 27244 49038 27300
rect 42130 27132 42140 27188
rect 42196 27132 43036 27188
rect 43092 27132 43102 27188
rect 44034 27132 44044 27188
rect 44100 27132 45836 27188
rect 45892 27132 45902 27188
rect 49074 27132 49084 27188
rect 49140 27132 50204 27188
rect 50260 27132 50428 27188
rect 50372 27076 50428 27132
rect 34850 27020 34860 27076
rect 34916 27020 35532 27076
rect 35588 27020 35598 27076
rect 47506 27020 47516 27076
rect 47572 27020 49532 27076
rect 49588 27020 49598 27076
rect 50372 27020 60396 27076
rect 60452 27020 60462 27076
rect 0 26964 800 26992
rect 68124 26964 68180 27580
rect 70690 27468 70700 27524
rect 70756 27468 76524 27524
rect 76580 27468 76590 27524
rect 76860 27412 76916 27580
rect 79200 27552 80000 27580
rect 70130 27356 70140 27412
rect 70196 27356 76916 27412
rect 71922 27244 71932 27300
rect 71988 27244 76860 27300
rect 76916 27244 76926 27300
rect 77186 27244 77196 27300
rect 77252 27244 77532 27300
rect 77588 27244 77598 27300
rect 72258 27132 72268 27188
rect 72324 27132 74620 27188
rect 74676 27132 74686 27188
rect 72706 27020 72716 27076
rect 72772 27020 73164 27076
rect 73220 27020 73230 27076
rect 73490 27020 73500 27076
rect 73556 27020 73566 27076
rect 74022 27020 74060 27076
rect 74116 27020 74126 27076
rect 74946 27020 74956 27076
rect 75012 27020 75292 27076
rect 75348 27020 75358 27076
rect 77410 27020 77420 27076
rect 77476 27020 77868 27076
rect 77924 27020 77934 27076
rect 0 26908 1708 26964
rect 1764 26908 2492 26964
rect 2548 26908 2558 26964
rect 40002 26908 40012 26964
rect 40068 26908 41692 26964
rect 41748 26908 41758 26964
rect 44930 26908 44940 26964
rect 44996 26908 47292 26964
rect 47348 26908 47358 26964
rect 49634 26908 49644 26964
rect 49700 26908 50652 26964
rect 50708 26908 68180 26964
rect 73500 26964 73556 27020
rect 73500 26908 74732 26964
rect 74788 26908 76188 26964
rect 76244 26908 76254 26964
rect 0 26880 800 26908
rect 36306 26796 36316 26852
rect 36372 26796 73948 26852
rect 74050 26796 74060 26852
rect 74116 26796 74956 26852
rect 75012 26796 75022 26852
rect 72706 26684 72716 26740
rect 72772 26684 72940 26740
rect 72996 26684 73006 26740
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 50546 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50830 26684
rect 73892 26628 73948 26796
rect 74274 26684 74284 26740
rect 74340 26684 77756 26740
rect 77812 26684 77822 26740
rect 73892 26572 74228 26628
rect 74610 26572 74620 26628
rect 74676 26572 76804 26628
rect 74172 26516 74228 26572
rect 76748 26516 76804 26572
rect 79200 26516 80000 26544
rect 33730 26460 33740 26516
rect 33796 26460 34300 26516
rect 34356 26460 35812 26516
rect 36978 26460 36988 26516
rect 37044 26460 41356 26516
rect 41412 26460 42364 26516
rect 42420 26460 42430 26516
rect 46050 26460 46060 26516
rect 46116 26460 46732 26516
rect 46788 26460 46798 26516
rect 48850 26460 48860 26516
rect 48916 26460 50092 26516
rect 50148 26460 50158 26516
rect 35756 26404 35812 26460
rect 50372 26404 50428 26516
rect 50484 26460 50494 26516
rect 64194 26460 64204 26516
rect 64260 26460 72492 26516
rect 72548 26460 72558 26516
rect 73266 26460 73276 26516
rect 73332 26460 73836 26516
rect 73892 26460 73902 26516
rect 74172 26460 74676 26516
rect 75842 26460 75852 26516
rect 75908 26460 76188 26516
rect 76244 26460 76254 26516
rect 76748 26460 80000 26516
rect 74620 26404 74676 26460
rect 79200 26432 80000 26460
rect 34850 26348 34860 26404
rect 34916 26348 35532 26404
rect 35588 26348 35598 26404
rect 35746 26348 35756 26404
rect 35812 26348 36428 26404
rect 36484 26348 36494 26404
rect 38210 26348 38220 26404
rect 38276 26348 39116 26404
rect 39172 26348 39182 26404
rect 46162 26348 46172 26404
rect 46228 26348 46844 26404
rect 46900 26348 47740 26404
rect 47796 26348 47806 26404
rect 49410 26348 49420 26404
rect 49476 26348 50428 26404
rect 74610 26348 74620 26404
rect 74676 26348 74686 26404
rect 35186 26236 35196 26292
rect 35252 26236 37212 26292
rect 37268 26236 37278 26292
rect 38770 26236 38780 26292
rect 38836 26236 40012 26292
rect 40068 26236 40078 26292
rect 41682 26236 41692 26292
rect 41748 26236 42028 26292
rect 42084 26236 42924 26292
rect 42980 26236 42990 26292
rect 45042 26236 45052 26292
rect 45108 26236 46396 26292
rect 46452 26236 46462 26292
rect 46610 26236 46620 26292
rect 46676 26236 48748 26292
rect 48804 26236 48814 26292
rect 49634 26236 49644 26292
rect 49700 26236 49980 26292
rect 50036 26236 50046 26292
rect 70914 26236 70924 26292
rect 70980 26236 73444 26292
rect 73826 26236 73836 26292
rect 73892 26236 77644 26292
rect 77700 26236 77710 26292
rect 34290 26124 34300 26180
rect 34356 26124 36988 26180
rect 37044 26124 37054 26180
rect 46946 26124 46956 26180
rect 47012 26124 47852 26180
rect 47908 26124 47918 26180
rect 49718 26124 49756 26180
rect 49812 26124 49822 26180
rect 58594 26124 58604 26180
rect 58660 26124 73164 26180
rect 73220 26124 73230 26180
rect 73388 26068 73444 26236
rect 74722 26124 74732 26180
rect 74788 26124 75852 26180
rect 75908 26124 75918 26180
rect 2034 26012 2044 26068
rect 2100 26012 44940 26068
rect 44996 26012 45500 26068
rect 45556 26012 45566 26068
rect 47506 26012 47516 26068
rect 47572 26012 49308 26068
rect 49364 26012 49374 26068
rect 73388 26012 77644 26068
rect 77700 26012 77710 26068
rect 72594 25900 72604 25956
rect 72660 25900 73500 25956
rect 73556 25900 73566 25956
rect 0 25844 800 25872
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 65906 25844 65916 25900
rect 65972 25844 66020 25900
rect 66076 25844 66124 25900
rect 66180 25844 66190 25900
rect 0 25788 1708 25844
rect 1764 25788 2492 25844
rect 2548 25788 2558 25844
rect 37314 25788 37324 25844
rect 37380 25788 50428 25844
rect 71362 25788 71372 25844
rect 71428 25788 72884 25844
rect 76962 25788 76972 25844
rect 77028 25788 77868 25844
rect 77924 25788 77934 25844
rect 0 25760 800 25788
rect 50372 25732 50428 25788
rect 72828 25732 72884 25788
rect 25554 25676 25564 25732
rect 25620 25676 26572 25732
rect 26628 25676 37660 25732
rect 37716 25676 37726 25732
rect 41906 25676 41916 25732
rect 41972 25676 43036 25732
rect 43092 25676 43484 25732
rect 43540 25676 45500 25732
rect 45556 25676 45566 25732
rect 50372 25676 71260 25732
rect 71316 25676 71326 25732
rect 72566 25676 72604 25732
rect 72660 25676 72670 25732
rect 72828 25676 78204 25732
rect 78260 25676 78270 25732
rect 2034 25564 2044 25620
rect 2100 25564 26908 25620
rect 37202 25564 37212 25620
rect 37268 25564 40460 25620
rect 40516 25564 42028 25620
rect 42084 25564 43708 25620
rect 43764 25564 43774 25620
rect 45826 25564 45836 25620
rect 45892 25564 46508 25620
rect 46564 25564 46574 25620
rect 50372 25564 72940 25620
rect 72996 25564 73006 25620
rect 26852 25396 26908 25564
rect 31826 25452 31836 25508
rect 31892 25452 36652 25508
rect 36708 25452 36718 25508
rect 37762 25452 37772 25508
rect 37828 25452 38332 25508
rect 38388 25452 38780 25508
rect 38836 25452 38846 25508
rect 41010 25452 41020 25508
rect 41076 25452 41356 25508
rect 41412 25452 41422 25508
rect 43362 25452 43372 25508
rect 43428 25452 44268 25508
rect 44324 25452 44940 25508
rect 44996 25452 45006 25508
rect 45602 25452 45612 25508
rect 45668 25452 46060 25508
rect 46116 25452 46126 25508
rect 26852 25340 46956 25396
rect 47012 25340 47516 25396
rect 47572 25340 47582 25396
rect 50372 25284 50428 25564
rect 64418 25452 64428 25508
rect 64484 25452 70924 25508
rect 70980 25452 70990 25508
rect 71922 25452 71932 25508
rect 71988 25452 75460 25508
rect 76514 25452 76524 25508
rect 76580 25452 77420 25508
rect 77476 25452 77486 25508
rect 75404 25396 75460 25452
rect 79200 25396 80000 25424
rect 70466 25340 70476 25396
rect 70532 25340 73948 25396
rect 75394 25340 75404 25396
rect 75460 25340 80000 25396
rect 73892 25284 73948 25340
rect 79200 25312 80000 25340
rect 34738 25228 34748 25284
rect 34804 25228 35532 25284
rect 35588 25228 35598 25284
rect 35970 25228 35980 25284
rect 36036 25228 36652 25284
rect 36708 25228 36718 25284
rect 37762 25228 37772 25284
rect 37828 25228 38220 25284
rect 38276 25228 38286 25284
rect 38658 25228 38668 25284
rect 38724 25228 39676 25284
rect 39732 25228 39742 25284
rect 42242 25228 42252 25284
rect 42308 25228 42812 25284
rect 42868 25228 44604 25284
rect 44660 25228 44670 25284
rect 45826 25228 45836 25284
rect 45892 25228 50428 25284
rect 71586 25228 71596 25284
rect 71652 25228 72940 25284
rect 72996 25228 73006 25284
rect 73892 25228 76188 25284
rect 76244 25228 76254 25284
rect 63186 25116 63196 25172
rect 63252 25116 71708 25172
rect 71764 25116 72156 25172
rect 72212 25116 72222 25172
rect 75730 25116 75740 25172
rect 75796 25116 77084 25172
rect 77140 25116 77150 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 50546 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50830 25116
rect 63298 25004 63308 25060
rect 63364 25004 64652 25060
rect 64708 25004 64718 25060
rect 70242 25004 70252 25060
rect 70308 25004 71036 25060
rect 71092 25004 71102 25060
rect 71782 25004 71820 25060
rect 71876 25004 71886 25060
rect 72230 25004 72268 25060
rect 72324 25004 72334 25060
rect 75618 25004 75628 25060
rect 75684 25004 76524 25060
rect 76580 25004 76590 25060
rect 32610 24892 32620 24948
rect 32676 24892 36876 24948
rect 36932 24892 36942 24948
rect 50372 24892 74060 24948
rect 74116 24892 74126 24948
rect 75618 24892 75628 24948
rect 75684 24892 77756 24948
rect 77812 24892 77822 24948
rect 35522 24780 35532 24836
rect 35588 24780 35980 24836
rect 36036 24780 36046 24836
rect 40338 24780 40348 24836
rect 40404 24780 41244 24836
rect 41300 24780 44828 24836
rect 44884 24780 45164 24836
rect 45220 24780 45230 24836
rect 0 24724 800 24752
rect 50372 24724 50428 24892
rect 73714 24780 73724 24836
rect 73780 24780 77700 24836
rect 77644 24724 77700 24780
rect 0 24668 1708 24724
rect 1764 24668 2492 24724
rect 2548 24668 2558 24724
rect 19730 24668 19740 24724
rect 19796 24668 19806 24724
rect 20290 24668 20300 24724
rect 20356 24668 21196 24724
rect 21252 24668 21262 24724
rect 34962 24668 34972 24724
rect 35028 24668 35308 24724
rect 35364 24668 50428 24724
rect 72706 24668 72716 24724
rect 72772 24668 73612 24724
rect 73668 24668 73678 24724
rect 75170 24668 75180 24724
rect 75236 24668 75628 24724
rect 75684 24668 75694 24724
rect 76486 24668 76524 24724
rect 76580 24668 76590 24724
rect 77634 24668 77644 24724
rect 77700 24668 77710 24724
rect 0 24640 800 24668
rect 19740 24612 19796 24668
rect 16370 24556 16380 24612
rect 16436 24556 19292 24612
rect 19348 24556 19796 24612
rect 24770 24556 24780 24612
rect 24836 24556 25676 24612
rect 25732 24556 25742 24612
rect 27682 24556 27692 24612
rect 27748 24556 30380 24612
rect 30436 24556 37884 24612
rect 37940 24556 37950 24612
rect 39666 24556 39676 24612
rect 39732 24556 41692 24612
rect 41748 24556 44604 24612
rect 44660 24556 45388 24612
rect 45444 24556 45454 24612
rect 50372 24556 63420 24612
rect 63476 24556 63486 24612
rect 71362 24556 71372 24612
rect 71428 24556 71438 24612
rect 73490 24556 73500 24612
rect 73556 24556 76468 24612
rect 50372 24500 50428 24556
rect 19730 24444 19740 24500
rect 19796 24444 21868 24500
rect 21924 24444 21934 24500
rect 37762 24444 37772 24500
rect 37828 24444 50428 24500
rect 71372 24500 71428 24556
rect 76412 24500 76468 24556
rect 71372 24444 75740 24500
rect 75796 24444 75806 24500
rect 76402 24444 76412 24500
rect 76468 24444 76478 24500
rect 76850 24444 76860 24500
rect 76916 24444 76926 24500
rect 76860 24388 76916 24444
rect 8306 24332 8316 24388
rect 8372 24332 14252 24388
rect 14308 24332 17500 24388
rect 17556 24332 18060 24388
rect 18116 24332 18126 24388
rect 40114 24332 40124 24388
rect 40180 24332 42700 24388
rect 42756 24332 42766 24388
rect 47954 24332 47964 24388
rect 48020 24332 48972 24388
rect 49028 24332 49038 24388
rect 70466 24332 70476 24388
rect 70532 24332 76916 24388
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 65906 24276 65916 24332
rect 65972 24276 66020 24332
rect 66076 24276 66124 24332
rect 66180 24276 66190 24332
rect 79200 24276 80000 24304
rect 37202 24220 37212 24276
rect 37268 24220 63532 24276
rect 63588 24220 63598 24276
rect 75730 24220 75740 24276
rect 75796 24220 78540 24276
rect 78596 24220 78606 24276
rect 78988 24220 80000 24276
rect 34066 24108 34076 24164
rect 34132 24108 35756 24164
rect 35812 24108 74060 24164
rect 74116 24108 74126 24164
rect 78988 24052 79044 24220
rect 79200 24192 80000 24220
rect 12674 23996 12684 24052
rect 12740 23996 23100 24052
rect 23156 23996 23166 24052
rect 36642 23996 36652 24052
rect 36708 23996 37660 24052
rect 37716 23996 37726 24052
rect 38108 23996 43428 24052
rect 43586 23996 43596 24052
rect 43652 23996 44940 24052
rect 44996 23996 45006 24052
rect 60162 23996 60172 24052
rect 60228 23996 63252 24052
rect 63410 23996 63420 24052
rect 63476 23996 64092 24052
rect 64148 23996 70812 24052
rect 70868 23996 70878 24052
rect 71036 23996 73164 24052
rect 73220 23996 73836 24052
rect 73892 23996 73902 24052
rect 74498 23996 74508 24052
rect 74564 23996 75292 24052
rect 75348 23996 75358 24052
rect 78988 23996 79268 24052
rect 2034 23884 2044 23940
rect 2100 23884 8428 23940
rect 21186 23884 21196 23940
rect 21252 23884 23996 23940
rect 24052 23884 24062 23940
rect 34514 23884 34524 23940
rect 34580 23884 37212 23940
rect 37268 23884 37278 23940
rect 8372 23828 8428 23884
rect 38108 23828 38164 23996
rect 43372 23940 43428 23996
rect 63196 23940 63252 23996
rect 71036 23940 71092 23996
rect 8372 23772 38164 23828
rect 38556 23884 40348 23940
rect 40404 23884 40414 23940
rect 43372 23884 44828 23940
rect 44884 23884 44894 23940
rect 45154 23884 45164 23940
rect 45220 23884 45724 23940
rect 45780 23884 45790 23940
rect 47282 23884 47292 23940
rect 47348 23884 48524 23940
rect 48580 23884 62188 23940
rect 63196 23884 71092 23940
rect 71810 23884 71820 23940
rect 71876 23884 72156 23940
rect 72212 23884 72222 23940
rect 72706 23884 72716 23940
rect 72772 23884 73276 23940
rect 73332 23884 73342 23940
rect 74386 23884 74396 23940
rect 74452 23884 74508 23940
rect 74564 23884 74574 23940
rect 38556 23716 38612 23884
rect 62132 23828 62188 23884
rect 40226 23772 40236 23828
rect 40292 23772 56812 23828
rect 56868 23772 56878 23828
rect 62132 23772 70588 23828
rect 70644 23772 70654 23828
rect 71586 23772 71596 23828
rect 71652 23772 72492 23828
rect 72548 23772 72558 23828
rect 76178 23772 76188 23828
rect 76244 23772 76748 23828
rect 76804 23772 76814 23828
rect 23314 23660 23324 23716
rect 23380 23660 27580 23716
rect 27636 23660 27646 23716
rect 35410 23660 35420 23716
rect 35476 23660 37772 23716
rect 37828 23660 37838 23716
rect 37996 23660 38612 23716
rect 45042 23660 45052 23716
rect 45108 23660 45388 23716
rect 45444 23660 45454 23716
rect 46050 23660 46060 23716
rect 46116 23660 47404 23716
rect 47460 23660 47470 23716
rect 48962 23660 48972 23716
rect 49028 23660 49308 23716
rect 49364 23660 49374 23716
rect 71026 23660 71036 23716
rect 71092 23660 77644 23716
rect 77700 23660 77710 23716
rect 0 23604 800 23632
rect 37996 23604 38052 23660
rect 0 23548 1708 23604
rect 1764 23548 2492 23604
rect 2548 23548 2558 23604
rect 17378 23548 17388 23604
rect 17444 23548 17454 23604
rect 21522 23548 21532 23604
rect 21588 23548 22316 23604
rect 22372 23548 23772 23604
rect 23828 23548 34860 23604
rect 34916 23548 38052 23604
rect 46386 23548 46396 23604
rect 46452 23548 47068 23604
rect 47124 23548 47134 23604
rect 68898 23548 68908 23604
rect 68964 23548 72380 23604
rect 72436 23548 72446 23604
rect 74946 23548 74956 23604
rect 75012 23548 77196 23604
rect 77252 23548 77262 23604
rect 0 23520 800 23548
rect 17388 23492 17444 23548
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 50546 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50830 23548
rect 79212 23492 79268 23996
rect 13458 23436 13468 23492
rect 13524 23436 14924 23492
rect 14980 23436 14990 23492
rect 16146 23436 16156 23492
rect 16212 23436 19292 23492
rect 19348 23436 19358 23492
rect 20290 23436 20300 23492
rect 20356 23436 36988 23492
rect 37044 23436 37054 23492
rect 50978 23436 50988 23492
rect 51044 23436 51548 23492
rect 51604 23436 51614 23492
rect 52770 23436 52780 23492
rect 52836 23436 53788 23492
rect 53844 23436 53854 23492
rect 76178 23436 76188 23492
rect 76244 23436 78316 23492
rect 78372 23436 79268 23492
rect 20300 23380 20356 23436
rect 17602 23324 17612 23380
rect 17668 23324 18396 23380
rect 18452 23324 20356 23380
rect 23650 23324 23660 23380
rect 23716 23324 23996 23380
rect 24052 23324 24332 23380
rect 24388 23324 25228 23380
rect 25284 23324 25294 23380
rect 26114 23324 26124 23380
rect 26180 23324 26572 23380
rect 26628 23324 28028 23380
rect 28084 23324 28094 23380
rect 34850 23324 34860 23380
rect 34916 23324 36204 23380
rect 36260 23324 36270 23380
rect 43698 23324 43708 23380
rect 43764 23324 44268 23380
rect 44324 23324 44334 23380
rect 46834 23324 46844 23380
rect 46900 23324 48972 23380
rect 49028 23324 49038 23380
rect 49522 23324 49532 23380
rect 49588 23324 49756 23380
rect 49812 23324 50764 23380
rect 50820 23324 50830 23380
rect 67778 23324 67788 23380
rect 67844 23324 71708 23380
rect 71764 23324 72156 23380
rect 72212 23324 72222 23380
rect 36306 23212 36316 23268
rect 36372 23212 36764 23268
rect 36820 23212 36830 23268
rect 38658 23212 38668 23268
rect 38724 23212 39676 23268
rect 39732 23212 40460 23268
rect 40516 23212 40526 23268
rect 45826 23212 45836 23268
rect 45892 23212 45902 23268
rect 47954 23212 47964 23268
rect 48020 23212 49420 23268
rect 49476 23212 49486 23268
rect 71810 23212 71820 23268
rect 71876 23212 73948 23268
rect 74004 23212 74014 23268
rect 45836 23156 45892 23212
rect 79200 23156 80000 23184
rect 14914 23100 14924 23156
rect 14980 23100 23548 23156
rect 23604 23100 24444 23156
rect 24500 23100 24510 23156
rect 25554 23100 25564 23156
rect 25620 23100 27356 23156
rect 27412 23100 27422 23156
rect 27794 23100 27804 23156
rect 27860 23100 31724 23156
rect 31780 23100 34076 23156
rect 34132 23100 34142 23156
rect 35746 23100 35756 23156
rect 35812 23100 37324 23156
rect 37380 23100 37390 23156
rect 39788 23100 45892 23156
rect 46274 23100 46284 23156
rect 46340 23100 47292 23156
rect 47348 23100 47358 23156
rect 47516 23100 61852 23156
rect 61908 23100 61918 23156
rect 72034 23100 72044 23156
rect 72100 23100 77644 23156
rect 77700 23100 77710 23156
rect 78194 23100 78204 23156
rect 78260 23100 80000 23156
rect 39788 23044 39844 23100
rect 47516 23044 47572 23100
rect 79200 23072 80000 23100
rect 1698 22988 1708 23044
rect 1764 22988 2492 23044
rect 2548 22988 2558 23044
rect 20066 22988 20076 23044
rect 20132 22988 20636 23044
rect 20692 22988 20702 23044
rect 27906 22988 27916 23044
rect 27972 22988 29148 23044
rect 29204 22988 29214 23044
rect 34962 22988 34972 23044
rect 35028 22988 36148 23044
rect 36306 22988 36316 23044
rect 36372 22988 39844 23044
rect 40002 22988 40012 23044
rect 40068 22988 47572 23044
rect 63746 22988 63756 23044
rect 63812 22988 76860 23044
rect 76916 22988 76926 23044
rect 36092 22932 36148 22988
rect 11442 22876 11452 22932
rect 11508 22876 14364 22932
rect 14420 22876 23996 22932
rect 24052 22876 25340 22932
rect 25396 22876 25406 22932
rect 34860 22876 36036 22932
rect 36092 22876 37324 22932
rect 37380 22876 37884 22932
rect 37940 22876 37950 22932
rect 38612 22876 39228 22932
rect 39284 22876 39294 22932
rect 46806 22876 46844 22932
rect 46900 22876 46910 22932
rect 47590 22876 47628 22932
rect 47684 22876 47694 22932
rect 49410 22876 49420 22932
rect 49476 22876 70700 22932
rect 70756 22876 70766 22932
rect 71026 22876 71036 22932
rect 71092 22876 74060 22932
rect 74116 22876 74126 22932
rect 34860 22820 34916 22876
rect 35980 22820 36036 22876
rect 38612 22820 38668 22876
rect 18498 22764 18508 22820
rect 18564 22764 20076 22820
rect 20132 22764 34860 22820
rect 34916 22764 34926 22820
rect 35980 22764 38668 22820
rect 43810 22764 43820 22820
rect 43876 22764 62188 22820
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 20402 22652 20412 22708
rect 20468 22652 21420 22708
rect 21476 22652 21486 22708
rect 21634 22652 21644 22708
rect 21700 22652 24668 22708
rect 24724 22652 24734 22708
rect 25554 22652 25564 22708
rect 25620 22652 27132 22708
rect 27188 22652 28364 22708
rect 28420 22652 29036 22708
rect 29092 22652 29102 22708
rect 36978 22652 36988 22708
rect 37044 22652 37548 22708
rect 37604 22652 40348 22708
rect 40404 22652 40414 22708
rect 47954 22652 47964 22708
rect 48020 22652 48030 22708
rect 51426 22652 51436 22708
rect 51492 22652 52556 22708
rect 52612 22652 52622 22708
rect 47964 22596 48020 22652
rect 62132 22596 62188 22764
rect 65906 22708 65916 22764
rect 65972 22708 66020 22764
rect 66076 22708 66124 22764
rect 66180 22708 66190 22764
rect 2034 22540 2044 22596
rect 2100 22540 46956 22596
rect 47012 22540 47022 22596
rect 47618 22540 47628 22596
rect 47684 22540 48020 22596
rect 48850 22540 48860 22596
rect 48916 22540 51772 22596
rect 51828 22540 51838 22596
rect 62132 22540 74284 22596
rect 74340 22540 74350 22596
rect 0 22484 800 22512
rect 0 22428 1708 22484
rect 1764 22428 1774 22484
rect 12898 22428 12908 22484
rect 12964 22428 14700 22484
rect 14756 22428 15596 22484
rect 15652 22428 15662 22484
rect 28354 22428 28364 22484
rect 28420 22428 29148 22484
rect 29204 22428 29214 22484
rect 34402 22428 34412 22484
rect 34468 22428 36316 22484
rect 36372 22428 36382 22484
rect 36540 22428 68908 22484
rect 68964 22428 68974 22484
rect 69234 22428 69244 22484
rect 69300 22428 71932 22484
rect 71988 22428 71998 22484
rect 0 22400 800 22428
rect 36540 22372 36596 22428
rect 16818 22316 16828 22372
rect 16884 22316 18844 22372
rect 18900 22316 18910 22372
rect 34850 22316 34860 22372
rect 34916 22316 35196 22372
rect 35252 22316 36596 22372
rect 37426 22316 37436 22372
rect 37492 22316 38332 22372
rect 38388 22316 38398 22372
rect 42018 22316 42028 22372
rect 42084 22316 42476 22372
rect 42532 22316 42542 22372
rect 45938 22316 45948 22372
rect 46004 22316 47068 22372
rect 47124 22316 47180 22372
rect 47236 22316 47246 22372
rect 48626 22316 48636 22372
rect 48692 22316 48972 22372
rect 49028 22316 49038 22372
rect 49382 22316 49420 22372
rect 49476 22316 49486 22372
rect 69458 22316 69468 22372
rect 69524 22316 74060 22372
rect 74116 22316 74126 22372
rect 17938 22204 17948 22260
rect 18004 22204 20412 22260
rect 20468 22204 20478 22260
rect 35858 22204 35868 22260
rect 35924 22204 36876 22260
rect 36932 22204 36942 22260
rect 43698 22204 43708 22260
rect 43764 22204 43774 22260
rect 50372 22204 67116 22260
rect 67172 22204 67182 22260
rect 70242 22204 70252 22260
rect 70308 22204 72268 22260
rect 72324 22204 72334 22260
rect 16706 22092 16716 22148
rect 16772 22092 18172 22148
rect 18228 22092 19852 22148
rect 19908 22092 19918 22148
rect 33954 22092 33964 22148
rect 34020 22092 35756 22148
rect 35812 22092 37212 22148
rect 37268 22092 37278 22148
rect 43708 22036 43764 22204
rect 46386 22092 46396 22148
rect 46452 22092 48076 22148
rect 48132 22092 48142 22148
rect 50372 22036 50428 22204
rect 77858 22092 77868 22148
rect 77924 22092 78652 22148
rect 78708 22092 78718 22148
rect 79200 22036 80000 22064
rect 38098 21980 38108 22036
rect 38164 21980 43764 22036
rect 43922 21980 43932 22036
rect 43988 21980 50428 22036
rect 75730 21980 75740 22036
rect 75796 21980 76300 22036
rect 76356 21980 76366 22036
rect 78418 21980 78428 22036
rect 78484 21980 80000 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 50546 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50830 21980
rect 79200 21952 80000 21980
rect 37202 21868 37212 21924
rect 37268 21868 37548 21924
rect 37604 21868 37614 21924
rect 45164 21868 46676 21924
rect 73378 21868 73388 21924
rect 73444 21868 77644 21924
rect 77700 21868 77710 21924
rect 45164 21812 45220 21868
rect 46620 21812 46676 21868
rect 9986 21756 9996 21812
rect 10052 21756 15484 21812
rect 15540 21756 15550 21812
rect 15810 21756 15820 21812
rect 15876 21756 17500 21812
rect 17556 21756 17566 21812
rect 17714 21756 17724 21812
rect 17780 21756 18508 21812
rect 18564 21756 18574 21812
rect 24658 21756 24668 21812
rect 24724 21756 37660 21812
rect 37716 21756 37726 21812
rect 38612 21756 45220 21812
rect 45378 21756 45388 21812
rect 45444 21756 46396 21812
rect 46452 21756 46462 21812
rect 46620 21756 48188 21812
rect 48244 21756 50204 21812
rect 50260 21756 50270 21812
rect 51538 21756 51548 21812
rect 51604 21756 53788 21812
rect 53844 21756 53854 21812
rect 54898 21756 54908 21812
rect 54964 21756 55804 21812
rect 55860 21756 55870 21812
rect 63634 21756 63644 21812
rect 63700 21756 77868 21812
rect 77924 21756 77934 21812
rect 38612 21700 38668 21756
rect 2034 21644 2044 21700
rect 2100 21644 38668 21700
rect 43250 21644 43260 21700
rect 43316 21644 44268 21700
rect 44324 21644 46004 21700
rect 46162 21644 46172 21700
rect 46228 21644 47404 21700
rect 47460 21644 47470 21700
rect 47618 21644 47628 21700
rect 47684 21644 47722 21700
rect 66434 21644 66444 21700
rect 66500 21644 71708 21700
rect 71764 21644 72156 21700
rect 72212 21644 72222 21700
rect 76066 21644 76076 21700
rect 76132 21644 76300 21700
rect 76356 21644 76636 21700
rect 76692 21644 76702 21700
rect 77718 21644 77756 21700
rect 77812 21644 77822 21700
rect 45948 21588 46004 21644
rect 33394 21532 33404 21588
rect 33460 21532 34972 21588
rect 35028 21532 35038 21588
rect 35410 21532 35420 21588
rect 35476 21532 35980 21588
rect 36036 21532 36046 21588
rect 36530 21532 36540 21588
rect 36596 21532 39116 21588
rect 39172 21532 39182 21588
rect 41346 21532 41356 21588
rect 41412 21532 42476 21588
rect 42532 21532 43036 21588
rect 43092 21532 43102 21588
rect 44034 21532 44044 21588
rect 44100 21532 45612 21588
rect 45668 21532 45678 21588
rect 45948 21532 46284 21588
rect 46340 21532 46350 21588
rect 47142 21532 47180 21588
rect 47236 21532 47246 21588
rect 49494 21532 49532 21588
rect 49588 21532 49598 21588
rect 51874 21532 51884 21588
rect 51940 21532 52668 21588
rect 52724 21532 52734 21588
rect 53330 21532 53340 21588
rect 53396 21532 54348 21588
rect 54404 21532 54414 21588
rect 68002 21532 68012 21588
rect 68068 21532 74956 21588
rect 75012 21532 75022 21588
rect 75394 21532 75404 21588
rect 75460 21532 75740 21588
rect 75796 21532 75806 21588
rect 15474 21420 15484 21476
rect 15540 21420 24668 21476
rect 24724 21420 25340 21476
rect 25396 21420 25406 21476
rect 34822 21420 34860 21476
rect 34916 21420 34926 21476
rect 42802 21420 42812 21476
rect 42868 21420 62636 21476
rect 62692 21420 62702 21476
rect 73490 21420 73500 21476
rect 73556 21420 75292 21476
rect 75348 21420 75358 21476
rect 0 21364 800 21392
rect 0 21308 1708 21364
rect 1764 21308 2492 21364
rect 2548 21308 2558 21364
rect 34738 21308 34748 21364
rect 34804 21308 36316 21364
rect 36372 21308 36382 21364
rect 42130 21308 42140 21364
rect 42196 21308 42924 21364
rect 42980 21308 42990 21364
rect 45490 21308 45500 21364
rect 45556 21308 50204 21364
rect 50260 21308 50764 21364
rect 50820 21308 52780 21364
rect 52836 21308 52846 21364
rect 0 21280 800 21308
rect 39218 21196 39228 21252
rect 39284 21196 61628 21252
rect 61684 21196 61694 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 65906 21140 65916 21196
rect 65972 21140 66020 21196
rect 66076 21140 66124 21196
rect 66180 21140 66190 21196
rect 42354 21084 42364 21140
rect 42420 21084 43260 21140
rect 43316 21084 46172 21140
rect 46228 21084 46238 21140
rect 48850 21084 48860 21140
rect 48916 21084 49532 21140
rect 49588 21084 49598 21140
rect 26852 20972 48188 21028
rect 48244 20972 48254 21028
rect 48402 20972 48412 21028
rect 48468 20972 51884 21028
rect 51940 20972 51950 21028
rect 73266 20972 73276 21028
rect 73332 20972 73948 21028
rect 75394 20972 75404 21028
rect 75460 20972 76524 21028
rect 76580 20972 76590 21028
rect 26852 20916 26908 20972
rect 73892 20916 73948 20972
rect 79200 20916 80000 20944
rect 2034 20860 2044 20916
rect 2100 20860 26908 20916
rect 33954 20860 33964 20916
rect 34020 20860 35084 20916
rect 35140 20860 35150 20916
rect 36418 20860 36428 20916
rect 36484 20860 37436 20916
rect 37492 20860 38108 20916
rect 38164 20860 38892 20916
rect 38948 20860 38958 20916
rect 39452 20860 41356 20916
rect 41412 20860 41422 20916
rect 55122 20860 55132 20916
rect 55188 20860 56924 20916
rect 56980 20860 56990 20916
rect 66546 20860 66556 20916
rect 66612 20860 71260 20916
rect 71316 20860 71326 20916
rect 73892 20860 77308 20916
rect 77364 20860 77374 20916
rect 77970 20860 77980 20916
rect 78036 20860 80000 20916
rect 39452 20804 39508 20860
rect 79200 20832 80000 20860
rect 34636 20748 35196 20804
rect 35252 20748 35532 20804
rect 35588 20748 35980 20804
rect 36036 20748 36046 20804
rect 37762 20748 37772 20804
rect 37828 20748 39452 20804
rect 39508 20748 39518 20804
rect 47058 20748 47068 20804
rect 47124 20748 47628 20804
rect 47684 20748 47852 20804
rect 47908 20748 47918 20804
rect 48962 20748 48972 20804
rect 49028 20748 50316 20804
rect 50372 20748 50382 20804
rect 54002 20748 54012 20804
rect 54068 20748 56476 20804
rect 56532 20748 56542 20804
rect 77522 20748 77532 20804
rect 77588 20748 78092 20804
rect 78148 20748 78158 20804
rect 34636 20692 34692 20748
rect 34626 20636 34636 20692
rect 34692 20636 34702 20692
rect 34850 20636 34860 20692
rect 34916 20636 35644 20692
rect 35700 20636 36092 20692
rect 36148 20636 36158 20692
rect 49970 20636 49980 20692
rect 50036 20636 50652 20692
rect 50708 20636 50988 20692
rect 51044 20636 51054 20692
rect 54338 20636 54348 20692
rect 54404 20636 55020 20692
rect 55076 20636 55086 20692
rect 70466 20636 70476 20692
rect 70532 20636 72268 20692
rect 72324 20636 72334 20692
rect 74050 20636 74060 20692
rect 74116 20636 74126 20692
rect 19618 20524 19628 20580
rect 19684 20524 20524 20580
rect 20580 20524 20590 20580
rect 23426 20524 23436 20580
rect 23492 20524 24108 20580
rect 24164 20524 25340 20580
rect 25396 20524 25406 20580
rect 25554 20524 25564 20580
rect 25620 20524 29484 20580
rect 29540 20524 29550 20580
rect 32918 20524 32956 20580
rect 33012 20524 33022 20580
rect 35746 20524 35756 20580
rect 35812 20524 37100 20580
rect 37156 20524 37166 20580
rect 38882 20524 38892 20580
rect 38948 20524 39900 20580
rect 39956 20524 40684 20580
rect 40740 20524 40750 20580
rect 48178 20524 48188 20580
rect 48244 20524 52780 20580
rect 52836 20524 52846 20580
rect 74060 20468 74116 20636
rect 22418 20412 22428 20468
rect 22484 20412 22988 20468
rect 23044 20412 24780 20468
rect 24836 20412 38444 20468
rect 38500 20412 38510 20468
rect 38658 20412 38668 20468
rect 38724 20412 40684 20468
rect 40740 20412 43148 20468
rect 43204 20412 43214 20468
rect 57250 20412 57260 20468
rect 57316 20412 74116 20468
rect 76374 20412 76412 20468
rect 76468 20412 76478 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 50546 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50830 20412
rect 2034 20300 2044 20356
rect 2100 20300 8428 20356
rect 0 20244 800 20272
rect 8372 20244 8428 20300
rect 26852 20300 31836 20356
rect 31892 20300 31902 20356
rect 34626 20300 34636 20356
rect 34692 20300 36540 20356
rect 36596 20300 37436 20356
rect 37492 20300 38780 20356
rect 38836 20300 39340 20356
rect 39396 20300 39406 20356
rect 48934 20300 48972 20356
rect 49028 20300 49038 20356
rect 53554 20300 53564 20356
rect 53620 20300 55468 20356
rect 55524 20300 55534 20356
rect 26852 20244 26908 20300
rect 0 20188 1708 20244
rect 1764 20188 2492 20244
rect 2548 20188 2558 20244
rect 8372 20188 26908 20244
rect 29698 20188 29708 20244
rect 29764 20188 32284 20244
rect 32340 20188 44156 20244
rect 44212 20188 44222 20244
rect 45042 20188 45052 20244
rect 45108 20188 46396 20244
rect 46452 20188 47124 20244
rect 47394 20188 47404 20244
rect 47460 20188 63532 20244
rect 63588 20188 63598 20244
rect 74722 20188 74732 20244
rect 74788 20188 76972 20244
rect 77028 20188 77038 20244
rect 0 20160 800 20188
rect 47068 20132 47124 20188
rect 17042 20076 17052 20132
rect 17108 20076 18620 20132
rect 18676 20076 18686 20132
rect 19058 20076 19068 20132
rect 19124 20076 20300 20132
rect 20356 20076 20366 20132
rect 20738 20076 20748 20132
rect 20804 20076 21756 20132
rect 21812 20076 21822 20132
rect 26674 20076 26684 20132
rect 26740 20076 29260 20132
rect 29316 20076 30156 20132
rect 30212 20076 30222 20132
rect 31266 20076 31276 20132
rect 31332 20076 33516 20132
rect 33572 20076 35700 20132
rect 40562 20076 40572 20132
rect 40628 20076 40908 20132
rect 40964 20076 40974 20132
rect 43474 20076 43484 20132
rect 43540 20076 44492 20132
rect 44548 20076 44558 20132
rect 47068 20076 47460 20132
rect 48514 20076 48524 20132
rect 48580 20076 49420 20132
rect 49476 20076 49486 20132
rect 51090 20076 51100 20132
rect 51156 20076 51324 20132
rect 51380 20076 53228 20132
rect 53284 20076 53452 20132
rect 53508 20076 53518 20132
rect 54226 20076 54236 20132
rect 54292 20076 57596 20132
rect 57652 20076 57662 20132
rect 72706 20076 72716 20132
rect 72772 20076 73948 20132
rect 75058 20076 75068 20132
rect 75124 20076 77644 20132
rect 77700 20076 77710 20132
rect 18620 19908 18676 20076
rect 18946 19964 18956 20020
rect 19012 19964 19516 20020
rect 19572 19964 19582 20020
rect 24210 19964 24220 20020
rect 24276 19964 25228 20020
rect 25284 19964 25294 20020
rect 32946 19964 32956 20020
rect 33012 19964 33740 20020
rect 33796 19964 33806 20020
rect 18620 19852 19628 19908
rect 19684 19852 19694 19908
rect 20962 19852 20972 19908
rect 21028 19852 35588 19908
rect 19058 19740 19068 19796
rect 19124 19740 22092 19796
rect 22148 19740 22158 19796
rect 26852 19740 34188 19796
rect 34244 19740 34254 19796
rect 19282 19628 19292 19684
rect 19348 19628 24108 19684
rect 24164 19628 24174 19684
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 26852 19572 26908 19740
rect 34066 19628 34076 19684
rect 34132 19628 34860 19684
rect 34916 19628 34926 19684
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 35532 19572 35588 19852
rect 35644 19796 35700 20076
rect 37874 19964 37884 20020
rect 37940 19964 39676 20020
rect 39732 19964 39742 20020
rect 40226 19964 40236 20020
rect 40292 19964 41132 20020
rect 41188 19964 41198 20020
rect 47404 19908 47460 20076
rect 73892 20020 73948 20076
rect 48066 19964 48076 20020
rect 48132 19964 48748 20020
rect 48804 19964 48814 20020
rect 49270 19964 49308 20020
rect 49364 19964 49374 20020
rect 51762 19964 51772 20020
rect 51828 19964 52108 20020
rect 52164 19964 52444 20020
rect 52500 19964 52510 20020
rect 52882 19964 52892 20020
rect 52948 19964 56700 20020
rect 56756 19964 56766 20020
rect 73892 19964 75740 20020
rect 75796 19964 75806 20020
rect 76374 19964 76412 20020
rect 76468 19964 76478 20020
rect 76850 19964 76860 20020
rect 76916 19964 77420 20020
rect 77476 19964 77486 20020
rect 47394 19852 47404 19908
rect 47460 19852 48524 19908
rect 48580 19852 48590 19908
rect 50866 19852 50876 19908
rect 50932 19852 56028 19908
rect 56084 19852 56094 19908
rect 75394 19852 75404 19908
rect 75460 19852 75964 19908
rect 76020 19852 76030 19908
rect 77606 19852 77644 19908
rect 77700 19852 77710 19908
rect 79200 19796 80000 19824
rect 35644 19740 47068 19796
rect 47124 19740 47134 19796
rect 52098 19740 52108 19796
rect 52164 19740 52444 19796
rect 52500 19740 52510 19796
rect 74834 19740 74844 19796
rect 74900 19740 80000 19796
rect 79200 19712 80000 19740
rect 37090 19628 37100 19684
rect 37156 19628 37996 19684
rect 38052 19628 38062 19684
rect 40562 19628 40572 19684
rect 40628 19628 41132 19684
rect 41188 19628 57260 19684
rect 57316 19628 57326 19684
rect 65906 19572 65916 19628
rect 65972 19572 66020 19628
rect 66076 19572 66124 19628
rect 66180 19572 66190 19628
rect 15092 19516 26908 19572
rect 35532 19516 39228 19572
rect 39284 19516 39294 19572
rect 45938 19516 45948 19572
rect 46004 19516 50204 19572
rect 50260 19516 50270 19572
rect 55346 19516 55356 19572
rect 55412 19516 56588 19572
rect 56644 19516 56654 19572
rect 15092 19348 15148 19516
rect 30146 19404 30156 19460
rect 30212 19404 34020 19460
rect 35634 19404 35644 19460
rect 35700 19404 36652 19460
rect 36708 19404 36718 19460
rect 37762 19404 37772 19460
rect 37828 19404 40012 19460
rect 40068 19404 40078 19460
rect 40786 19404 40796 19460
rect 40852 19404 41244 19460
rect 41300 19404 41310 19460
rect 41570 19404 41580 19460
rect 41636 19404 70476 19460
rect 70532 19404 70542 19460
rect 33964 19348 34020 19404
rect 7522 19292 7532 19348
rect 7588 19292 15148 19348
rect 25900 19292 26572 19348
rect 26628 19292 26638 19348
rect 33964 19292 37100 19348
rect 37156 19292 37166 19348
rect 37874 19292 37884 19348
rect 37940 19292 38332 19348
rect 38388 19292 38668 19348
rect 39218 19292 39228 19348
rect 39284 19292 43036 19348
rect 43092 19292 43102 19348
rect 46722 19292 46732 19348
rect 46788 19292 48524 19348
rect 48580 19292 48590 19348
rect 48748 19292 73836 19348
rect 73892 19292 73902 19348
rect 76066 19292 76076 19348
rect 76132 19292 76524 19348
rect 76580 19292 76590 19348
rect 25900 19236 25956 19292
rect 38612 19236 38668 19292
rect 21746 19180 21756 19236
rect 21812 19180 25564 19236
rect 25620 19180 25956 19236
rect 26114 19180 26124 19236
rect 26180 19180 26908 19236
rect 26964 19180 26974 19236
rect 27570 19180 27580 19236
rect 27636 19180 29932 19236
rect 29988 19180 29998 19236
rect 30482 19180 30492 19236
rect 30548 19180 31276 19236
rect 31332 19180 31342 19236
rect 34962 19180 34972 19236
rect 35028 19180 35644 19236
rect 35700 19180 35710 19236
rect 36418 19180 36428 19236
rect 36484 19180 37996 19236
rect 38052 19180 38062 19236
rect 38612 19180 39116 19236
rect 39172 19180 39182 19236
rect 39554 19180 39564 19236
rect 39620 19180 41020 19236
rect 41076 19180 41086 19236
rect 46274 19180 46284 19236
rect 46340 19180 46620 19236
rect 46676 19180 46956 19236
rect 47012 19180 47022 19236
rect 0 19124 800 19152
rect 48748 19124 48804 19292
rect 48934 19180 48972 19236
rect 49028 19180 49038 19236
rect 49298 19180 49308 19236
rect 49364 19180 50428 19236
rect 50484 19180 50494 19236
rect 51762 19180 51772 19236
rect 51828 19180 51996 19236
rect 52052 19180 52668 19236
rect 52724 19180 52734 19236
rect 78194 19180 78204 19236
rect 78260 19180 78428 19236
rect 78484 19180 78494 19236
rect 0 19068 1708 19124
rect 1764 19068 2492 19124
rect 2548 19068 2558 19124
rect 17938 19068 17948 19124
rect 18004 19068 18956 19124
rect 19012 19068 19022 19124
rect 19618 19068 19628 19124
rect 19684 19068 21532 19124
rect 21588 19068 22764 19124
rect 22820 19068 22830 19124
rect 23314 19068 23324 19124
rect 23380 19068 23996 19124
rect 24052 19068 24062 19124
rect 24434 19068 24444 19124
rect 24500 19068 25452 19124
rect 25508 19068 26236 19124
rect 26292 19068 26302 19124
rect 29698 19068 29708 19124
rect 29764 19068 30604 19124
rect 30660 19068 33404 19124
rect 33460 19068 33470 19124
rect 34290 19068 34300 19124
rect 34356 19068 35308 19124
rect 35364 19068 35374 19124
rect 35858 19068 35868 19124
rect 35924 19068 37100 19124
rect 37156 19068 37660 19124
rect 37716 19068 37726 19124
rect 38658 19068 38668 19124
rect 38724 19068 39340 19124
rect 39396 19068 39406 19124
rect 39778 19068 39788 19124
rect 39844 19068 40460 19124
rect 40516 19068 40526 19124
rect 41346 19068 41356 19124
rect 41412 19068 42140 19124
rect 42196 19068 48804 19124
rect 75954 19068 75964 19124
rect 76020 19068 76524 19124
rect 76580 19068 76590 19124
rect 77522 19068 77532 19124
rect 77588 19068 77980 19124
rect 78036 19068 78046 19124
rect 0 19040 800 19068
rect 19506 18956 19516 19012
rect 19572 18956 23548 19012
rect 23604 18956 23614 19012
rect 24098 18956 24108 19012
rect 24164 18956 24174 19012
rect 26562 18956 26572 19012
rect 26628 18956 29484 19012
rect 29540 18956 29550 19012
rect 30706 18956 30716 19012
rect 30772 18956 30782 19012
rect 32274 18956 32284 19012
rect 32340 18956 33852 19012
rect 33908 18956 33918 19012
rect 39106 18956 39116 19012
rect 39172 18956 41804 19012
rect 41860 18956 41870 19012
rect 46610 18956 46620 19012
rect 46676 18956 64652 19012
rect 64708 18956 64718 19012
rect 67106 18956 67116 19012
rect 67172 18956 75404 19012
rect 75460 18956 75470 19012
rect 76738 18956 76748 19012
rect 76804 18956 77868 19012
rect 77924 18956 77934 19012
rect 24108 18900 24164 18956
rect 30716 18900 30772 18956
rect 24108 18844 30772 18900
rect 31826 18844 31836 18900
rect 31892 18844 36316 18900
rect 36372 18844 36382 18900
rect 40002 18844 40012 18900
rect 40068 18844 40460 18900
rect 40516 18844 41580 18900
rect 41636 18844 41646 18900
rect 47170 18844 47180 18900
rect 47236 18844 48524 18900
rect 48580 18844 48590 18900
rect 56354 18844 56364 18900
rect 56420 18844 68572 18900
rect 68628 18844 68638 18900
rect 74274 18844 74284 18900
rect 74340 18844 76636 18900
rect 76692 18844 76702 18900
rect 77186 18844 77196 18900
rect 77252 18844 78204 18900
rect 78260 18844 78270 18900
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 50546 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50830 18844
rect 21522 18732 21532 18788
rect 21588 18732 23660 18788
rect 23716 18732 24332 18788
rect 24388 18732 24398 18788
rect 27346 18732 27356 18788
rect 27412 18732 27916 18788
rect 27972 18732 28476 18788
rect 28532 18732 33012 18788
rect 33394 18732 33404 18788
rect 33460 18732 45052 18788
rect 45108 18732 45118 18788
rect 48290 18732 48300 18788
rect 48356 18732 48972 18788
rect 49028 18732 49038 18788
rect 32956 18676 33012 18732
rect 79200 18676 80000 18704
rect 6290 18620 6300 18676
rect 6356 18620 32732 18676
rect 32788 18620 32798 18676
rect 32956 18620 46620 18676
rect 46676 18620 46686 18676
rect 76738 18620 76748 18676
rect 76804 18620 77532 18676
rect 77588 18620 77598 18676
rect 78194 18620 78204 18676
rect 78260 18620 80000 18676
rect 79200 18592 80000 18620
rect 25564 18508 26012 18564
rect 26068 18508 26078 18564
rect 39106 18508 39116 18564
rect 39172 18508 39900 18564
rect 39956 18508 39966 18564
rect 46274 18508 46284 18564
rect 46340 18508 49420 18564
rect 49476 18508 50988 18564
rect 51044 18508 51054 18564
rect 53218 18508 53228 18564
rect 53284 18508 54124 18564
rect 54180 18508 54190 18564
rect 55122 18508 55132 18564
rect 55188 18508 56140 18564
rect 56196 18508 57092 18564
rect 76514 18508 76524 18564
rect 76580 18508 77420 18564
rect 77476 18508 77486 18564
rect 25564 18452 25620 18508
rect 57036 18452 57092 18508
rect 22194 18396 22204 18452
rect 22260 18396 25340 18452
rect 25396 18396 25620 18452
rect 25778 18396 25788 18452
rect 25844 18396 26348 18452
rect 26404 18396 26908 18452
rect 28130 18396 28140 18452
rect 28196 18396 31948 18452
rect 32004 18396 33628 18452
rect 33684 18396 33694 18452
rect 38546 18396 38556 18452
rect 38612 18396 39340 18452
rect 39396 18396 39406 18452
rect 39666 18396 39676 18452
rect 39732 18396 41244 18452
rect 41300 18396 41310 18452
rect 41906 18396 41916 18452
rect 41972 18396 42588 18452
rect 42644 18396 42654 18452
rect 45602 18396 45612 18452
rect 45668 18396 50428 18452
rect 54898 18396 54908 18452
rect 54964 18396 56700 18452
rect 56756 18396 56766 18452
rect 57036 18396 58828 18452
rect 58884 18396 58894 18452
rect 77746 18396 77756 18452
rect 77812 18396 77980 18452
rect 78036 18396 78046 18452
rect 26852 18340 26908 18396
rect 2034 18284 2044 18340
rect 2100 18284 8428 18340
rect 24658 18284 24668 18340
rect 24724 18284 25900 18340
rect 25956 18284 25966 18340
rect 26852 18284 28700 18340
rect 28756 18284 28766 18340
rect 35186 18284 35196 18340
rect 35252 18284 38220 18340
rect 38276 18284 40572 18340
rect 40628 18284 40638 18340
rect 43138 18284 43148 18340
rect 43204 18284 45500 18340
rect 45556 18284 45566 18340
rect 48738 18284 48748 18340
rect 48804 18284 49084 18340
rect 49140 18284 49150 18340
rect 8372 18228 8428 18284
rect 50372 18228 50428 18396
rect 53330 18284 53340 18340
rect 53396 18284 57148 18340
rect 57204 18284 57214 18340
rect 8372 18172 36540 18228
rect 36596 18172 36606 18228
rect 39442 18172 39452 18228
rect 39508 18172 41244 18228
rect 41300 18172 41310 18228
rect 41906 18172 41916 18228
rect 41972 18172 44716 18228
rect 44772 18172 44782 18228
rect 50372 18172 52556 18228
rect 52612 18172 55916 18228
rect 55972 18172 55982 18228
rect 77746 18172 77756 18228
rect 77812 18172 77822 18228
rect 77756 18116 77812 18172
rect 39106 18060 39116 18116
rect 39172 18060 43372 18116
rect 43428 18060 43438 18116
rect 74610 18060 74620 18116
rect 74676 18060 77812 18116
rect 0 18004 800 18032
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 65906 18004 65916 18060
rect 65972 18004 66020 18060
rect 66076 18004 66124 18060
rect 66180 18004 66190 18060
rect 0 17948 1708 18004
rect 1764 17948 2492 18004
rect 2548 17948 2558 18004
rect 23986 17948 23996 18004
rect 24052 17948 25116 18004
rect 25172 17948 32788 18004
rect 40114 17948 40124 18004
rect 40180 17948 43932 18004
rect 43988 17948 43998 18004
rect 47730 17948 47740 18004
rect 47796 17948 64540 18004
rect 64596 17948 64606 18004
rect 0 17920 800 17948
rect 32732 17892 32788 17948
rect 2034 17836 2044 17892
rect 2100 17836 26908 17892
rect 32732 17836 41076 17892
rect 44034 17836 44044 17892
rect 44100 17836 45388 17892
rect 45444 17836 45454 17892
rect 45612 17836 70588 17892
rect 70644 17836 70654 17892
rect 26852 17780 26908 17836
rect 16930 17724 16940 17780
rect 16996 17724 17724 17780
rect 17780 17724 18732 17780
rect 18788 17724 18798 17780
rect 21634 17724 21644 17780
rect 21700 17724 22316 17780
rect 22372 17724 25004 17780
rect 25060 17724 25070 17780
rect 26852 17724 35420 17780
rect 35476 17724 35486 17780
rect 35634 17724 35644 17780
rect 35700 17724 36092 17780
rect 36148 17724 37212 17780
rect 37268 17724 37278 17780
rect 38612 17724 39116 17780
rect 39172 17724 39182 17780
rect 38612 17668 38668 17724
rect 41020 17668 41076 17836
rect 45612 17780 45668 17836
rect 43026 17724 43036 17780
rect 43092 17724 43820 17780
rect 43876 17724 43886 17780
rect 44930 17724 44940 17780
rect 44996 17724 45668 17780
rect 46722 17724 46732 17780
rect 46788 17724 61740 17780
rect 61796 17724 61806 17780
rect 32946 17612 32956 17668
rect 33012 17612 38668 17668
rect 39302 17612 39340 17668
rect 39396 17612 39406 17668
rect 39974 17612 40012 17668
rect 40068 17612 40348 17668
rect 40404 17612 40414 17668
rect 40646 17612 40684 17668
rect 40740 17612 40750 17668
rect 41010 17612 41020 17668
rect 41076 17612 43148 17668
rect 43204 17612 43214 17668
rect 45042 17612 45052 17668
rect 45108 17612 46956 17668
rect 47012 17612 47022 17668
rect 53442 17612 53452 17668
rect 53508 17612 54012 17668
rect 54068 17612 54078 17668
rect 55234 17612 55244 17668
rect 55300 17612 56812 17668
rect 56868 17612 56878 17668
rect 57138 17612 57148 17668
rect 57204 17612 58716 17668
rect 58772 17612 58782 17668
rect 77634 17612 77644 17668
rect 77700 17612 78204 17668
rect 78260 17612 78270 17668
rect 79200 17556 80000 17584
rect 28690 17500 28700 17556
rect 28756 17500 29596 17556
rect 29652 17500 29662 17556
rect 33842 17500 33852 17556
rect 33908 17500 35308 17556
rect 35364 17500 35374 17556
rect 76962 17500 76972 17556
rect 77028 17500 77532 17556
rect 77588 17500 80000 17556
rect 79200 17472 80000 17500
rect 1698 17388 1708 17444
rect 1764 17388 2492 17444
rect 2548 17388 2558 17444
rect 17826 17388 17836 17444
rect 17892 17388 19404 17444
rect 19460 17388 19470 17444
rect 19730 17388 19740 17444
rect 19796 17388 20412 17444
rect 20468 17388 20478 17444
rect 26852 17388 28476 17444
rect 28532 17388 39396 17444
rect 39554 17388 39564 17444
rect 39620 17388 41356 17444
rect 41412 17388 41422 17444
rect 43596 17388 49308 17444
rect 49364 17388 50876 17444
rect 50932 17388 50942 17444
rect 51762 17388 51772 17444
rect 51828 17388 52780 17444
rect 52836 17388 52846 17444
rect 75282 17388 75292 17444
rect 75348 17388 78204 17444
rect 78260 17388 78270 17444
rect 26338 17276 26348 17332
rect 26404 17276 26796 17332
rect 26852 17276 26908 17388
rect 32946 17276 32956 17332
rect 33012 17276 33022 17332
rect 35410 17276 35420 17332
rect 35476 17276 37100 17332
rect 37156 17276 37166 17332
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 32956 17220 33012 17276
rect 39340 17220 39396 17388
rect 43596 17220 43652 17388
rect 53442 17276 53452 17332
rect 53508 17276 55132 17332
rect 55188 17276 55198 17332
rect 77298 17276 77308 17332
rect 77364 17276 77588 17332
rect 77858 17276 77868 17332
rect 77924 17276 78652 17332
rect 78708 17276 78718 17332
rect 50546 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50830 17276
rect 77532 17220 77588 17276
rect 20402 17164 20412 17220
rect 20468 17164 21644 17220
rect 21700 17164 33012 17220
rect 37202 17164 37212 17220
rect 37268 17164 38892 17220
rect 38948 17164 38958 17220
rect 39340 17164 43652 17220
rect 43810 17164 43820 17220
rect 43876 17164 44940 17220
rect 44996 17164 45006 17220
rect 77522 17164 77532 17220
rect 77588 17164 77598 17220
rect 29362 17052 29372 17108
rect 29428 17052 32508 17108
rect 32564 17052 34524 17108
rect 34580 17052 34590 17108
rect 34748 17052 50988 17108
rect 51044 17052 51054 17108
rect 34748 16996 34804 17052
rect 30146 16940 30156 16996
rect 30212 16940 32060 16996
rect 32116 16940 34804 16996
rect 37090 16940 37100 16996
rect 37156 16940 37268 16996
rect 38882 16940 38892 16996
rect 38948 16940 39900 16996
rect 39956 16940 39966 16996
rect 42690 16940 42700 16996
rect 42756 16940 45612 16996
rect 45668 16940 45678 16996
rect 45836 16940 72156 16996
rect 72212 16940 72222 16996
rect 75618 16940 75628 16996
rect 75684 16940 77308 16996
rect 77364 16940 77374 16996
rect 0 16884 800 16912
rect 37212 16884 37268 16940
rect 45836 16884 45892 16940
rect 0 16828 1708 16884
rect 1764 16828 1774 16884
rect 25890 16828 25900 16884
rect 25956 16828 27132 16884
rect 27188 16828 27198 16884
rect 33506 16828 33516 16884
rect 33572 16828 34580 16884
rect 34738 16828 34748 16884
rect 34804 16828 36988 16884
rect 37044 16828 37054 16884
rect 37212 16828 37772 16884
rect 37828 16828 37838 16884
rect 38658 16828 38668 16884
rect 38724 16828 40012 16884
rect 40068 16828 40124 16884
rect 40180 16828 40190 16884
rect 41458 16828 41468 16884
rect 41524 16828 41916 16884
rect 41972 16828 45892 16884
rect 47030 16828 47068 16884
rect 47124 16828 47134 16884
rect 48066 16828 48076 16884
rect 48132 16828 48748 16884
rect 48804 16828 48814 16884
rect 51874 16828 51884 16884
rect 51940 16828 52668 16884
rect 52724 16828 52734 16884
rect 77186 16828 77196 16884
rect 77252 16828 78092 16884
rect 78148 16828 78372 16884
rect 0 16800 800 16828
rect 34524 16772 34580 16828
rect 34524 16716 34636 16772
rect 34692 16716 34702 16772
rect 36530 16716 36540 16772
rect 36596 16716 37436 16772
rect 37492 16716 37502 16772
rect 39750 16716 39788 16772
rect 39844 16716 39854 16772
rect 47170 16716 47180 16772
rect 47236 16716 47740 16772
rect 47796 16716 47806 16772
rect 77410 16716 77420 16772
rect 77476 16716 77756 16772
rect 77812 16716 77822 16772
rect 38098 16604 38108 16660
rect 38164 16604 43372 16660
rect 43428 16604 43438 16660
rect 43670 16604 43708 16660
rect 43764 16604 43774 16660
rect 42354 16492 42364 16548
rect 42420 16492 45500 16548
rect 45556 16492 46060 16548
rect 46116 16492 46126 16548
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 65906 16436 65916 16492
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 66180 16436 66190 16492
rect 78316 16436 78372 16828
rect 79200 16436 80000 16464
rect 42578 16380 42588 16436
rect 42644 16380 54572 16436
rect 54628 16380 54638 16436
rect 78316 16380 80000 16436
rect 79200 16352 80000 16380
rect 2034 16268 2044 16324
rect 2100 16268 36092 16324
rect 36148 16268 36988 16324
rect 37044 16268 37054 16324
rect 37986 16268 37996 16324
rect 38052 16268 39340 16324
rect 39396 16268 39406 16324
rect 43586 16268 43596 16324
rect 43652 16268 45388 16324
rect 45444 16268 45454 16324
rect 45826 16268 45836 16324
rect 45892 16268 71036 16324
rect 71092 16268 71102 16324
rect 8372 16156 33516 16212
rect 33572 16156 33582 16212
rect 37884 16156 39676 16212
rect 39732 16156 39742 16212
rect 41458 16156 41468 16212
rect 41524 16156 42924 16212
rect 42980 16156 42990 16212
rect 43474 16156 43484 16212
rect 43540 16156 44268 16212
rect 44324 16156 70252 16212
rect 70308 16156 70318 16212
rect 8372 16100 8428 16156
rect 2146 16044 2156 16100
rect 2212 16044 8428 16100
rect 31490 16044 31500 16100
rect 31556 16044 32172 16100
rect 32228 16044 32238 16100
rect 37884 15988 37940 16156
rect 41234 16044 41244 16100
rect 41300 16044 43036 16100
rect 43092 16044 43708 16100
rect 43764 16044 43774 16100
rect 51426 16044 51436 16100
rect 51492 16044 52668 16100
rect 52724 16044 52734 16100
rect 27346 15932 27356 15988
rect 27412 15932 28364 15988
rect 28420 15932 31444 15988
rect 34626 15932 34636 15988
rect 34692 15932 37884 15988
rect 37940 15932 37950 15988
rect 38612 15932 46284 15988
rect 46340 15932 46350 15988
rect 31388 15876 31444 15932
rect 38612 15876 38668 15932
rect 23762 15820 23772 15876
rect 23828 15820 26908 15876
rect 26964 15820 27244 15876
rect 27300 15820 27310 15876
rect 28130 15820 28140 15876
rect 28196 15820 29596 15876
rect 29652 15820 29662 15876
rect 31388 15820 38668 15876
rect 40114 15820 40124 15876
rect 40180 15820 42252 15876
rect 42308 15820 42588 15876
rect 42644 15820 42654 15876
rect 44034 15820 44044 15876
rect 44100 15820 45836 15876
rect 45892 15820 45902 15876
rect 46386 15820 46396 15876
rect 46452 15820 48076 15876
rect 48132 15820 51436 15876
rect 51492 15820 54684 15876
rect 54740 15820 54750 15876
rect 77634 15820 77644 15876
rect 77700 15820 78204 15876
rect 78260 15820 78270 15876
rect 0 15764 800 15792
rect 0 15708 1708 15764
rect 1764 15708 2492 15764
rect 2548 15708 2558 15764
rect 34962 15708 34972 15764
rect 35028 15708 35644 15764
rect 35700 15708 35710 15764
rect 45714 15708 45724 15764
rect 45780 15708 47852 15764
rect 47908 15708 50316 15764
rect 50372 15708 50382 15764
rect 0 15680 800 15708
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 50546 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50830 15708
rect 20178 15596 20188 15652
rect 20244 15596 34076 15652
rect 34132 15596 34142 15652
rect 42690 15596 42700 15652
rect 42756 15596 43260 15652
rect 43316 15596 43326 15652
rect 46386 15596 46396 15652
rect 46452 15596 47740 15652
rect 47796 15596 48188 15652
rect 48244 15596 50428 15652
rect 8372 15484 23548 15540
rect 8372 15428 8428 15484
rect 2034 15372 2044 15428
rect 2100 15372 8428 15428
rect 23492 15428 23548 15484
rect 26852 15484 38892 15540
rect 38948 15484 39452 15540
rect 39508 15484 39518 15540
rect 26852 15428 26908 15484
rect 50372 15428 50428 15596
rect 23492 15372 26908 15428
rect 33394 15372 33404 15428
rect 33460 15372 35420 15428
rect 35476 15372 47292 15428
rect 47348 15372 47358 15428
rect 50372 15372 50652 15428
rect 50708 15372 50718 15428
rect 79200 15316 80000 15344
rect 9986 15260 9996 15316
rect 10052 15260 20188 15316
rect 20244 15260 20254 15316
rect 46834 15260 46844 15316
rect 46900 15260 48972 15316
rect 49028 15260 49038 15316
rect 51986 15260 51996 15316
rect 52052 15260 54236 15316
rect 54292 15260 54302 15316
rect 78194 15260 78204 15316
rect 78260 15260 80000 15316
rect 79200 15232 80000 15260
rect 5842 15148 5852 15204
rect 5908 15148 32508 15204
rect 32564 15148 33852 15204
rect 33908 15148 33918 15204
rect 39218 15148 39228 15204
rect 39284 15148 41692 15204
rect 41748 15148 42028 15204
rect 42084 15148 42094 15204
rect 51650 15148 51660 15204
rect 51716 15148 53676 15204
rect 53732 15148 53742 15204
rect 55234 15148 55244 15204
rect 55300 15148 69692 15204
rect 69748 15148 69758 15204
rect 34850 15036 34860 15092
rect 34916 15036 48300 15092
rect 48356 15036 50876 15092
rect 50932 15036 50942 15092
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 65906 14868 65916 14924
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 66180 14868 66190 14924
rect 38546 14812 38556 14868
rect 38612 14812 38622 14868
rect 49410 14812 49420 14868
rect 49476 14812 51324 14868
rect 51380 14812 51390 14868
rect 0 14644 800 14672
rect 38556 14644 38612 14812
rect 42690 14700 42700 14756
rect 42756 14700 45164 14756
rect 45220 14700 54460 14756
rect 54516 14700 54526 14756
rect 74582 14700 74620 14756
rect 74676 14700 74686 14756
rect 0 14588 1708 14644
rect 1764 14588 2492 14644
rect 2548 14588 2558 14644
rect 8306 14588 8316 14644
rect 8372 14588 38612 14644
rect 47058 14588 47068 14644
rect 47124 14588 50092 14644
rect 50148 14588 50158 14644
rect 50306 14588 50316 14644
rect 50372 14588 55468 14644
rect 55524 14588 55534 14644
rect 0 14560 800 14588
rect 3332 14476 31948 14532
rect 32004 14476 32014 14532
rect 34066 14476 34076 14532
rect 34132 14476 35420 14532
rect 35476 14476 35486 14532
rect 35858 14476 35868 14532
rect 35924 14476 37436 14532
rect 37492 14476 48748 14532
rect 48804 14476 48814 14532
rect 50418 14476 50428 14532
rect 50484 14476 51324 14532
rect 51380 14476 52668 14532
rect 52724 14476 52734 14532
rect 3332 14420 3388 14476
rect 1586 14364 1596 14420
rect 1652 14364 3388 14420
rect 26786 14364 26796 14420
rect 26852 14364 28252 14420
rect 28308 14364 29148 14420
rect 29204 14364 29214 14420
rect 32050 14364 32060 14420
rect 32116 14364 33404 14420
rect 33460 14364 33470 14420
rect 37202 14364 37212 14420
rect 37268 14364 42924 14420
rect 42980 14364 42990 14420
rect 52770 14364 52780 14420
rect 52836 14364 71372 14420
rect 71428 14364 71438 14420
rect 77298 14364 77308 14420
rect 77364 14364 77868 14420
rect 77924 14364 77934 14420
rect 26562 14252 26572 14308
rect 26628 14252 27244 14308
rect 27300 14252 27310 14308
rect 28578 14252 28588 14308
rect 28644 14252 29484 14308
rect 29540 14252 34412 14308
rect 34468 14252 34478 14308
rect 38434 14252 38444 14308
rect 38500 14252 45500 14308
rect 45556 14252 45566 14308
rect 79200 14196 80000 14224
rect 29362 14140 29372 14196
rect 29428 14140 30156 14196
rect 30212 14140 30828 14196
rect 30884 14140 49420 14196
rect 49476 14140 49486 14196
rect 77634 14140 77644 14196
rect 77700 14140 78204 14196
rect 78260 14140 80000 14196
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 50546 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50830 14140
rect 79200 14112 80000 14140
rect 26852 14028 34636 14084
rect 34692 14028 34702 14084
rect 39330 14028 39340 14084
rect 39396 14028 40292 14084
rect 41458 14028 41468 14084
rect 41524 14028 50316 14084
rect 50372 14028 50382 14084
rect 2034 13916 2044 13972
rect 2100 13916 3388 13972
rect 3332 13860 3388 13916
rect 26852 13860 26908 14028
rect 40236 13972 40292 14028
rect 33394 13916 33404 13972
rect 33460 13916 34188 13972
rect 34244 13916 34860 13972
rect 34916 13916 34926 13972
rect 37650 13916 37660 13972
rect 37716 13916 39676 13972
rect 39732 13916 39742 13972
rect 40226 13916 40236 13972
rect 40292 13916 42476 13972
rect 42532 13916 42542 13972
rect 76290 13916 76300 13972
rect 76356 13916 77084 13972
rect 77140 13916 77150 13972
rect 3332 13804 26908 13860
rect 33618 13804 33628 13860
rect 33684 13804 34748 13860
rect 34804 13804 36092 13860
rect 36148 13804 36158 13860
rect 40002 13804 40012 13860
rect 40068 13804 41580 13860
rect 41636 13804 54796 13860
rect 54852 13804 54862 13860
rect 21410 13692 21420 13748
rect 21476 13692 23436 13748
rect 23492 13692 23502 13748
rect 26562 13692 26572 13748
rect 26628 13692 27356 13748
rect 27412 13692 27804 13748
rect 27860 13692 27870 13748
rect 34402 13692 34412 13748
rect 34468 13692 37884 13748
rect 37940 13692 39004 13748
rect 39060 13692 39070 13748
rect 42690 13692 42700 13748
rect 42756 13692 45388 13748
rect 45444 13692 51324 13748
rect 51380 13692 51390 13748
rect 16594 13580 16604 13636
rect 16660 13580 18620 13636
rect 18676 13580 19628 13636
rect 19684 13580 19694 13636
rect 0 13524 800 13552
rect 0 13468 1708 13524
rect 1764 13468 2492 13524
rect 2548 13468 2558 13524
rect 26674 13468 26684 13524
rect 26740 13468 29596 13524
rect 29652 13468 29662 13524
rect 35746 13468 35756 13524
rect 35812 13468 38444 13524
rect 38500 13468 38510 13524
rect 39778 13468 39788 13524
rect 39844 13468 40796 13524
rect 40852 13468 40862 13524
rect 45266 13468 45276 13524
rect 45332 13468 46956 13524
rect 47012 13468 47022 13524
rect 76066 13468 76076 13524
rect 76132 13468 77812 13524
rect 78082 13468 78092 13524
rect 78148 13468 78158 13524
rect 0 13440 800 13468
rect 21746 13356 21756 13412
rect 21812 13356 22988 13412
rect 23044 13356 25004 13412
rect 25060 13356 25070 13412
rect 49858 13356 49868 13412
rect 49924 13356 58156 13412
rect 58212 13356 58222 13412
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 65906 13300 65916 13356
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 66180 13300 66190 13356
rect 25442 13244 25452 13300
rect 25508 13244 26124 13300
rect 26180 13244 26190 13300
rect 77756 13188 77812 13468
rect 3332 13132 32956 13188
rect 33012 13132 33022 13188
rect 35074 13132 35084 13188
rect 35140 13132 37436 13188
rect 37492 13132 39228 13188
rect 39284 13132 39294 13188
rect 77746 13132 77756 13188
rect 77812 13132 77822 13188
rect 3332 13076 3388 13132
rect 78092 13076 78148 13468
rect 79200 13076 80000 13104
rect 1922 13020 1932 13076
rect 1988 13020 3388 13076
rect 11666 13020 11676 13076
rect 11732 13020 19572 13076
rect 21410 13020 21420 13076
rect 21476 13020 22540 13076
rect 22596 13020 22606 13076
rect 23762 13020 23772 13076
rect 23828 13020 26572 13076
rect 26628 13020 26638 13076
rect 78092 13020 80000 13076
rect 19516 12964 19572 13020
rect 79200 12992 80000 13020
rect 19506 12908 19516 12964
rect 19572 12908 20972 12964
rect 21028 12908 25676 12964
rect 25732 12908 25742 12964
rect 33170 12908 33180 12964
rect 33236 12908 33852 12964
rect 33908 12908 34412 12964
rect 34468 12908 34478 12964
rect 34738 12908 34748 12964
rect 34804 12908 35420 12964
rect 35476 12908 35486 12964
rect 36194 12908 36204 12964
rect 36260 12908 42364 12964
rect 42420 12908 42430 12964
rect 2034 12796 2044 12852
rect 2100 12796 8316 12852
rect 8372 12796 8382 12852
rect 19516 12516 19572 12908
rect 27122 12796 27132 12852
rect 27188 12796 27916 12852
rect 27972 12796 29148 12852
rect 29204 12796 29214 12852
rect 41990 12796 42028 12852
rect 42084 12796 42094 12852
rect 43138 12796 43148 12852
rect 43204 12796 59500 12852
rect 59556 12796 59566 12852
rect 20178 12684 20188 12740
rect 20244 12684 21420 12740
rect 21476 12684 21486 12740
rect 31378 12684 31388 12740
rect 31444 12684 73052 12740
rect 73108 12684 73118 12740
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 50546 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50830 12572
rect 19506 12460 19516 12516
rect 19572 12460 19582 12516
rect 28242 12460 28252 12516
rect 28308 12460 33964 12516
rect 34020 12460 34030 12516
rect 37986 12460 37996 12516
rect 38052 12460 39564 12516
rect 39620 12460 39630 12516
rect 40898 12460 40908 12516
rect 40964 12460 40974 12516
rect 0 12404 800 12432
rect 40908 12404 40964 12460
rect 0 12348 1708 12404
rect 1764 12348 2492 12404
rect 2548 12348 2558 12404
rect 8306 12348 8316 12404
rect 8372 12348 42364 12404
rect 42420 12348 42430 12404
rect 75170 12348 75180 12404
rect 75236 12348 75964 12404
rect 76020 12348 76030 12404
rect 0 12320 800 12348
rect 19842 12236 19852 12292
rect 19908 12236 20412 12292
rect 20468 12236 20478 12292
rect 24546 12236 24556 12292
rect 24612 12236 25452 12292
rect 25508 12236 25518 12292
rect 31490 12236 31500 12292
rect 31556 12236 32060 12292
rect 32116 12236 36988 12292
rect 37044 12236 37054 12292
rect 26338 12124 26348 12180
rect 26404 12124 33068 12180
rect 33124 12124 33134 12180
rect 36866 12124 36876 12180
rect 36932 12124 37324 12180
rect 37380 12124 37390 12180
rect 40674 12124 40684 12180
rect 40740 12124 41580 12180
rect 41636 12124 41646 12180
rect 9426 12012 9436 12068
rect 9492 12012 10332 12068
rect 10388 12012 10398 12068
rect 17938 12012 17948 12068
rect 18004 12012 19292 12068
rect 19348 12012 19358 12068
rect 22530 12012 22540 12068
rect 22596 12012 25340 12068
rect 25396 12012 25406 12068
rect 33954 12012 33964 12068
rect 34020 12012 36988 12068
rect 37044 12012 37054 12068
rect 39218 12012 39228 12068
rect 39284 12012 41468 12068
rect 41524 12012 41534 12068
rect 79200 11956 80000 11984
rect 31714 11900 31724 11956
rect 31780 11900 37436 11956
rect 37492 11900 37502 11956
rect 77634 11900 77644 11956
rect 77700 11900 78204 11956
rect 78260 11900 80000 11956
rect 79200 11872 80000 11900
rect 16034 11788 16044 11844
rect 16100 11788 20300 11844
rect 20356 11788 20366 11844
rect 24322 11788 24332 11844
rect 24388 11788 27244 11844
rect 27300 11788 27310 11844
rect 27458 11788 27468 11844
rect 27524 11788 33852 11844
rect 33908 11788 33918 11844
rect 45602 11788 45612 11844
rect 45668 11788 48860 11844
rect 48916 11788 48926 11844
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 65906 11732 65916 11788
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 66180 11732 66190 11788
rect 14578 11676 14588 11732
rect 14644 11676 16380 11732
rect 16436 11676 16446 11732
rect 24098 11676 24108 11732
rect 24164 11676 25228 11732
rect 25284 11676 25676 11732
rect 25732 11676 26684 11732
rect 26740 11676 26750 11732
rect 37202 11676 37212 11732
rect 37268 11676 56588 11732
rect 56644 11676 56654 11732
rect 33282 11564 33292 11620
rect 33348 11564 53900 11620
rect 53956 11564 53966 11620
rect 11666 11452 11676 11508
rect 11732 11452 12460 11508
rect 12516 11452 12526 11508
rect 19842 11452 19852 11508
rect 19908 11452 20636 11508
rect 20692 11452 21532 11508
rect 21588 11452 21598 11508
rect 25890 11452 25900 11508
rect 25956 11452 28252 11508
rect 28308 11452 28318 11508
rect 31826 11452 31836 11508
rect 31892 11452 55020 11508
rect 55076 11452 55086 11508
rect 19058 11340 19068 11396
rect 19124 11340 22092 11396
rect 22148 11340 22158 11396
rect 32386 11340 32396 11396
rect 32452 11340 35980 11396
rect 36036 11340 36046 11396
rect 38210 11340 38220 11396
rect 38276 11340 39676 11396
rect 39732 11340 39742 11396
rect 40338 11340 40348 11396
rect 40404 11340 41692 11396
rect 41748 11340 41758 11396
rect 75506 11340 75516 11396
rect 75572 11340 76412 11396
rect 76468 11340 76478 11396
rect 0 11284 800 11312
rect 0 11228 1708 11284
rect 1764 11228 1774 11284
rect 2034 11228 2044 11284
rect 2100 11228 8316 11284
rect 8372 11228 8382 11284
rect 9538 11228 9548 11284
rect 9604 11228 11564 11284
rect 11620 11228 11630 11284
rect 24882 11228 24892 11284
rect 24948 11228 26124 11284
rect 26180 11228 26190 11284
rect 30034 11228 30044 11284
rect 30100 11228 31388 11284
rect 31444 11228 31454 11284
rect 31938 11228 31948 11284
rect 32004 11228 32620 11284
rect 32676 11228 32686 11284
rect 46498 11228 46508 11284
rect 46564 11228 67452 11284
rect 67508 11228 67518 11284
rect 0 11200 800 11228
rect 1708 11172 1764 11228
rect 1708 11116 2492 11172
rect 2548 11116 2558 11172
rect 18610 11116 18620 11172
rect 18676 11116 19740 11172
rect 19796 11116 19806 11172
rect 22082 11116 22092 11172
rect 22148 11116 24780 11172
rect 24836 11116 24846 11172
rect 26898 11116 26908 11172
rect 26964 11116 32508 11172
rect 32564 11116 36428 11172
rect 36484 11116 38668 11172
rect 38724 11116 38734 11172
rect 45154 11116 45164 11172
rect 45220 11116 54908 11172
rect 54964 11116 54974 11172
rect 31266 11004 31276 11060
rect 31332 11004 32172 11060
rect 32228 11004 32238 11060
rect 33730 11004 33740 11060
rect 33796 11004 34132 11060
rect 38546 11004 38556 11060
rect 38612 11004 47348 11060
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 34076 10948 34132 11004
rect 47292 10948 47348 11004
rect 50546 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50830 11004
rect 33170 10892 33180 10948
rect 33236 10892 33852 10948
rect 33908 10892 33918 10948
rect 34076 10892 38668 10948
rect 39554 10892 39564 10948
rect 39620 10892 40348 10948
rect 40404 10892 40414 10948
rect 47282 10892 47292 10948
rect 47348 10892 47358 10948
rect 38612 10836 38668 10892
rect 79200 10836 80000 10864
rect 11106 10780 11116 10836
rect 11172 10780 11564 10836
rect 11620 10780 14924 10836
rect 14980 10780 14990 10836
rect 24994 10780 25004 10836
rect 25060 10780 25788 10836
rect 25844 10780 25854 10836
rect 30930 10780 30940 10836
rect 30996 10780 31500 10836
rect 31556 10780 31566 10836
rect 38612 10780 52556 10836
rect 52612 10780 52622 10836
rect 77634 10780 77644 10836
rect 77700 10780 78204 10836
rect 78260 10780 80000 10836
rect 79200 10752 80000 10780
rect 2034 10668 2044 10724
rect 2100 10668 27972 10724
rect 28130 10668 28140 10724
rect 28196 10668 29484 10724
rect 29540 10668 33292 10724
rect 33348 10668 33358 10724
rect 27916 10612 27972 10668
rect 12674 10556 12684 10612
rect 12740 10556 15372 10612
rect 15428 10556 15438 10612
rect 24770 10556 24780 10612
rect 24836 10556 25228 10612
rect 25284 10556 26236 10612
rect 26292 10556 26302 10612
rect 8194 10444 8204 10500
rect 8260 10444 11452 10500
rect 11508 10444 11518 10500
rect 18274 10444 18284 10500
rect 18340 10444 19516 10500
rect 19572 10444 19582 10500
rect 22530 10444 22540 10500
rect 22596 10444 24220 10500
rect 24276 10444 24286 10500
rect 26852 10388 26908 10612
rect 26964 10556 26974 10612
rect 27916 10556 30156 10612
rect 30212 10556 30222 10612
rect 29474 10444 29484 10500
rect 29540 10444 31388 10500
rect 31444 10444 31454 10500
rect 2370 10332 2380 10388
rect 2436 10332 9996 10388
rect 10052 10332 10062 10388
rect 22754 10332 22764 10388
rect 22820 10332 26908 10388
rect 20962 10220 20972 10276
rect 21028 10220 31780 10276
rect 42354 10220 42364 10276
rect 42420 10220 45164 10276
rect 45220 10220 45230 10276
rect 0 10164 800 10192
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 31724 10164 31780 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 65906 10164 65916 10220
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 66180 10164 66190 10220
rect 0 10108 1708 10164
rect 1764 10108 2492 10164
rect 2548 10108 2558 10164
rect 28018 10108 28028 10164
rect 28084 10108 29820 10164
rect 29876 10108 29886 10164
rect 31714 10108 31724 10164
rect 31780 10108 31790 10164
rect 0 10080 800 10108
rect 11218 9996 11228 10052
rect 11284 9996 12236 10052
rect 12292 9996 12302 10052
rect 14914 9996 14924 10052
rect 14980 9996 24668 10052
rect 24724 9996 24734 10052
rect 31826 9996 31836 10052
rect 31892 9996 37996 10052
rect 38052 9996 38062 10052
rect 38210 9996 38220 10052
rect 38276 9996 38780 10052
rect 38836 9996 38846 10052
rect 42578 9996 42588 10052
rect 42644 9996 42654 10052
rect 43362 9996 43372 10052
rect 43428 9996 60172 10052
rect 60228 9996 60238 10052
rect 42588 9940 42644 9996
rect 8418 9884 8428 9940
rect 8484 9884 13468 9940
rect 13524 9884 13534 9940
rect 13906 9884 13916 9940
rect 13972 9884 14476 9940
rect 14532 9884 15484 9940
rect 15540 9884 15550 9940
rect 20178 9884 20188 9940
rect 20244 9884 20748 9940
rect 20804 9884 22764 9940
rect 22820 9884 22830 9940
rect 30146 9884 30156 9940
rect 30212 9884 34860 9940
rect 34916 9884 34926 9940
rect 37538 9884 37548 9940
rect 37604 9884 41580 9940
rect 41636 9884 41646 9940
rect 41794 9884 41804 9940
rect 41860 9884 42364 9940
rect 42420 9884 42430 9940
rect 42588 9884 60060 9940
rect 60116 9884 60126 9940
rect 11890 9772 11900 9828
rect 11956 9772 12572 9828
rect 12628 9772 13244 9828
rect 13300 9772 14028 9828
rect 14084 9772 14094 9828
rect 14252 9772 28812 9828
rect 28868 9772 28878 9828
rect 36866 9772 36876 9828
rect 36932 9772 38220 9828
rect 38276 9772 38286 9828
rect 39778 9772 39788 9828
rect 39844 9772 42588 9828
rect 42644 9772 42654 9828
rect 45826 9772 45836 9828
rect 45892 9772 64764 9828
rect 64820 9772 64830 9828
rect 14252 9716 14308 9772
rect 79200 9716 80000 9744
rect 8082 9660 8092 9716
rect 8148 9660 9324 9716
rect 9380 9660 9390 9716
rect 9986 9660 9996 9716
rect 10052 9660 14308 9716
rect 14466 9660 14476 9716
rect 14532 9660 21140 9716
rect 23538 9660 23548 9716
rect 23604 9660 25340 9716
rect 25396 9660 26124 9716
rect 26180 9660 26190 9716
rect 31686 9660 31724 9716
rect 31780 9660 31790 9716
rect 32274 9660 32284 9716
rect 32340 9660 33740 9716
rect 33796 9660 33806 9716
rect 37314 9660 37324 9716
rect 37380 9660 37660 9716
rect 37716 9660 37726 9716
rect 38994 9660 39004 9716
rect 39060 9660 39452 9716
rect 39508 9660 40908 9716
rect 40964 9660 57036 9716
rect 57092 9660 57102 9716
rect 77634 9660 77644 9716
rect 77700 9660 78204 9716
rect 78260 9660 80000 9716
rect 1698 9548 1708 9604
rect 1764 9548 2492 9604
rect 2548 9548 2558 9604
rect 11330 9548 11340 9604
rect 11396 9548 12012 9604
rect 12068 9548 13468 9604
rect 13524 9548 14140 9604
rect 14196 9548 14206 9604
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 21084 9380 21140 9660
rect 79200 9632 80000 9660
rect 26852 9548 33292 9604
rect 33348 9548 33358 9604
rect 37986 9548 37996 9604
rect 38052 9548 42140 9604
rect 42196 9548 42206 9604
rect 43138 9548 43148 9604
rect 43204 9548 43932 9604
rect 43988 9548 43998 9604
rect 47954 9548 47964 9604
rect 48020 9548 51716 9604
rect 51874 9548 51884 9604
rect 51940 9548 59612 9604
rect 59668 9548 59678 9604
rect 75282 9548 75292 9604
rect 75348 9548 78092 9604
rect 78148 9548 78158 9604
rect 26852 9492 26908 9548
rect 25666 9436 25676 9492
rect 25732 9436 26908 9492
rect 38546 9436 38556 9492
rect 38612 9436 43372 9492
rect 43428 9436 43438 9492
rect 50546 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50830 9436
rect 51660 9380 51716 9548
rect 18694 9324 18732 9380
rect 18788 9324 18798 9380
rect 21084 9324 29036 9380
rect 29092 9324 29102 9380
rect 31266 9324 31276 9380
rect 31332 9324 38668 9380
rect 51660 9324 52052 9380
rect 53666 9324 53676 9380
rect 53732 9324 69804 9380
rect 69860 9324 69870 9380
rect 75282 9324 75292 9380
rect 75348 9324 76188 9380
rect 76244 9324 76254 9380
rect 38612 9268 38668 9324
rect 51996 9268 52052 9324
rect 13794 9212 13804 9268
rect 13860 9212 14252 9268
rect 14308 9212 14924 9268
rect 14980 9212 14990 9268
rect 18274 9212 18284 9268
rect 18340 9212 19180 9268
rect 19236 9212 19246 9268
rect 19590 9212 19628 9268
rect 19684 9212 19694 9268
rect 24658 9212 24668 9268
rect 24724 9212 25452 9268
rect 25508 9212 32396 9268
rect 32452 9212 32844 9268
rect 32900 9212 34076 9268
rect 34132 9212 34142 9268
rect 38612 9212 51772 9268
rect 51828 9212 51838 9268
rect 51996 9212 67116 9268
rect 67172 9212 67182 9268
rect 26562 9100 26572 9156
rect 26628 9100 34524 9156
rect 34580 9100 34590 9156
rect 38658 9100 38668 9156
rect 38724 9100 39788 9156
rect 39844 9100 39854 9156
rect 48402 9100 48412 9156
rect 48468 9100 63868 9156
rect 63924 9100 63934 9156
rect 0 9044 800 9072
rect 0 8988 1708 9044
rect 1764 8988 1774 9044
rect 18834 8988 18844 9044
rect 18900 8988 19516 9044
rect 19572 8988 21644 9044
rect 21700 8988 22764 9044
rect 22820 8988 23548 9044
rect 23604 8988 23614 9044
rect 24994 8988 25004 9044
rect 25060 8988 29260 9044
rect 29316 8988 29326 9044
rect 0 8960 800 8988
rect 8866 8876 8876 8932
rect 8932 8876 10332 8932
rect 10388 8876 10398 8932
rect 12450 8876 12460 8932
rect 12516 8876 13244 8932
rect 13300 8876 13310 8932
rect 16258 8876 16268 8932
rect 16324 8876 18172 8932
rect 18228 8876 18238 8932
rect 19170 8876 19180 8932
rect 19236 8876 20300 8932
rect 20356 8876 20366 8932
rect 26898 8876 26908 8932
rect 26964 8876 27580 8932
rect 27636 8876 27646 8932
rect 29026 8876 29036 8932
rect 29092 8876 32732 8932
rect 32788 8876 32798 8932
rect 33506 8876 33516 8932
rect 33572 8876 34748 8932
rect 34804 8876 34814 8932
rect 43922 8876 43932 8932
rect 43988 8876 45276 8932
rect 45332 8876 57148 8932
rect 57204 8876 57214 8932
rect 77858 8876 77868 8932
rect 77924 8876 78428 8932
rect 78484 8876 78494 8932
rect 8978 8764 8988 8820
rect 9044 8764 12124 8820
rect 12180 8764 12190 8820
rect 20626 8764 20636 8820
rect 20692 8764 29484 8820
rect 29540 8764 29550 8820
rect 34290 8764 34300 8820
rect 34356 8764 36876 8820
rect 36932 8764 36942 8820
rect 23090 8652 23100 8708
rect 23156 8652 27244 8708
rect 27300 8652 27310 8708
rect 28242 8652 28252 8708
rect 28308 8652 28700 8708
rect 28756 8652 28766 8708
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 65906 8596 65916 8652
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 66180 8596 66190 8652
rect 79200 8596 80000 8624
rect 16818 8540 16828 8596
rect 16884 8540 28196 8596
rect 78082 8540 78092 8596
rect 78148 8540 80000 8596
rect 28140 8484 28196 8540
rect 79200 8512 80000 8540
rect 20626 8428 20636 8484
rect 20692 8428 22204 8484
rect 22260 8428 22270 8484
rect 26786 8428 26796 8484
rect 26852 8428 27972 8484
rect 28130 8428 28140 8484
rect 28196 8428 28206 8484
rect 28364 8428 29036 8484
rect 29092 8428 29102 8484
rect 30370 8428 30380 8484
rect 30436 8428 50988 8484
rect 51044 8428 51884 8484
rect 51940 8428 51950 8484
rect 27916 8372 27972 8428
rect 28364 8372 28420 8428
rect 15586 8316 15596 8372
rect 15652 8316 18172 8372
rect 18228 8316 18238 8372
rect 19954 8316 19964 8372
rect 20020 8316 20748 8372
rect 20804 8316 22540 8372
rect 22596 8316 22606 8372
rect 26898 8316 26908 8372
rect 26964 8316 27356 8372
rect 27412 8316 27422 8372
rect 27916 8316 28420 8372
rect 28802 8316 28812 8372
rect 28868 8316 73612 8372
rect 73668 8316 73678 8372
rect 76850 8316 76860 8372
rect 76916 8316 77196 8372
rect 77252 8316 77262 8372
rect 17714 8204 17724 8260
rect 17780 8204 18284 8260
rect 18340 8204 18350 8260
rect 19618 8204 19628 8260
rect 19684 8204 19796 8260
rect 19740 8148 19796 8204
rect 26852 8204 29260 8260
rect 29316 8204 29820 8260
rect 29876 8204 31276 8260
rect 31332 8204 31342 8260
rect 37314 8204 37324 8260
rect 37380 8204 38332 8260
rect 38388 8204 38398 8260
rect 38612 8204 38892 8260
rect 38948 8204 38958 8260
rect 39778 8204 39788 8260
rect 39844 8204 39854 8260
rect 43026 8204 43036 8260
rect 43092 8204 44716 8260
rect 44772 8204 44782 8260
rect 46162 8204 46172 8260
rect 46228 8204 75628 8260
rect 75684 8204 76188 8260
rect 76244 8204 76254 8260
rect 76514 8204 76524 8260
rect 76580 8204 77868 8260
rect 77924 8204 77934 8260
rect 19282 8092 19292 8148
rect 19348 8092 19740 8148
rect 19796 8092 19806 8148
rect 26852 8036 26908 8204
rect 38612 8148 38668 8204
rect 32834 8092 32844 8148
rect 32900 8092 38668 8148
rect 39788 8036 39844 8204
rect 40898 8092 40908 8148
rect 40964 8092 42364 8148
rect 42420 8092 43596 8148
rect 43652 8092 43662 8148
rect 44370 8092 44380 8148
rect 44436 8092 45052 8148
rect 45108 8092 45118 8148
rect 74050 8092 74060 8148
rect 74116 8092 76412 8148
rect 76468 8092 76478 8148
rect 25778 7980 25788 8036
rect 25844 7980 26908 8036
rect 28466 7980 28476 8036
rect 28532 7980 33292 8036
rect 33348 7980 33358 8036
rect 37090 7980 37100 8036
rect 37156 7980 39844 8036
rect 43922 7980 43932 8036
rect 43988 7980 45948 8036
rect 46004 7980 49532 8036
rect 49588 7980 49598 8036
rect 49746 7980 49756 8036
rect 49812 7980 62188 8036
rect 62244 7980 62254 8036
rect 0 7924 800 7952
rect 0 7868 1708 7924
rect 1764 7868 2492 7924
rect 2548 7868 2558 7924
rect 26236 7868 28140 7924
rect 28196 7868 28206 7924
rect 29026 7868 29036 7924
rect 29092 7868 30044 7924
rect 30100 7868 30110 7924
rect 31612 7868 37660 7924
rect 37716 7868 38668 7924
rect 0 7840 800 7868
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 18386 7756 18396 7812
rect 18452 7756 19180 7812
rect 19236 7756 19246 7812
rect 26236 7700 26292 7868
rect 31612 7812 31668 7868
rect 27234 7756 27244 7812
rect 27300 7756 31668 7812
rect 31826 7756 31836 7812
rect 31892 7756 35308 7812
rect 35364 7756 35374 7812
rect 2034 7644 2044 7700
rect 2100 7644 5852 7700
rect 5908 7644 5918 7700
rect 13122 7644 13132 7700
rect 13188 7644 13580 7700
rect 13636 7644 14364 7700
rect 14420 7644 14430 7700
rect 16930 7644 16940 7700
rect 16996 7644 17836 7700
rect 17892 7644 17902 7700
rect 19954 7644 19964 7700
rect 20020 7644 20412 7700
rect 20468 7644 20860 7700
rect 20916 7644 22204 7700
rect 22260 7644 23100 7700
rect 23156 7644 23166 7700
rect 24770 7644 24780 7700
rect 24836 7644 26236 7700
rect 26292 7644 26302 7700
rect 26572 7644 27020 7700
rect 27076 7644 27086 7700
rect 27794 7644 27804 7700
rect 27860 7644 28812 7700
rect 28868 7644 28878 7700
rect 29474 7644 29484 7700
rect 29540 7644 30044 7700
rect 30100 7644 30110 7700
rect 33954 7644 33964 7700
rect 34020 7644 34972 7700
rect 35028 7644 35038 7700
rect 17836 7588 17892 7644
rect 26572 7588 26628 7644
rect 13794 7532 13804 7588
rect 13860 7532 14588 7588
rect 14644 7532 14654 7588
rect 15092 7532 15596 7588
rect 15652 7532 15662 7588
rect 17836 7532 18508 7588
rect 18564 7532 18574 7588
rect 25778 7532 25788 7588
rect 25844 7532 26012 7588
rect 26068 7532 26572 7588
rect 26628 7532 26638 7588
rect 15092 7476 15148 7532
rect 27804 7476 27860 7644
rect 28242 7532 28252 7588
rect 28308 7532 30380 7588
rect 30436 7532 33236 7588
rect 33842 7532 33852 7588
rect 33908 7532 37324 7588
rect 37380 7532 37390 7588
rect 38612 7532 38668 7868
rect 38892 7812 38948 7980
rect 50546 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50830 7868
rect 38882 7756 38892 7812
rect 38948 7756 38958 7812
rect 41010 7756 41020 7812
rect 41076 7756 41244 7812
rect 41300 7756 42476 7812
rect 42532 7756 46732 7812
rect 46788 7756 46798 7812
rect 55234 7756 55244 7812
rect 55300 7756 71708 7812
rect 71764 7756 72380 7812
rect 72436 7756 72446 7812
rect 39106 7644 39116 7700
rect 39172 7644 39676 7700
rect 39732 7644 40908 7700
rect 40964 7644 44940 7700
rect 44996 7644 45006 7700
rect 57698 7644 57708 7700
rect 57764 7644 74732 7700
rect 74788 7644 75292 7700
rect 75348 7644 75358 7700
rect 38724 7532 38734 7588
rect 41458 7532 41468 7588
rect 41524 7532 44044 7588
rect 44100 7532 44492 7588
rect 44548 7532 44558 7588
rect 49970 7532 49980 7588
rect 50036 7532 66668 7588
rect 66724 7532 66734 7588
rect 29260 7476 29316 7532
rect 33180 7476 33236 7532
rect 79200 7476 80000 7504
rect 11106 7420 11116 7476
rect 11172 7420 15148 7476
rect 17714 7420 17724 7476
rect 17780 7420 19628 7476
rect 19684 7420 19694 7476
rect 22530 7420 22540 7476
rect 22596 7420 25340 7476
rect 25396 7420 27860 7476
rect 28550 7420 28588 7476
rect 28644 7420 28654 7476
rect 29250 7420 29260 7476
rect 29316 7420 29326 7476
rect 33170 7420 33180 7476
rect 33236 7420 33246 7476
rect 33730 7420 33740 7476
rect 33796 7420 34412 7476
rect 34468 7420 34478 7476
rect 36418 7420 36428 7476
rect 36484 7420 37772 7476
rect 37828 7420 37838 7476
rect 41346 7420 41356 7476
rect 41412 7420 43036 7476
rect 43092 7420 43102 7476
rect 77522 7420 77532 7476
rect 77588 7420 80000 7476
rect 79200 7392 80000 7420
rect 1698 7308 1708 7364
rect 1764 7308 2492 7364
rect 2548 7308 2558 7364
rect 11218 7308 11228 7364
rect 11284 7308 13468 7364
rect 13524 7308 13534 7364
rect 15810 7308 15820 7364
rect 15876 7308 18508 7364
rect 18564 7308 18574 7364
rect 23762 7308 23772 7364
rect 23828 7308 25788 7364
rect 25844 7308 25854 7364
rect 30902 7308 30940 7364
rect 30996 7308 31006 7364
rect 33058 7308 33068 7364
rect 33124 7308 46508 7364
rect 46564 7308 47068 7364
rect 47124 7308 53452 7364
rect 53508 7308 53518 7364
rect 27458 7196 27468 7252
rect 27524 7196 27860 7252
rect 28130 7196 28140 7252
rect 28196 7196 28588 7252
rect 28644 7196 38668 7252
rect 27804 7140 27860 7196
rect 9538 7084 9548 7140
rect 9604 7084 19516 7140
rect 19572 7084 19582 7140
rect 21746 7084 21756 7140
rect 21812 7084 27580 7140
rect 27636 7084 27646 7140
rect 27804 7084 30604 7140
rect 30660 7084 33068 7140
rect 33124 7084 33134 7140
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 6066 6972 6076 7028
rect 6132 6972 13916 7028
rect 13972 6972 13982 7028
rect 17714 6972 17724 7028
rect 17780 6972 19068 7028
rect 19124 6972 19134 7028
rect 24434 6972 24444 7028
rect 24500 6972 25340 7028
rect 25396 6972 25406 7028
rect 26338 6972 26348 7028
rect 26404 6972 26796 7028
rect 26852 6972 26862 7028
rect 28914 6972 28924 7028
rect 28980 6972 31500 7028
rect 31556 6972 31566 7028
rect 38612 6916 38668 7196
rect 65906 7028 65916 7084
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 66180 7028 66190 7084
rect 39218 6972 39228 7028
rect 39284 6972 40124 7028
rect 40180 6972 44268 7028
rect 44324 6972 44334 7028
rect 8194 6860 8204 6916
rect 8260 6860 8652 6916
rect 8708 6860 8876 6916
rect 8932 6860 8942 6916
rect 12338 6860 12348 6916
rect 12404 6860 13468 6916
rect 13524 6860 14252 6916
rect 14308 6860 14318 6916
rect 20178 6860 20188 6916
rect 20244 6860 20972 6916
rect 21028 6860 21038 6916
rect 24322 6860 24332 6916
rect 24388 6860 27916 6916
rect 27972 6860 28140 6916
rect 28196 6860 28206 6916
rect 29586 6860 29596 6916
rect 29652 6860 30044 6916
rect 30100 6860 30110 6916
rect 30790 6860 30828 6916
rect 30884 6860 30894 6916
rect 31164 6860 32172 6916
rect 32228 6860 32238 6916
rect 34402 6860 34412 6916
rect 34468 6860 36428 6916
rect 36484 6860 36494 6916
rect 38612 6860 40292 6916
rect 75170 6860 75180 6916
rect 75236 6860 77196 6916
rect 77252 6860 77262 6916
rect 0 6804 800 6832
rect 0 6748 1708 6804
rect 1764 6748 1774 6804
rect 2146 6748 2156 6804
rect 2212 6748 7532 6804
rect 7588 6748 7598 6804
rect 10770 6748 10780 6804
rect 10836 6748 13580 6804
rect 13636 6748 13646 6804
rect 13794 6748 13804 6804
rect 13860 6748 13870 6804
rect 21858 6748 21868 6804
rect 21924 6748 22540 6804
rect 22596 6748 22606 6804
rect 23314 6748 23324 6804
rect 23380 6748 26236 6804
rect 26292 6748 26302 6804
rect 26898 6748 26908 6804
rect 26964 6748 27804 6804
rect 27860 6748 27870 6804
rect 28242 6748 28252 6804
rect 28308 6748 29260 6804
rect 29316 6748 30268 6804
rect 30324 6748 30884 6804
rect 0 6720 800 6748
rect 13804 6692 13860 6748
rect 30828 6692 30884 6748
rect 12114 6636 12124 6692
rect 12180 6636 12796 6692
rect 12852 6636 13860 6692
rect 14242 6636 14252 6692
rect 14308 6636 15932 6692
rect 15988 6636 15998 6692
rect 18834 6636 18844 6692
rect 18900 6636 19628 6692
rect 19684 6636 19694 6692
rect 19842 6636 19852 6692
rect 19908 6636 27916 6692
rect 27972 6636 27982 6692
rect 28550 6636 28588 6692
rect 28644 6636 28654 6692
rect 30818 6636 30828 6692
rect 30884 6636 30894 6692
rect 31164 6580 31220 6860
rect 31462 6748 31500 6804
rect 31556 6748 31566 6804
rect 31826 6748 31836 6804
rect 31892 6748 32732 6804
rect 32788 6748 32798 6804
rect 33282 6748 33292 6804
rect 33348 6748 34636 6804
rect 34692 6748 34702 6804
rect 34860 6748 38444 6804
rect 38500 6748 38510 6804
rect 32610 6636 32620 6692
rect 32676 6636 34188 6692
rect 34244 6636 34254 6692
rect 34860 6580 34916 6748
rect 40236 6692 40292 6860
rect 43026 6748 43036 6804
rect 43092 6748 45724 6804
rect 45780 6748 45790 6804
rect 75282 6748 75292 6804
rect 75348 6748 76412 6804
rect 76468 6748 77532 6804
rect 77588 6748 78092 6804
rect 78148 6748 78158 6804
rect 36530 6636 36540 6692
rect 36596 6636 39564 6692
rect 39620 6636 39630 6692
rect 40236 6636 49980 6692
rect 50036 6636 50046 6692
rect 51426 6636 51436 6692
rect 51492 6636 69524 6692
rect 69682 6636 69692 6692
rect 69748 6636 71260 6692
rect 71316 6636 71326 6692
rect 69468 6580 69524 6636
rect 4274 6524 4284 6580
rect 4340 6524 9436 6580
rect 9492 6524 9502 6580
rect 14018 6524 14028 6580
rect 14084 6524 15148 6580
rect 15204 6524 21532 6580
rect 21588 6524 21868 6580
rect 21924 6524 21934 6580
rect 25890 6524 25900 6580
rect 25956 6524 26348 6580
rect 26404 6524 26414 6580
rect 28130 6524 28140 6580
rect 28196 6524 28476 6580
rect 28532 6524 30156 6580
rect 30212 6524 30222 6580
rect 31154 6524 31164 6580
rect 31220 6524 31230 6580
rect 33170 6524 33180 6580
rect 33236 6524 34916 6580
rect 50530 6524 50540 6580
rect 50596 6524 51324 6580
rect 51380 6524 69244 6580
rect 69300 6524 69310 6580
rect 69468 6524 74956 6580
rect 75012 6524 75022 6580
rect 76850 6524 76860 6580
rect 76916 6524 77700 6580
rect 4946 6412 4956 6468
rect 5012 6412 8652 6468
rect 8708 6412 8718 6468
rect 8978 6412 8988 6468
rect 9044 6412 9660 6468
rect 9716 6412 9996 6468
rect 10052 6412 10062 6468
rect 12898 6412 12908 6468
rect 12964 6412 13916 6468
rect 13972 6412 14364 6468
rect 14420 6412 14430 6468
rect 14690 6412 14700 6468
rect 14756 6412 15148 6468
rect 18610 6412 18620 6468
rect 18676 6412 18956 6468
rect 19012 6412 19022 6468
rect 19394 6412 19404 6468
rect 19460 6412 19964 6468
rect 20020 6412 20030 6468
rect 21410 6412 21420 6468
rect 21476 6412 23100 6468
rect 23156 6412 23166 6468
rect 28690 6412 28700 6468
rect 28756 6412 30044 6468
rect 30100 6412 40684 6468
rect 40740 6412 40750 6468
rect 47282 6412 47292 6468
rect 47348 6412 56028 6468
rect 56084 6412 56924 6468
rect 56980 6412 56990 6468
rect 60050 6412 60060 6468
rect 60116 6412 61516 6468
rect 61572 6412 61582 6468
rect 62738 6412 62748 6468
rect 62804 6412 64428 6468
rect 64484 6412 64494 6468
rect 67554 6412 67564 6468
rect 67620 6412 69356 6468
rect 69412 6412 69422 6468
rect 70466 6412 70476 6468
rect 70532 6412 72268 6468
rect 72324 6412 72334 6468
rect 75506 6412 75516 6468
rect 75572 6412 77420 6468
rect 77476 6412 77486 6468
rect 14364 6356 14420 6412
rect 15092 6356 15148 6412
rect 77644 6356 77700 6524
rect 79200 6356 80000 6384
rect 14364 6300 14812 6356
rect 14868 6300 14878 6356
rect 15092 6300 18508 6356
rect 18564 6300 18574 6356
rect 26450 6300 26460 6356
rect 26516 6300 29036 6356
rect 29092 6300 29102 6356
rect 30818 6300 30828 6356
rect 30884 6300 31164 6356
rect 31220 6300 31230 6356
rect 62178 6300 62188 6356
rect 62244 6300 67900 6356
rect 67956 6300 67966 6356
rect 69234 6300 69244 6356
rect 69300 6300 76860 6356
rect 76916 6300 76926 6356
rect 77644 6300 80000 6356
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 50546 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50830 6300
rect 79200 6272 80000 6300
rect 7858 6188 7868 6244
rect 7924 6188 8372 6244
rect 12674 6188 12684 6244
rect 12740 6188 14140 6244
rect 14196 6188 16716 6244
rect 16772 6188 16782 6244
rect 22978 6188 22988 6244
rect 23044 6188 27020 6244
rect 27076 6188 27086 6244
rect 30594 6188 30604 6244
rect 30660 6188 31500 6244
rect 31556 6188 31566 6244
rect 39778 6188 39788 6244
rect 39844 6188 44380 6244
rect 44436 6188 44446 6244
rect 58146 6188 58156 6244
rect 58212 6188 67340 6244
rect 67396 6188 68460 6244
rect 68516 6188 68526 6244
rect 73602 6188 73612 6244
rect 73668 6188 75516 6244
rect 75572 6188 75582 6244
rect 8316 6132 8372 6188
rect 3602 6076 3612 6132
rect 3668 6076 7980 6132
rect 8036 6076 8046 6132
rect 8306 6076 8316 6132
rect 8372 6076 8988 6132
rect 9044 6076 9054 6132
rect 13458 6076 13468 6132
rect 13524 6076 15148 6132
rect 15204 6076 15242 6132
rect 17388 6076 18284 6132
rect 18340 6076 18732 6132
rect 18788 6076 18798 6132
rect 22306 6076 22316 6132
rect 22372 6076 24332 6132
rect 24388 6076 24398 6132
rect 26338 6076 26348 6132
rect 26404 6076 27132 6132
rect 27188 6076 27198 6132
rect 29922 6076 29932 6132
rect 29988 6076 35644 6132
rect 35700 6076 35710 6132
rect 46050 6076 46060 6132
rect 46116 6076 47964 6132
rect 48020 6076 48030 6132
rect 48626 6076 48636 6132
rect 48692 6076 49644 6132
rect 49700 6076 49710 6132
rect 49970 6076 49980 6132
rect 50036 6076 50764 6132
rect 50820 6076 52332 6132
rect 52388 6076 52398 6132
rect 68562 6076 68572 6132
rect 68628 6076 77308 6132
rect 77364 6076 78204 6132
rect 78260 6076 78270 6132
rect 17388 6020 17444 6076
rect 2370 5964 2380 6020
rect 2436 5964 6300 6020
rect 6356 5964 6366 6020
rect 6626 5964 6636 6020
rect 6692 5964 8428 6020
rect 8484 5964 8494 6020
rect 13682 5964 13692 6020
rect 13748 5964 17444 6020
rect 18386 5964 18396 6020
rect 18452 5964 22036 6020
rect 23986 5964 23996 6020
rect 24052 5964 29036 6020
rect 29092 5964 29102 6020
rect 30828 5964 34300 6020
rect 34356 5964 34366 6020
rect 42242 5964 42252 6020
rect 42308 5964 45164 6020
rect 45220 5964 45612 6020
rect 45668 5964 45678 6020
rect 48850 5964 48860 6020
rect 48916 5964 63196 6020
rect 63252 5964 63262 6020
rect 21980 5908 22036 5964
rect 30828 5908 30884 5964
rect 5618 5852 5628 5908
rect 5684 5852 8092 5908
rect 8148 5852 8158 5908
rect 10210 5852 10220 5908
rect 10276 5852 12572 5908
rect 12628 5852 12638 5908
rect 14018 5852 14028 5908
rect 14084 5852 14094 5908
rect 14690 5852 14700 5908
rect 14756 5852 17388 5908
rect 17444 5852 17454 5908
rect 18610 5852 18620 5908
rect 18676 5852 21756 5908
rect 21812 5852 21822 5908
rect 21980 5852 25564 5908
rect 25620 5852 25630 5908
rect 29250 5852 29260 5908
rect 29316 5852 30044 5908
rect 30100 5852 30110 5908
rect 30818 5852 30828 5908
rect 30884 5852 30894 5908
rect 32162 5852 32172 5908
rect 32228 5852 33516 5908
rect 33572 5852 33582 5908
rect 33842 5852 33852 5908
rect 33908 5852 37548 5908
rect 37604 5852 37614 5908
rect 41794 5852 41804 5908
rect 41860 5852 42476 5908
rect 42532 5852 44268 5908
rect 44324 5852 44828 5908
rect 44884 5852 44894 5908
rect 47506 5852 47516 5908
rect 47572 5852 49868 5908
rect 49924 5852 49934 5908
rect 55346 5852 55356 5908
rect 55412 5852 71708 5908
rect 71764 5852 72268 5908
rect 72324 5852 72334 5908
rect 14028 5796 14084 5852
rect 6850 5740 6860 5796
rect 6916 5740 11004 5796
rect 11060 5740 11070 5796
rect 12002 5740 12012 5796
rect 12068 5740 14084 5796
rect 15586 5740 15596 5796
rect 15652 5740 16828 5796
rect 16884 5740 16894 5796
rect 19618 5740 19628 5796
rect 19684 5740 21084 5796
rect 21140 5740 21150 5796
rect 21970 5740 21980 5796
rect 22036 5740 26292 5796
rect 26898 5740 26908 5796
rect 26964 5740 27244 5796
rect 27300 5740 27310 5796
rect 30930 5740 30940 5796
rect 30996 5740 34300 5796
rect 34356 5740 34366 5796
rect 38098 5740 38108 5796
rect 38164 5740 40012 5796
rect 40068 5740 50092 5796
rect 50148 5740 50158 5796
rect 54338 5740 54348 5796
rect 54404 5740 70476 5796
rect 70532 5740 70542 5796
rect 72818 5740 72828 5796
rect 72884 5740 75628 5796
rect 75684 5740 75694 5796
rect 0 5684 800 5712
rect 26236 5684 26292 5740
rect 0 5628 1708 5684
rect 1764 5628 2492 5684
rect 2548 5628 2558 5684
rect 11218 5628 11228 5684
rect 11284 5628 13804 5684
rect 13860 5628 13870 5684
rect 21186 5628 21196 5684
rect 21252 5628 23660 5684
rect 23716 5628 23726 5684
rect 25106 5628 25116 5684
rect 25172 5628 25788 5684
rect 25844 5628 25854 5684
rect 26226 5628 26236 5684
rect 26292 5628 26302 5684
rect 26674 5628 26684 5684
rect 26740 5628 32620 5684
rect 32676 5628 32686 5684
rect 33842 5628 33852 5684
rect 33908 5628 36764 5684
rect 36820 5628 36830 5684
rect 56690 5628 56700 5684
rect 56756 5628 57932 5684
rect 57988 5628 57998 5684
rect 59378 5628 59388 5684
rect 59444 5628 60844 5684
rect 60900 5628 60910 5684
rect 70802 5628 70812 5684
rect 70868 5628 73276 5684
rect 73332 5628 73342 5684
rect 0 5600 800 5628
rect 4834 5516 4844 5572
rect 4900 5516 8652 5572
rect 8708 5516 8718 5572
rect 9986 5516 9996 5572
rect 10052 5516 13468 5572
rect 13524 5516 13534 5572
rect 13906 5516 13916 5572
rect 13972 5516 14028 5572
rect 14084 5516 14094 5572
rect 14354 5516 14364 5572
rect 14420 5516 21924 5572
rect 22642 5516 22652 5572
rect 22708 5516 28028 5572
rect 28084 5516 28094 5572
rect 33282 5516 33292 5572
rect 33348 5516 33740 5572
rect 33796 5516 33806 5572
rect 45154 5516 45164 5572
rect 45220 5516 47628 5572
rect 47684 5516 47694 5572
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 21868 5460 21924 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 65906 5460 65916 5516
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 66180 5460 66190 5516
rect 6290 5404 6300 5460
rect 6356 5404 10556 5460
rect 10612 5404 10622 5460
rect 13906 5404 13916 5460
rect 13972 5404 20412 5460
rect 20468 5404 20478 5460
rect 21858 5404 21868 5460
rect 21924 5404 21934 5460
rect 25778 5404 25788 5460
rect 25844 5404 26572 5460
rect 26628 5404 26796 5460
rect 26852 5404 26862 5460
rect 27234 5404 27244 5460
rect 27300 5404 29260 5460
rect 29316 5404 29326 5460
rect 48066 5404 48076 5460
rect 48132 5404 50428 5460
rect 75058 5404 75068 5460
rect 75124 5404 77588 5460
rect 50372 5348 50428 5404
rect 7634 5292 7644 5348
rect 7700 5292 8988 5348
rect 9044 5292 9054 5348
rect 11442 5292 11452 5348
rect 11508 5292 14812 5348
rect 14868 5292 14878 5348
rect 16594 5292 16604 5348
rect 16660 5292 18284 5348
rect 18340 5292 18350 5348
rect 19394 5292 19404 5348
rect 19460 5292 20748 5348
rect 20804 5292 21420 5348
rect 21476 5292 21486 5348
rect 22306 5292 22316 5348
rect 22372 5292 23604 5348
rect 24658 5292 24668 5348
rect 24724 5292 24734 5348
rect 27794 5292 27804 5348
rect 27860 5292 31612 5348
rect 31668 5292 31678 5348
rect 31826 5292 31836 5348
rect 31892 5292 36540 5348
rect 36596 5292 36606 5348
rect 38322 5292 38332 5348
rect 38388 5292 39452 5348
rect 39508 5292 39518 5348
rect 45938 5292 45948 5348
rect 46004 5292 49196 5348
rect 49252 5292 49756 5348
rect 49812 5292 49822 5348
rect 50372 5292 50540 5348
rect 50596 5292 51212 5348
rect 51268 5292 51278 5348
rect 66322 5292 66332 5348
rect 66388 5292 69356 5348
rect 69412 5292 69422 5348
rect 70466 5292 70476 5348
rect 70532 5292 75180 5348
rect 75236 5292 75246 5348
rect 23548 5236 23604 5292
rect 24668 5236 24724 5292
rect 77532 5236 77588 5404
rect 79200 5236 80000 5264
rect 8306 5180 8316 5236
rect 8372 5180 12460 5236
rect 12516 5180 12526 5236
rect 13458 5180 13468 5236
rect 13524 5180 14420 5236
rect 16706 5180 16716 5236
rect 16772 5180 17388 5236
rect 17444 5180 17454 5236
rect 18694 5180 18732 5236
rect 18788 5180 18798 5236
rect 21186 5180 21196 5236
rect 21252 5180 22988 5236
rect 23044 5180 23054 5236
rect 23538 5180 23548 5236
rect 23604 5180 23614 5236
rect 24668 5180 27580 5236
rect 27636 5180 27646 5236
rect 27906 5180 27916 5236
rect 27972 5180 28700 5236
rect 28756 5180 28924 5236
rect 28980 5180 29596 5236
rect 29652 5180 29662 5236
rect 31378 5180 31388 5236
rect 31444 5180 31724 5236
rect 31780 5180 33852 5236
rect 33908 5180 33918 5236
rect 34066 5180 34076 5236
rect 34132 5180 40516 5236
rect 42130 5180 42140 5236
rect 42196 5180 43260 5236
rect 43316 5180 45500 5236
rect 45556 5180 45566 5236
rect 47954 5180 47964 5236
rect 48020 5180 48748 5236
rect 48804 5180 48814 5236
rect 54002 5180 54012 5236
rect 54068 5180 55244 5236
rect 55300 5180 55310 5236
rect 56130 5180 56140 5236
rect 56196 5180 58156 5236
rect 58212 5180 58222 5236
rect 60722 5180 60732 5236
rect 60788 5180 64428 5236
rect 64484 5180 64494 5236
rect 64642 5180 64652 5236
rect 64708 5180 66444 5236
rect 66500 5180 66510 5236
rect 68114 5180 68124 5236
rect 68180 5180 72268 5236
rect 72324 5180 72334 5236
rect 73490 5180 73500 5236
rect 73556 5180 76300 5236
rect 76356 5180 76366 5236
rect 77532 5180 78092 5236
rect 78148 5180 80000 5236
rect 6066 5068 6076 5124
rect 6132 5068 7980 5124
rect 8036 5068 8046 5124
rect 8866 5068 8876 5124
rect 8932 5068 11676 5124
rect 11732 5068 11742 5124
rect 13010 5068 13020 5124
rect 13076 5068 14196 5124
rect 14140 5012 14196 5068
rect 14364 5012 14420 5180
rect 40460 5124 40516 5180
rect 79200 5152 80000 5180
rect 14578 5068 14588 5124
rect 14644 5068 15932 5124
rect 15988 5068 15998 5124
rect 16482 5068 16492 5124
rect 16548 5068 19404 5124
rect 19460 5068 19470 5124
rect 20066 5068 20076 5124
rect 20132 5068 22484 5124
rect 22866 5068 22876 5124
rect 22932 5068 25228 5124
rect 25284 5068 25294 5124
rect 27122 5068 27132 5124
rect 27188 5068 28028 5124
rect 28084 5068 28094 5124
rect 29474 5068 29484 5124
rect 29540 5068 30604 5124
rect 30660 5068 30670 5124
rect 32274 5068 32284 5124
rect 32340 5068 33180 5124
rect 33236 5068 33246 5124
rect 33506 5068 33516 5124
rect 33572 5068 37324 5124
rect 37380 5068 37390 5124
rect 37874 5068 37884 5124
rect 37940 5068 39676 5124
rect 39732 5068 40012 5124
rect 40068 5068 40078 5124
rect 40450 5068 40460 5124
rect 40516 5068 40526 5124
rect 41794 5068 41804 5124
rect 41860 5068 46396 5124
rect 46452 5068 46844 5124
rect 46900 5068 46910 5124
rect 48178 5068 48188 5124
rect 48244 5068 48972 5124
rect 49028 5068 49038 5124
rect 63746 5068 63756 5124
rect 63812 5068 65548 5124
rect 65604 5068 65614 5124
rect 66770 5068 66780 5124
rect 66836 5068 67788 5124
rect 67844 5068 67854 5124
rect 72146 5068 72156 5124
rect 72212 5068 73948 5124
rect 74004 5068 74014 5124
rect 76962 5068 76972 5124
rect 77028 5068 78316 5124
rect 78372 5068 78382 5124
rect 17948 5012 18004 5068
rect 22428 5012 22484 5068
rect 1586 4956 1596 5012
rect 1652 4956 2716 5012
rect 2772 4956 2782 5012
rect 6738 4956 6748 5012
rect 6804 4956 7308 5012
rect 7364 4956 7374 5012
rect 14130 4956 14140 5012
rect 14196 4956 14206 5012
rect 14364 4956 14700 5012
rect 14756 4956 14766 5012
rect 17938 4956 17948 5012
rect 18004 4956 18014 5012
rect 22418 4956 22428 5012
rect 22484 4956 22494 5012
rect 28802 4956 28812 5012
rect 28868 4956 29932 5012
rect 29988 4956 29998 5012
rect 30258 4956 30268 5012
rect 30324 4956 35308 5012
rect 35364 4956 35374 5012
rect 40226 4956 40236 5012
rect 40292 4956 42476 5012
rect 42532 4956 42542 5012
rect 55010 4956 55020 5012
rect 55076 4956 55916 5012
rect 55972 4956 55982 5012
rect 6178 4844 6188 4900
rect 6244 4844 6524 4900
rect 6580 4844 6590 4900
rect 6850 4844 6860 4900
rect 6916 4844 7644 4900
rect 7700 4844 7710 4900
rect 13794 4844 13804 4900
rect 13860 4844 14252 4900
rect 14308 4844 14924 4900
rect 14980 4844 15260 4900
rect 15316 4844 15326 4900
rect 27122 4844 27132 4900
rect 27188 4844 33292 4900
rect 33348 4844 33358 4900
rect 39778 4844 39788 4900
rect 39844 4844 41580 4900
rect 41636 4844 45388 4900
rect 45444 4844 45454 4900
rect 46610 4844 46620 4900
rect 46676 4844 49868 4900
rect 49924 4844 49934 4900
rect 58706 4844 58716 4900
rect 58772 4844 61516 4900
rect 61572 4844 61582 4900
rect 14326 4732 14364 4788
rect 14420 4732 14430 4788
rect 25442 4732 25452 4788
rect 25508 4732 30716 4788
rect 30772 4732 30782 4788
rect 30930 4732 30940 4788
rect 30996 4732 36428 4788
rect 36484 4732 36494 4788
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 30940 4676 30996 4732
rect 50546 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50830 4732
rect 7074 4620 7084 4676
rect 7140 4620 7150 4676
rect 8530 4620 8540 4676
rect 8596 4620 14924 4676
rect 14980 4620 14990 4676
rect 15138 4620 15148 4676
rect 15204 4620 16044 4676
rect 16100 4620 16110 4676
rect 23762 4620 23772 4676
rect 23828 4620 29820 4676
rect 29876 4620 29886 4676
rect 30258 4620 30268 4676
rect 30324 4620 30996 4676
rect 33394 4620 33404 4676
rect 33460 4620 34524 4676
rect 34580 4620 34590 4676
rect 46620 4620 47404 4676
rect 47460 4620 47470 4676
rect 0 4564 800 4592
rect 7084 4564 7140 4620
rect 46620 4564 46676 4620
rect 0 4508 1708 4564
rect 1764 4508 2492 4564
rect 2548 4508 2558 4564
rect 7084 4508 8764 4564
rect 8820 4508 14252 4564
rect 14308 4508 14318 4564
rect 19954 4508 19964 4564
rect 20020 4508 20300 4564
rect 20356 4508 20366 4564
rect 20626 4508 20636 4564
rect 20692 4508 21308 4564
rect 21364 4508 21868 4564
rect 21924 4508 22876 4564
rect 22932 4508 22942 4564
rect 32386 4508 32396 4564
rect 32452 4508 34188 4564
rect 34244 4508 34254 4564
rect 36082 4508 36092 4564
rect 36148 4508 43708 4564
rect 43764 4508 43774 4564
rect 45602 4508 45612 4564
rect 45668 4508 46620 4564
rect 46676 4508 46686 4564
rect 47170 4508 47180 4564
rect 47236 4508 48748 4564
rect 48804 4508 48814 4564
rect 53778 4508 53788 4564
rect 53844 4508 71708 4564
rect 71764 4508 72268 4564
rect 72324 4508 72334 4564
rect 0 4480 800 4508
rect 7634 4396 7644 4452
rect 7700 4396 10892 4452
rect 10948 4396 10958 4452
rect 12226 4396 12236 4452
rect 12292 4396 17724 4452
rect 17780 4396 17790 4452
rect 18274 4396 18284 4452
rect 18340 4396 20412 4452
rect 20468 4396 20478 4452
rect 21746 4396 21756 4452
rect 21812 4396 23100 4452
rect 23156 4396 23166 4452
rect 23986 4396 23996 4452
rect 24052 4396 28812 4452
rect 28868 4396 28878 4452
rect 30034 4396 30044 4452
rect 30100 4396 31108 4452
rect 32722 4396 32732 4452
rect 32788 4396 36652 4452
rect 36708 4396 36718 4452
rect 61618 4396 61628 4452
rect 61684 4396 62524 4452
rect 62580 4396 62590 4452
rect 31052 4340 31108 4396
rect 4498 4284 4508 4340
rect 4564 4284 6636 4340
rect 6692 4284 6702 4340
rect 10210 4284 10220 4340
rect 10276 4284 13692 4340
rect 13748 4284 14588 4340
rect 14644 4284 14654 4340
rect 15026 4284 15036 4340
rect 15092 4284 18956 4340
rect 19012 4284 19022 4340
rect 19394 4284 19404 4340
rect 19460 4284 22876 4340
rect 22932 4284 22942 4340
rect 25778 4284 25788 4340
rect 25844 4284 30828 4340
rect 30884 4284 30894 4340
rect 31052 4284 32956 4340
rect 33012 4284 33022 4340
rect 33170 4284 33180 4340
rect 33236 4284 33274 4340
rect 33394 4284 33404 4340
rect 33460 4284 36540 4340
rect 36596 4284 36606 4340
rect 42690 4284 42700 4340
rect 42756 4284 48524 4340
rect 48580 4284 48590 4340
rect 49074 4284 49084 4340
rect 49140 4284 52556 4340
rect 52612 4284 52622 4340
rect 56578 4284 56588 4340
rect 56644 4284 58044 4340
rect 58100 4284 58110 4340
rect 64530 4284 64540 4340
rect 64596 4284 65660 4340
rect 65716 4284 65726 4340
rect 1810 4172 1820 4228
rect 1876 4172 2492 4228
rect 2548 4172 2558 4228
rect 4610 4172 4620 4228
rect 4676 4172 6188 4228
rect 6244 4172 6254 4228
rect 6402 4172 6412 4228
rect 6468 4172 7364 4228
rect 8194 4172 8204 4228
rect 8260 4172 11004 4228
rect 11060 4172 11070 4228
rect 11890 4172 11900 4228
rect 11956 4172 14476 4228
rect 14532 4172 14542 4228
rect 16034 4172 16044 4228
rect 16100 4172 21196 4228
rect 21252 4172 21262 4228
rect 21746 4172 21756 4228
rect 21812 4172 26012 4228
rect 26068 4172 26078 4228
rect 30258 4172 30268 4228
rect 30324 4172 34972 4228
rect 35028 4172 35038 4228
rect 35522 4172 35532 4228
rect 35588 4172 43148 4228
rect 43204 4172 43214 4228
rect 46610 4172 46620 4228
rect 46676 4172 48972 4228
rect 49028 4172 49038 4228
rect 52210 4172 52220 4228
rect 52276 4172 70532 4228
rect 73042 4172 73052 4228
rect 73108 4172 74172 4228
rect 74228 4172 74238 4228
rect 7308 4116 7364 4172
rect 6290 4060 6300 4116
rect 6356 4060 6972 4116
rect 7028 4060 7038 4116
rect 7298 4060 7308 4116
rect 7364 4060 9268 4116
rect 9650 4060 9660 4116
rect 9716 4060 10220 4116
rect 10276 4060 13580 4116
rect 13636 4060 13646 4116
rect 15092 4060 16268 4116
rect 16324 4060 16334 4116
rect 17490 4060 17500 4116
rect 17556 4060 17948 4116
rect 18004 4060 18014 4116
rect 18582 4060 18620 4116
rect 18676 4060 18686 4116
rect 19170 4060 19180 4116
rect 19236 4060 19964 4116
rect 20020 4060 20030 4116
rect 20738 4060 20748 4116
rect 20804 4060 22988 4116
rect 23044 4060 23054 4116
rect 24322 4060 24332 4116
rect 24388 4060 26348 4116
rect 26404 4060 26414 4116
rect 29922 4060 29932 4116
rect 29988 4060 33180 4116
rect 33236 4060 33246 4116
rect 34738 4060 34748 4116
rect 34804 4060 40572 4116
rect 40628 4060 40638 4116
rect 40786 4060 40796 4116
rect 40852 4060 41244 4116
rect 41300 4060 48860 4116
rect 48916 4060 48926 4116
rect 49298 4060 49308 4116
rect 49364 4060 50540 4116
rect 50596 4060 50606 4116
rect 52658 4060 52668 4116
rect 52724 4060 53900 4116
rect 53956 4060 53966 4116
rect 57362 4060 57372 4116
rect 57428 4060 59724 4116
rect 59780 4060 59790 4116
rect 64082 4060 64092 4116
rect 64148 4060 68348 4116
rect 68404 4060 68414 4116
rect 9212 4004 9268 4060
rect 15092 4004 15148 4060
rect 17500 4004 17556 4060
rect 70476 4004 70532 4172
rect 79200 4116 80000 4144
rect 71474 4060 71484 4116
rect 71540 4060 76188 4116
rect 76244 4060 76254 4116
rect 78418 4060 78428 4116
rect 78484 4060 80000 4116
rect 79200 4032 80000 4060
rect 6514 3948 6524 4004
rect 6580 3948 8988 4004
rect 9044 3948 9054 4004
rect 9212 3948 11452 4004
rect 11508 3948 11518 4004
rect 11676 3948 15148 4004
rect 15698 3948 15708 4004
rect 15764 3948 17556 4004
rect 17826 3948 17836 4004
rect 17892 3948 20524 4004
rect 20580 3948 21756 4004
rect 21812 3948 21822 4004
rect 22418 3948 22428 4004
rect 22484 3948 27020 4004
rect 27076 3948 27086 4004
rect 39330 3948 39340 4004
rect 39396 3948 43036 4004
rect 43092 3948 43102 4004
rect 43922 3948 43932 4004
rect 43988 3948 48972 4004
rect 49028 3948 49038 4004
rect 50082 3948 50092 4004
rect 50148 3948 53564 4004
rect 53620 3948 53630 4004
rect 70466 3948 70476 4004
rect 70532 3948 74060 4004
rect 74116 3948 74126 4004
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 11676 3892 11732 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 65906 3892 65916 3948
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 66180 3892 66190 3948
rect 5394 3836 5404 3892
rect 5460 3836 6972 3892
rect 7028 3836 7038 3892
rect 7410 3836 7420 3892
rect 7476 3836 9996 3892
rect 10052 3836 10062 3892
rect 10322 3836 10332 3892
rect 10388 3836 10780 3892
rect 10836 3836 11732 3892
rect 14130 3836 14140 3892
rect 14196 3836 19068 3892
rect 19124 3836 19134 3892
rect 21074 3836 21084 3892
rect 21140 3836 27692 3892
rect 27748 3836 27758 3892
rect 28578 3836 28588 3892
rect 28644 3836 34860 3892
rect 34916 3836 34926 3892
rect 36306 3836 36316 3892
rect 36372 3836 36876 3892
rect 36932 3836 36942 3892
rect 38612 3836 41132 3892
rect 41188 3836 41198 3892
rect 41906 3836 41916 3892
rect 41972 3836 48748 3892
rect 48804 3836 51100 3892
rect 51156 3836 51166 3892
rect 61394 3836 61404 3892
rect 61460 3836 65548 3892
rect 65604 3836 65614 3892
rect 68786 3836 68796 3892
rect 68852 3836 73276 3892
rect 73332 3836 73342 3892
rect 38612 3780 38668 3836
rect 4722 3724 4732 3780
rect 4788 3724 5068 3780
rect 5124 3724 9548 3780
rect 9604 3724 9614 3780
rect 13458 3724 13468 3780
rect 13524 3724 18396 3780
rect 18452 3724 18462 3780
rect 22978 3724 22988 3780
rect 23044 3724 25956 3780
rect 26114 3724 26124 3780
rect 26180 3724 31836 3780
rect 31892 3724 31902 3780
rect 34962 3724 34972 3780
rect 35028 3724 35868 3780
rect 35924 3724 38668 3780
rect 42578 3724 42588 3780
rect 42644 3724 49420 3780
rect 49476 3724 51548 3780
rect 51604 3724 51614 3780
rect 51986 3724 51996 3780
rect 52052 3724 53228 3780
rect 53284 3724 53676 3780
rect 53732 3724 53742 3780
rect 62066 3724 62076 3780
rect 62132 3724 67452 3780
rect 67508 3724 67518 3780
rect 69458 3724 69468 3780
rect 69524 3724 75068 3780
rect 75124 3724 75134 3780
rect 25900 3668 25956 3724
rect 5842 3612 5852 3668
rect 5908 3612 10332 3668
rect 10388 3612 10398 3668
rect 14802 3612 14812 3668
rect 14868 3612 19404 3668
rect 19460 3612 19470 3668
rect 19954 3612 19964 3668
rect 20020 3612 25676 3668
rect 25732 3612 25742 3668
rect 25900 3612 26404 3668
rect 26898 3612 26908 3668
rect 26964 3612 32508 3668
rect 32564 3612 32574 3668
rect 33730 3612 33740 3668
rect 33796 3612 39900 3668
rect 39956 3612 39966 3668
rect 40226 3612 40236 3668
rect 40292 3612 42308 3668
rect 44594 3612 44604 3668
rect 44660 3612 50092 3668
rect 50148 3612 50158 3668
rect 50372 3612 50652 3668
rect 50708 3612 50718 3668
rect 51314 3612 51324 3668
rect 51380 3612 53004 3668
rect 53060 3612 53070 3668
rect 53330 3612 53340 3668
rect 53396 3612 56028 3668
rect 56084 3612 56094 3668
rect 59042 3612 59052 3668
rect 59108 3612 59118 3668
rect 71250 3612 71260 3668
rect 71316 3612 71326 3668
rect 26348 3556 26404 3612
rect 42252 3556 42308 3612
rect 50372 3556 50428 3612
rect 53004 3556 53060 3612
rect 59052 3556 59108 3612
rect 1810 3500 1820 3556
rect 1876 3500 1886 3556
rect 3378 3500 3388 3556
rect 3444 3500 5628 3556
rect 5684 3500 5694 3556
rect 6514 3500 6524 3556
rect 6580 3500 7196 3556
rect 7252 3500 8260 3556
rect 9650 3500 9660 3556
rect 9716 3500 10444 3556
rect 10500 3500 10510 3556
rect 11666 3500 11676 3556
rect 11732 3500 17052 3556
rect 17108 3500 17118 3556
rect 18498 3500 18508 3556
rect 18564 3500 19180 3556
rect 19236 3500 19246 3556
rect 19506 3500 19516 3556
rect 19572 3500 24780 3556
rect 24836 3500 24846 3556
rect 25330 3500 25340 3556
rect 25396 3500 26124 3556
rect 26180 3500 26190 3556
rect 26348 3500 28476 3556
rect 28532 3500 28542 3556
rect 32386 3500 32396 3556
rect 32452 3500 32462 3556
rect 34514 3500 34524 3556
rect 34580 3500 40572 3556
rect 40628 3500 40638 3556
rect 42242 3500 42252 3556
rect 42308 3500 45276 3556
rect 45332 3500 45342 3556
rect 49522 3500 49532 3556
rect 49588 3500 50428 3556
rect 50866 3500 50876 3556
rect 50932 3500 52332 3556
rect 52388 3500 52398 3556
rect 53004 3500 54236 3556
rect 54292 3500 54302 3556
rect 55346 3500 55356 3556
rect 55412 3500 59108 3556
rect 65426 3500 65436 3556
rect 65492 3500 68908 3556
rect 68964 3500 68974 3556
rect 0 3444 800 3472
rect 1820 3444 1876 3500
rect 8204 3444 8260 3500
rect 32396 3444 32452 3500
rect 71260 3444 71316 3612
rect 0 3388 1876 3444
rect 3938 3388 3948 3444
rect 4004 3388 4172 3444
rect 4228 3388 7532 3444
rect 7588 3388 7598 3444
rect 8204 3388 11004 3444
rect 11060 3388 11070 3444
rect 12562 3388 12572 3444
rect 12628 3388 21644 3444
rect 21700 3388 21710 3444
rect 22642 3388 22652 3444
rect 22708 3388 28700 3444
rect 28756 3388 28766 3444
rect 32396 3388 38556 3444
rect 38612 3388 38622 3444
rect 43026 3388 43036 3444
rect 43092 3388 45388 3444
rect 45444 3388 45454 3444
rect 49970 3388 49980 3444
rect 50036 3388 51212 3444
rect 51268 3388 51660 3444
rect 51716 3388 51726 3444
rect 51874 3388 51884 3444
rect 51940 3388 52780 3444
rect 52836 3388 52846 3444
rect 54674 3388 54684 3444
rect 54740 3388 57596 3444
rect 57652 3388 57662 3444
rect 58034 3388 58044 3444
rect 58100 3388 63868 3444
rect 63924 3388 63934 3444
rect 64754 3388 64764 3444
rect 64820 3388 71316 3444
rect 73602 3388 73612 3444
rect 73668 3388 74844 3444
rect 74900 3388 74910 3444
rect 0 3360 800 3388
rect 6738 3276 6748 3332
rect 6804 3276 8428 3332
rect 9986 3276 9996 3332
rect 10052 3276 15372 3332
rect 15428 3276 15438 3332
rect 18834 3276 18844 3332
rect 18900 3276 27356 3332
rect 27412 3276 27422 3332
rect 30930 3276 30940 3332
rect 30996 3276 38668 3332
rect 38724 3276 38734 3332
rect 8372 2772 8428 3276
rect 8754 3164 8764 3220
rect 8820 3164 17388 3220
rect 17444 3164 17454 3220
rect 22306 3164 22316 3220
rect 22372 3164 23324 3220
rect 23380 3164 23390 3220
rect 26852 3164 30604 3220
rect 30660 3164 30670 3220
rect 35074 3164 35084 3220
rect 35140 3164 42476 3220
rect 42532 3164 42542 3220
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 26852 3108 26908 3164
rect 50546 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50830 3164
rect 10434 3052 10444 3108
rect 10500 3052 15708 3108
rect 15764 3052 15774 3108
rect 24098 3052 24108 3108
rect 24164 3052 26908 3108
rect 28914 3052 28924 3108
rect 28980 3052 37436 3108
rect 37492 3052 37502 3108
rect 79200 2996 80000 3024
rect 11890 2940 11900 2996
rect 11956 2940 22204 2996
rect 22260 2940 22270 2996
rect 27794 2940 27804 2996
rect 27860 2940 36988 2996
rect 37044 2940 37054 2996
rect 74050 2940 74060 2996
rect 74116 2940 80000 2996
rect 79200 2912 80000 2940
rect 9874 2828 9884 2884
rect 9940 2828 23212 2884
rect 23268 2828 23278 2884
rect 23436 2828 26236 2884
rect 26292 2828 26302 2884
rect 33058 2828 33068 2884
rect 33124 2828 39228 2884
rect 39284 2828 39294 2884
rect 23436 2772 23492 2828
rect 8372 2716 15260 2772
rect 15316 2716 15326 2772
rect 16370 2716 16380 2772
rect 16436 2716 23492 2772
rect 24658 2716 24668 2772
rect 24724 2716 33516 2772
rect 33572 2716 33582 2772
rect 7074 2604 7084 2660
rect 7140 2604 12348 2660
rect 12404 2604 12414 2660
rect 23314 2604 23324 2660
rect 23380 2604 29148 2660
rect 29204 2604 29214 2660
rect 7746 2492 7756 2548
rect 7812 2492 13020 2548
rect 13076 2492 13086 2548
rect 10546 2380 10556 2436
rect 10612 2380 20860 2436
rect 20916 2380 20926 2436
rect 23426 2380 23436 2436
rect 23492 2380 35980 2436
rect 36036 2380 36046 2436
rect 0 2324 800 2352
rect 0 2268 2380 2324
rect 2436 2268 2446 2324
rect 8082 2268 8092 2324
rect 8148 2268 17276 2324
rect 17332 2268 17342 2324
rect 27570 2268 27580 2324
rect 27636 2268 34524 2324
rect 34580 2268 34590 2324
rect 0 2240 800 2268
rect 30594 2156 30604 2212
rect 30660 2156 37212 2212
rect 37268 2156 37278 2212
rect 79200 1876 80000 1904
rect 29250 1820 29260 1876
rect 29316 1820 35868 1876
rect 35924 1820 35934 1876
rect 75506 1820 75516 1876
rect 75572 1820 80000 1876
rect 79200 1792 80000 1820
rect 31490 1708 31500 1764
rect 31556 1708 37884 1764
rect 37940 1708 37950 1764
rect 21298 1596 21308 1652
rect 21364 1596 38892 1652
rect 38948 1596 38958 1652
rect 31602 1484 31612 1540
rect 31668 1484 39004 1540
rect 39060 1484 39070 1540
rect 22754 1372 22764 1428
rect 22820 1372 33628 1428
rect 33684 1372 33694 1428
rect 74610 924 74620 980
rect 74676 924 74686 980
rect 74620 756 74676 924
rect 79200 756 80000 784
rect 74620 700 80000 756
rect 79200 672 80000 700
<< via3 >>
rect 19836 76804 19892 76860
rect 19940 76804 19996 76860
rect 20044 76804 20100 76860
rect 50556 76804 50612 76860
rect 50660 76804 50716 76860
rect 50764 76804 50820 76860
rect 76076 76524 76132 76580
rect 47068 76300 47124 76356
rect 4476 76020 4532 76076
rect 4580 76020 4636 76076
rect 4684 76020 4740 76076
rect 35196 76020 35252 76076
rect 35300 76020 35356 76076
rect 35404 76020 35460 76076
rect 65916 76020 65972 76076
rect 66020 76020 66076 76076
rect 66124 76020 66180 76076
rect 19836 75236 19892 75292
rect 19940 75236 19996 75292
rect 20044 75236 20100 75292
rect 50556 75236 50612 75292
rect 50660 75236 50716 75292
rect 50764 75236 50820 75292
rect 4476 74452 4532 74508
rect 4580 74452 4636 74508
rect 4684 74452 4740 74508
rect 35196 74452 35252 74508
rect 35300 74452 35356 74508
rect 35404 74452 35460 74508
rect 65916 74452 65972 74508
rect 66020 74452 66076 74508
rect 66124 74452 66180 74508
rect 19836 73668 19892 73724
rect 19940 73668 19996 73724
rect 20044 73668 20100 73724
rect 50556 73668 50612 73724
rect 50660 73668 50716 73724
rect 50764 73668 50820 73724
rect 4476 72884 4532 72940
rect 4580 72884 4636 72940
rect 4684 72884 4740 72940
rect 35196 72884 35252 72940
rect 35300 72884 35356 72940
rect 35404 72884 35460 72940
rect 65916 72884 65972 72940
rect 66020 72884 66076 72940
rect 66124 72884 66180 72940
rect 19836 72100 19892 72156
rect 19940 72100 19996 72156
rect 20044 72100 20100 72156
rect 50556 72100 50612 72156
rect 50660 72100 50716 72156
rect 50764 72100 50820 72156
rect 4476 71316 4532 71372
rect 4580 71316 4636 71372
rect 4684 71316 4740 71372
rect 35196 71316 35252 71372
rect 35300 71316 35356 71372
rect 35404 71316 35460 71372
rect 65916 71316 65972 71372
rect 66020 71316 66076 71372
rect 66124 71316 66180 71372
rect 19836 70532 19892 70588
rect 19940 70532 19996 70588
rect 20044 70532 20100 70588
rect 50556 70532 50612 70588
rect 50660 70532 50716 70588
rect 50764 70532 50820 70588
rect 4476 69748 4532 69804
rect 4580 69748 4636 69804
rect 4684 69748 4740 69804
rect 35196 69748 35252 69804
rect 35300 69748 35356 69804
rect 35404 69748 35460 69804
rect 65916 69748 65972 69804
rect 66020 69748 66076 69804
rect 66124 69748 66180 69804
rect 19836 68964 19892 69020
rect 19940 68964 19996 69020
rect 20044 68964 20100 69020
rect 50556 68964 50612 69020
rect 50660 68964 50716 69020
rect 50764 68964 50820 69020
rect 4476 68180 4532 68236
rect 4580 68180 4636 68236
rect 4684 68180 4740 68236
rect 35196 68180 35252 68236
rect 35300 68180 35356 68236
rect 35404 68180 35460 68236
rect 65916 68180 65972 68236
rect 66020 68180 66076 68236
rect 66124 68180 66180 68236
rect 76300 67788 76356 67844
rect 19836 67396 19892 67452
rect 19940 67396 19996 67452
rect 20044 67396 20100 67452
rect 50556 67396 50612 67452
rect 50660 67396 50716 67452
rect 50764 67396 50820 67452
rect 75852 67116 75908 67172
rect 4476 66612 4532 66668
rect 4580 66612 4636 66668
rect 4684 66612 4740 66668
rect 35196 66612 35252 66668
rect 35300 66612 35356 66668
rect 35404 66612 35460 66668
rect 65916 66612 65972 66668
rect 66020 66612 66076 66668
rect 66124 66612 66180 66668
rect 19836 65828 19892 65884
rect 19940 65828 19996 65884
rect 20044 65828 20100 65884
rect 50556 65828 50612 65884
rect 50660 65828 50716 65884
rect 50764 65828 50820 65884
rect 4476 65044 4532 65100
rect 4580 65044 4636 65100
rect 4684 65044 4740 65100
rect 35196 65044 35252 65100
rect 35300 65044 35356 65100
rect 35404 65044 35460 65100
rect 65916 65044 65972 65100
rect 66020 65044 66076 65100
rect 66124 65044 66180 65100
rect 19836 64260 19892 64316
rect 19940 64260 19996 64316
rect 20044 64260 20100 64316
rect 50556 64260 50612 64316
rect 50660 64260 50716 64316
rect 50764 64260 50820 64316
rect 4476 63476 4532 63532
rect 4580 63476 4636 63532
rect 4684 63476 4740 63532
rect 35196 63476 35252 63532
rect 35300 63476 35356 63532
rect 35404 63476 35460 63532
rect 65916 63476 65972 63532
rect 66020 63476 66076 63532
rect 66124 63476 66180 63532
rect 19836 62692 19892 62748
rect 19940 62692 19996 62748
rect 20044 62692 20100 62748
rect 50556 62692 50612 62748
rect 50660 62692 50716 62748
rect 50764 62692 50820 62748
rect 76412 62188 76468 62244
rect 4476 61908 4532 61964
rect 4580 61908 4636 61964
rect 4684 61908 4740 61964
rect 35196 61908 35252 61964
rect 35300 61908 35356 61964
rect 35404 61908 35460 61964
rect 65916 61908 65972 61964
rect 66020 61908 66076 61964
rect 66124 61908 66180 61964
rect 76972 61292 77028 61348
rect 19836 61124 19892 61180
rect 19940 61124 19996 61180
rect 20044 61124 20100 61180
rect 50556 61124 50612 61180
rect 50660 61124 50716 61180
rect 50764 61124 50820 61180
rect 4476 60340 4532 60396
rect 4580 60340 4636 60396
rect 4684 60340 4740 60396
rect 35196 60340 35252 60396
rect 35300 60340 35356 60396
rect 35404 60340 35460 60396
rect 65916 60340 65972 60396
rect 66020 60340 66076 60396
rect 66124 60340 66180 60396
rect 19836 59556 19892 59612
rect 19940 59556 19996 59612
rect 20044 59556 20100 59612
rect 50556 59556 50612 59612
rect 50660 59556 50716 59612
rect 50764 59556 50820 59612
rect 4476 58772 4532 58828
rect 4580 58772 4636 58828
rect 4684 58772 4740 58828
rect 35196 58772 35252 58828
rect 35300 58772 35356 58828
rect 35404 58772 35460 58828
rect 65916 58772 65972 58828
rect 66020 58772 66076 58828
rect 66124 58772 66180 58828
rect 19836 57988 19892 58044
rect 19940 57988 19996 58044
rect 20044 57988 20100 58044
rect 50556 57988 50612 58044
rect 50660 57988 50716 58044
rect 50764 57988 50820 58044
rect 4476 57204 4532 57260
rect 4580 57204 4636 57260
rect 4684 57204 4740 57260
rect 35196 57204 35252 57260
rect 35300 57204 35356 57260
rect 35404 57204 35460 57260
rect 65916 57204 65972 57260
rect 66020 57204 66076 57260
rect 66124 57204 66180 57260
rect 74060 56588 74116 56644
rect 19836 56420 19892 56476
rect 19940 56420 19996 56476
rect 20044 56420 20100 56476
rect 50556 56420 50612 56476
rect 50660 56420 50716 56476
rect 50764 56420 50820 56476
rect 4476 55636 4532 55692
rect 4580 55636 4636 55692
rect 4684 55636 4740 55692
rect 35196 55636 35252 55692
rect 35300 55636 35356 55692
rect 35404 55636 35460 55692
rect 65916 55636 65972 55692
rect 66020 55636 66076 55692
rect 66124 55636 66180 55692
rect 19836 54852 19892 54908
rect 19940 54852 19996 54908
rect 20044 54852 20100 54908
rect 50556 54852 50612 54908
rect 50660 54852 50716 54908
rect 50764 54852 50820 54908
rect 4476 54068 4532 54124
rect 4580 54068 4636 54124
rect 4684 54068 4740 54124
rect 35196 54068 35252 54124
rect 35300 54068 35356 54124
rect 35404 54068 35460 54124
rect 65916 54068 65972 54124
rect 66020 54068 66076 54124
rect 66124 54068 66180 54124
rect 19836 53284 19892 53340
rect 19940 53284 19996 53340
rect 20044 53284 20100 53340
rect 50556 53284 50612 53340
rect 50660 53284 50716 53340
rect 50764 53284 50820 53340
rect 4476 52500 4532 52556
rect 4580 52500 4636 52556
rect 4684 52500 4740 52556
rect 35196 52500 35252 52556
rect 35300 52500 35356 52556
rect 35404 52500 35460 52556
rect 65916 52500 65972 52556
rect 66020 52500 66076 52556
rect 66124 52500 66180 52556
rect 19836 51716 19892 51772
rect 19940 51716 19996 51772
rect 20044 51716 20100 51772
rect 50556 51716 50612 51772
rect 50660 51716 50716 51772
rect 50764 51716 50820 51772
rect 4476 50932 4532 50988
rect 4580 50932 4636 50988
rect 4684 50932 4740 50988
rect 35196 50932 35252 50988
rect 35300 50932 35356 50988
rect 35404 50932 35460 50988
rect 65916 50932 65972 50988
rect 66020 50932 66076 50988
rect 66124 50932 66180 50988
rect 19836 50148 19892 50204
rect 19940 50148 19996 50204
rect 20044 50148 20100 50204
rect 50556 50148 50612 50204
rect 50660 50148 50716 50204
rect 50764 50148 50820 50204
rect 4476 49364 4532 49420
rect 4580 49364 4636 49420
rect 4684 49364 4740 49420
rect 35196 49364 35252 49420
rect 35300 49364 35356 49420
rect 35404 49364 35460 49420
rect 65916 49364 65972 49420
rect 66020 49364 66076 49420
rect 66124 49364 66180 49420
rect 19836 48580 19892 48636
rect 19940 48580 19996 48636
rect 20044 48580 20100 48636
rect 50556 48580 50612 48636
rect 50660 48580 50716 48636
rect 50764 48580 50820 48636
rect 4476 47796 4532 47852
rect 4580 47796 4636 47852
rect 4684 47796 4740 47852
rect 35196 47796 35252 47852
rect 35300 47796 35356 47852
rect 35404 47796 35460 47852
rect 65916 47796 65972 47852
rect 66020 47796 66076 47852
rect 66124 47796 66180 47852
rect 19836 47012 19892 47068
rect 19940 47012 19996 47068
rect 20044 47012 20100 47068
rect 50556 47012 50612 47068
rect 50660 47012 50716 47068
rect 50764 47012 50820 47068
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 65916 46228 65972 46284
rect 66020 46228 66076 46284
rect 66124 46228 66180 46284
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 50556 45444 50612 45500
rect 50660 45444 50716 45500
rect 50764 45444 50820 45500
rect 72604 45052 72660 45108
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 65916 44660 65972 44716
rect 66020 44660 66076 44716
rect 66124 44660 66180 44716
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 50556 43876 50612 43932
rect 50660 43876 50716 43932
rect 50764 43876 50820 43932
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 65916 43092 65972 43148
rect 66020 43092 66076 43148
rect 66124 43092 66180 43148
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 50556 42308 50612 42364
rect 50660 42308 50716 42364
rect 50764 42308 50820 42364
rect 65772 42140 65828 42196
rect 76188 41916 76244 41972
rect 74620 41580 74676 41636
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 65916 41524 65972 41580
rect 66020 41524 66076 41580
rect 66124 41524 66180 41580
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 50556 40740 50612 40796
rect 50660 40740 50716 40796
rect 50764 40740 50820 40796
rect 75068 40572 75124 40628
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 65916 39956 65972 40012
rect 66020 39956 66076 40012
rect 66124 39956 66180 40012
rect 72828 39564 72884 39620
rect 65772 39452 65828 39508
rect 75068 39340 75124 39396
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 50556 39172 50612 39228
rect 50660 39172 50716 39228
rect 50764 39172 50820 39228
rect 72716 39116 72772 39172
rect 73724 38780 73780 38836
rect 75068 38780 75124 38836
rect 72828 38556 72884 38612
rect 73388 38556 73444 38612
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 65916 38388 65972 38444
rect 66020 38388 66076 38444
rect 66124 38388 66180 38444
rect 76188 38220 76244 38276
rect 72604 38108 72660 38164
rect 72940 38108 72996 38164
rect 73948 37660 74004 37716
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 50556 37604 50612 37660
rect 50660 37604 50716 37660
rect 50764 37604 50820 37660
rect 74396 37436 74452 37492
rect 73388 37324 73444 37380
rect 73724 37212 73780 37268
rect 75964 37212 76020 37268
rect 76636 37212 76692 37268
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 65916 36820 65972 36876
rect 66020 36820 66076 36876
rect 66124 36820 66180 36876
rect 72940 36764 72996 36820
rect 73276 36316 73332 36372
rect 73948 36316 74004 36372
rect 74396 36316 74452 36372
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 50556 36036 50612 36092
rect 50660 36036 50716 36092
rect 50764 36036 50820 36092
rect 77868 35868 77924 35924
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 65916 35252 65972 35308
rect 66020 35252 66076 35308
rect 66124 35252 66180 35308
rect 72268 35196 72324 35252
rect 72716 35196 72772 35252
rect 72940 35084 72996 35140
rect 77868 35084 77924 35140
rect 74956 34860 75012 34916
rect 70812 34636 70868 34692
rect 72380 34636 72436 34692
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 50556 34468 50612 34524
rect 50660 34468 50716 34524
rect 50764 34468 50820 34524
rect 75964 34300 76020 34356
rect 76188 34300 76244 34356
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 65916 33684 65972 33740
rect 66020 33684 66076 33740
rect 66124 33684 66180 33740
rect 76636 33404 76692 33460
rect 72604 33292 72660 33348
rect 72940 33292 72996 33348
rect 77084 33180 77140 33236
rect 75628 33068 75684 33124
rect 74508 32956 74564 33012
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 50556 32900 50612 32956
rect 50660 32900 50716 32956
rect 50764 32900 50820 32956
rect 72380 32620 72436 32676
rect 71596 32396 71652 32452
rect 72604 32396 72660 32452
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 65916 32116 65972 32172
rect 66020 32116 66076 32172
rect 66124 32116 66180 32172
rect 77084 31948 77140 32004
rect 72380 31836 72436 31892
rect 75068 31724 75124 31780
rect 76300 31724 76356 31780
rect 72492 31388 72548 31444
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 50556 31332 50612 31388
rect 50660 31332 50716 31388
rect 50764 31332 50820 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 65916 30548 65972 30604
rect 66020 30548 66076 30604
rect 66124 30548 66180 30604
rect 71820 30492 71876 30548
rect 76860 30156 76916 30212
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 50556 29764 50612 29820
rect 50660 29764 50716 29820
rect 50764 29764 50820 29820
rect 49756 29372 49812 29428
rect 72268 29372 72324 29428
rect 75852 29372 75908 29428
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 65916 28980 65972 29036
rect 66020 28980 66076 29036
rect 66124 28980 66180 29036
rect 72716 28924 72772 28980
rect 76860 28588 76916 28644
rect 72380 28476 72436 28532
rect 76524 28476 76580 28532
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 50556 28196 50612 28252
rect 50660 28196 50716 28252
rect 50764 28196 50820 28252
rect 40124 27804 40180 27860
rect 75628 27916 75684 27972
rect 71932 27804 71988 27860
rect 72268 27692 72324 27748
rect 73724 27692 73780 27748
rect 40124 27580 40180 27636
rect 74060 27580 74116 27636
rect 76972 27580 77028 27636
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 65916 27412 65972 27468
rect 66020 27412 66076 27468
rect 66124 27412 66180 27468
rect 71932 27244 71988 27300
rect 74060 27020 74116 27076
rect 74956 26796 75012 26852
rect 72716 26684 72772 26740
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 50556 26628 50612 26684
rect 50660 26628 50716 26684
rect 50764 26628 50820 26684
rect 75852 26460 75908 26516
rect 73836 26236 73892 26292
rect 49756 26124 49812 26180
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 65916 25844 65972 25900
rect 66020 25844 66076 25900
rect 66124 25844 66180 25900
rect 72604 25676 72660 25732
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 50556 25060 50612 25116
rect 50660 25060 50716 25116
rect 50764 25060 50820 25116
rect 71820 25004 71876 25060
rect 72268 25004 72324 25060
rect 75628 25004 75684 25060
rect 76524 24668 76580 24724
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 65916 24276 65972 24332
rect 66020 24276 66076 24332
rect 66124 24276 66180 24332
rect 70812 23996 70868 24052
rect 73276 23884 73332 23940
rect 74508 23884 74564 23940
rect 71596 23772 71652 23828
rect 49308 23660 49364 23716
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 50556 23492 50612 23548
rect 50660 23492 50716 23548
rect 50764 23492 50820 23548
rect 49532 23324 49588 23380
rect 46844 22876 46900 22932
rect 47628 22876 47684 22932
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 65916 22708 65972 22764
rect 66020 22708 66076 22764
rect 66124 22708 66180 22764
rect 34860 22316 34916 22372
rect 42028 22316 42084 22372
rect 47180 22316 47236 22372
rect 49420 22316 49476 22372
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 50556 21924 50612 21980
rect 50660 21924 50716 21980
rect 50764 21924 50820 21980
rect 77644 21868 77700 21924
rect 47628 21644 47684 21700
rect 77756 21644 77812 21700
rect 47180 21532 47236 21588
rect 49532 21532 49588 21588
rect 75404 21532 75460 21588
rect 34860 21420 34916 21476
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 65916 21140 65972 21196
rect 66020 21140 66076 21196
rect 66124 21140 66180 21196
rect 32956 20524 33012 20580
rect 40684 20524 40740 20580
rect 38444 20412 38500 20468
rect 38668 20412 38724 20468
rect 76412 20412 76468 20468
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 50556 20356 50612 20412
rect 50660 20356 50716 20412
rect 50764 20356 50820 20412
rect 48972 20300 49028 20356
rect 32956 19964 33012 20020
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 49308 19964 49364 20020
rect 76412 19964 76468 20020
rect 77644 19852 77700 19908
rect 65916 19572 65972 19628
rect 66020 19572 66076 19628
rect 66124 19572 66180 19628
rect 48972 19180 49028 19236
rect 39788 19068 39844 19124
rect 75404 18956 75460 19012
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 50556 18788 50612 18844
rect 50660 18788 50716 18844
rect 50764 18788 50820 18844
rect 49420 18508 49476 18564
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 65916 18004 65972 18060
rect 66020 18004 66076 18060
rect 66124 18004 66180 18060
rect 39340 17612 39396 17668
rect 40012 17612 40068 17668
rect 40684 17612 40740 17668
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 50556 17220 50612 17276
rect 50660 17220 50716 17276
rect 50764 17220 50820 17276
rect 40012 16828 40068 16884
rect 47068 16828 47124 16884
rect 39788 16716 39844 16772
rect 77756 16716 77812 16772
rect 43708 16604 43764 16660
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 65916 16436 65972 16492
rect 66020 16436 66076 16492
rect 66124 16436 66180 16492
rect 39340 16268 39396 16324
rect 43708 16044 43764 16100
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 50556 15652 50612 15708
rect 50660 15652 50716 15708
rect 50764 15652 50820 15708
rect 20188 15596 20244 15652
rect 20188 15260 20244 15316
rect 46844 15260 46900 15316
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 65916 14868 65972 14924
rect 66020 14868 66076 14924
rect 66124 14868 66180 14924
rect 74620 14700 74676 14756
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 50556 14084 50612 14140
rect 50660 14084 50716 14140
rect 50764 14084 50820 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 65916 13300 65972 13356
rect 66020 13300 66076 13356
rect 66124 13300 66180 13356
rect 32956 13132 33012 13188
rect 42028 12796 42084 12852
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 50556 12516 50612 12572
rect 50660 12516 50716 12572
rect 50764 12516 50820 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 65916 11732 65972 11788
rect 66020 11732 66076 11788
rect 66124 11732 66180 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 50556 10948 50612 11004
rect 50660 10948 50716 11004
rect 50764 10948 50820 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 65916 10164 65972 10220
rect 66020 10164 66076 10220
rect 66124 10164 66180 10220
rect 31724 10108 31780 10164
rect 38220 9996 38276 10052
rect 38220 9772 38276 9828
rect 31724 9660 31780 9716
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 50556 9380 50612 9436
rect 50660 9380 50716 9436
rect 50764 9380 50820 9436
rect 18732 9324 18788 9380
rect 19628 9212 19684 9268
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 65916 8596 65972 8652
rect 66020 8596 66076 8652
rect 66124 8596 66180 8652
rect 19628 8204 19684 8260
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 50556 7812 50612 7868
rect 50660 7812 50716 7868
rect 50764 7812 50820 7868
rect 28588 7420 28644 7476
rect 33180 7420 33236 7476
rect 30940 7308 30996 7364
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 13916 6972 13972 7028
rect 65916 7028 65972 7084
rect 66020 7028 66076 7084
rect 66124 7028 66180 7084
rect 30828 6860 30884 6916
rect 28588 6636 28644 6692
rect 31500 6748 31556 6804
rect 15148 6524 15204 6580
rect 33180 6524 33236 6580
rect 18620 6412 18676 6468
rect 30828 6300 30884 6356
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 50556 6244 50612 6300
rect 50660 6244 50716 6300
rect 50764 6244 50820 6300
rect 31500 6188 31556 6244
rect 15148 6076 15204 6132
rect 18732 6076 18788 6132
rect 9996 5516 10052 5572
rect 13916 5516 13972 5572
rect 14364 5516 14420 5572
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 65916 5460 65972 5516
rect 66020 5460 66076 5516
rect 66124 5460 66180 5516
rect 18732 5180 18788 5236
rect 14364 4732 14420 4788
rect 30940 4732 30996 4788
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 50556 4676 50612 4732
rect 50660 4676 50716 4732
rect 50764 4676 50820 4732
rect 33180 4284 33236 4340
rect 18620 4060 18676 4116
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 65916 3892 65972 3948
rect 66020 3892 66076 3948
rect 66124 3892 66180 3948
rect 9996 3836 10052 3892
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
rect 50556 3108 50612 3164
rect 50660 3108 50716 3164
rect 50764 3108 50820 3164
<< metal4 >>
rect 4448 76076 4768 76892
rect 4448 76020 4476 76076
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4740 76020 4768 76076
rect 4448 74508 4768 76020
rect 4448 74452 4476 74508
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4740 74452 4768 74508
rect 4448 72940 4768 74452
rect 4448 72884 4476 72940
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4740 72884 4768 72940
rect 4448 71372 4768 72884
rect 4448 71316 4476 71372
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4740 71316 4768 71372
rect 4448 69804 4768 71316
rect 4448 69748 4476 69804
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4740 69748 4768 69804
rect 4448 68236 4768 69748
rect 4448 68180 4476 68236
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4740 68180 4768 68236
rect 4448 66668 4768 68180
rect 4448 66612 4476 66668
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4740 66612 4768 66668
rect 4448 65100 4768 66612
rect 4448 65044 4476 65100
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4740 65044 4768 65100
rect 4448 63532 4768 65044
rect 4448 63476 4476 63532
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4740 63476 4768 63532
rect 4448 61964 4768 63476
rect 4448 61908 4476 61964
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4740 61908 4768 61964
rect 4448 60396 4768 61908
rect 4448 60340 4476 60396
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4740 60340 4768 60396
rect 4448 58828 4768 60340
rect 4448 58772 4476 58828
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4740 58772 4768 58828
rect 4448 57260 4768 58772
rect 4448 57204 4476 57260
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4740 57204 4768 57260
rect 4448 55692 4768 57204
rect 4448 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4768 55692
rect 4448 54124 4768 55636
rect 4448 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4768 54124
rect 4448 52556 4768 54068
rect 4448 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4768 52556
rect 4448 50988 4768 52500
rect 4448 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4768 50988
rect 4448 49420 4768 50932
rect 4448 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4768 49420
rect 4448 47852 4768 49364
rect 4448 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4768 47852
rect 4448 46284 4768 47796
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 19808 76860 20128 76892
rect 19808 76804 19836 76860
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 20100 76804 20128 76860
rect 19808 75292 20128 76804
rect 19808 75236 19836 75292
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 20100 75236 20128 75292
rect 19808 73724 20128 75236
rect 19808 73668 19836 73724
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 20100 73668 20128 73724
rect 19808 72156 20128 73668
rect 19808 72100 19836 72156
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 20100 72100 20128 72156
rect 19808 70588 20128 72100
rect 19808 70532 19836 70588
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 20100 70532 20128 70588
rect 19808 69020 20128 70532
rect 19808 68964 19836 69020
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 20100 68964 20128 69020
rect 19808 67452 20128 68964
rect 19808 67396 19836 67452
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 20100 67396 20128 67452
rect 19808 65884 20128 67396
rect 19808 65828 19836 65884
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 20100 65828 20128 65884
rect 19808 64316 20128 65828
rect 19808 64260 19836 64316
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 20100 64260 20128 64316
rect 19808 62748 20128 64260
rect 19808 62692 19836 62748
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 20100 62692 20128 62748
rect 19808 61180 20128 62692
rect 19808 61124 19836 61180
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 20100 61124 20128 61180
rect 19808 59612 20128 61124
rect 19808 59556 19836 59612
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 20100 59556 20128 59612
rect 19808 58044 20128 59556
rect 19808 57988 19836 58044
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 20100 57988 20128 58044
rect 19808 56476 20128 57988
rect 19808 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20128 56476
rect 19808 54908 20128 56420
rect 19808 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20128 54908
rect 19808 53340 20128 54852
rect 19808 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20128 53340
rect 19808 51772 20128 53284
rect 19808 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20128 51772
rect 19808 50204 20128 51716
rect 19808 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20128 50204
rect 19808 48636 20128 50148
rect 19808 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20128 48636
rect 19808 47068 20128 48580
rect 19808 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20128 47068
rect 19808 45500 20128 47012
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 19808 43932 20128 45444
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 19808 42364 20128 43876
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 35168 76076 35488 76892
rect 50528 76860 50848 76892
rect 50528 76804 50556 76860
rect 50612 76804 50660 76860
rect 50716 76804 50764 76860
rect 50820 76804 50848 76860
rect 35168 76020 35196 76076
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35460 76020 35488 76076
rect 35168 74508 35488 76020
rect 35168 74452 35196 74508
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35460 74452 35488 74508
rect 35168 72940 35488 74452
rect 35168 72884 35196 72940
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35460 72884 35488 72940
rect 35168 71372 35488 72884
rect 35168 71316 35196 71372
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35460 71316 35488 71372
rect 35168 69804 35488 71316
rect 35168 69748 35196 69804
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35460 69748 35488 69804
rect 35168 68236 35488 69748
rect 35168 68180 35196 68236
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35460 68180 35488 68236
rect 35168 66668 35488 68180
rect 35168 66612 35196 66668
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35460 66612 35488 66668
rect 35168 65100 35488 66612
rect 35168 65044 35196 65100
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35460 65044 35488 65100
rect 35168 63532 35488 65044
rect 35168 63476 35196 63532
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35460 63476 35488 63532
rect 35168 61964 35488 63476
rect 35168 61908 35196 61964
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35460 61908 35488 61964
rect 35168 60396 35488 61908
rect 35168 60340 35196 60396
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35460 60340 35488 60396
rect 35168 58828 35488 60340
rect 35168 58772 35196 58828
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35460 58772 35488 58828
rect 35168 57260 35488 58772
rect 35168 57204 35196 57260
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35460 57204 35488 57260
rect 35168 55692 35488 57204
rect 35168 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35488 55692
rect 35168 54124 35488 55636
rect 35168 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35488 54124
rect 35168 52556 35488 54068
rect 35168 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35488 52556
rect 35168 50988 35488 52500
rect 35168 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35488 50988
rect 35168 49420 35488 50932
rect 35168 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35488 49420
rect 35168 47852 35488 49364
rect 35168 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35488 47852
rect 35168 46284 35488 47796
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 47068 76356 47124 76366
rect 40124 27860 40180 27870
rect 40124 27636 40180 27804
rect 40124 27570 40180 27580
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 34860 22372 34916 22382
rect 34860 21476 34916 22316
rect 34860 21410 34916 21420
rect 35168 21196 35488 22708
rect 46844 22932 46900 22942
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 32956 20580 33012 20590
rect 32956 20020 33012 20524
rect 19808 14140 20128 15652
rect 20188 15652 20244 15662
rect 20188 15316 20244 15596
rect 20188 15250 20244 15260
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 32956 13188 33012 19964
rect 32956 13122 33012 13132
rect 35168 19628 35488 21140
rect 42028 22372 42084 22382
rect 40684 20580 40740 20590
rect 38444 20468 38500 20478
rect 38668 20468 38724 20478
rect 38500 20412 38668 20458
rect 38444 20402 38724 20412
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 39788 19124 39844 19134
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 39340 17668 39396 17678
rect 39340 16324 39396 17612
rect 39788 16772 39844 19068
rect 40012 17668 40068 17678
rect 40012 16884 40068 17612
rect 40684 17668 40740 20524
rect 40684 17602 40740 17612
rect 40012 16818 40068 16828
rect 39788 16706 39844 16716
rect 39340 16258 39396 16268
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 35168 11788 35488 13300
rect 42028 12852 42084 22316
rect 43708 16660 43764 16670
rect 43708 16100 43764 16604
rect 43708 16034 43764 16044
rect 46844 15316 46900 22876
rect 47068 16884 47124 76300
rect 50528 75292 50848 76804
rect 50528 75236 50556 75292
rect 50612 75236 50660 75292
rect 50716 75236 50764 75292
rect 50820 75236 50848 75292
rect 50528 73724 50848 75236
rect 50528 73668 50556 73724
rect 50612 73668 50660 73724
rect 50716 73668 50764 73724
rect 50820 73668 50848 73724
rect 50528 72156 50848 73668
rect 50528 72100 50556 72156
rect 50612 72100 50660 72156
rect 50716 72100 50764 72156
rect 50820 72100 50848 72156
rect 50528 70588 50848 72100
rect 50528 70532 50556 70588
rect 50612 70532 50660 70588
rect 50716 70532 50764 70588
rect 50820 70532 50848 70588
rect 50528 69020 50848 70532
rect 50528 68964 50556 69020
rect 50612 68964 50660 69020
rect 50716 68964 50764 69020
rect 50820 68964 50848 69020
rect 50528 67452 50848 68964
rect 50528 67396 50556 67452
rect 50612 67396 50660 67452
rect 50716 67396 50764 67452
rect 50820 67396 50848 67452
rect 50528 65884 50848 67396
rect 50528 65828 50556 65884
rect 50612 65828 50660 65884
rect 50716 65828 50764 65884
rect 50820 65828 50848 65884
rect 50528 64316 50848 65828
rect 50528 64260 50556 64316
rect 50612 64260 50660 64316
rect 50716 64260 50764 64316
rect 50820 64260 50848 64316
rect 50528 62748 50848 64260
rect 50528 62692 50556 62748
rect 50612 62692 50660 62748
rect 50716 62692 50764 62748
rect 50820 62692 50848 62748
rect 50528 61180 50848 62692
rect 50528 61124 50556 61180
rect 50612 61124 50660 61180
rect 50716 61124 50764 61180
rect 50820 61124 50848 61180
rect 50528 59612 50848 61124
rect 50528 59556 50556 59612
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50820 59556 50848 59612
rect 50528 58044 50848 59556
rect 50528 57988 50556 58044
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50820 57988 50848 58044
rect 50528 56476 50848 57988
rect 50528 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50848 56476
rect 50528 54908 50848 56420
rect 50528 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50848 54908
rect 50528 53340 50848 54852
rect 50528 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50848 53340
rect 50528 51772 50848 53284
rect 50528 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50848 51772
rect 50528 50204 50848 51716
rect 50528 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50848 50204
rect 50528 48636 50848 50148
rect 50528 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50848 48636
rect 50528 47068 50848 48580
rect 50528 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50848 47068
rect 50528 45500 50848 47012
rect 50528 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50848 45500
rect 50528 43932 50848 45444
rect 50528 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50848 43932
rect 50528 42364 50848 43876
rect 50528 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50848 42364
rect 50528 40796 50848 42308
rect 65888 76076 66208 76892
rect 65888 76020 65916 76076
rect 65972 76020 66020 76076
rect 66076 76020 66124 76076
rect 66180 76020 66208 76076
rect 65888 74508 66208 76020
rect 65888 74452 65916 74508
rect 65972 74452 66020 74508
rect 66076 74452 66124 74508
rect 66180 74452 66208 74508
rect 65888 72940 66208 74452
rect 65888 72884 65916 72940
rect 65972 72884 66020 72940
rect 66076 72884 66124 72940
rect 66180 72884 66208 72940
rect 65888 71372 66208 72884
rect 65888 71316 65916 71372
rect 65972 71316 66020 71372
rect 66076 71316 66124 71372
rect 66180 71316 66208 71372
rect 65888 69804 66208 71316
rect 65888 69748 65916 69804
rect 65972 69748 66020 69804
rect 66076 69748 66124 69804
rect 66180 69748 66208 69804
rect 65888 68236 66208 69748
rect 65888 68180 65916 68236
rect 65972 68180 66020 68236
rect 66076 68180 66124 68236
rect 66180 68180 66208 68236
rect 65888 66668 66208 68180
rect 76076 76580 76132 76590
rect 65888 66612 65916 66668
rect 65972 66612 66020 66668
rect 66076 66612 66124 66668
rect 66180 66612 66208 66668
rect 65888 65100 66208 66612
rect 65888 65044 65916 65100
rect 65972 65044 66020 65100
rect 66076 65044 66124 65100
rect 66180 65044 66208 65100
rect 65888 63532 66208 65044
rect 65888 63476 65916 63532
rect 65972 63476 66020 63532
rect 66076 63476 66124 63532
rect 66180 63476 66208 63532
rect 65888 61964 66208 63476
rect 65888 61908 65916 61964
rect 65972 61908 66020 61964
rect 66076 61908 66124 61964
rect 66180 61908 66208 61964
rect 65888 60396 66208 61908
rect 65888 60340 65916 60396
rect 65972 60340 66020 60396
rect 66076 60340 66124 60396
rect 66180 60340 66208 60396
rect 65888 58828 66208 60340
rect 65888 58772 65916 58828
rect 65972 58772 66020 58828
rect 66076 58772 66124 58828
rect 66180 58772 66208 58828
rect 65888 57260 66208 58772
rect 65888 57204 65916 57260
rect 65972 57204 66020 57260
rect 66076 57204 66124 57260
rect 66180 57204 66208 57260
rect 65888 55692 66208 57204
rect 75852 67172 75908 67182
rect 65888 55636 65916 55692
rect 65972 55636 66020 55692
rect 66076 55636 66124 55692
rect 66180 55636 66208 55692
rect 65888 54124 66208 55636
rect 65888 54068 65916 54124
rect 65972 54068 66020 54124
rect 66076 54068 66124 54124
rect 66180 54068 66208 54124
rect 65888 52556 66208 54068
rect 65888 52500 65916 52556
rect 65972 52500 66020 52556
rect 66076 52500 66124 52556
rect 66180 52500 66208 52556
rect 65888 50988 66208 52500
rect 65888 50932 65916 50988
rect 65972 50932 66020 50988
rect 66076 50932 66124 50988
rect 66180 50932 66208 50988
rect 65888 49420 66208 50932
rect 65888 49364 65916 49420
rect 65972 49364 66020 49420
rect 66076 49364 66124 49420
rect 66180 49364 66208 49420
rect 65888 47852 66208 49364
rect 65888 47796 65916 47852
rect 65972 47796 66020 47852
rect 66076 47796 66124 47852
rect 66180 47796 66208 47852
rect 65888 46284 66208 47796
rect 65888 46228 65916 46284
rect 65972 46228 66020 46284
rect 66076 46228 66124 46284
rect 66180 46228 66208 46284
rect 65888 44716 66208 46228
rect 74060 56644 74116 56654
rect 65888 44660 65916 44716
rect 65972 44660 66020 44716
rect 66076 44660 66124 44716
rect 66180 44660 66208 44716
rect 65888 43148 66208 44660
rect 65888 43092 65916 43148
rect 65972 43092 66020 43148
rect 66076 43092 66124 43148
rect 66180 43092 66208 43148
rect 50528 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50848 40796
rect 50528 39228 50848 40740
rect 65772 42196 65828 42206
rect 65772 39508 65828 42140
rect 65772 39442 65828 39452
rect 65888 41580 66208 43092
rect 65888 41524 65916 41580
rect 65972 41524 66020 41580
rect 66076 41524 66124 41580
rect 66180 41524 66208 41580
rect 65888 40012 66208 41524
rect 65888 39956 65916 40012
rect 65972 39956 66020 40012
rect 66076 39956 66124 40012
rect 66180 39956 66208 40012
rect 50528 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50848 39228
rect 50528 37660 50848 39172
rect 50528 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50848 37660
rect 50528 36092 50848 37604
rect 50528 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50848 36092
rect 50528 34524 50848 36036
rect 50528 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50848 34524
rect 50528 32956 50848 34468
rect 50528 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50848 32956
rect 50528 31388 50848 32900
rect 50528 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50848 31388
rect 50528 29820 50848 31332
rect 50528 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50848 29820
rect 49756 29428 49812 29438
rect 49756 26180 49812 29372
rect 49756 26114 49812 26124
rect 50528 28252 50848 29764
rect 50528 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50848 28252
rect 50528 26684 50848 28196
rect 50528 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50848 26684
rect 50528 25116 50848 26628
rect 50528 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50848 25116
rect 49308 23716 49364 23726
rect 47628 22932 47684 22942
rect 47180 22372 47236 22382
rect 47180 21588 47236 22316
rect 47628 21700 47684 22876
rect 47628 21634 47684 21644
rect 47180 21522 47236 21532
rect 48972 20356 49028 20366
rect 48972 19236 49028 20300
rect 49308 20020 49364 23660
rect 50528 23548 50848 25060
rect 50528 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50848 23548
rect 49532 23380 49588 23390
rect 49308 19954 49364 19964
rect 49420 22372 49476 22382
rect 48972 19170 49028 19180
rect 49420 18564 49476 22316
rect 49532 21588 49588 23324
rect 49532 21522 49588 21532
rect 50528 21980 50848 23492
rect 50528 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50848 21980
rect 49420 18498 49476 18508
rect 50528 20412 50848 21924
rect 50528 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50848 20412
rect 50528 18844 50848 20356
rect 50528 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50848 18844
rect 47068 16818 47124 16828
rect 50528 17276 50848 18788
rect 50528 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50848 17276
rect 46844 15250 46900 15260
rect 50528 15708 50848 17220
rect 50528 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50848 15708
rect 42028 12786 42084 12796
rect 50528 14140 50848 15652
rect 50528 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50848 14140
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 31724 10164 31780 10174
rect 31724 9716 31780 10108
rect 31724 9650 31780 9660
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 18732 9380 18788 9390
rect 4448 5516 4768 7028
rect 13916 7028 13972 7038
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 9996 5572 10052 5582
rect 9996 3892 10052 5516
rect 13916 5572 13972 6972
rect 15148 6580 15204 6590
rect 15148 6132 15204 6524
rect 15148 6066 15204 6076
rect 18620 6468 18676 6478
rect 13916 5506 13972 5516
rect 14364 5572 14420 5582
rect 14364 4788 14420 5516
rect 14364 4722 14420 4732
rect 18620 4116 18676 6412
rect 18732 6132 18788 9324
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19628 9268 19684 9278
rect 19628 8260 19684 9212
rect 19628 8194 19684 8204
rect 18732 5236 18788 6076
rect 18732 5170 18788 5180
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 35168 8652 35488 10164
rect 50528 12572 50848 14084
rect 50528 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50848 12572
rect 50528 11004 50848 12516
rect 50528 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50848 11004
rect 38220 10052 38276 10062
rect 38220 9828 38276 9996
rect 38220 9762 38276 9772
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 28588 7476 28644 7486
rect 28588 6692 28644 7420
rect 33180 7476 33236 7486
rect 30940 7364 30996 7374
rect 28588 6626 28644 6636
rect 30828 6916 30884 6926
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 30828 6356 30884 6860
rect 30828 6290 30884 6300
rect 18620 4050 18676 4060
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 30940 4788 30996 7308
rect 31500 6804 31556 6814
rect 31500 6244 31556 6748
rect 31500 6178 31556 6188
rect 33180 6580 33236 7420
rect 30940 4722 30996 4732
rect 9996 3826 10052 3836
rect 19808 3164 20128 4676
rect 33180 4340 33236 6524
rect 33180 4274 33236 4284
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
rect 50528 9436 50848 10948
rect 50528 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50848 9436
rect 50528 7868 50848 9380
rect 50528 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50848 7868
rect 50528 6300 50848 7812
rect 50528 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50848 6300
rect 50528 4732 50848 6244
rect 50528 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50848 4732
rect 50528 3164 50848 4676
rect 50528 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50848 3164
rect 50528 3076 50848 3108
rect 65888 38444 66208 39956
rect 72604 45108 72660 45118
rect 72604 38668 72660 45052
rect 72828 39620 72884 39630
rect 65888 38388 65916 38444
rect 65972 38388 66020 38444
rect 66076 38388 66124 38444
rect 66180 38388 66208 38444
rect 65888 36876 66208 38388
rect 65888 36820 65916 36876
rect 65972 36820 66020 36876
rect 66076 36820 66124 36876
rect 66180 36820 66208 36876
rect 65888 35308 66208 36820
rect 65888 35252 65916 35308
rect 65972 35252 66020 35308
rect 66076 35252 66124 35308
rect 66180 35252 66208 35308
rect 72492 38612 72660 38668
rect 72716 39172 72772 39182
rect 65888 33740 66208 35252
rect 72268 35252 72324 35262
rect 65888 33684 65916 33740
rect 65972 33684 66020 33740
rect 66076 33684 66124 33740
rect 66180 33684 66208 33740
rect 65888 32172 66208 33684
rect 65888 32116 65916 32172
rect 65972 32116 66020 32172
rect 66076 32116 66124 32172
rect 66180 32116 66208 32172
rect 65888 30604 66208 32116
rect 65888 30548 65916 30604
rect 65972 30548 66020 30604
rect 66076 30548 66124 30604
rect 66180 30548 66208 30604
rect 65888 29036 66208 30548
rect 65888 28980 65916 29036
rect 65972 28980 66020 29036
rect 66076 28980 66124 29036
rect 66180 28980 66208 29036
rect 65888 27468 66208 28980
rect 65888 27412 65916 27468
rect 65972 27412 66020 27468
rect 66076 27412 66124 27468
rect 66180 27412 66208 27468
rect 65888 25900 66208 27412
rect 65888 25844 65916 25900
rect 65972 25844 66020 25900
rect 66076 25844 66124 25900
rect 66180 25844 66208 25900
rect 65888 24332 66208 25844
rect 65888 24276 65916 24332
rect 65972 24276 66020 24332
rect 66076 24276 66124 24332
rect 66180 24276 66208 24332
rect 65888 22764 66208 24276
rect 70812 34692 70868 34702
rect 70812 24052 70868 34636
rect 70812 23986 70868 23996
rect 71596 32452 71652 32462
rect 71596 23828 71652 32396
rect 71820 30548 71876 30558
rect 71820 25060 71876 30492
rect 72268 29428 72324 35196
rect 72380 34692 72436 34702
rect 72380 32676 72436 34636
rect 72380 32610 72436 32620
rect 72268 29362 72324 29372
rect 72380 31892 72436 31902
rect 72380 28532 72436 31836
rect 72492 31444 72548 38612
rect 72604 38164 72660 38174
rect 72604 33348 72660 38108
rect 72716 35252 72772 39116
rect 72828 38612 72884 39564
rect 73724 38836 73780 38846
rect 72828 38546 72884 38556
rect 73388 38612 73444 38622
rect 72940 38164 72996 38174
rect 72940 36820 72996 38108
rect 73388 37380 73444 38556
rect 73388 37314 73444 37324
rect 73724 37268 73780 38780
rect 73724 37202 73780 37212
rect 73948 37716 74004 37726
rect 72940 36754 72996 36764
rect 72716 35186 72772 35196
rect 73276 36372 73332 36382
rect 72604 33282 72660 33292
rect 72940 35140 72996 35150
rect 72940 33348 72996 35084
rect 72940 33282 72996 33292
rect 72492 31378 72548 31388
rect 72604 32452 72660 32462
rect 72380 28466 72436 28476
rect 71932 27860 71988 27870
rect 71932 27300 71988 27804
rect 71932 27234 71988 27244
rect 72268 27748 72324 27758
rect 71820 24994 71876 25004
rect 72268 25060 72324 27692
rect 72604 25732 72660 32396
rect 72716 28980 72772 28990
rect 72716 26740 72772 28924
rect 72716 26674 72772 26684
rect 72604 25666 72660 25676
rect 72268 24994 72324 25004
rect 73276 23940 73332 36316
rect 73948 36372 74004 37660
rect 73948 36306 74004 36316
rect 73724 27748 73780 27758
rect 73724 26908 73780 27692
rect 74060 27636 74116 56588
rect 74620 41636 74676 41646
rect 74396 37492 74452 37502
rect 74396 36372 74452 37436
rect 74396 36306 74452 36316
rect 74060 27076 74116 27580
rect 74060 27010 74116 27020
rect 74508 33012 74564 33022
rect 73724 26852 73892 26908
rect 73836 26292 73892 26852
rect 73836 26226 73892 26236
rect 73276 23874 73332 23884
rect 74508 23940 74564 32956
rect 74508 23874 74564 23884
rect 71596 23762 71652 23772
rect 65888 22708 65916 22764
rect 65972 22708 66020 22764
rect 66076 22708 66124 22764
rect 66180 22708 66208 22764
rect 65888 21196 66208 22708
rect 65888 21140 65916 21196
rect 65972 21140 66020 21196
rect 66076 21140 66124 21196
rect 66180 21140 66208 21196
rect 65888 19628 66208 21140
rect 65888 19572 65916 19628
rect 65972 19572 66020 19628
rect 66076 19572 66124 19628
rect 66180 19572 66208 19628
rect 65888 18060 66208 19572
rect 65888 18004 65916 18060
rect 65972 18004 66020 18060
rect 66076 18004 66124 18060
rect 66180 18004 66208 18060
rect 65888 16492 66208 18004
rect 65888 16436 65916 16492
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 66180 16436 66208 16492
rect 65888 14924 66208 16436
rect 65888 14868 65916 14924
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 66180 14868 66208 14924
rect 65888 13356 66208 14868
rect 74620 14756 74676 41580
rect 75068 40628 75124 40638
rect 75068 39396 75124 40572
rect 75068 39330 75124 39340
rect 75068 38836 75124 38846
rect 74956 34916 75012 34926
rect 74956 26852 75012 34860
rect 75068 31780 75124 38780
rect 75068 31714 75124 31724
rect 75628 33124 75684 33134
rect 74956 26786 75012 26796
rect 75628 27972 75684 33068
rect 75628 25060 75684 27916
rect 75852 29428 75908 67116
rect 76076 55468 76132 76524
rect 75964 55412 76132 55468
rect 76300 67844 76356 67854
rect 75964 37268 76020 55412
rect 75964 34356 76020 37212
rect 75964 34290 76020 34300
rect 76188 41972 76244 41982
rect 76188 38276 76244 41916
rect 76188 34356 76244 38220
rect 76188 34290 76244 34300
rect 76300 31780 76356 67788
rect 76412 62244 76468 62254
rect 76412 38668 76468 62188
rect 76972 61348 77028 61358
rect 76412 38612 76916 38668
rect 76636 37268 76692 37278
rect 76636 33460 76692 37212
rect 76636 33394 76692 33404
rect 76300 31714 76356 31724
rect 75852 26516 75908 29372
rect 76860 30212 76916 38612
rect 76860 28644 76916 30156
rect 76860 28578 76916 28588
rect 75852 26450 75908 26460
rect 76524 28532 76580 28542
rect 75628 24994 75684 25004
rect 76524 24724 76580 28476
rect 76972 27636 77028 61292
rect 77868 35924 77924 35934
rect 77868 35140 77924 35868
rect 77868 35074 77924 35084
rect 77084 33236 77140 33246
rect 77084 32004 77140 33180
rect 77084 31938 77140 31948
rect 76972 27570 77028 27580
rect 76524 24658 76580 24668
rect 77644 21924 77700 21934
rect 75404 21588 75460 21598
rect 75404 19012 75460 21532
rect 76412 20468 76468 20478
rect 76412 20020 76468 20412
rect 76412 19954 76468 19964
rect 77644 19908 77700 21868
rect 77644 19842 77700 19852
rect 77756 21700 77812 21710
rect 75404 18946 75460 18956
rect 77756 16772 77812 21644
rect 77756 16706 77812 16716
rect 74620 14690 74676 14700
rect 65888 13300 65916 13356
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 66180 13300 66208 13356
rect 65888 11788 66208 13300
rect 65888 11732 65916 11788
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 66180 11732 66208 11788
rect 65888 10220 66208 11732
rect 65888 10164 65916 10220
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 66180 10164 66208 10220
rect 65888 8652 66208 10164
rect 65888 8596 65916 8652
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 66180 8596 66208 8652
rect 65888 7084 66208 8596
rect 65888 7028 65916 7084
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 66180 7028 66208 7084
rect 65888 5516 66208 7028
rect 65888 5460 65916 5516
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 66180 5460 66208 5516
rect 65888 3948 66208 5460
rect 65888 3892 65916 3948
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 66180 3892 66208 3948
rect 65888 3076 66208 3892
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0663_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 48384 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0664_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 48832 0 1 6272
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _0665_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 48272 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0666_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 41440 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0667_
timestamp 1698431365
transform -1 0 44464 0 1 4704
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0668_
timestamp 1698431365
transform 1 0 36400 0 -1 4704
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0669_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 43232 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0670_
timestamp 1698431365
transform 1 0 34944 0 -1 6272
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0671_
timestamp 1698431365
transform -1 0 36624 0 1 4704
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0672_
timestamp 1698431365
transform -1 0 32704 0 -1 4704
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _0673_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 33488 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0674_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 40320 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0675_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 33376 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0676_
timestamp 1698431365
transform 1 0 35840 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0677_
timestamp 1698431365
transform 1 0 42448 0 -1 6272
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0678_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 42896 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0679_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 40208 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _0680_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 38416 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _0681_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 39872 0 1 4704
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or4_2  _0682_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 42448 0 -1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _0683_
timestamp 1698431365
transform -1 0 40544 0 -1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0684_
timestamp 1698431365
transform 1 0 42336 0 -1 4704
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0685_
timestamp 1698431365
transform -1 0 44240 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0686_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 47488 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0687_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 45248 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0688_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 43232 0 1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0689_
timestamp 1698431365
transform -1 0 46928 0 -1 17248
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _0690_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 47040 0 -1 18816
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0691_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 40768 0 -1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0692_
timestamp 1698431365
transform 1 0 39424 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0693_
timestamp 1698431365
transform 1 0 43456 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0694_
timestamp 1698431365
transform 1 0 41776 0 -1 7840
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0695_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 42560 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0696_
timestamp 1698431365
transform 1 0 70784 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0697_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 72464 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0698_
timestamp 1698431365
transform 1 0 73920 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0699_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 50736 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0700_
timestamp 1698431365
transform 1 0 49840 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0701_
timestamp 1698431365
transform -1 0 46816 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _0702_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 70784 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0703_
timestamp 1698431365
transform 1 0 74032 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0704_
timestamp 1698431365
transform 1 0 74816 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0705_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 40544 0 1 7840
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0706_
timestamp 1698431365
transform -1 0 41664 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0707_
timestamp 1698431365
transform 1 0 69888 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0708_
timestamp 1698431365
transform -1 0 68432 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0709_
timestamp 1698431365
transform -1 0 60816 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0710_
timestamp 1698431365
transform -1 0 58688 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0711_
timestamp 1698431365
transform 1 0 54992 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0712_
timestamp 1698431365
transform 1 0 55328 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0713_
timestamp 1698431365
transform 1 0 55216 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0714_
timestamp 1698431365
transform 1 0 56448 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0715_
timestamp 1698431365
transform -1 0 57344 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0716_
timestamp 1698431365
transform 1 0 56560 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0717_
timestamp 1698431365
transform -1 0 58240 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0718_
timestamp 1698431365
transform 1 0 57456 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0719_
timestamp 1698431365
transform 1 0 44688 0 1 4704
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0720_
timestamp 1698431365
transform 1 0 72240 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0721_
timestamp 1698431365
transform 1 0 73472 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0722_
timestamp 1698431365
transform 1 0 75040 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0723_
timestamp 1698431365
transform 1 0 74816 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0724_
timestamp 1698431365
transform -1 0 76720 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0725_
timestamp 1698431365
transform 1 0 76944 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0726_
timestamp 1698431365
transform 1 0 77728 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0727_
timestamp 1698431365
transform 1 0 74816 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0728_
timestamp 1698431365
transform -1 0 77728 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0729_
timestamp 1698431365
transform 1 0 76048 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0730_
timestamp 1698431365
transform -1 0 76720 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0731_
timestamp 1698431365
transform 1 0 31472 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0732_
timestamp 1698431365
transform -1 0 42896 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0733_
timestamp 1698431365
transform -1 0 43568 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _0734_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 37968 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0735_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 74704 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0736_
timestamp 1698431365
transform 1 0 75600 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0737_
timestamp 1698431365
transform -1 0 77392 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0738_
timestamp 1698431365
transform -1 0 76160 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0739_
timestamp 1698431365
transform 1 0 44016 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0740_
timestamp 1698431365
transform -1 0 62720 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0741_
timestamp 1698431365
transform -1 0 62496 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0742_
timestamp 1698431365
transform -1 0 60144 0 1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0743_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 73360 0 -1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0744_
timestamp 1698431365
transform -1 0 39872 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0745_
timestamp 1698431365
transform -1 0 36512 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0746_
timestamp 1698431365
transform 1 0 33712 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0747_
timestamp 1698431365
transform 1 0 39872 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0748_
timestamp 1698431365
transform -1 0 40432 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0749_
timestamp 1698431365
transform -1 0 36624 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0750_
timestamp 1698431365
transform 1 0 34832 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0751_
timestamp 1698431365
transform 1 0 36064 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0752_
timestamp 1698431365
transform -1 0 41440 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0753_
timestamp 1698431365
transform -1 0 34496 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0754_
timestamp 1698431365
transform -1 0 42560 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0755_
timestamp 1698431365
transform -1 0 35392 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0756_
timestamp 1698431365
transform 1 0 34832 0 1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0757_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 36960 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0758_
timestamp 1698431365
transform -1 0 26880 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0759_
timestamp 1698431365
transform -1 0 74704 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0760_
timestamp 1698431365
transform -1 0 75824 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0761_
timestamp 1698431365
transform -1 0 61824 0 1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0762_
timestamp 1698431365
transform 1 0 73248 0 1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0763_
timestamp 1698431365
transform 1 0 33152 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0764_
timestamp 1698431365
transform 1 0 34944 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0765_
timestamp 1698431365
transform 1 0 35504 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0766_
timestamp 1698431365
transform -1 0 35168 0 1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0767_
timestamp 1698431365
transform 1 0 35392 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0768_
timestamp 1698431365
transform 1 0 30128 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0769_
timestamp 1698431365
transform -1 0 73808 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0770_
timestamp 1698431365
transform 1 0 73472 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0771_
timestamp 1698431365
transform 1 0 75488 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0772_
timestamp 1698431365
transform 1 0 59696 0 -1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0773_
timestamp 1698431365
transform 1 0 73808 0 -1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0774_
timestamp 1698431365
transform 1 0 34048 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0775_
timestamp 1698431365
transform 1 0 34160 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0776_
timestamp 1698431365
transform 1 0 35056 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0777_
timestamp 1698431365
transform 1 0 35280 0 -1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0778_
timestamp 1698431365
transform 1 0 35616 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0779_
timestamp 1698431365
transform 1 0 29008 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0780_
timestamp 1698431365
transform -1 0 73024 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0781_
timestamp 1698431365
transform -1 0 71680 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0782_
timestamp 1698431365
transform 1 0 76048 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0783_
timestamp 1698431365
transform 1 0 61376 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0784_
timestamp 1698431365
transform -1 0 63280 0 1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0785_
timestamp 1698431365
transform 1 0 72128 0 -1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0786_
timestamp 1698431365
transform 1 0 33600 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0787_
timestamp 1698431365
transform 1 0 35056 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0788_
timestamp 1698431365
transform -1 0 35504 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0789_
timestamp 1698431365
transform 1 0 35168 0 1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0790_
timestamp 1698431365
transform 1 0 35728 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0791_
timestamp 1698431365
transform 1 0 19824 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _0792_
timestamp 1698431365
transform -1 0 39760 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0793_
timestamp 1698431365
transform 1 0 71680 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0794_
timestamp 1698431365
transform 1 0 76608 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0795_
timestamp 1698431365
transform 1 0 77392 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0796_
timestamp 1698431365
transform -1 0 64064 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0797_
timestamp 1698431365
transform 1 0 62496 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0798_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 63840 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0799_
timestamp 1698431365
transform 1 0 34496 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0800_
timestamp 1698431365
transform 1 0 33600 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0801_
timestamp 1698431365
transform -1 0 37632 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0802_
timestamp 1698431365
transform 1 0 35168 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0803_
timestamp 1698431365
transform 1 0 36960 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0804_
timestamp 1698431365
transform 1 0 36848 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0805_
timestamp 1698431365
transform 1 0 37072 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0806_
timestamp 1698431365
transform -1 0 39088 0 -1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0807_
timestamp 1698431365
transform 1 0 37968 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0808_
timestamp 1698431365
transform 1 0 23296 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0809_
timestamp 1698431365
transform -1 0 73472 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0810_
timestamp 1698431365
transform -1 0 77392 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0811_
timestamp 1698431365
transform 1 0 62496 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0812_
timestamp 1698431365
transform -1 0 63728 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0813_
timestamp 1698431365
transform 1 0 34048 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0814_
timestamp 1698431365
transform 1 0 35168 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0815_
timestamp 1698431365
transform 1 0 37520 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0816_
timestamp 1698431365
transform -1 0 39200 0 1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0817_
timestamp 1698431365
transform 1 0 38080 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0818_
timestamp 1698431365
transform 1 0 19600 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0819_
timestamp 1698431365
transform 1 0 71680 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0820_
timestamp 1698431365
transform 1 0 71008 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0821_
timestamp 1698431365
transform 1 0 71568 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0822_
timestamp 1698431365
transform 1 0 77392 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0823_
timestamp 1698431365
transform -1 0 64736 0 1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0824_
timestamp 1698431365
transform 1 0 71008 0 1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0825_
timestamp 1698431365
transform 1 0 34496 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0826_
timestamp 1698431365
transform 1 0 36848 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0827_
timestamp 1698431365
transform -1 0 36064 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0828_
timestamp 1698431365
transform 1 0 37968 0 1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0829_
timestamp 1698431365
transform 1 0 36960 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0830_
timestamp 1698431365
transform 1 0 24416 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0831_
timestamp 1698431365
transform -1 0 73696 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0832_
timestamp 1698431365
transform 1 0 72128 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0833_
timestamp 1698431365
transform 1 0 77392 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0834_
timestamp 1698431365
transform 1 0 64288 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0835_
timestamp 1698431365
transform 1 0 64288 0 -1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0836_
timestamp 1698431365
transform 1 0 72688 0 1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0837_
timestamp 1698431365
transform 1 0 34944 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0838_
timestamp 1698431365
transform 1 0 35616 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0839_
timestamp 1698431365
transform 1 0 36064 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0840_
timestamp 1698431365
transform -1 0 40432 0 -1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0841_
timestamp 1698431365
transform -1 0 40544 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0842_
timestamp 1698431365
transform -1 0 21504 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _0843_
timestamp 1698431365
transform 1 0 41216 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0844_
timestamp 1698431365
transform -1 0 71904 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0845_
timestamp 1698431365
transform -1 0 76608 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0846_
timestamp 1698431365
transform 1 0 75264 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0847_
timestamp 1698431365
transform 1 0 64512 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0848_
timestamp 1698431365
transform -1 0 66976 0 1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0849_
timestamp 1698431365
transform 1 0 71344 0 1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0850_
timestamp 1698431365
transform 1 0 38752 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0851_
timestamp 1698431365
transform -1 0 41216 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0852_
timestamp 1698431365
transform -1 0 40880 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0853_
timestamp 1698431365
transform -1 0 39312 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0854_
timestamp 1698431365
transform 1 0 39760 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0855_
timestamp 1698431365
transform 1 0 42224 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0856_
timestamp 1698431365
transform 1 0 40320 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0857_
timestamp 1698431365
transform 1 0 40768 0 -1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0858_
timestamp 1698431365
transform 1 0 40768 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0859_
timestamp 1698431365
transform 1 0 21168 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0860_
timestamp 1698431365
transform 1 0 72128 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0861_
timestamp 1698431365
transform -1 0 75824 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0862_
timestamp 1698431365
transform -1 0 66864 0 1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0863_
timestamp 1698431365
transform 1 0 72128 0 -1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0864_
timestamp 1698431365
transform 1 0 38192 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0865_
timestamp 1698431365
transform 1 0 39312 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0866_
timestamp 1698431365
transform 1 0 41216 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0867_
timestamp 1698431365
transform -1 0 40880 0 1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0868_
timestamp 1698431365
transform 1 0 40880 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0869_
timestamp 1698431365
transform 1 0 24640 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0870_
timestamp 1698431365
transform 1 0 72352 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0871_
timestamp 1698431365
transform -1 0 73360 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0872_
timestamp 1698431365
transform 1 0 77280 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0873_
timestamp 1698431365
transform -1 0 67200 0 -1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0874_
timestamp 1698431365
transform -1 0 75488 0 -1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0875_
timestamp 1698431365
transform 1 0 37744 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0876_
timestamp 1698431365
transform 1 0 39312 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0877_
timestamp 1698431365
transform 1 0 41104 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0878_
timestamp 1698431365
transform 1 0 40768 0 -1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0879_
timestamp 1698431365
transform 1 0 40880 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0880_
timestamp 1698431365
transform 1 0 24304 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0881_
timestamp 1698431365
transform 1 0 74928 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0882_
timestamp 1698431365
transform -1 0 76720 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0883_
timestamp 1698431365
transform 1 0 72800 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0884_
timestamp 1698431365
transform 1 0 76384 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0885_
timestamp 1698431365
transform 1 0 69216 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0886_
timestamp 1698431365
transform -1 0 67984 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0887_
timestamp 1698431365
transform 1 0 66080 0 -1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0888_
timestamp 1698431365
transform 1 0 73024 0 1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0889_
timestamp 1698431365
transform 1 0 38752 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0890_
timestamp 1698431365
transform 1 0 39424 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0891_
timestamp 1698431365
transform 1 0 40320 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0892_
timestamp 1698431365
transform 1 0 40880 0 1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0893_
timestamp 1698431365
transform 1 0 40880 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0894_
timestamp 1698431365
transform -1 0 28784 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _0895_
timestamp 1698431365
transform 1 0 42336 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0896_
timestamp 1698431365
transform 1 0 72688 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0897_
timestamp 1698431365
transform 1 0 76496 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0898_
timestamp 1698431365
transform 1 0 77056 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0899_
timestamp 1698431365
transform 1 0 65184 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0900_
timestamp 1698431365
transform -1 0 68992 0 -1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0901_
timestamp 1698431365
transform 1 0 72128 0 -1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0902_
timestamp 1698431365
transform 1 0 37296 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0903_
timestamp 1698431365
transform 1 0 36848 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0904_
timestamp 1698431365
transform 1 0 37968 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0905_
timestamp 1698431365
transform 1 0 38752 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0906_
timestamp 1698431365
transform 1 0 41664 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0907_
timestamp 1698431365
transform 1 0 41216 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0908_
timestamp 1698431365
transform 1 0 43568 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0909_
timestamp 1698431365
transform -1 0 43568 0 1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0910_
timestamp 1698431365
transform 1 0 44352 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0911_
timestamp 1698431365
transform 1 0 32928 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0912_
timestamp 1698431365
transform 1 0 73584 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0913_
timestamp 1698431365
transform 1 0 77280 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0914_
timestamp 1698431365
transform -1 0 69664 0 1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0915_
timestamp 1698431365
transform 1 0 72016 0 1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0916_
timestamp 1698431365
transform 1 0 37744 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0917_
timestamp 1698431365
transform 1 0 37968 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0918_
timestamp 1698431365
transform 1 0 43232 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0919_
timestamp 1698431365
transform -1 0 44352 0 -1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0920_
timestamp 1698431365
transform 1 0 44688 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0921_
timestamp 1698431365
transform 1 0 33040 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0922_
timestamp 1698431365
transform 1 0 74928 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0923_
timestamp 1698431365
transform -1 0 75376 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0924_
timestamp 1698431365
transform 1 0 76608 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0925_
timestamp 1698431365
transform -1 0 69664 0 1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0926_
timestamp 1698431365
transform 1 0 73808 0 -1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0927_
timestamp 1698431365
transform 1 0 37296 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0928_
timestamp 1698431365
transform -1 0 40208 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0929_
timestamp 1698431365
transform 1 0 43792 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0930_
timestamp 1698431365
transform -1 0 44800 0 -1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0931_
timestamp 1698431365
transform 1 0 44688 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0932_
timestamp 1698431365
transform 1 0 32256 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0933_
timestamp 1698431365
transform 1 0 76272 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0934_
timestamp 1698431365
transform 1 0 76944 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0935_
timestamp 1698431365
transform -1 0 77056 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0936_
timestamp 1698431365
transform 1 0 68544 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0937_
timestamp 1698431365
transform 1 0 68432 0 -1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0938_
timestamp 1698431365
transform 1 0 74032 0 1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0939_
timestamp 1698431365
transform 1 0 36176 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0940_
timestamp 1698431365
transform 1 0 37856 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0941_
timestamp 1698431365
transform 1 0 43568 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0942_
timestamp 1698431365
transform 1 0 44688 0 1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0943_
timestamp 1698431365
transform -1 0 47040 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0944_
timestamp 1698431365
transform -1 0 37744 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0945_
timestamp 1698431365
transform 1 0 45248 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _0946_
timestamp 1698431365
transform -1 0 48160 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0947_
timestamp 1698431365
transform 1 0 76496 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0948_
timestamp 1698431365
transform 1 0 76048 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0949_
timestamp 1698431365
transform -1 0 77616 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0950_
timestamp 1698431365
transform 1 0 77392 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0951_
timestamp 1698431365
transform 1 0 69664 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0952_
timestamp 1698431365
transform 1 0 70448 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0953_
timestamp 1698431365
transform 1 0 69888 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0954_
timestamp 1698431365
transform -1 0 71120 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0955_
timestamp 1698431365
transform 1 0 46256 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0956_
timestamp 1698431365
transform 1 0 45696 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0957_
timestamp 1698431365
transform -1 0 48384 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0958_
timestamp 1698431365
transform 1 0 45024 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0959_
timestamp 1698431365
transform 1 0 46592 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0960_
timestamp 1698431365
transform -1 0 47936 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0961_
timestamp 1698431365
transform 1 0 47712 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0962_
timestamp 1698431365
transform 1 0 45024 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0963_
timestamp 1698431365
transform -1 0 45808 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0964_
timestamp 1698431365
transform 1 0 45920 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0965_
timestamp 1698431365
transform -1 0 47936 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0966_
timestamp 1698431365
transform -1 0 47264 0 1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0967_
timestamp 1698431365
transform 1 0 46256 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0968_
timestamp 1698431365
transform 1 0 38192 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0969_
timestamp 1698431365
transform 1 0 76496 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0970_
timestamp 1698431365
transform -1 0 77392 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0971_
timestamp 1698431365
transform 1 0 70784 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0972_
timestamp 1698431365
transform 1 0 70336 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0973_
timestamp 1698431365
transform -1 0 48384 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0974_
timestamp 1698431365
transform -1 0 46592 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0975_
timestamp 1698431365
transform 1 0 47152 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0976_
timestamp 1698431365
transform 1 0 47264 0 1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0977_
timestamp 1698431365
transform -1 0 48384 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0978_
timestamp 1698431365
transform 1 0 34384 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0979_
timestamp 1698431365
transform 1 0 74256 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0980_
timestamp 1698431365
transform 1 0 76048 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0981_
timestamp 1698431365
transform 1 0 77392 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0982_
timestamp 1698431365
transform 1 0 70224 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0983_
timestamp 1698431365
transform 1 0 69888 0 1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0984_
timestamp 1698431365
transform -1 0 47040 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0985_
timestamp 1698431365
transform -1 0 46592 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0986_
timestamp 1698431365
transform 1 0 46592 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0987_
timestamp 1698431365
transform -1 0 48384 0 -1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0988_
timestamp 1698431365
transform 1 0 48608 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0989_
timestamp 1698431365
transform 1 0 35168 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0990_
timestamp 1698431365
transform -1 0 76944 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0991_
timestamp 1698431365
transform 1 0 76048 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0992_
timestamp 1698431365
transform -1 0 75824 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0993_
timestamp 1698431365
transform 1 0 70448 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0994_
timestamp 1698431365
transform -1 0 71792 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0995_
timestamp 1698431365
transform 1 0 73472 0 -1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0996_
timestamp 1698431365
transform 1 0 44912 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0997_
timestamp 1698431365
transform 1 0 45696 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0998_
timestamp 1698431365
transform 1 0 47264 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0999_
timestamp 1698431365
transform 1 0 48608 0 -1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1000_
timestamp 1698431365
transform -1 0 50176 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1001_
timestamp 1698431365
transform -1 0 28784 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1002_
timestamp 1698431365
transform 1 0 50176 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1003_
timestamp 1698431365
transform 1 0 75376 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1004_
timestamp 1698431365
transform -1 0 78064 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1005_
timestamp 1698431365
transform -1 0 77392 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1006_
timestamp 1698431365
transform 1 0 72016 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1007_
timestamp 1698431365
transform 1 0 72128 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1008_
timestamp 1698431365
transform 1 0 71680 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1009_
timestamp 1698431365
transform 1 0 45696 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1010_
timestamp 1698431365
transform 1 0 46816 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1011_
timestamp 1698431365
transform 1 0 46144 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1012_
timestamp 1698431365
transform 1 0 47264 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1013_
timestamp 1698431365
transform 1 0 49168 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1014_
timestamp 1698431365
transform 1 0 50064 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1015_
timestamp 1698431365
transform 1 0 47936 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1016_
timestamp 1698431365
transform 1 0 48720 0 1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1017_
timestamp 1698431365
transform 1 0 48608 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1018_
timestamp 1698431365
transform 1 0 31584 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1019_
timestamp 1698431365
transform 1 0 75376 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1020_
timestamp 1698431365
transform 1 0 77392 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1021_
timestamp 1698431365
transform 1 0 73024 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1022_
timestamp 1698431365
transform 1 0 72576 0 1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1023_
timestamp 1698431365
transform 1 0 44800 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1024_
timestamp 1698431365
transform 1 0 46368 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1025_
timestamp 1698431365
transform 1 0 48608 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1026_
timestamp 1698431365
transform 1 0 48608 0 -1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1027_
timestamp 1698431365
transform 1 0 48720 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1028_
timestamp 1698431365
transform 1 0 28112 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1029_
timestamp 1698431365
transform 1 0 75152 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1030_
timestamp 1698431365
transform 1 0 76048 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1031_
timestamp 1698431365
transform 1 0 77392 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1032_
timestamp 1698431365
transform 1 0 72688 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1033_
timestamp 1698431365
transform -1 0 74144 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1034_
timestamp 1698431365
transform 1 0 44688 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1035_
timestamp 1698431365
transform 1 0 47264 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1036_
timestamp 1698431365
transform 1 0 49392 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1037_
timestamp 1698431365
transform 1 0 50176 0 1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1038_
timestamp 1698431365
transform 1 0 48720 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1039_
timestamp 1698431365
transform -1 0 31136 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1040_
timestamp 1698431365
transform 1 0 76944 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1041_
timestamp 1698431365
transform 1 0 76384 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1042_
timestamp 1698431365
transform 1 0 77392 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1043_
timestamp 1698431365
transform 1 0 71120 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1044_
timestamp 1698431365
transform -1 0 74480 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1045_
timestamp 1698431365
transform -1 0 74480 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1046_
timestamp 1698431365
transform 1 0 44912 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1047_
timestamp 1698431365
transform 1 0 46368 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1048_
timestamp 1698431365
transform 1 0 48832 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1049_
timestamp 1698431365
transform 1 0 48832 0 1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1050_
timestamp 1698431365
transform 1 0 48720 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1051_
timestamp 1698431365
transform -1 0 41888 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1052_
timestamp 1698431365
transform 1 0 51072 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1053_
timestamp 1698431365
transform 1 0 77056 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1054_
timestamp 1698431365
transform -1 0 78064 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1055_
timestamp 1698431365
transform -1 0 75152 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1056_
timestamp 1698431365
transform 1 0 74144 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1057_
timestamp 1698431365
transform 1 0 74480 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1058_
timestamp 1698431365
transform 1 0 74144 0 1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1059_
timestamp 1698431365
transform 1 0 46592 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1060_
timestamp 1698431365
transform 1 0 44688 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1061_
timestamp 1698431365
transform 1 0 45024 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1062_
timestamp 1698431365
transform -1 0 47488 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1063_
timestamp 1698431365
transform 1 0 50736 0 1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1064_
timestamp 1698431365
transform 1 0 50624 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1065_
timestamp 1698431365
transform 1 0 51296 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1066_
timestamp 1698431365
transform -1 0 51968 0 -1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1067_
timestamp 1698431365
transform 1 0 52528 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1068_
timestamp 1698431365
transform 1 0 45136 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1069_
timestamp 1698431365
transform 1 0 76160 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1070_
timestamp 1698431365
transform 1 0 77392 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1071_
timestamp 1698431365
transform 1 0 74704 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1072_
timestamp 1698431365
transform -1 0 75600 0 -1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1073_
timestamp 1698431365
transform 1 0 44240 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1074_
timestamp 1698431365
transform 1 0 45696 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1075_
timestamp 1698431365
transform 1 0 52304 0 -1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1076_
timestamp 1698431365
transform 1 0 52528 0 1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1077_
timestamp 1698431365
transform -1 0 54208 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1078_
timestamp 1698431365
transform 1 0 44912 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1079_
timestamp 1698431365
transform 1 0 75600 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1080_
timestamp 1698431365
transform 1 0 76384 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1081_
timestamp 1698431365
transform -1 0 77280 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1082_
timestamp 1698431365
transform 1 0 76048 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1083_
timestamp 1698431365
transform 1 0 76048 0 1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1084_
timestamp 1698431365
transform 1 0 45136 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1085_
timestamp 1698431365
transform 1 0 45696 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1086_
timestamp 1698431365
transform 1 0 51296 0 -1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1087_
timestamp 1698431365
transform 1 0 51968 0 -1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1088_
timestamp 1698431365
transform 1 0 52192 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1089_
timestamp 1698431365
transform 1 0 42000 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1090_
timestamp 1698431365
transform 1 0 74704 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1091_
timestamp 1698431365
transform -1 0 76720 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1092_
timestamp 1698431365
transform 1 0 75152 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1093_
timestamp 1698431365
transform 1 0 69104 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1094_
timestamp 1698431365
transform 1 0 76048 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1095_
timestamp 1698431365
transform 1 0 76048 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1096_
timestamp 1698431365
transform 1 0 44688 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1097_
timestamp 1698431365
transform 1 0 45696 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1098_
timestamp 1698431365
transform 1 0 51296 0 1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1099_
timestamp 1698431365
transform -1 0 52640 0 -1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1100_
timestamp 1698431365
transform 1 0 52304 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1101_
timestamp 1698431365
transform 1 0 41440 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1102_
timestamp 1698431365
transform 1 0 52528 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1103_
timestamp 1698431365
transform -1 0 76720 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1104_
timestamp 1698431365
transform 1 0 77280 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1105_
timestamp 1698431365
transform -1 0 75152 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1106_
timestamp 1698431365
transform 1 0 73472 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1107_
timestamp 1698431365
transform 1 0 76944 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1108_
timestamp 1698431365
transform -1 0 78400 0 -1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1109_
timestamp 1698431365
transform -1 0 46928 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1110_
timestamp 1698431365
transform 1 0 44240 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1111_
timestamp 1698431365
transform 1 0 45584 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1112_
timestamp 1698431365
transform 1 0 45360 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1113_
timestamp 1698431365
transform 1 0 52864 0 -1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1114_
timestamp 1698431365
transform 1 0 52640 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1115_
timestamp 1698431365
transform 1 0 54880 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1116_
timestamp 1698431365
transform 1 0 53424 0 -1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1117_
timestamp 1698431365
transform 1 0 52864 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1118_
timestamp 1698431365
transform 1 0 44688 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1119_
timestamp 1698431365
transform -1 0 77840 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1120_
timestamp 1698431365
transform 1 0 77728 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1121_
timestamp 1698431365
transform 1 0 77056 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1122_
timestamp 1698431365
transform 1 0 76720 0 -1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1123_
timestamp 1698431365
transform 1 0 44688 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1124_
timestamp 1698431365
transform 1 0 45360 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1125_
timestamp 1698431365
transform -1 0 54320 0 1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1126_
timestamp 1698431365
transform 1 0 53312 0 1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1127_
timestamp 1698431365
transform 1 0 52640 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1128_
timestamp 1698431365
transform 1 0 40656 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1129_
timestamp 1698431365
transform 1 0 74928 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1130_
timestamp 1698431365
transform 1 0 77728 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1131_
timestamp 1698431365
transform 1 0 76832 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1132_
timestamp 1698431365
transform -1 0 77728 0 1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1133_
timestamp 1698431365
transform 1 0 44464 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1134_
timestamp 1698431365
transform 1 0 45360 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1135_
timestamp 1698431365
transform 1 0 54096 0 -1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1136_
timestamp 1698431365
transform -1 0 56224 0 1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1137_
timestamp 1698431365
transform 1 0 54208 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1138_
timestamp 1698431365
transform 1 0 44912 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1139_
timestamp 1698431365
transform -1 0 73808 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1140_
timestamp 1698431365
transform 1 0 74816 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1141_
timestamp 1698431365
transform 1 0 73136 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1142_
timestamp 1698431365
transform 1 0 72688 0 1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1143_
timestamp 1698431365
transform 1 0 44688 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1144_
timestamp 1698431365
transform -1 0 47152 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1145_
timestamp 1698431365
transform 1 0 54320 0 1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1146_
timestamp 1698431365
transform -1 0 55664 0 -1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1147_
timestamp 1698431365
transform 1 0 56448 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1148_
timestamp 1698431365
transform -1 0 42784 0 -1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1149_
timestamp 1698431365
transform -1 0 41776 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1150_
timestamp 1698431365
transform 1 0 42784 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1151_
timestamp 1698431365
transform -1 0 42896 0 1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1152_
timestamp 1698431365
transform 1 0 74928 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1153_
timestamp 1698431365
transform -1 0 78400 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1154_
timestamp 1698431365
transform 1 0 40320 0 1 6272
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1155_
timestamp 1698431365
transform 1 0 29120 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1156_
timestamp 1698431365
transform -1 0 28448 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1157_
timestamp 1698431365
transform -1 0 15792 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1158_
timestamp 1698431365
transform -1 0 14448 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1159_
timestamp 1698431365
transform 1 0 29792 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1160_
timestamp 1698431365
transform -1 0 28672 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1161_
timestamp 1698431365
transform 1 0 17584 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1162_
timestamp 1698431365
transform 1 0 21728 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1163_
timestamp 1698431365
transform -1 0 20160 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1164_
timestamp 1698431365
transform 1 0 17920 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1165_
timestamp 1698431365
transform -1 0 16464 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1166_
timestamp 1698431365
transform 1 0 15344 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1167_
timestamp 1698431365
transform 1 0 17920 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1168_
timestamp 1698431365
transform -1 0 15792 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1169_
timestamp 1698431365
transform -1 0 11424 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1170_
timestamp 1698431365
transform 1 0 18256 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1171_
timestamp 1698431365
transform -1 0 16016 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1172_
timestamp 1698431365
transform -1 0 15120 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1173_
timestamp 1698431365
transform 1 0 17920 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1174_
timestamp 1698431365
transform -1 0 17920 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1175_
timestamp 1698431365
transform -1 0 17024 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1176_
timestamp 1698431365
transform -1 0 17696 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1177_
timestamp 1698431365
transform -1 0 19824 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1178_
timestamp 1698431365
transform -1 0 20608 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1179_
timestamp 1698431365
transform 1 0 19040 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1180_
timestamp 1698431365
transform -1 0 18144 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1181_
timestamp 1698431365
transform -1 0 15904 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1182_
timestamp 1698431365
transform 1 0 19824 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1183_
timestamp 1698431365
transform 1 0 19936 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1184_
timestamp 1698431365
transform 1 0 19264 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1185_
timestamp 1698431365
transform 1 0 19488 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1186_
timestamp 1698431365
transform -1 0 18592 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1187_
timestamp 1698431365
transform -1 0 18144 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1188_
timestamp 1698431365
transform 1 0 19600 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1189_
timestamp 1698431365
transform -1 0 19488 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1190_
timestamp 1698431365
transform -1 0 30576 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1191_
timestamp 1698431365
transform 1 0 20160 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1192_
timestamp 1698431365
transform 1 0 22848 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1193_
timestamp 1698431365
transform -1 0 28672 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1194_
timestamp 1698431365
transform -1 0 27104 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1195_
timestamp 1698431365
transform -1 0 27552 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1196_
timestamp 1698431365
transform 1 0 25984 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1197_
timestamp 1698431365
transform -1 0 22176 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1198_
timestamp 1698431365
transform -1 0 21504 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1199_
timestamp 1698431365
transform 1 0 25984 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1200_
timestamp 1698431365
transform -1 0 23520 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1201_
timestamp 1698431365
transform -1 0 22736 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1202_
timestamp 1698431365
transform 1 0 25536 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1203_
timestamp 1698431365
transform -1 0 23968 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1204_
timestamp 1698431365
transform -1 0 22176 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1205_
timestamp 1698431365
transform -1 0 27216 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1206_
timestamp 1698431365
transform 1 0 27216 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1207_
timestamp 1698431365
transform -1 0 20160 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1208_
timestamp 1698431365
transform -1 0 20944 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1209_
timestamp 1698431365
transform -1 0 27440 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1210_
timestamp 1698431365
transform 1 0 13776 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1211_
timestamp 1698431365
transform -1 0 25760 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1212_
timestamp 1698431365
transform 1 0 23968 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1213_
timestamp 1698431365
transform -1 0 22736 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1214_
timestamp 1698431365
transform 1 0 21392 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1215_
timestamp 1698431365
transform 1 0 25536 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1216_
timestamp 1698431365
transform -1 0 25200 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1217_
timestamp 1698431365
transform -1 0 19488 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1218_
timestamp 1698431365
transform 1 0 25088 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1219_
timestamp 1698431365
transform -1 0 22624 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1220_
timestamp 1698431365
transform 1 0 21280 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1221_
timestamp 1698431365
transform -1 0 26880 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1222_
timestamp 1698431365
transform -1 0 23968 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1223_
timestamp 1698431365
transform -1 0 33488 0 -1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1224_
timestamp 1698431365
transform -1 0 27440 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1225_
timestamp 1698431365
transform -1 0 26768 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1226_
timestamp 1698431365
transform 1 0 30464 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1227_
timestamp 1698431365
transform -1 0 32032 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1228_
timestamp 1698431365
transform -1 0 34272 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1229_
timestamp 1698431365
transform 1 0 31472 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1230_
timestamp 1698431365
transform -1 0 30464 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1231_
timestamp 1698431365
transform -1 0 25984 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1232_
timestamp 1698431365
transform 1 0 32032 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1233_
timestamp 1698431365
transform 1 0 32928 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1234_
timestamp 1698431365
transform 1 0 27104 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1235_
timestamp 1698431365
transform 1 0 31136 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1236_
timestamp 1698431365
transform -1 0 30240 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1237_
timestamp 1698431365
transform -1 0 25312 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1238_
timestamp 1698431365
transform 1 0 31136 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1239_
timestamp 1698431365
transform -1 0 29680 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1240_
timestamp 1698431365
transform -1 0 29456 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1241_
timestamp 1698431365
transform -1 0 28784 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1242_
timestamp 1698431365
transform 1 0 32032 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1243_
timestamp 1698431365
transform 1 0 32480 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1244_
timestamp 1698431365
transform 1 0 33936 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1245_
timestamp 1698431365
transform -1 0 33824 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1246_
timestamp 1698431365
transform -1 0 29792 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1247_
timestamp 1698431365
transform 1 0 34048 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1248_
timestamp 1698431365
transform -1 0 31136 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1249_
timestamp 1698431365
transform -1 0 28112 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1250_
timestamp 1698431365
transform 1 0 32480 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1251_
timestamp 1698431365
transform -1 0 32032 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1252_
timestamp 1698431365
transform 1 0 31360 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1253_
timestamp 1698431365
transform -1 0 34272 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1254_
timestamp 1698431365
transform 1 0 34832 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1255_
timestamp 1698431365
transform -1 0 29120 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1256_
timestamp 1698431365
transform -1 0 26096 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1257_
timestamp 1698431365
transform 1 0 25648 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1258_
timestamp 1698431365
transform -1 0 24864 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1259_
timestamp 1698431365
transform -1 0 24416 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1260_
timestamp 1698431365
transform 1 0 25088 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1261_
timestamp 1698431365
transform -1 0 28224 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1262_
timestamp 1698431365
transform 1 0 24192 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1263_
timestamp 1698431365
transform -1 0 25984 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1264_
timestamp 1698431365
transform -1 0 23856 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1265_
timestamp 1698431365
transform -1 0 28224 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1266_
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1267_
timestamp 1698431365
transform -1 0 26768 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1268_
timestamp 1698431365
transform -1 0 20944 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1269_
timestamp 1698431365
transform -1 0 19824 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1270_
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1271_
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1272_
timestamp 1698431365
transform 1 0 19488 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1273_
timestamp 1698431365
transform 1 0 21168 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1274_
timestamp 1698431365
transform -1 0 16352 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1275_
timestamp 1698431365
transform -1 0 18144 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1276_
timestamp 1698431365
transform 1 0 19824 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1277_
timestamp 1698431365
transform -1 0 22064 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1278_
timestamp 1698431365
transform -1 0 22064 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1279_
timestamp 1698431365
transform -1 0 19600 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1280_
timestamp 1698431365
transform 1 0 19376 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1281_
timestamp 1698431365
transform 1 0 19264 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1282_
timestamp 1698431365
transform -1 0 18144 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1283_
timestamp 1698431365
transform -1 0 20160 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1284_
timestamp 1698431365
transform 1 0 18704 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1285_
timestamp 1698431365
transform 1 0 22960 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1286_
timestamp 1698431365
transform 1 0 18816 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1287_
timestamp 1698431365
transform -1 0 22960 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1288_
timestamp 1698431365
transform 1 0 26432 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1289_
timestamp 1698431365
transform 1 0 25088 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1290_
timestamp 1698431365
transform 1 0 25648 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1291_
timestamp 1698431365
transform -1 0 27776 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1292_
timestamp 1698431365
transform 1 0 26096 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1293_
timestamp 1698431365
transform -1 0 30128 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1294_
timestamp 1698431365
transform -1 0 24640 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1295_
timestamp 1698431365
transform 1 0 30128 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1296_
timestamp 1698431365
transform 1 0 25088 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1297_
timestamp 1698431365
transform -1 0 30128 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1298_
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1299_
timestamp 1698431365
transform 1 0 34272 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1300_
timestamp 1698431365
transform 1 0 27776 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1301_
timestamp 1698431365
transform -1 0 34272 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1302_
timestamp 1698431365
transform 1 0 33712 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1303_
timestamp 1698431365
transform -1 0 36288 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1304_
timestamp 1698431365
transform 1 0 34272 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1305_
timestamp 1698431365
transform -1 0 36176 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1306_
timestamp 1698431365
transform -1 0 33376 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1307_
timestamp 1698431365
transform -1 0 33824 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1308_
timestamp 1698431365
transform -1 0 32816 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1309_
timestamp 1698431365
transform -1 0 33824 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1310_
timestamp 1698431365
transform -1 0 28784 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1311_
timestamp 1698431365
transform -1 0 28336 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1312_
timestamp 1698431365
transform -1 0 27552 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1313_
timestamp 1698431365
transform 1 0 26432 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1314_
timestamp 1698431365
transform 1 0 27664 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1315_
timestamp 1698431365
transform 1 0 29008 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1316_
timestamp 1698431365
transform -1 0 26432 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1317_
timestamp 1698431365
transform -1 0 26992 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1318_
timestamp 1698431365
transform 1 0 26432 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1319_
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1320_
timestamp 1698431365
transform 1 0 38864 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1321_
timestamp 1698431365
transform 1 0 36848 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1322_
timestamp 1698431365
transform 1 0 37744 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1323_
timestamp 1698431365
transform -1 0 40432 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1324_
timestamp 1698431365
transform -1 0 36736 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1325_
timestamp 1698431365
transform -1 0 43232 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1326_
timestamp 1698431365
transform 1 0 36736 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1327_
timestamp 1698431365
transform 1 0 42336 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1328_
timestamp 1698431365
transform 1 0 37184 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1329_
timestamp 1698431365
transform -1 0 40544 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1330_
timestamp 1698431365
transform 1 0 38304 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1331_
timestamp 1698431365
transform 1 0 36848 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1332_
timestamp 1698431365
transform 1 0 38528 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1333_
timestamp 1698431365
transform -1 0 39984 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1334_
timestamp 1698431365
transform 1 0 37520 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1335_
timestamp 1698431365
transform -1 0 42784 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1336_
timestamp 1698431365
transform 1 0 38640 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1337_
timestamp 1698431365
transform 1 0 38528 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1338_
timestamp 1698431365
transform 1 0 38080 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1339_
timestamp 1698431365
transform 1 0 42784 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1340_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 37856 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1341_
timestamp 1698431365
transform -1 0 38416 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1342_
timestamp 1698431365
transform -1 0 29568 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1343_
timestamp 1698431365
transform -1 0 9184 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1344_
timestamp 1698431365
transform 1 0 9072 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1345_
timestamp 1698431365
transform -1 0 30016 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1346_
timestamp 1698431365
transform -1 0 14672 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1347_
timestamp 1698431365
transform -1 0 14000 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1348_
timestamp 1698431365
transform 1 0 11872 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1349_
timestamp 1698431365
transform -1 0 9184 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1350_
timestamp 1698431365
transform -1 0 8400 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1351_
timestamp 1698431365
transform 1 0 11200 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1352_
timestamp 1698431365
transform -1 0 8400 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1353_
timestamp 1698431365
transform -1 0 9072 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1354_
timestamp 1698431365
transform 1 0 11312 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1355_
timestamp 1698431365
transform -1 0 9744 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1356_
timestamp 1698431365
transform -1 0 8848 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1357_
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1358_
timestamp 1698431365
transform -1 0 14000 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1359_
timestamp 1698431365
transform -1 0 9856 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1360_
timestamp 1698431365
transform -1 0 7168 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1361_
timestamp 1698431365
transform -1 0 14784 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1362_
timestamp 1698431365
transform -1 0 15344 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1363_
timestamp 1698431365
transform 1 0 13216 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1364_
timestamp 1698431365
transform -1 0 11424 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1365_
timestamp 1698431365
transform -1 0 6496 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1366_
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1367_
timestamp 1698431365
transform -1 0 10976 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1368_
timestamp 1698431365
transform -1 0 7840 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1369_
timestamp 1698431365
transform 1 0 12208 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1370_
timestamp 1698431365
transform -1 0 8512 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1371_
timestamp 1698431365
transform -1 0 9184 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1372_
timestamp 1698431365
transform 1 0 13776 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1373_
timestamp 1698431365
transform -1 0 12208 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1374_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15232 0 1 10976
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1375_
timestamp 1698431365
transform 1 0 14448 0 1 7840
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1376_
timestamp 1698431365
transform 1 0 14784 0 1 6272
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1377_
timestamp 1698431365
transform 1 0 15792 0 1 4704
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1378_
timestamp 1698431365
transform 1 0 16352 0 1 12544
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1379_
timestamp 1698431365
transform 1 0 19488 0 -1 14112
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1380_
timestamp 1698431365
transform 1 0 18592 0 -1 10976
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1381_
timestamp 1698431365
transform 1 0 19376 0 -1 9408
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1382_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25088 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1383_
timestamp 1698431365
transform 1 0 22736 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1384_
timestamp 1698431365
transform 1 0 22512 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1385_
timestamp 1698431365
transform 1 0 25984 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1386_
timestamp 1698431365
transform 1 0 21504 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1387_
timestamp 1698431365
transform 1 0 25200 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1388_
timestamp 1698431365
transform 1 0 21504 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1389_
timestamp 1698431365
transform 1 0 22736 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1390_
timestamp 1698431365
transform 1 0 29232 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1391_
timestamp 1698431365
transform 1 0 32928 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1392_
timestamp 1698431365
transform 1 0 29008 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1393_
timestamp 1698431365
transform 1 0 27888 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1394_
timestamp 1698431365
transform 1 0 33824 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1395_
timestamp 1698431365
transform 1 0 33376 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1396_
timestamp 1698431365
transform 1 0 29456 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1397_
timestamp 1698431365
transform 1 0 34272 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1398_
timestamp 1698431365
transform 1 0 28224 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1399_
timestamp 1698431365
transform 1 0 23856 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1400_
timestamp 1698431365
transform 1 0 26880 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1401_
timestamp 1698431365
transform 1 0 25312 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1402_
timestamp 1698431365
transform 1 0 16576 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1403_
timestamp 1698431365
transform 1 0 20048 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1404_
timestamp 1698431365
transform 1 0 16352 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1405_
timestamp 1698431365
transform 1 0 21168 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1406_
timestamp 1698431365
transform 1 0 18704 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1407_
timestamp 1698431365
transform 1 0 18368 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1408_
timestamp 1698431365
transform 1 0 21616 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1409_
timestamp 1698431365
transform 1 0 21504 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1410_
timestamp 1698431365
transform 1 0 26208 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1411_
timestamp 1698431365
transform 1 0 29120 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1412_
timestamp 1698431365
transform 1 0 29456 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1413_
timestamp 1698431365
transform 1 0 29008 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1414_
timestamp 1698431365
transform 1 0 35056 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1415_
timestamp 1698431365
transform 1 0 34944 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1416_
timestamp 1698431365
transform 1 0 31136 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1417_
timestamp 1698431365
transform 1 0 31920 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1418_
timestamp 1698431365
transform 1 0 25536 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1419_
timestamp 1698431365
transform 1 0 28336 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1420_
timestamp 1698431365
transform 1 0 24864 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1421_
timestamp 1698431365
transform 1 0 28224 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1422_
timestamp 1698431365
transform 1 0 38976 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1423_
timestamp 1698431365
transform 1 0 41888 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1424_
timestamp 1698431365
transform 1 0 41552 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1425_
timestamp 1698431365
transform 1 0 39088 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1426_
timestamp 1698431365
transform 1 0 37296 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1427_
timestamp 1698431365
transform 1 0 41216 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1428_
timestamp 1698431365
transform 1 0 37296 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1429_
timestamp 1698431365
transform 1 0 41664 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1430_
timestamp 1698431365
transform 1 0 40768 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1431_
timestamp 1698431365
transform 1 0 37072 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1432_
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1433_
timestamp 1698431365
transform 1 0 8400 0 1 9408
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1434_
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1435_
timestamp 1698431365
transform 1 0 12432 0 -1 10976
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1436_
timestamp 1698431365
transform 1 0 9632 0 1 7840
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1437_
timestamp 1698431365
transform 1 0 9744 0 -1 6272
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1438_
timestamp 1698431365
transform 1 0 10080 0 -1 4704
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1439_
timestamp 1698431365
transform 1 0 13552 0 -1 4704
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1456_
timestamp 1698431365
transform -1 0 3248 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1457_
timestamp 1698431365
transform -1 0 2576 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1458_
timestamp 1698431365
transform -1 0 2576 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1459_
timestamp 1698431365
transform -1 0 3920 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1460_
timestamp 1698431365
transform -1 0 2576 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1461_
timestamp 1698431365
transform -1 0 3248 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1462_
timestamp 1698431365
transform -1 0 3920 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1463_
timestamp 1698431365
transform -1 0 3360 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1464_
timestamp 1698431365
transform -1 0 4032 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1465_
timestamp 1698431365
transform 1 0 2688 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1466_
timestamp 1698431365
transform -1 0 4032 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1467_
timestamp 1698431365
transform -1 0 2576 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1468_
timestamp 1698431365
transform 1 0 3248 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1469_
timestamp 1698431365
transform -1 0 5152 0 1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1470_
timestamp 1698431365
transform -1 0 2576 0 -1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1471_
timestamp 1698431365
transform -1 0 3248 0 -1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1472_
timestamp 1698431365
transform -1 0 2576 0 1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1473_
timestamp 1698431365
transform -1 0 3920 0 1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1474_
timestamp 1698431365
transform 1 0 2688 0 -1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1475_
timestamp 1698431365
transform -1 0 4032 0 -1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1476_
timestamp 1698431365
transform -1 0 2576 0 -1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1477_
timestamp 1698431365
transform 1 0 2576 0 -1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1478_
timestamp 1698431365
transform -1 0 4592 0 -1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1479_
timestamp 1698431365
transform -1 0 2576 0 1 68992
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1480_
timestamp 1698431365
transform -1 0 3248 0 1 68992
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1481_
timestamp 1698431365
transform 1 0 2688 0 -1 72128
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1482_
timestamp 1698431365
transform -1 0 4032 0 -1 72128
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1483_
timestamp 1698431365
transform -1 0 5152 0 -1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1484_
timestamp 1698431365
transform -1 0 5152 0 1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1485_
timestamp 1698431365
transform -1 0 5152 0 -1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1486_
timestamp 1698431365
transform -1 0 5152 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1487_
timestamp 1698431365
transform -1 0 5152 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 27776 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0674__I
timestamp 1698431365
transform -1 0 40096 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0678__I
timestamp 1698431365
transform 1 0 44912 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0681__A2
timestamp 1698431365
transform 1 0 37072 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0689__A1
timestamp 1698431365
transform -1 0 41552 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0689__A3
timestamp 1698431365
transform 1 0 46928 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0690__A1
timestamp 1698431365
transform -1 0 52640 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0690__B
timestamp 1698431365
transform 1 0 43008 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0694__A2
timestamp 1698431365
transform 1 0 45920 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0696__I
timestamp 1698431365
transform 1 0 70560 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0697__I
timestamp 1698431365
transform 1 0 71680 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0699__I
timestamp 1698431365
transform 1 0 51856 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0700__I
timestamp 1698431365
transform 1 0 50736 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0701__I
timestamp 1698431365
transform 1 0 47040 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0702__A1
timestamp 1698431365
transform -1 0 71232 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0702__A2
timestamp 1698431365
transform -1 0 70784 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0702__A3
timestamp 1698431365
transform 1 0 70112 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0702__A4
timestamp 1698431365
transform -1 0 70336 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0707__I
timestamp 1698431365
transform -1 0 69888 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0708__I
timestamp 1698431365
transform 1 0 67536 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0711__A1
timestamp 1698431365
transform -1 0 54992 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0713__A1
timestamp 1698431365
transform 1 0 54992 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0715__A1
timestamp 1698431365
transform 1 0 56336 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0717__A1
timestamp 1698431365
transform 1 0 57120 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0720__I
timestamp 1698431365
transform -1 0 72576 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0723__A1
timestamp 1698431365
transform 1 0 74592 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0723__A2
timestamp 1698431365
transform 1 0 75936 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0725__A1
timestamp 1698431365
transform 1 0 78176 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0725__A2
timestamp 1698431365
transform -1 0 77280 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0727__A1
timestamp 1698431365
transform -1 0 74816 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0727__A2
timestamp 1698431365
transform 1 0 76272 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0729__A1
timestamp 1698431365
transform 1 0 75600 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0729__A2
timestamp 1698431365
transform 1 0 78064 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0736__I
timestamp 1698431365
transform 1 0 75376 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0738__A1
timestamp 1698431365
transform -1 0 71456 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0740__I
timestamp 1698431365
transform 1 0 61824 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0742__A1
timestamp 1698431365
transform 1 0 61040 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0743__B
timestamp 1698431365
transform 1 0 73136 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0744__I
timestamp 1698431365
transform 1 0 41664 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0746__I
timestamp 1698431365
transform 1 0 32256 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0747__I
timestamp 1698431365
transform 1 0 42784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0751__A1
timestamp 1698431365
transform -1 0 36960 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0756__A2
timestamp 1698431365
transform -1 0 34832 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0761__A1
timestamp 1698431365
transform 1 0 61824 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0762__B
timestamp 1698431365
transform -1 0 72800 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0763__I
timestamp 1698431365
transform 1 0 32704 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0765__A1
timestamp 1698431365
transform -1 0 34160 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0766__A2
timestamp 1698431365
transform 1 0 35056 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0772__A1
timestamp 1698431365
transform -1 0 61376 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0773__B
timestamp 1698431365
transform -1 0 73248 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0774__I
timestamp 1698431365
transform -1 0 34160 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0776__A1
timestamp 1698431365
transform -1 0 35056 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0777__A2
timestamp 1698431365
transform 1 0 36960 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0781__A1
timestamp 1698431365
transform -1 0 71904 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0784__A1
timestamp 1698431365
transform -1 0 61600 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0785__B
timestamp 1698431365
transform 1 0 71680 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0786__I
timestamp 1698431365
transform -1 0 33040 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0788__A1
timestamp 1698431365
transform -1 0 34944 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0789__A2
timestamp 1698431365
transform 1 0 37072 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0793__A1
timestamp 1698431365
transform -1 0 73472 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0797__A1
timestamp 1698431365
transform 1 0 62272 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0798__A1
timestamp 1698431365
transform 1 0 64064 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0798__B
timestamp 1698431365
transform -1 0 62944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0800__I
timestamp 1698431365
transform 1 0 32480 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0803__A1
timestamp 1698431365
transform -1 0 34608 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0806__A2
timestamp 1698431365
transform 1 0 37408 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0807__A1
timestamp 1698431365
transform -1 0 37296 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0809__A1
timestamp 1698431365
transform -1 0 73920 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0811__A1
timestamp 1698431365
transform 1 0 63392 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0812__A1
timestamp 1698431365
transform -1 0 64736 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0813__I
timestamp 1698431365
transform 1 0 34048 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0815__A1
timestamp 1698431365
transform -1 0 35504 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0816__A2
timestamp 1698431365
transform 1 0 39312 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0817__A1
timestamp 1698431365
transform 1 0 34832 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0819__I
timestamp 1698431365
transform 1 0 71456 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0821__A1
timestamp 1698431365
transform 1 0 72688 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0823__A1
timestamp 1698431365
transform 1 0 64960 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0824__B
timestamp 1698431365
transform -1 0 71008 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0825__I
timestamp 1698431365
transform -1 0 33600 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0827__A1
timestamp 1698431365
transform -1 0 34048 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0828__A2
timestamp 1698431365
transform 1 0 39648 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0829__A1
timestamp 1698431365
transform 1 0 34720 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0832__A1
timestamp 1698431365
transform -1 0 73472 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0835__A1
timestamp 1698431365
transform 1 0 65856 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0836__B
timestamp 1698431365
transform 1 0 72464 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0837__I
timestamp 1698431365
transform -1 0 34944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0839__A1
timestamp 1698431365
transform -1 0 34496 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0840__A2
timestamp 1698431365
transform 1 0 40096 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0844__A1
timestamp 1698431365
transform -1 0 72128 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0848__A1
timestamp 1698431365
transform 1 0 65408 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0849__B
timestamp 1698431365
transform -1 0 71344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0851__I
timestamp 1698431365
transform 1 0 42336 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0854__A1
timestamp 1698431365
transform -1 0 40544 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0857__A2
timestamp 1698431365
transform 1 0 40320 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0858__A1
timestamp 1698431365
transform -1 0 39312 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0860__A1
timestamp 1698431365
transform -1 0 73248 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0862__A1
timestamp 1698431365
transform 1 0 67088 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0863__B
timestamp 1698431365
transform 1 0 71680 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0864__I
timestamp 1698431365
transform 1 0 38528 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0866__A1
timestamp 1698431365
transform -1 0 42000 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0867__A2
timestamp 1698431365
transform 1 0 42560 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0868__A1
timestamp 1698431365
transform 1 0 39088 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0871__A1
timestamp 1698431365
transform -1 0 73584 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0873__A1
timestamp 1698431365
transform 1 0 67424 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0874__B
timestamp 1698431365
transform -1 0 75152 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0875__I
timestamp 1698431365
transform 1 0 39648 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0877__A1
timestamp 1698431365
transform -1 0 42224 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0878__A2
timestamp 1698431365
transform 1 0 42448 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0879__A1
timestamp 1698431365
transform -1 0 40992 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0881__I
timestamp 1698431365
transform 1 0 75152 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0883__A1
timestamp 1698431365
transform -1 0 72800 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0885__I
timestamp 1698431365
transform 1 0 68992 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0887__A1
timestamp 1698431365
transform 1 0 69664 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0888__B
timestamp 1698431365
transform -1 0 73024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0889__I
timestamp 1698431365
transform 1 0 39424 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0891__A1
timestamp 1698431365
transform -1 0 41216 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0892__A2
timestamp 1698431365
transform 1 0 43008 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0893__A1
timestamp 1698431365
transform 1 0 40656 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0896__A1
timestamp 1698431365
transform -1 0 74144 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0900__A1
timestamp 1698431365
transform 1 0 69216 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0901__B
timestamp 1698431365
transform 1 0 71680 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0903__I
timestamp 1698431365
transform -1 0 36176 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0906__A1
timestamp 1698431365
transform -1 0 42672 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0909__A2
timestamp 1698431365
transform 1 0 44576 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0910__A1
timestamp 1698431365
transform 1 0 48496 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0912__A1
timestamp 1698431365
transform -1 0 74816 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0914__A1
timestamp 1698431365
transform -1 0 68208 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0915__B
timestamp 1698431365
transform -1 0 72016 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0916__I
timestamp 1698431365
transform 1 0 37072 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0918__A1
timestamp 1698431365
transform -1 0 44016 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0919__A2
timestamp 1698431365
transform 1 0 44912 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0920__A1
timestamp 1698431365
transform -1 0 44464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0923__A1
timestamp 1698431365
transform -1 0 76608 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0925__A1
timestamp 1698431365
transform 1 0 71904 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0926__B
timestamp 1698431365
transform 1 0 72128 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0927__I
timestamp 1698431365
transform -1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0929__A1
timestamp 1698431365
transform -1 0 45808 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0930__A2
timestamp 1698431365
transform 1 0 45808 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0931__A1
timestamp 1698431365
transform 1 0 48496 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0934__A1
timestamp 1698431365
transform -1 0 71904 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0937__A1
timestamp 1698431365
transform 1 0 71344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0938__B
timestamp 1698431365
transform -1 0 74032 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0939__I
timestamp 1698431365
transform 1 0 36288 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0941__A1
timestamp 1698431365
transform -1 0 44352 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0942__A2
timestamp 1698431365
transform 1 0 46592 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0947__A1
timestamp 1698431365
transform -1 0 70224 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0948__I
timestamp 1698431365
transform -1 0 70560 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0951__I
timestamp 1698431365
transform 1 0 70560 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0953__A1
timestamp 1698431365
transform 1 0 71344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0955__I
timestamp 1698431365
transform 1 0 45360 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0957__I
timestamp 1698431365
transform 1 0 52752 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0961__A1
timestamp 1698431365
transform -1 0 49504 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0966__A2
timestamp 1698431365
transform 1 0 50288 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0969__A1
timestamp 1698431365
transform -1 0 71904 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0971__A1
timestamp 1698431365
transform 1 0 72352 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0973__I
timestamp 1698431365
transform 1 0 49728 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0975__A1
timestamp 1698431365
transform 1 0 48496 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0976__A2
timestamp 1698431365
transform 1 0 51856 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0980__A1
timestamp 1698431365
transform -1 0 71456 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0982__A1
timestamp 1698431365
transform -1 0 71344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0984__I
timestamp 1698431365
transform 1 0 47040 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0986__A1
timestamp 1698431365
transform -1 0 49056 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0987__A2
timestamp 1698431365
transform 1 0 50064 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0988__A1
timestamp 1698431365
transform -1 0 48384 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0991__A1
timestamp 1698431365
transform -1 0 77392 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0994__A1
timestamp 1698431365
transform -1 0 72016 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0996__I
timestamp 1698431365
transform 1 0 45360 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0998__A1
timestamp 1698431365
transform 1 0 48048 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0999__A2
timestamp 1698431365
transform 1 0 48944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1003__A1
timestamp 1698431365
transform -1 0 76496 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1007__A1
timestamp 1698431365
transform 1 0 73248 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1010__I
timestamp 1698431365
transform 1 0 47488 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1013__A1
timestamp 1698431365
transform -1 0 50624 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1016__A2
timestamp 1698431365
transform 1 0 51744 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1017__A1
timestamp 1698431365
transform -1 0 49056 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1019__A1
timestamp 1698431365
transform -1 0 76272 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1021__A1
timestamp 1698431365
transform -1 0 73024 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1023__I
timestamp 1698431365
transform 1 0 45472 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1025__A1
timestamp 1698431365
transform -1 0 50176 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1026__A2
timestamp 1698431365
transform 1 0 50736 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1027__A1
timestamp 1698431365
transform -1 0 50736 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1029__I
timestamp 1698431365
transform 1 0 74704 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1030__A1
timestamp 1698431365
transform -1 0 72800 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1032__A1
timestamp 1698431365
transform 1 0 75600 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1034__I
timestamp 1698431365
transform 1 0 45360 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1036__A1
timestamp 1698431365
transform 1 0 50624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1037__A2
timestamp 1698431365
transform 1 0 53760 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1038__A1
timestamp 1698431365
transform -1 0 49616 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1041__A1
timestamp 1698431365
transform -1 0 78288 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1044__A1
timestamp 1698431365
transform -1 0 74480 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1046__I
timestamp 1698431365
transform 1 0 44688 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1048__A1
timestamp 1698431365
transform 1 0 50176 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1049__A2
timestamp 1698431365
transform 1 0 50288 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1050__A1
timestamp 1698431365
transform -1 0 49504 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1053__A1
timestamp 1698431365
transform -1 0 71456 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1057__A1
timestamp 1698431365
transform -1 0 74032 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1060__I
timestamp 1698431365
transform -1 0 44688 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1063__A1
timestamp 1698431365
transform 1 0 51968 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1066__A2
timestamp 1698431365
transform 1 0 56000 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1069__A1
timestamp 1698431365
transform -1 0 77392 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1071__A1
timestamp 1698431365
transform -1 0 76048 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1073__I
timestamp 1698431365
transform -1 0 44240 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1075__A1
timestamp 1698431365
transform -1 0 53760 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1076__A2
timestamp 1698431365
transform 1 0 57120 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1079__I
timestamp 1698431365
transform 1 0 76048 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1080__A1
timestamp 1698431365
transform -1 0 77728 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1082__A1
timestamp 1698431365
transform 1 0 78176 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1084__I
timestamp 1698431365
transform -1 0 45136 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1086__A1
timestamp 1698431365
transform -1 0 52976 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1087__A2
timestamp 1698431365
transform 1 0 56672 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1090__I
timestamp 1698431365
transform 1 0 75600 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1091__A1
timestamp 1698431365
transform -1 0 76608 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1093__I
timestamp 1698431365
transform -1 0 69104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1094__A1
timestamp 1698431365
transform 1 0 78064 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1096__I
timestamp 1698431365
transform -1 0 44464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1098__A1
timestamp 1698431365
transform 1 0 52752 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1099__A2
timestamp 1698431365
transform 1 0 52752 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1103__A1
timestamp 1698431365
transform -1 0 73024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1107__A1
timestamp 1698431365
transform -1 0 78288 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1110__I
timestamp 1698431365
transform -1 0 44240 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1113__A1
timestamp 1698431365
transform -1 0 54096 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1116__A2
timestamp 1698431365
transform 1 0 57568 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1117__A1
timestamp 1698431365
transform 1 0 56672 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1119__A1
timestamp 1698431365
transform 1 0 78176 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1121__A1
timestamp 1698431365
transform 1 0 78176 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1123__I
timestamp 1698431365
transform -1 0 44464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1125__A1
timestamp 1698431365
transform 1 0 54320 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1126__A2
timestamp 1698431365
transform 1 0 56448 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1127__A1
timestamp 1698431365
transform 1 0 56672 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1129__A1
timestamp 1698431365
transform -1 0 73472 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1131__A1
timestamp 1698431365
transform -1 0 75824 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1133__I
timestamp 1698431365
transform 1 0 44240 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1135__A1
timestamp 1698431365
transform -1 0 55552 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1136__A2
timestamp 1698431365
transform 1 0 56896 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1137__A1
timestamp 1698431365
transform 1 0 57120 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1139__A1
timestamp 1698431365
transform 1 0 74592 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1141__A1
timestamp 1698431365
transform 1 0 74032 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1143__I
timestamp 1698431365
transform 1 0 45360 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1145__A1
timestamp 1698431365
transform 1 0 55552 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1146__A2
timestamp 1698431365
transform 1 0 55888 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1147__A1
timestamp 1698431365
transform 1 0 57120 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1147__B1
timestamp 1698431365
transform -1 0 56560 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1148__A1
timestamp 1698431365
transform 1 0 43568 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1149__A1
timestamp 1698431365
transform -1 0 41216 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1150__A1
timestamp 1698431365
transform 1 0 44016 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1151__A1
timestamp 1698431365
transform 1 0 43232 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1152__A1
timestamp 1698431365
transform -1 0 74816 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1156__A1
timestamp 1698431365
transform -1 0 26320 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1160__A1
timestamp 1698431365
transform -1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1162__I
timestamp 1698431365
transform 1 0 21504 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1163__I
timestamp 1698431365
transform -1 0 19488 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1164__A1
timestamp 1698431365
transform -1 0 19264 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1167__A1
timestamp 1698431365
transform 1 0 17696 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1170__A1
timestamp 1698431365
transform -1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1173__A1
timestamp 1698431365
transform -1 0 13776 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1178__I
timestamp 1698431365
transform 1 0 20832 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1179__A1
timestamp 1698431365
transform -1 0 21056 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1182__A1
timestamp 1698431365
transform 1 0 21392 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1185__A1
timestamp 1698431365
transform 1 0 20608 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1188__A1
timestamp 1698431365
transform 1 0 20720 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1190__A1
timestamp 1698431365
transform -1 0 27888 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1193__A1
timestamp 1698431365
transform -1 0 24416 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1195__I
timestamp 1698431365
transform 1 0 23072 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1210__I
timestamp 1698431365
transform -1 0 13776 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1211__I
timestamp 1698431365
transform 1 0 24640 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1223__A1
timestamp 1698431365
transform 1 0 32256 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1226__A1
timestamp 1698431365
transform -1 0 27552 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1228__I
timestamp 1698431365
transform -1 0 32928 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1243__I
timestamp 1698431365
transform 1 0 32256 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1255__A1
timestamp 1698431365
transform 1 0 25312 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1260__A1
timestamp 1698431365
transform 1 0 23968 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1262__A1
timestamp 1698431365
transform 1 0 23520 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1264__A1
timestamp 1698431365
transform 1 0 23072 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1266__A1
timestamp 1698431365
transform 1 0 24640 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1270__A1
timestamp 1698431365
transform 1 0 18032 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1271__A1
timestamp 1698431365
transform 1 0 18368 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1272__A1
timestamp 1698431365
transform 1 0 19264 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1273__A1
timestamp 1698431365
transform 1 0 22288 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1274__A1
timestamp 1698431365
transform 1 0 15568 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1275__A1
timestamp 1698431365
transform -1 0 18592 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1276__A1
timestamp 1698431365
transform 1 0 20608 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1280__A1
timestamp 1698431365
transform 1 0 18592 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1281__A1
timestamp 1698431365
transform -1 0 20608 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1282__A1
timestamp 1698431365
transform 1 0 18144 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1283__A1
timestamp 1698431365
transform 1 0 20384 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1284__A1
timestamp 1698431365
transform 1 0 17696 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1285__A1
timestamp 1698431365
transform 1 0 23968 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1286__A1
timestamp 1698431365
transform 1 0 20160 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1287__A1
timestamp 1698431365
transform 1 0 22960 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1290__A1
timestamp 1698431365
transform 1 0 25984 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1291__A1
timestamp 1698431365
transform -1 0 28000 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1292__A1
timestamp 1698431365
transform 1 0 25312 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1293__A1
timestamp 1698431365
transform -1 0 30576 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1294__A1
timestamp 1698431365
transform 1 0 23632 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1295__A1
timestamp 1698431365
transform 1 0 31248 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1296__A1
timestamp 1698431365
transform 1 0 24080 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1307__A1
timestamp 1698431365
transform -1 0 34272 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1313__A1
timestamp 1698431365
transform -1 0 26432 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1315__A1
timestamp 1698431365
transform 1 0 30128 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1317__A1
timestamp 1698431365
transform 1 0 27216 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1319__A1
timestamp 1698431365
transform 1 0 30128 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1333__A1
timestamp 1698431365
transform -1 0 40432 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1335__A1
timestamp 1698431365
transform -1 0 41888 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1337__A1
timestamp 1698431365
transform 1 0 39424 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1339__A1
timestamp 1698431365
transform 1 0 43904 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1340__S
timestamp 1698431365
transform -1 0 37744 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1342__A1
timestamp 1698431365
transform -1 0 25872 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1343__I
timestamp 1698431365
transform 1 0 8288 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1345__A1
timestamp 1698431365
transform 1 0 31248 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1347__I
timestamp 1698431365
transform 1 0 14896 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1348__A1
timestamp 1698431365
transform -1 0 13328 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1351__A1
timestamp 1698431365
transform -1 0 11200 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1354__A1
timestamp 1698431365
transform 1 0 12432 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1357__A1
timestamp 1698431365
transform 1 0 14448 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1359__I
timestamp 1698431365
transform -1 0 8064 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1362__I
timestamp 1698431365
transform -1 0 13776 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1363__A1
timestamp 1698431365
transform -1 0 13216 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1366__A1
timestamp 1698431365
transform -1 0 12208 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1369__A1
timestamp 1698431365
transform -1 0 10304 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1372__A1
timestamp 1698431365
transform -1 0 12656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1411__CLK
timestamp 1698431365
transform 1 0 32480 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1412__CLK
timestamp 1698431365
transform 1 0 32368 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1416__CLK
timestamp 1698431365
transform 1 0 34496 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1417__CLK
timestamp 1698431365
transform 1 0 35168 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1430__CLK
timestamp 1698431365
transform 1 0 40992 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1471__I
timestamp 1698431365
transform 1 0 3472 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698431365
transform -1 0 31472 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_0__f_clk_I
timestamp 1698431365
transform -1 0 20832 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_1__f_clk_I
timestamp 1698431365
transform 1 0 26768 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_2__f_clk_I
timestamp 1698431365
transform 1 0 23744 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_3__f_clk_I
timestamp 1698431365
transform 1 0 27552 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_4__f_clk_I
timestamp 1698431365
transform 1 0 32480 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_5__f_clk_I
timestamp 1698431365
transform 1 0 36400 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_6__f_clk_I
timestamp 1698431365
transform 1 0 28112 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_7__f_clk_I
timestamp 1698431365
transform -1 0 32032 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout331_I
timestamp 1698431365
transform -1 0 4368 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout332_I
timestamp 1698431365
transform 1 0 4480 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout334_I
timestamp 1698431365
transform -1 0 2016 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout335_I
timestamp 1698431365
transform 1 0 4928 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout336_I
timestamp 1698431365
transform -1 0 4368 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout338_I
timestamp 1698431365
transform 1 0 2912 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout341_I
timestamp 1698431365
transform -1 0 2016 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout342_I
timestamp 1698431365
transform 1 0 5376 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform -1 0 23968 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform -1 0 28336 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform -1 0 31360 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform -1 0 27888 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform -1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform -1 0 30128 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform -1 0 31024 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698431365
transform -1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698431365
transform -1 0 30912 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698431365
transform -1 0 33600 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698431365
transform -1 0 32480 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698431365
transform -1 0 20160 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698431365
transform -1 0 33376 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1698431365
transform -1 0 33376 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1698431365
transform -1 0 35952 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1698431365
transform 1 0 51072 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1698431365
transform 1 0 51520 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1698431365
transform 1 0 45472 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1698431365
transform 1 0 52528 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1698431365
transform 1 0 53536 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1698431365
transform -1 0 47712 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input22_I
timestamp 1698431365
transform 1 0 49728 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input23_I
timestamp 1698431365
transform -1 0 19712 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input24_I
timestamp 1698431365
transform 1 0 49056 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input25_I
timestamp 1698431365
transform -1 0 49728 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input26_I
timestamp 1698431365
transform -1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input27_I
timestamp 1698431365
transform -1 0 21504 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input28_I
timestamp 1698431365
transform -1 0 21280 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input29_I
timestamp 1698431365
transform -1 0 30576 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input30_I
timestamp 1698431365
transform -1 0 24416 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input31_I
timestamp 1698431365
transform -1 0 25424 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input32_I
timestamp 1698431365
transform -1 0 22848 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input33_I
timestamp 1698431365
transform 1 0 51184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input34_I
timestamp 1698431365
transform -1 0 3808 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input35_I
timestamp 1698431365
transform -1 0 6272 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input36_I
timestamp 1698431365
transform -1 0 6720 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input37_I
timestamp 1698431365
transform -1 0 7728 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input38_I
timestamp 1698431365
transform -1 0 10304 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input39_I
timestamp 1698431365
transform -1 0 7168 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input40_I
timestamp 1698431365
transform -1 0 6720 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input41_I
timestamp 1698431365
transform -1 0 10304 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input42_I
timestamp 1698431365
transform -1 0 10976 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input43_I
timestamp 1698431365
transform -1 0 11760 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input44_I
timestamp 1698431365
transform -1 0 11872 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input45_I
timestamp 1698431365
transform -1 0 3360 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input46_I
timestamp 1698431365
transform -1 0 12768 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input47_I
timestamp 1698431365
transform -1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input48_I
timestamp 1698431365
transform -1 0 11536 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input49_I
timestamp 1698431365
transform -1 0 16576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input50_I
timestamp 1698431365
transform -1 0 15344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input51_I
timestamp 1698431365
transform -1 0 20608 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input52_I
timestamp 1698431365
transform -1 0 19040 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input53_I
timestamp 1698431365
transform -1 0 14784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input54_I
timestamp 1698431365
transform -1 0 21952 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input55_I
timestamp 1698431365
transform -1 0 23520 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input56_I
timestamp 1698431365
transform -1 0 4816 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input57_I
timestamp 1698431365
transform -1 0 22400 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input58_I
timestamp 1698431365
transform -1 0 19264 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input59_I
timestamp 1698431365
transform -1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input60_I
timestamp 1698431365
transform -1 0 4368 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input61_I
timestamp 1698431365
transform -1 0 7616 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input62_I
timestamp 1698431365
transform -1 0 6272 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input63_I
timestamp 1698431365
transform -1 0 5376 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input64_I
timestamp 1698431365
transform -1 0 5824 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input65_I
timestamp 1698431365
transform -1 0 7168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input66_I
timestamp 1698431365
transform 1 0 51632 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input67_I
timestamp 1698431365
transform -1 0 52192 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input68_I
timestamp 1698431365
transform 1 0 54208 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input69_I
timestamp 1698431365
transform -1 0 53312 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input70_I
timestamp 1698431365
transform -1 0 2240 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input71_I
timestamp 1698431365
transform 1 0 2464 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input72_I
timestamp 1698431365
transform 1 0 2464 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input73_I
timestamp 1698431365
transform 1 0 2464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input74_I
timestamp 1698431365
transform 1 0 2464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input75_I
timestamp 1698431365
transform 1 0 2464 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input76_I
timestamp 1698431365
transform 1 0 2464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input77_I
timestamp 1698431365
transform 1 0 2464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input78_I
timestamp 1698431365
transform 1 0 2464 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input79_I
timestamp 1698431365
transform 1 0 2464 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input80_I
timestamp 1698431365
transform 1 0 2464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input81_I
timestamp 1698431365
transform 1 0 2464 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input82_I
timestamp 1698431365
transform 1 0 2464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input83_I
timestamp 1698431365
transform 1 0 2464 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input84_I
timestamp 1698431365
transform 1 0 2464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input85_I
timestamp 1698431365
transform 1 0 2464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input86_I
timestamp 1698431365
transform 1 0 2464 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input87_I
timestamp 1698431365
transform 1 0 2464 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input88_I
timestamp 1698431365
transform 1 0 2464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input89_I
timestamp 1698431365
transform 1 0 2464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input90_I
timestamp 1698431365
transform 1 0 2464 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input91_I
timestamp 1698431365
transform 1 0 2464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input92_I
timestamp 1698431365
transform 1 0 2464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input93_I
timestamp 1698431365
transform 1 0 2464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input94_I
timestamp 1698431365
transform 1 0 2464 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input95_I
timestamp 1698431365
transform 1 0 2464 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input96_I
timestamp 1698431365
transform 1 0 2464 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input97_I
timestamp 1698431365
transform 1 0 2464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input98_I
timestamp 1698431365
transform 1 0 2464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input99_I
timestamp 1698431365
transform 1 0 2464 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input100_I
timestamp 1698431365
transform 1 0 2464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input101_I
timestamp 1698431365
transform 1 0 2464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input102_I
timestamp 1698431365
transform -1 0 73696 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input103_I
timestamp 1698431365
transform -1 0 78400 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input104_I
timestamp 1698431365
transform -1 0 77728 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input105_I
timestamp 1698431365
transform -1 0 77504 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input106_I
timestamp 1698431365
transform -1 0 77728 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input107_I
timestamp 1698431365
transform -1 0 77728 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input108_I
timestamp 1698431365
transform -1 0 77504 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input109_I
timestamp 1698431365
transform -1 0 77728 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input110_I
timestamp 1698431365
transform -1 0 77728 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input111_I
timestamp 1698431365
transform -1 0 77504 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input112_I
timestamp 1698431365
transform -1 0 77728 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input113_I
timestamp 1698431365
transform -1 0 77504 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input114_I
timestamp 1698431365
transform -1 0 77728 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input115_I
timestamp 1698431365
transform -1 0 77504 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input116_I
timestamp 1698431365
transform -1 0 77728 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input117_I
timestamp 1698431365
transform -1 0 77504 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input118_I
timestamp 1698431365
transform -1 0 77728 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input119_I
timestamp 1698431365
transform -1 0 77504 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input120_I
timestamp 1698431365
transform -1 0 77728 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input121_I
timestamp 1698431365
transform -1 0 77728 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input122_I
timestamp 1698431365
transform -1 0 77504 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input123_I
timestamp 1698431365
transform -1 0 75376 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input124_I
timestamp 1698431365
transform -1 0 74144 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input125_I
timestamp 1698431365
transform -1 0 77728 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input126_I
timestamp 1698431365
transform -1 0 77056 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input127_I
timestamp 1698431365
transform 1 0 77952 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input128_I
timestamp 1698431365
transform -1 0 77728 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input129_I
timestamp 1698431365
transform -1 0 77728 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input130_I
timestamp 1698431365
transform -1 0 77728 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input131_I
timestamp 1698431365
transform -1 0 77728 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input132_I
timestamp 1698431365
transform -1 0 77728 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input133_I
timestamp 1698431365
transform -1 0 77728 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input134_I
timestamp 1698431365
transform -1 0 77728 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input135_I
timestamp 1698431365
transform -1 0 77280 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input136_I
timestamp 1698431365
transform -1 0 74928 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input137_I
timestamp 1698431365
transform -1 0 77280 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input138_I
timestamp 1698431365
transform -1 0 77056 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input139_I
timestamp 1698431365
transform -1 0 77728 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input140_I
timestamp 1698431365
transform -1 0 75152 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input141_I
timestamp 1698431365
transform -1 0 76832 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input142_I
timestamp 1698431365
transform -1 0 77280 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input143_I
timestamp 1698431365
transform -1 0 78400 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input144_I
timestamp 1698431365
transform -1 0 78400 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input145_I
timestamp 1698431365
transform -1 0 71904 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input146_I
timestamp 1698431365
transform -1 0 72352 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input147_I
timestamp 1698431365
transform -1 0 77280 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input148_I
timestamp 1698431365
transform -1 0 71456 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input149_I
timestamp 1698431365
transform -1 0 72688 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input150_I
timestamp 1698431365
transform -1 0 76608 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input151_I
timestamp 1698431365
transform -1 0 75152 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input152_I
timestamp 1698431365
transform -1 0 74928 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input153_I
timestamp 1698431365
transform -1 0 71008 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input154_I
timestamp 1698431365
transform -1 0 73472 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input155_I
timestamp 1698431365
transform -1 0 74704 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input156_I
timestamp 1698431365
transform -1 0 77728 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input157_I
timestamp 1698431365
transform -1 0 72576 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input158_I
timestamp 1698431365
transform -1 0 77280 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input159_I
timestamp 1698431365
transform -1 0 77392 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input160_I
timestamp 1698431365
transform -1 0 77056 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input161_I
timestamp 1698431365
transform -1 0 75376 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input162_I
timestamp 1698431365
transform -1 0 77728 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input163_I
timestamp 1698431365
transform -1 0 77728 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input164_I
timestamp 1698431365
transform -1 0 77728 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input165_I
timestamp 1698431365
transform -1 0 77728 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input166_I
timestamp 1698431365
transform -1 0 77728 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input167_I
timestamp 1698431365
transform -1 0 77728 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input168_I
timestamp 1698431365
transform -1 0 34160 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input169_I
timestamp 1698431365
transform 1 0 42000 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input170_I
timestamp 1698431365
transform -1 0 41552 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input171_I
timestamp 1698431365
transform 1 0 42448 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input172_I
timestamp 1698431365
transform -1 0 43456 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input173_I
timestamp 1698431365
transform -1 0 44016 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input174_I
timestamp 1698431365
transform 1 0 46032 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input175_I
timestamp 1698431365
transform -1 0 44464 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input176_I
timestamp 1698431365
transform 1 0 46480 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input177_I
timestamp 1698431365
transform 1 0 48048 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input178_I
timestamp 1698431365
transform -1 0 46928 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input179_I
timestamp 1698431365
transform -1 0 34832 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input180_I
timestamp 1698431365
transform 1 0 48496 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input181_I
timestamp 1698431365
transform -1 0 49168 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input182_I
timestamp 1698431365
transform 1 0 50736 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input183_I
timestamp 1698431365
transform -1 0 49616 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input184_I
timestamp 1698431365
transform 1 0 51184 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input185_I
timestamp 1698431365
transform -1 0 51856 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input186_I
timestamp 1698431365
transform -1 0 52864 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input187_I
timestamp 1698431365
transform -1 0 52304 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input188_I
timestamp 1698431365
transform 1 0 55104 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input189_I
timestamp 1698431365
transform -1 0 53648 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input190_I
timestamp 1698431365
transform -1 0 35504 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input191_I
timestamp 1698431365
transform -1 0 54544 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input192_I
timestamp 1698431365
transform -1 0 55440 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input193_I
timestamp 1698431365
transform 1 0 36400 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input194_I
timestamp 1698431365
transform 1 0 37296 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input195_I
timestamp 1698431365
transform -1 0 37520 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input196_I
timestamp 1698431365
transform 1 0 38864 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input197_I
timestamp 1698431365
transform -1 0 37968 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input198_I
timestamp 1698431365
transform 1 0 39984 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input199_I
timestamp 1698431365
transform 1 0 40880 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input200_I
timestamp 1698431365
transform -1 0 32816 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input201_I
timestamp 1698431365
transform -1 0 59248 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input202_I
timestamp 1698431365
transform -1 0 65072 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input203_I
timestamp 1698431365
transform 1 0 66416 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input204_I
timestamp 1698431365
transform -1 0 67088 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input205_I
timestamp 1698431365
transform -1 0 67648 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input206_I
timestamp 1698431365
transform 1 0 68432 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input207_I
timestamp 1698431365
transform -1 0 69104 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input208_I
timestamp 1698431365
transform -1 0 70112 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input209_I
timestamp 1698431365
transform -1 0 70784 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input210_I
timestamp 1698431365
transform -1 0 71456 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input211_I
timestamp 1698431365
transform -1 0 72016 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input212_I
timestamp 1698431365
transform 1 0 61264 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input213_I
timestamp 1698431365
transform 1 0 73360 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input214_I
timestamp 1698431365
transform -1 0 72464 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input215_I
timestamp 1698431365
transform -1 0 74032 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input216_I
timestamp 1698431365
transform -1 0 74592 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input217_I
timestamp 1698431365
transform -1 0 75152 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input218_I
timestamp 1698431365
transform -1 0 75824 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input219_I
timestamp 1698431365
transform -1 0 75040 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input220_I
timestamp 1698431365
transform -1 0 74592 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input221_I
timestamp 1698431365
transform -1 0 76160 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input222_I
timestamp 1698431365
transform -1 0 76608 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input223_I
timestamp 1698431365
transform 1 0 62608 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input224_I
timestamp 1698431365
transform -1 0 76496 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input225_I
timestamp 1698431365
transform -1 0 75488 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input226_I
timestamp 1698431365
transform 1 0 61712 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input227_I
timestamp 1698431365
transform 1 0 62160 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input228_I
timestamp 1698431365
transform 1 0 63056 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input229_I
timestamp 1698431365
transform 1 0 63504 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input230_I
timestamp 1698431365
transform 1 0 63952 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input231_I
timestamp 1698431365
transform -1 0 64624 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input232_I
timestamp 1698431365
transform 1 0 65968 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output233_I
timestamp 1698431365
transform 1 0 14336 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output234_I
timestamp 1698431365
transform -1 0 18032 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output235_I
timestamp 1698431365
transform 1 0 19824 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output236_I
timestamp 1698431365
transform 1 0 19376 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output237_I
timestamp 1698431365
transform 1 0 22960 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output238_I
timestamp 1698431365
transform 1 0 24752 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output239_I
timestamp 1698431365
transform 1 0 25200 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output240_I
timestamp 1698431365
transform 1 0 14112 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output241_I
timestamp 1698431365
transform 1 0 13552 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output242_I
timestamp 1698431365
transform -1 0 14336 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output243_I
timestamp 1698431365
transform -1 0 13440 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output244_I
timestamp 1698431365
transform -1 0 14112 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output245_I
timestamp 1698431365
transform -1 0 14784 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output246_I
timestamp 1698431365
transform 1 0 18032 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output247_I
timestamp 1698431365
transform -1 0 17248 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output248_I
timestamp 1698431365
transform 1 0 18256 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output249_I
timestamp 1698431365
transform 1 0 52528 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output250_I
timestamp 1698431365
transform 1 0 59472 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output251_I
timestamp 1698431365
transform -1 0 60144 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output252_I
timestamp 1698431365
transform -1 0 63280 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output253_I
timestamp 1698431365
transform 1 0 65632 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output254_I
timestamp 1698431365
transform 1 0 66416 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output255_I
timestamp 1698431365
transform -1 0 63280 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output256_I
timestamp 1698431365
transform 1 0 63840 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output257_I
timestamp 1698431365
transform 1 0 67424 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output258_I
timestamp 1698431365
transform -1 0 69888 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output259_I
timestamp 1698431365
transform -1 0 67200 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output260_I
timestamp 1698431365
transform 1 0 55888 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output261_I
timestamp 1698431365
transform 1 0 67312 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output262_I
timestamp 1698431365
transform 1 0 66640 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output263_I
timestamp 1698431365
transform -1 0 67984 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output264_I
timestamp 1698431365
transform -1 0 71120 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output265_I
timestamp 1698431365
transform 1 0 71680 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output266_I
timestamp 1698431365
transform 1 0 70448 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output267_I
timestamp 1698431365
transform -1 0 71120 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output268_I
timestamp 1698431365
transform 1 0 71680 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output269_I
timestamp 1698431365
transform 1 0 70448 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output270_I
timestamp 1698431365
transform 1 0 71680 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output271_I
timestamp 1698431365
transform 1 0 53872 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output272_I
timestamp 1698431365
transform 1 0 78176 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output273_I
timestamp 1698431365
transform -1 0 74816 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output274_I
timestamp 1698431365
transform 1 0 58016 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output275_I
timestamp 1698431365
transform 1 0 61824 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output276_I
timestamp 1698431365
transform 1 0 56784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output277_I
timestamp 1698431365
transform 1 0 56000 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output278_I
timestamp 1698431365
transform 1 0 62496 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output279_I
timestamp 1698431365
transform 1 0 63504 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output280_I
timestamp 1698431365
transform 1 0 60144 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output281_I
timestamp 1698431365
transform 1 0 50624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output283_I
timestamp 1698431365
transform 1 0 4704 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output284_I
timestamp 1698431365
transform 1 0 4704 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output285_I
timestamp 1698431365
transform 1 0 4704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output324_I
timestamp 1698431365
transform 1 0 35728 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output325_I
timestamp 1698431365
transform 1 0 58464 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output326_I
timestamp 1698431365
transform 1 0 59472 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output327_I
timestamp 1698431365
transform 1 0 57456 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output328_I
timestamp 1698431365
transform 1 0 60816 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 31024 0 -1 15680
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_0__f_clk
timestamp 1698431365
transform -1 0 20384 0 1 9408
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_1__f_clk
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_2__f_clk
timestamp 1698431365
transform -1 0 23744 0 -1 18816
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_3__f_clk
timestamp 1698431365
transform -1 0 27440 0 1 17248
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_4__f_clk
timestamp 1698431365
transform -1 0 38528 0 -1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_5__f_clk
timestamp 1698431365
transform 1 0 38640 0 1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_6__f_clk
timestamp 1698431365
transform -1 0 34832 0 1 17248
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_7__f_clk
timestamp 1698431365
transform 1 0 33040 0 -1 18816
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout329
timestamp 1698431365
transform 1 0 2016 0 -1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout330
timestamp 1698431365
transform 1 0 3248 0 -1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout331
timestamp 1698431365
transform 1 0 2576 0 1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout332
timestamp 1698431365
transform -1 0 4256 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout333
timestamp 1698431365
transform -1 0 3248 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout334
timestamp 1698431365
transform 1 0 2016 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout335
timestamp 1698431365
transform -1 0 3360 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout336
timestamp 1698431365
transform 1 0 2576 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout337
timestamp 1698431365
transform 1 0 2016 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout338
timestamp 1698431365
transform -1 0 2688 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout339
timestamp 1698431365
transform -1 0 5152 0 1 72128
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout340
timestamp 1698431365
transform -1 0 6048 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout341
timestamp 1698431365
transform 1 0 2016 0 -1 72128
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout342
timestamp 1698431365
transform -1 0 2464 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_14 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2912 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_36
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_70
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_104
timestamp 1698431365
transform 1 0 12992 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_138
timestamp 1698431365
transform 1 0 16800 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_172
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_200
timestamp 1698431365
transform 1 0 23744 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_206
timestamp 1698431365
transform 1 0 24416 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_240
timestamp 1698431365
transform 1 0 28224 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_274
timestamp 1698431365
transform 1 0 32032 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_438
timestamp 1698431365
transform 1 0 50400 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_470
timestamp 1698431365
transform 1 0 53984 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_474
timestamp 1698431365
transform 1 0 54432 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_504
timestamp 1698431365
transform 1 0 57792 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_508
timestamp 1698431365
transform 1 0 58240 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_538
timestamp 1698431365
transform 1 0 61600 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_542
timestamp 1698431365
transform 1 0 62048 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_572
timestamp 1698431365
transform 1 0 65408 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_576
timestamp 1698431365
transform 1 0 65856 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_606 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 69216 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_640
timestamp 1698431365
transform 1 0 73024 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_674
timestamp 1698431365
transform 1 0 76832 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_678
timestamp 1698431365
transform 1 0 77280 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_2
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_8
timestamp 1698431365
transform 1 0 2240 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_12
timestamp 1698431365
transform 1 0 2688 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_18
timestamp 1698431365
transform 1 0 3360 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_142
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_241
timestamp 1698431365
transform 1 0 28336 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_419 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 48272 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_428
timestamp 1698431365
transform 1 0 49280 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_455
timestamp 1698431365
transform 1 0 52304 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_485
timestamp 1698431365
transform 1 0 55664 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_489
timestamp 1698431365
transform 1 0 56112 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_544
timestamp 1698431365
transform 1 0 62272 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_548
timestamp 1698431365
transform 1 0 62720 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_550
timestamp 1698431365
transform 1 0 62944 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_553
timestamp 1698431365
transform 1 0 63280 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_557
timestamp 1698431365
transform 1 0 63728 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_559
timestamp 1698431365
transform 1 0 63952 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_614
timestamp 1698431365
transform 1 0 70112 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_616
timestamp 1698431365
transform 1 0 70336 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_619
timestamp 1698431365
transform 1 0 70672 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_623
timestamp 1698431365
transform 1 0 71120 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_627
timestamp 1698431365
transform 1 0 71568 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_684
timestamp 1698431365
transform 1 0 77952 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_8
timestamp 1698431365
transform 1 0 2240 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_12 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2688 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_20
timestamp 1698431365
transform 1 0 3584 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_24
timestamp 1698431365
transform 1 0 4032 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_27
timestamp 1698431365
transform 1 0 4368 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_31
timestamp 1698431365
transform 1 0 4816 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_41
timestamp 1698431365
transform 1 0 5936 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_50
timestamp 1698431365
transform 1 0 6944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_76
timestamp 1698431365
transform 1 0 9856 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_86
timestamp 1698431365
transform 1 0 10976 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_88
timestamp 1698431365
transform 1 0 11200 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_107
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_166
timestamp 1698431365
transform 1 0 19936 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_168
timestamp 1698431365
transform 1 0 20160 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_177
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_220
timestamp 1698431365
transform 1 0 25984 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_247
timestamp 1698431365
transform 1 0 29008 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_274
timestamp 1698431365
transform 1 0 32032 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_430
timestamp 1698431365
transform 1 0 49504 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_442
timestamp 1698431365
transform 1 0 50848 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_446
timestamp 1698431365
transform 1 0 51296 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_450
timestamp 1698431365
transform 1 0 51744 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_454
timestamp 1698431365
transform 1 0 52192 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_457
timestamp 1698431365
transform 1 0 52528 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_461
timestamp 1698431365
transform 1 0 52976 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_464
timestamp 1698431365
transform 1 0 53312 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_468
timestamp 1698431365
transform 1 0 53760 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_470
timestamp 1698431365
transform 1 0 53984 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_523
timestamp 1698431365
transform 1 0 59920 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_579
timestamp 1698431365
transform 1 0 66192 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_583
timestamp 1698431365
transform 1 0 66640 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_585
timestamp 1698431365
transform 1 0 66864 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_588
timestamp 1698431365
transform 1 0 67200 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_592
timestamp 1698431365
transform 1 0 67648 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_594
timestamp 1698431365
transform 1 0 67872 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_649
timestamp 1698431365
transform 1 0 74032 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_653
timestamp 1698431365
transform 1 0 74480 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_656
timestamp 1698431365
transform 1 0 74816 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_673
timestamp 1698431365
transform 1 0 76720 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_675
timestamp 1698431365
transform 1 0 76944 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_8
timestamp 1698431365
transform 1 0 2240 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_12 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2688 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_28
timestamp 1698431365
transform 1 0 4480 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_32
timestamp 1698431365
transform 1 0 4928 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_36
timestamp 1698431365
transform 1 0 5376 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_40
timestamp 1698431365
transform 1 0 5824 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_44
timestamp 1698431365
transform 1 0 6272 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_48
timestamp 1698431365
transform 1 0 6720 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_52
timestamp 1698431365
transform 1 0 7168 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_56
timestamp 1698431365
transform 1 0 7616 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_60
timestamp 1698431365
transform 1 0 8064 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_74
timestamp 1698431365
transform 1 0 9632 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_106
timestamp 1698431365
transform 1 0 13216 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_108
timestamp 1698431365
transform 1 0 13440 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_131
timestamp 1698431365
transform 1 0 16016 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_133
timestamp 1698431365
transform 1 0 16240 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_156
timestamp 1698431365
transform 1 0 18816 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_160
timestamp 1698431365
transform 1 0 19264 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_164
timestamp 1698431365
transform 1 0 19712 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_168
timestamp 1698431365
transform 1 0 20160 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_172
timestamp 1698431365
transform 1 0 20608 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_184
timestamp 1698431365
transform 1 0 21952 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_212
timestamp 1698431365
transform 1 0 25088 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_228
timestamp 1698431365
transform 1 0 26880 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_244
timestamp 1698431365
transform 1 0 28672 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_282
timestamp 1698431365
transform 1 0 32928 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_352
timestamp 1698431365
transform 1 0 40768 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_418
timestamp 1698431365
transform 1 0 48160 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_428
timestamp 1698431365
transform 1 0 49280 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_436
timestamp 1698431365
transform 1 0 50176 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_440
timestamp 1698431365
transform 1 0 50624 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_443
timestamp 1698431365
transform 1 0 50960 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_447
timestamp 1698431365
transform 1 0 51408 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_451
timestamp 1698431365
transform 1 0 51856 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_455
timestamp 1698431365
transform 1 0 52304 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_459
timestamp 1698431365
transform 1 0 52752 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_467
timestamp 1698431365
transform 1 0 53648 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_471
timestamp 1698431365
transform 1 0 54096 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_487
timestamp 1698431365
transform 1 0 55888 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_492
timestamp 1698431365
transform 1 0 56448 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_494
timestamp 1698431365
transform 1 0 56672 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_547
timestamp 1698431365
transform 1 0 62608 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_553
timestamp 1698431365
transform 1 0 63280 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_557
timestamp 1698431365
transform 1 0 63728 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_614
timestamp 1698431365
transform 1 0 70112 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_616
timestamp 1698431365
transform 1 0 70336 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_619
timestamp 1698431365
transform 1 0 70672 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_623
timestamp 1698431365
transform 1 0 71120 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_627
timestamp 1698431365
transform 1 0 71568 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_684
timestamp 1698431365
transform 1 0 77952 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_45
timestamp 1698431365
transform 1 0 6384 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_48
timestamp 1698431365
transform 1 0 6720 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_52
timestamp 1698431365
transform 1 0 7168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_54
timestamp 1698431365
transform 1 0 7392 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_75
timestamp 1698431365
transform 1 0 9744 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_77
timestamp 1698431365
transform 1 0 9968 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_80
timestamp 1698431365
transform 1 0 10304 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_86
timestamp 1698431365
transform 1 0 10976 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_90
timestamp 1698431365
transform 1 0 11424 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_93
timestamp 1698431365
transform 1 0 11760 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_97
timestamp 1698431365
transform 1 0 12208 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_101
timestamp 1698431365
transform 1 0 12656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_115
timestamp 1698431365
transform 1 0 14224 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_117
timestamp 1698431365
transform 1 0 14448 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_151
timestamp 1698431365
transform 1 0 18256 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_155
timestamp 1698431365
transform 1 0 18704 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_158
timestamp 1698431365
transform 1 0 19040 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_168
timestamp 1698431365
transform 1 0 20160 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_172
timestamp 1698431365
transform 1 0 20608 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_177
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_179
timestamp 1698431365
transform 1 0 21392 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_188
timestamp 1698431365
transform 1 0 22400 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_218
timestamp 1698431365
transform 1 0 25760 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_234
timestamp 1698431365
transform 1 0 27552 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_244
timestamp 1698431365
transform 1 0 28672 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_247
timestamp 1698431365
transform 1 0 29008 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_274
timestamp 1698431365
transform 1 0 32032 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_317
timestamp 1698431365
transform 1 0 36848 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_424
timestamp 1698431365
transform 1 0 48832 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_428
timestamp 1698431365
transform 1 0 49280 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_432
timestamp 1698431365
transform 1 0 49728 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_449
timestamp 1698431365
transform 1 0 51632 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_453
timestamp 1698431365
transform 1 0 52080 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_457
timestamp 1698431365
transform 1 0 52528 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_489
timestamp 1698431365
transform 1 0 56112 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_493
timestamp 1698431365
transform 1 0 56560 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_497
timestamp 1698431365
transform 1 0 57008 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_513
timestamp 1698431365
transform 1 0 58800 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_517
timestamp 1698431365
transform 1 0 59248 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_521
timestamp 1698431365
transform 1 0 59696 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_579
timestamp 1698431365
transform 1 0 66192 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_587
timestamp 1698431365
transform 1 0 67088 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_591
timestamp 1698431365
transform 1 0 67536 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_649
timestamp 1698431365
transform 1 0 74032 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_653
timestamp 1698431365
transform 1 0 74480 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_664
timestamp 1698431365
transform 1 0 75712 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_683
timestamp 1698431365
transform 1 0 77840 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_687
timestamp 1698431365
transform 1 0 78288 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_8
timestamp 1698431365
transform 1 0 2240 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_12
timestamp 1698431365
transform 1 0 2688 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_44
timestamp 1698431365
transform 1 0 6272 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_60
timestamp 1698431365
transform 1 0 8064 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_67
timestamp 1698431365
transform 1 0 8848 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_69
timestamp 1698431365
transform 1 0 9072 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_76
timestamp 1698431365
transform 1 0 9856 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_80
timestamp 1698431365
transform 1 0 10304 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_90
timestamp 1698431365
transform 1 0 11424 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_94
timestamp 1698431365
transform 1 0 11872 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_98
timestamp 1698431365
transform 1 0 12320 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_102
timestamp 1698431365
transform 1 0 12768 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_120
timestamp 1698431365
transform 1 0 14784 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_122
timestamp 1698431365
transform 1 0 15008 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_131
timestamp 1698431365
transform 1 0 16016 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_133
timestamp 1698431365
transform 1 0 16240 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_136
timestamp 1698431365
transform 1 0 16576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_142
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_144
timestamp 1698431365
transform 1 0 17472 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_165
timestamp 1698431365
transform 1 0 19824 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_172
timestamp 1698431365
transform 1 0 20608 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_176
timestamp 1698431365
transform 1 0 21056 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_180
timestamp 1698431365
transform 1 0 21504 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_184
timestamp 1698431365
transform 1 0 21952 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_188
timestamp 1698431365
transform 1 0 22400 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_192
timestamp 1698431365
transform 1 0 22848 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_202
timestamp 1698431365
transform 1 0 23968 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_206
timestamp 1698431365
transform 1 0 24416 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_212
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_230
timestamp 1698431365
transform 1 0 27104 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_234
timestamp 1698431365
transform 1 0 27552 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_238
timestamp 1698431365
transform 1 0 28000 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_267
timestamp 1698431365
transform 1 0 31248 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_282
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_323
timestamp 1698431365
transform 1 0 37520 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_325
timestamp 1698431365
transform 1 0 37744 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_347
timestamp 1698431365
transform 1 0 40208 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_349
timestamp 1698431365
transform 1 0 40432 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_406
timestamp 1698431365
transform 1 0 46816 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_410
timestamp 1698431365
transform 1 0 47264 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_414
timestamp 1698431365
transform 1 0 47712 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_418
timestamp 1698431365
transform 1 0 48160 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_422 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 48608 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_486
timestamp 1698431365
transform 1 0 55776 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_492
timestamp 1698431365
transform 1 0 56448 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_524
timestamp 1698431365
transform 1 0 60032 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_527
timestamp 1698431365
transform 1 0 60368 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_559
timestamp 1698431365
transform 1 0 63952 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_562
timestamp 1698431365
transform 1 0 64288 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_578
timestamp 1698431365
transform 1 0 66080 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_582
timestamp 1698431365
transform 1 0 66528 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_611
timestamp 1698431365
transform 1 0 69776 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_627
timestamp 1698431365
transform 1 0 71568 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_632
timestamp 1698431365
transform 1 0 72128 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_685
timestamp 1698431365
transform 1 0 78064 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_687
timestamp 1698431365
transform 1 0 78288 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_8
timestamp 1698431365
transform 1 0 2240 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_12
timestamp 1698431365
transform 1 0 2688 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_28
timestamp 1698431365
transform 1 0 4480 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_32
timestamp 1698431365
transform 1 0 4928 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_69
timestamp 1698431365
transform 1 0 9072 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_73
timestamp 1698431365
transform 1 0 9520 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_107
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_162
timestamp 1698431365
transform 1 0 19488 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_171
timestamp 1698431365
transform 1 0 20496 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_177
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_179
timestamp 1698431365
transform 1 0 21392 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_209
timestamp 1698431365
transform 1 0 24752 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_215
timestamp 1698431365
transform 1 0 25424 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_219
timestamp 1698431365
transform 1 0 25872 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_242
timestamp 1698431365
transform 1 0 28448 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_244
timestamp 1698431365
transform 1 0 28672 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_252
timestamp 1698431365
transform 1 0 29568 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_260
timestamp 1698431365
transform 1 0 30464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_264
timestamp 1698431365
transform 1 0 30912 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_274
timestamp 1698431365
transform 1 0 32032 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_284
timestamp 1698431365
transform 1 0 33152 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_288
timestamp 1698431365
transform 1 0 33600 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_290
timestamp 1698431365
transform 1 0 33824 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_305
timestamp 1698431365
transform 1 0 35504 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_309
timestamp 1698431365
transform 1 0 35952 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_313
timestamp 1698431365
transform 1 0 36400 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_317
timestamp 1698431365
transform 1 0 36848 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_321
timestamp 1698431365
transform 1 0 37296 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_331
timestamp 1698431365
transform 1 0 38416 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_374
timestamp 1698431365
transform 1 0 43232 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_376
timestamp 1698431365
transform 1 0 43456 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_383
timestamp 1698431365
transform 1 0 44240 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_392
timestamp 1698431365
transform 1 0 45248 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_396
timestamp 1698431365
transform 1 0 45696 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_400
timestamp 1698431365
transform 1 0 46144 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_432
timestamp 1698431365
transform 1 0 49728 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_448
timestamp 1698431365
transform 1 0 51520 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_452
timestamp 1698431365
transform 1 0 51968 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_454
timestamp 1698431365
transform 1 0 52192 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_457
timestamp 1698431365
transform 1 0 52528 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_521
timestamp 1698431365
transform 1 0 59696 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_527
timestamp 1698431365
transform 1 0 60368 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_591
timestamp 1698431365
transform 1 0 67536 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_597
timestamp 1698431365
transform 1 0 68208 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_629
timestamp 1698431365
transform 1 0 71792 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_637
timestamp 1698431365
transform 1 0 72688 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_667
timestamp 1698431365
transform 1 0 76048 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_669
timestamp 1698431365
transform 1 0 76272 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_34
timestamp 1698431365
transform 1 0 5152 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_50
timestamp 1698431365
transform 1 0 6944 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_58
timestamp 1698431365
transform 1 0 7840 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_62
timestamp 1698431365
transform 1 0 8288 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_103
timestamp 1698431365
transform 1 0 12880 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_119
timestamp 1698431365
transform 1 0 14672 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_135
timestamp 1698431365
transform 1 0 16464 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_139
timestamp 1698431365
transform 1 0 16912 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_142
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_156
timestamp 1698431365
transform 1 0 18816 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_160
timestamp 1698431365
transform 1 0 19264 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_192
timestamp 1698431365
transform 1 0 22848 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_198
timestamp 1698431365
transform 1 0 23520 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_202
timestamp 1698431365
transform 1 0 23968 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_206
timestamp 1698431365
transform 1 0 24416 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_218
timestamp 1698431365
transform 1 0 25760 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_278
timestamp 1698431365
transform 1 0 32480 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_282
timestamp 1698431365
transform 1 0 32928 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_319
timestamp 1698431365
transform 1 0 37072 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_395
timestamp 1698431365
transform 1 0 45584 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_411
timestamp 1698431365
transform 1 0 47376 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_419
timestamp 1698431365
transform 1 0 48272 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_422
timestamp 1698431365
transform 1 0 48608 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_486
timestamp 1698431365
transform 1 0 55776 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_492
timestamp 1698431365
transform 1 0 56448 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_556
timestamp 1698431365
transform 1 0 63616 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_562
timestamp 1698431365
transform 1 0 64288 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_626
timestamp 1698431365
transform 1 0 71456 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_632
timestamp 1698431365
transform 1 0 72128 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_8
timestamp 1698431365
transform 1 0 2240 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_12
timestamp 1698431365
transform 1 0 2688 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_28
timestamp 1698431365
transform 1 0 4480 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_32
timestamp 1698431365
transform 1 0 4928 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_53
timestamp 1698431365
transform 1 0 7280 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_102
timestamp 1698431365
transform 1 0 12768 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_104
timestamp 1698431365
transform 1 0 12992 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_115
timestamp 1698431365
transform 1 0 14224 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_119
timestamp 1698431365
transform 1 0 14672 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_170
timestamp 1698431365
transform 1 0 20384 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_174
timestamp 1698431365
transform 1 0 20832 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_233
timestamp 1698431365
transform 1 0 27440 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_237
timestamp 1698431365
transform 1 0 27888 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_241
timestamp 1698431365
transform 1 0 28336 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_253
timestamp 1698431365
transform 1 0 29680 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_257
timestamp 1698431365
transform 1 0 30128 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_261
timestamp 1698431365
transform 1 0 30576 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_265
timestamp 1698431365
transform 1 0 31024 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_277
timestamp 1698431365
transform 1 0 32368 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_279
timestamp 1698431365
transform 1 0 32592 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_294
timestamp 1698431365
transform 1 0 34272 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_304
timestamp 1698431365
transform 1 0 35392 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_312
timestamp 1698431365
transform 1 0 36288 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_314
timestamp 1698431365
transform 1 0 36512 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_338
timestamp 1698431365
transform 1 0 39200 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_342
timestamp 1698431365
transform 1 0 39648 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_346
timestamp 1698431365
transform 1 0 40096 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_350
timestamp 1698431365
transform 1 0 40544 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_357
timestamp 1698431365
transform 1 0 41328 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_359
timestamp 1698431365
transform 1 0 41552 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_378
timestamp 1698431365
transform 1 0 43680 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_382
timestamp 1698431365
transform 1 0 44128 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_384
timestamp 1698431365
transform 1 0 44352 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_387
timestamp 1698431365
transform 1 0 44688 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_451
timestamp 1698431365
transform 1 0 51856 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_457
timestamp 1698431365
transform 1 0 52528 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_521
timestamp 1698431365
transform 1 0 59696 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_527
timestamp 1698431365
transform 1 0 60368 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_591
timestamp 1698431365
transform 1 0 67536 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_597
timestamp 1698431365
transform 1 0 68208 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_629
timestamp 1698431365
transform 1 0 71792 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_645
timestamp 1698431365
transform 1 0 73584 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_653
timestamp 1698431365
transform 1 0 74480 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_657
timestamp 1698431365
transform 1 0 74928 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_661
timestamp 1698431365
transform 1 0 75376 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_667
timestamp 1698431365
transform 1 0 76048 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_671
timestamp 1698431365
transform 1 0 76496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_675
timestamp 1698431365
transform 1 0 76944 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_678
timestamp 1698431365
transform 1 0 77280 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_8
timestamp 1698431365
transform 1 0 2240 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_12
timestamp 1698431365
transform 1 0 2688 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_44
timestamp 1698431365
transform 1 0 6272 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_60
timestamp 1698431365
transform 1 0 8064 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_68
timestamp 1698431365
transform 1 0 8960 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_72
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_80
timestamp 1698431365
transform 1 0 10304 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_84
timestamp 1698431365
transform 1 0 10752 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_96
timestamp 1698431365
transform 1 0 12096 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_98
timestamp 1698431365
transform 1 0 12320 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_130
timestamp 1698431365
transform 1 0 15904 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_138
timestamp 1698431365
transform 1 0 16800 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_146
timestamp 1698431365
transform 1 0 17696 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_191
timestamp 1698431365
transform 1 0 22736 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_199
timestamp 1698431365
transform 1 0 23632 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_201
timestamp 1698431365
transform 1 0 23856 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_212
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_224
timestamp 1698431365
transform 1 0 26432 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_226
timestamp 1698431365
transform 1 0 26656 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_229
timestamp 1698431365
transform 1 0 26992 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_233
timestamp 1698431365
transform 1 0 27440 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_274
timestamp 1698431365
transform 1 0 32032 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_345
timestamp 1698431365
transform 1 0 39984 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_349
timestamp 1698431365
transform 1 0 40432 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_352
timestamp 1698431365
transform 1 0 40768 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_385
timestamp 1698431365
transform 1 0 44464 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_417
timestamp 1698431365
transform 1 0 48048 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_419
timestamp 1698431365
transform 1 0 48272 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_422
timestamp 1698431365
transform 1 0 48608 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_486
timestamp 1698431365
transform 1 0 55776 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_492
timestamp 1698431365
transform 1 0 56448 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_556
timestamp 1698431365
transform 1 0 63616 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_562
timestamp 1698431365
transform 1 0 64288 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_626
timestamp 1698431365
transform 1 0 71456 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_632
timestamp 1698431365
transform 1 0 72128 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_648
timestamp 1698431365
transform 1 0 73920 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_656
timestamp 1698431365
transform 1 0 74816 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_660
timestamp 1698431365
transform 1 0 75264 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_8
timestamp 1698431365
transform 1 0 2240 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_12
timestamp 1698431365
transform 1 0 2688 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_28
timestamp 1698431365
transform 1 0 4480 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_32
timestamp 1698431365
transform 1 0 4928 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698431365
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_37
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_75
timestamp 1698431365
transform 1 0 9744 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_83
timestamp 1698431365
transform 1 0 10640 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_87
timestamp 1698431365
transform 1 0 11088 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_97
timestamp 1698431365
transform 1 0 12208 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698431365
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_113
timestamp 1698431365
transform 1 0 14000 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_121
timestamp 1698431365
transform 1 0 14896 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_123
timestamp 1698431365
transform 1 0 15120 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_155
timestamp 1698431365
transform 1 0 18704 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_159
timestamp 1698431365
transform 1 0 19152 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_161
timestamp 1698431365
transform 1 0 19376 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_170
timestamp 1698431365
transform 1 0 20384 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_174
timestamp 1698431365
transform 1 0 20832 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_177
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_181
timestamp 1698431365
transform 1 0 21616 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_183
timestamp 1698431365
transform 1 0 21840 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_190
timestamp 1698431365
transform 1 0 22624 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_206
timestamp 1698431365
transform 1 0 24416 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_242
timestamp 1698431365
transform 1 0 28448 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_244
timestamp 1698431365
transform 1 0 28672 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_247
timestamp 1698431365
transform 1 0 29008 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_251
timestamp 1698431365
transform 1 0 29456 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_258
timestamp 1698431365
transform 1 0 30240 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_311
timestamp 1698431365
transform 1 0 36176 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_323
timestamp 1698431365
transform 1 0 37520 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_330
timestamp 1698431365
transform 1 0 38304 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_332
timestamp 1698431365
transform 1 0 38528 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_383
timestamp 1698431365
transform 1 0 44240 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_393
timestamp 1698431365
transform 1 0 45360 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_425
timestamp 1698431365
transform 1 0 48944 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_441
timestamp 1698431365
transform 1 0 50736 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_449
timestamp 1698431365
transform 1 0 51632 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_453
timestamp 1698431365
transform 1 0 52080 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_457
timestamp 1698431365
transform 1 0 52528 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_521
timestamp 1698431365
transform 1 0 59696 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_527
timestamp 1698431365
transform 1 0 60368 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_591
timestamp 1698431365
transform 1 0 67536 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_597
timestamp 1698431365
transform 1 0 68208 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_661
timestamp 1698431365
transform 1 0 75376 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_673
timestamp 1698431365
transform 1 0 76720 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_675
timestamp 1698431365
transform 1 0 76944 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_678
timestamp 1698431365
transform 1 0 77280 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698431365
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_103
timestamp 1698431365
transform 1 0 12880 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_135
timestamp 1698431365
transform 1 0 16464 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_139
timestamp 1698431365
transform 1 0 16912 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_150
timestamp 1698431365
transform 1 0 18144 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_172
timestamp 1698431365
transform 1 0 20608 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_176
timestamp 1698431365
transform 1 0 21056 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_209
timestamp 1698431365
transform 1 0 24752 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_220
timestamp 1698431365
transform 1 0 25984 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_242
timestamp 1698431365
transform 1 0 28448 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_246
timestamp 1698431365
transform 1 0 28896 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698431365
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_282
timestamp 1698431365
transform 1 0 32928 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_286
timestamp 1698431365
transform 1 0 33376 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_294
timestamp 1698431365
transform 1 0 34272 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_310
timestamp 1698431365
transform 1 0 36064 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_356
timestamp 1698431365
transform 1 0 41216 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_364
timestamp 1698431365
transform 1 0 42112 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_368
timestamp 1698431365
transform 1 0 42560 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_400
timestamp 1698431365
transform 1 0 46144 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_416
timestamp 1698431365
transform 1 0 47936 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_422
timestamp 1698431365
transform 1 0 48608 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_486
timestamp 1698431365
transform 1 0 55776 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_492
timestamp 1698431365
transform 1 0 56448 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_556
timestamp 1698431365
transform 1 0 63616 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_562
timestamp 1698431365
transform 1 0 64288 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_626
timestamp 1698431365
transform 1 0 71456 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_632
timestamp 1698431365
transform 1 0 72128 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_648
timestamp 1698431365
transform 1 0 73920 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_652
timestamp 1698431365
transform 1 0 74368 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_664
timestamp 1698431365
transform 1 0 75712 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_668
timestamp 1698431365
transform 1 0 76160 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_676
timestamp 1698431365
transform 1 0 77056 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_8
timestamp 1698431365
transform 1 0 2240 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_12
timestamp 1698431365
transform 1 0 2688 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_28
timestamp 1698431365
transform 1 0 4480 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_32
timestamp 1698431365
transform 1 0 4928 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698431365
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698431365
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_107
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_123
timestamp 1698431365
transform 1 0 15120 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_131
timestamp 1698431365
transform 1 0 16016 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_133
timestamp 1698431365
transform 1 0 16240 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_173
timestamp 1698431365
transform 1 0 20720 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_177
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_181
timestamp 1698431365
transform 1 0 21616 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_189
timestamp 1698431365
transform 1 0 22512 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_228
timestamp 1698431365
transform 1 0 26880 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_232
timestamp 1698431365
transform 1 0 27328 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_234
timestamp 1698431365
transform 1 0 27552 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698431365
transform 1 0 28336 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_253
timestamp 1698431365
transform 1 0 29680 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_269
timestamp 1698431365
transform 1 0 31472 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_273
timestamp 1698431365
transform 1 0 31920 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_275
timestamp 1698431365
transform 1 0 32144 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_286
timestamp 1698431365
transform 1 0 33376 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_288
timestamp 1698431365
transform 1 0 33600 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_299
timestamp 1698431365
transform 1 0 34832 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698431365
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_317
timestamp 1698431365
transform 1 0 36848 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_319
timestamp 1698431365
transform 1 0 37072 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_325
timestamp 1698431365
transform 1 0 37744 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_329
timestamp 1698431365
transform 1 0 38192 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_365
timestamp 1698431365
transform 1 0 42224 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_374
timestamp 1698431365
transform 1 0 43232 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_382
timestamp 1698431365
transform 1 0 44128 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_384
timestamp 1698431365
transform 1 0 44352 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_387
timestamp 1698431365
transform 1 0 44688 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_451
timestamp 1698431365
transform 1 0 51856 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_457
timestamp 1698431365
transform 1 0 52528 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_521
timestamp 1698431365
transform 1 0 59696 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_527
timestamp 1698431365
transform 1 0 60368 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_591
timestamp 1698431365
transform 1 0 67536 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_597
timestamp 1698431365
transform 1 0 68208 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_661
timestamp 1698431365
transform 1 0 75376 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_667
timestamp 1698431365
transform 1 0 76048 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_683
timestamp 1698431365
transform 1 0 77840 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_687
timestamp 1698431365
transform 1 0 78288 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_8
timestamp 1698431365
transform 1 0 2240 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_12
timestamp 1698431365
transform 1 0 2688 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_44
timestamp 1698431365
transform 1 0 6272 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_60
timestamp 1698431365
transform 1 0 8064 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_68
timestamp 1698431365
transform 1 0 8960 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698431365
transform 1 0 16576 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_142
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_158
timestamp 1698431365
transform 1 0 19040 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_193
timestamp 1698431365
transform 1 0 22960 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_195
timestamp 1698431365
transform 1 0 23184 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_202
timestamp 1698431365
transform 1 0 23968 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_212
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_216
timestamp 1698431365
transform 1 0 25536 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_218
timestamp 1698431365
transform 1 0 25760 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_234
timestamp 1698431365
transform 1 0 27552 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_269
timestamp 1698431365
transform 1 0 31472 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_277
timestamp 1698431365
transform 1 0 32368 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_279
timestamp 1698431365
transform 1 0 32592 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_290
timestamp 1698431365
transform 1 0 33824 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_333
timestamp 1698431365
transform 1 0 38640 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_349
timestamp 1698431365
transform 1 0 40432 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_352
timestamp 1698431365
transform 1 0 40768 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_395
timestamp 1698431365
transform 1 0 45584 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_403
timestamp 1698431365
transform 1 0 46480 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_409
timestamp 1698431365
transform 1 0 47152 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_417
timestamp 1698431365
transform 1 0 48048 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_422
timestamp 1698431365
transform 1 0 48608 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_426
timestamp 1698431365
transform 1 0 49056 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_430
timestamp 1698431365
transform 1 0 49504 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_438
timestamp 1698431365
transform 1 0 50400 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_472
timestamp 1698431365
transform 1 0 54208 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_488
timestamp 1698431365
transform 1 0 56000 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_492
timestamp 1698431365
transform 1 0 56448 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_556
timestamp 1698431365
transform 1 0 63616 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_562
timestamp 1698431365
transform 1 0 64288 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_626
timestamp 1698431365
transform 1 0 71456 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_632
timestamp 1698431365
transform 1 0 72128 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_664
timestamp 1698431365
transform 1 0 75712 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698431365
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698431365
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_107
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_171
timestamp 1698431365
transform 1 0 20496 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_177
timestamp 1698431365
transform 1 0 21168 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_209
timestamp 1698431365
transform 1 0 24752 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_217
timestamp 1698431365
transform 1 0 25648 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_229
timestamp 1698431365
transform 1 0 26992 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_233
timestamp 1698431365
transform 1 0 27440 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_237
timestamp 1698431365
transform 1 0 27888 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_255
timestamp 1698431365
transform 1 0 29904 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_259
timestamp 1698431365
transform 1 0 30352 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_301
timestamp 1698431365
transform 1 0 35056 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_303
timestamp 1698431365
transform 1 0 35280 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_312
timestamp 1698431365
transform 1 0 36288 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_314
timestamp 1698431365
transform 1 0 36512 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_317
timestamp 1698431365
transform 1 0 36848 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_333
timestamp 1698431365
transform 1 0 38640 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_374
timestamp 1698431365
transform 1 0 43232 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_378
timestamp 1698431365
transform 1 0 43680 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_381
timestamp 1698431365
transform 1 0 44016 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_387
timestamp 1698431365
transform 1 0 44688 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_393
timestamp 1698431365
transform 1 0 45360 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_397
timestamp 1698431365
transform 1 0 45808 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_433
timestamp 1698431365
transform 1 0 49840 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_437
timestamp 1698431365
transform 1 0 50288 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_441
timestamp 1698431365
transform 1 0 50736 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_443
timestamp 1698431365
transform 1 0 50960 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_454
timestamp 1698431365
transform 1 0 52192 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_467
timestamp 1698431365
transform 1 0 53648 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_499
timestamp 1698431365
transform 1 0 57232 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_515
timestamp 1698431365
transform 1 0 59024 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_523
timestamp 1698431365
transform 1 0 59920 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_527
timestamp 1698431365
transform 1 0 60368 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_591
timestamp 1698431365
transform 1 0 67536 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_597
timestamp 1698431365
transform 1 0 68208 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_661
timestamp 1698431365
transform 1 0 75376 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_667
timestamp 1698431365
transform 1 0 76048 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_675
timestamp 1698431365
transform 1 0 76944 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_679
timestamp 1698431365
transform 1 0 77392 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_8
timestamp 1698431365
transform 1 0 2240 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_12
timestamp 1698431365
transform 1 0 2688 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_44
timestamp 1698431365
transform 1 0 6272 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_60
timestamp 1698431365
transform 1 0 8064 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_68
timestamp 1698431365
transform 1 0 8960 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_72
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_136
timestamp 1698431365
transform 1 0 16576 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_142
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_206
timestamp 1698431365
transform 1 0 24416 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_212
timestamp 1698431365
transform 1 0 25088 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_214
timestamp 1698431365
transform 1 0 25312 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_265
timestamp 1698431365
transform 1 0 31024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_269
timestamp 1698431365
transform 1 0 31472 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_277
timestamp 1698431365
transform 1 0 32368 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_290
timestamp 1698431365
transform 1 0 33824 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_294
timestamp 1698431365
transform 1 0 34272 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_298
timestamp 1698431365
transform 1 0 34720 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_300
timestamp 1698431365
transform 1 0 34944 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_330
timestamp 1698431365
transform 1 0 38304 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_338
timestamp 1698431365
transform 1 0 39200 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_352
timestamp 1698431365
transform 1 0 40768 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_356
timestamp 1698431365
transform 1 0 41216 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_358
timestamp 1698431365
transform 1 0 41440 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_486
timestamp 1698431365
transform 1 0 55776 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_492
timestamp 1698431365
transform 1 0 56448 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_556
timestamp 1698431365
transform 1 0 63616 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_562
timestamp 1698431365
transform 1 0 64288 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_626
timestamp 1698431365
transform 1 0 71456 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_632
timestamp 1698431365
transform 1 0 72128 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_664
timestamp 1698431365
transform 1 0 75712 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_680
timestamp 1698431365
transform 1 0 77504 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_8
timestamp 1698431365
transform 1 0 2240 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_12
timestamp 1698431365
transform 1 0 2688 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_28
timestamp 1698431365
transform 1 0 4480 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_32
timestamp 1698431365
transform 1 0 4928 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698431365
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698431365
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_107
timestamp 1698431365
transform 1 0 13328 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_171
timestamp 1698431365
transform 1 0 20496 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_177
timestamp 1698431365
transform 1 0 21168 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_193
timestamp 1698431365
transform 1 0 22960 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_197
timestamp 1698431365
transform 1 0 23408 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_199
timestamp 1698431365
transform 1 0 23632 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_202
timestamp 1698431365
transform 1 0 23968 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_255
timestamp 1698431365
transform 1 0 29904 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_259
timestamp 1698431365
transform 1 0 30352 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_267
timestamp 1698431365
transform 1 0 31248 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_271
timestamp 1698431365
transform 1 0 31696 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_306
timestamp 1698431365
transform 1 0 35616 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_308
timestamp 1698431365
transform 1 0 35840 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_311
timestamp 1698431365
transform 1 0 36176 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_333
timestamp 1698431365
transform 1 0 38640 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_340
timestamp 1698431365
transform 1 0 39424 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_344
timestamp 1698431365
transform 1 0 39872 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_350
timestamp 1698431365
transform 1 0 40544 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_354
timestamp 1698431365
transform 1 0 40992 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_356
timestamp 1698431365
transform 1 0 41216 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_359
timestamp 1698431365
transform 1 0 41552 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_369
timestamp 1698431365
transform 1 0 42672 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_371
timestamp 1698431365
transform 1 0 42896 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_384
timestamp 1698431365
transform 1 0 44352 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_387
timestamp 1698431365
transform 1 0 44688 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_391
timestamp 1698431365
transform 1 0 45136 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_454
timestamp 1698431365
transform 1 0 52192 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_489
timestamp 1698431365
transform 1 0 56112 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_493
timestamp 1698431365
transform 1 0 56560 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_527
timestamp 1698431365
transform 1 0 60368 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_591
timestamp 1698431365
transform 1 0 67536 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_597
timestamp 1698431365
transform 1 0 68208 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_661
timestamp 1698431365
transform 1 0 75376 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_667
timestamp 1698431365
transform 1 0 76048 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_675
timestamp 1698431365
transform 1 0 76944 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_679
timestamp 1698431365
transform 1 0 77392 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698431365
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_72
timestamp 1698431365
transform 1 0 9408 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_136
timestamp 1698431365
transform 1 0 16576 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_142
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_150
timestamp 1698431365
transform 1 0 18144 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_212
timestamp 1698431365
transform 1 0 25088 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_220
timestamp 1698431365
transform 1 0 25984 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_232
timestamp 1698431365
transform 1 0 27328 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_236
timestamp 1698431365
transform 1 0 27776 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_238
timestamp 1698431365
transform 1 0 28000 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_276
timestamp 1698431365
transform 1 0 32256 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_282
timestamp 1698431365
transform 1 0 32928 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_300
timestamp 1698431365
transform 1 0 34944 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_304
timestamp 1698431365
transform 1 0 35392 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_314
timestamp 1698431365
transform 1 0 36512 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_318
timestamp 1698431365
transform 1 0 36960 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_329
timestamp 1698431365
transform 1 0 38192 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_339
timestamp 1698431365
transform 1 0 39312 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_348
timestamp 1698431365
transform 1 0 40320 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_352
timestamp 1698431365
transform 1 0 40768 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_361
timestamp 1698431365
transform 1 0 41776 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_365
timestamp 1698431365
transform 1 0 42224 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_369
timestamp 1698431365
transform 1 0 42672 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_422
timestamp 1698431365
transform 1 0 48608 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_487
timestamp 1698431365
transform 1 0 55888 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_489
timestamp 1698431365
transform 1 0 56112 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_492
timestamp 1698431365
transform 1 0 56448 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_496
timestamp 1698431365
transform 1 0 56896 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_500
timestamp 1698431365
transform 1 0 57344 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_532
timestamp 1698431365
transform 1 0 60928 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_548
timestamp 1698431365
transform 1 0 62720 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_556
timestamp 1698431365
transform 1 0 63616 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_562
timestamp 1698431365
transform 1 0 64288 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_626
timestamp 1698431365
transform 1 0 71456 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_632
timestamp 1698431365
transform 1 0 72128 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_664
timestamp 1698431365
transform 1 0 75712 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_672
timestamp 1698431365
transform 1 0 76608 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_678
timestamp 1698431365
transform 1 0 77280 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_8
timestamp 1698431365
transform 1 0 2240 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_12
timestamp 1698431365
transform 1 0 2688 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_28
timestamp 1698431365
transform 1 0 4480 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_32
timestamp 1698431365
transform 1 0 4928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698431365
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698431365
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_107
timestamp 1698431365
transform 1 0 13328 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_139
timestamp 1698431365
transform 1 0 16912 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_143
timestamp 1698431365
transform 1 0 17360 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_145
timestamp 1698431365
transform 1 0 17584 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_148
timestamp 1698431365
transform 1 0 17920 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_152
timestamp 1698431365
transform 1 0 18368 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_154
timestamp 1698431365
transform 1 0 18592 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_168
timestamp 1698431365
transform 1 0 20160 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_172
timestamp 1698431365
transform 1 0 20608 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_174
timestamp 1698431365
transform 1 0 20832 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_233
timestamp 1698431365
transform 1 0 27440 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_235
timestamp 1698431365
transform 1 0 27664 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_238
timestamp 1698431365
transform 1 0 28000 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_247
timestamp 1698431365
transform 1 0 29008 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_299
timestamp 1698431365
transform 1 0 34832 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_301
timestamp 1698431365
transform 1 0 35056 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_310
timestamp 1698431365
transform 1 0 36064 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_314
timestamp 1698431365
transform 1 0 36512 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_325
timestamp 1698431365
transform 1 0 37744 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_335
timestamp 1698431365
transform 1 0 38864 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_419
timestamp 1698431365
transform 1 0 48272 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_457
timestamp 1698431365
transform 1 0 52528 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_459
timestamp 1698431365
transform 1 0 52752 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_524
timestamp 1698431365
transform 1 0 60032 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_527
timestamp 1698431365
transform 1 0 60368 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_591
timestamp 1698431365
transform 1 0 67536 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_597
timestamp 1698431365
transform 1 0 68208 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_661
timestamp 1698431365
transform 1 0 75376 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_667
timestamp 1698431365
transform 1 0 76048 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_671
timestamp 1698431365
transform 1 0 76496 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_673
timestamp 1698431365
transform 1 0 76720 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_8
timestamp 1698431365
transform 1 0 2240 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_12
timestamp 1698431365
transform 1 0 2688 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_44
timestamp 1698431365
transform 1 0 6272 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_60
timestamp 1698431365
transform 1 0 8064 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_68
timestamp 1698431365
transform 1 0 8960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_72
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_136
timestamp 1698431365
transform 1 0 16576 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_142
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_144
timestamp 1698431365
transform 1 0 17472 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_200
timestamp 1698431365
transform 1 0 23744 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_212
timestamp 1698431365
transform 1 0 25088 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_245
timestamp 1698431365
transform 1 0 28784 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_247
timestamp 1698431365
transform 1 0 29008 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_277
timestamp 1698431365
transform 1 0 32368 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_279
timestamp 1698431365
transform 1 0 32592 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_282
timestamp 1698431365
transform 1 0 32928 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_333
timestamp 1698431365
transform 1 0 38640 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_347
timestamp 1698431365
transform 1 0 40208 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_349
timestamp 1698431365
transform 1 0 40432 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_352
timestamp 1698431365
transform 1 0 40768 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_354
timestamp 1698431365
transform 1 0 40992 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_418
timestamp 1698431365
transform 1 0 48160 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_454
timestamp 1698431365
transform 1 0 52192 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_492
timestamp 1698431365
transform 1 0 56448 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_496
timestamp 1698431365
transform 1 0 56896 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_500
timestamp 1698431365
transform 1 0 57344 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_532
timestamp 1698431365
transform 1 0 60928 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_548
timestamp 1698431365
transform 1 0 62720 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_556
timestamp 1698431365
transform 1 0 63616 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_562
timestamp 1698431365
transform 1 0 64288 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_594
timestamp 1698431365
transform 1 0 67872 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_610
timestamp 1698431365
transform 1 0 69664 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_626
timestamp 1698431365
transform 1 0 71456 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_632
timestamp 1698431365
transform 1 0 72128 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_664
timestamp 1698431365
transform 1 0 75712 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_674
timestamp 1698431365
transform 1 0 76832 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_684
timestamp 1698431365
transform 1 0 77952 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_8
timestamp 1698431365
transform 1 0 2240 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_12
timestamp 1698431365
transform 1 0 2688 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_28
timestamp 1698431365
transform 1 0 4480 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_32
timestamp 1698431365
transform 1 0 4928 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698431365
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698431365
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_107
timestamp 1698431365
transform 1 0 13328 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_139
timestamp 1698431365
transform 1 0 16912 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_155
timestamp 1698431365
transform 1 0 18704 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_163
timestamp 1698431365
transform 1 0 19600 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_171
timestamp 1698431365
transform 1 0 20496 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_177
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_201
timestamp 1698431365
transform 1 0 23856 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_214
timestamp 1698431365
transform 1 0 25312 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_226
timestamp 1698431365
transform 1 0 26656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_236
timestamp 1698431365
transform 1 0 27776 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_238
timestamp 1698431365
transform 1 0 28000 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_247
timestamp 1698431365
transform 1 0 29008 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_265
timestamp 1698431365
transform 1 0 31024 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_269
timestamp 1698431365
transform 1 0 31472 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_271
timestamp 1698431365
transform 1 0 31696 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_274
timestamp 1698431365
transform 1 0 32032 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_278
timestamp 1698431365
transform 1 0 32480 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_288
timestamp 1698431365
transform 1 0 33600 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_293
timestamp 1698431365
transform 1 0 34160 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_295
timestamp 1698431365
transform 1 0 34384 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_310
timestamp 1698431365
transform 1 0 36064 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_317
timestamp 1698431365
transform 1 0 36848 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_324
timestamp 1698431365
transform 1 0 37632 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_342
timestamp 1698431365
transform 1 0 39648 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_419
timestamp 1698431365
transform 1 0 48272 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_470
timestamp 1698431365
transform 1 0 53984 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_504
timestamp 1698431365
transform 1 0 57792 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_520
timestamp 1698431365
transform 1 0 59584 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_524
timestamp 1698431365
transform 1 0 60032 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_527
timestamp 1698431365
transform 1 0 60368 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_591
timestamp 1698431365
transform 1 0 67536 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_597
timestamp 1698431365
transform 1 0 68208 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_629
timestamp 1698431365
transform 1 0 71792 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_645
timestamp 1698431365
transform 1 0 73584 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_653
timestamp 1698431365
transform 1 0 74480 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_659
timestamp 1698431365
transform 1 0 75152 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_663
timestamp 1698431365
transform 1 0 75600 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_667
timestamp 1698431365
transform 1 0 76048 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_669
timestamp 1698431365
transform 1 0 76272 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698431365
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_72
timestamp 1698431365
transform 1 0 9408 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_136
timestamp 1698431365
transform 1 0 16576 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_142
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_150
timestamp 1698431365
transform 1 0 18144 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_166
timestamp 1698431365
transform 1 0 19936 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_170
timestamp 1698431365
transform 1 0 20384 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_209
timestamp 1698431365
transform 1 0 24752 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_218
timestamp 1698431365
transform 1 0 25760 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_282
timestamp 1698431365
transform 1 0 32928 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_296
timestamp 1698431365
transform 1 0 34496 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_298
timestamp 1698431365
transform 1 0 34720 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_347
timestamp 1698431365
transform 1 0 40208 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_349
timestamp 1698431365
transform 1 0 40432 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_435
timestamp 1698431365
transform 1 0 50064 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_486
timestamp 1698431365
transform 1 0 55776 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_492
timestamp 1698431365
transform 1 0 56448 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_496
timestamp 1698431365
transform 1 0 56896 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_500
timestamp 1698431365
transform 1 0 57344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_504
timestamp 1698431365
transform 1 0 57792 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_536
timestamp 1698431365
transform 1 0 61376 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_552
timestamp 1698431365
transform 1 0 63168 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_562
timestamp 1698431365
transform 1 0 64288 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_626
timestamp 1698431365
transform 1 0 71456 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_632
timestamp 1698431365
transform 1 0 72128 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_636
timestamp 1698431365
transform 1 0 72576 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_640
timestamp 1698431365
transform 1 0 73024 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_644
timestamp 1698431365
transform 1 0 73472 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_646
timestamp 1698431365
transform 1 0 73696 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_649
timestamp 1698431365
transform 1 0 74032 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_653
timestamp 1698431365
transform 1 0 74480 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_684
timestamp 1698431365
transform 1 0 77952 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_8
timestamp 1698431365
transform 1 0 2240 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_12
timestamp 1698431365
transform 1 0 2688 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_28
timestamp 1698431365
transform 1 0 4480 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_32
timestamp 1698431365
transform 1 0 4928 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698431365
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698431365
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_107
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_139
timestamp 1698431365
transform 1 0 16912 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_155
timestamp 1698431365
transform 1 0 18704 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_159
timestamp 1698431365
transform 1 0 19152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_168
timestamp 1698431365
transform 1 0 20160 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_172
timestamp 1698431365
transform 1 0 20608 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_174
timestamp 1698431365
transform 1 0 20832 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_177
timestamp 1698431365
transform 1 0 21168 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_195
timestamp 1698431365
transform 1 0 23184 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_201
timestamp 1698431365
transform 1 0 23856 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_211
timestamp 1698431365
transform 1 0 24976 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_222
timestamp 1698431365
transform 1 0 26208 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_230
timestamp 1698431365
transform 1 0 27104 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_238
timestamp 1698431365
transform 1 0 28000 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_242
timestamp 1698431365
transform 1 0 28448 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_244
timestamp 1698431365
transform 1 0 28672 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_247
timestamp 1698431365
transform 1 0 29008 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_257
timestamp 1698431365
transform 1 0 30128 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_261
timestamp 1698431365
transform 1 0 30576 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_279
timestamp 1698431365
transform 1 0 32592 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_289
timestamp 1698431365
transform 1 0 33712 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_317
timestamp 1698431365
transform 1 0 36848 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_349
timestamp 1698431365
transform 1 0 40432 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_387
timestamp 1698431365
transform 1 0 44688 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_449
timestamp 1698431365
transform 1 0 51632 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_453
timestamp 1698431365
transform 1 0 52080 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_457
timestamp 1698431365
transform 1 0 52528 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_461
timestamp 1698431365
transform 1 0 52976 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_463
timestamp 1698431365
transform 1 0 53200 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_490
timestamp 1698431365
transform 1 0 56224 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_494
timestamp 1698431365
transform 1 0 56672 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_498
timestamp 1698431365
transform 1 0 57120 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_514
timestamp 1698431365
transform 1 0 58912 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_522
timestamp 1698431365
transform 1 0 59808 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_524
timestamp 1698431365
transform 1 0 60032 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_527
timestamp 1698431365
transform 1 0 60368 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_591
timestamp 1698431365
transform 1 0 67536 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_597
timestamp 1698431365
transform 1 0 68208 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_613
timestamp 1698431365
transform 1 0 70000 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_621
timestamp 1698431365
transform 1 0 70896 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_655
timestamp 1698431365
transform 1 0 74704 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_667
timestamp 1698431365
transform 1 0 76048 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_669
timestamp 1698431365
transform 1 0 76272 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_8
timestamp 1698431365
transform 1 0 2240 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_12
timestamp 1698431365
transform 1 0 2688 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_44
timestamp 1698431365
transform 1 0 6272 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_60
timestamp 1698431365
transform 1 0 8064 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_68
timestamp 1698431365
transform 1 0 8960 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_72
timestamp 1698431365
transform 1 0 9408 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_136
timestamp 1698431365
transform 1 0 16576 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_150
timestamp 1698431365
transform 1 0 18144 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_154
timestamp 1698431365
transform 1 0 18592 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_184
timestamp 1698431365
transform 1 0 21952 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_206
timestamp 1698431365
transform 1 0 24416 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_217
timestamp 1698431365
transform 1 0 25648 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_227
timestamp 1698431365
transform 1 0 26768 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_243
timestamp 1698431365
transform 1 0 28560 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_282
timestamp 1698431365
transform 1 0 32928 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_314
timestamp 1698431365
transform 1 0 36512 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_352
timestamp 1698431365
transform 1 0 40768 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_443
timestamp 1698431365
transform 1 0 50960 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_466
timestamp 1698431365
transform 1 0 53536 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_470
timestamp 1698431365
transform 1 0 53984 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_485
timestamp 1698431365
transform 1 0 55664 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_489
timestamp 1698431365
transform 1 0 56112 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_492
timestamp 1698431365
transform 1 0 56448 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_556
timestamp 1698431365
transform 1 0 63616 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_562
timestamp 1698431365
transform 1 0 64288 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_626
timestamp 1698431365
transform 1 0 71456 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_662
timestamp 1698431365
transform 1 0 75488 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_669
timestamp 1698431365
transform 1 0 76272 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_677
timestamp 1698431365
transform 1 0 77168 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_685
timestamp 1698431365
transform 1 0 78064 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_687
timestamp 1698431365
transform 1 0 78288 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698431365
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698431365
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_107
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_123
timestamp 1698431365
transform 1 0 15120 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_212
timestamp 1698431365
transform 1 0 25088 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_243
timestamp 1698431365
transform 1 0 28560 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_253
timestamp 1698431365
transform 1 0 29680 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_285
timestamp 1698431365
transform 1 0 33264 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_289
timestamp 1698431365
transform 1 0 33712 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_292
timestamp 1698431365
transform 1 0 34048 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_296
timestamp 1698431365
transform 1 0 34496 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_359
timestamp 1698431365
transform 1 0 41552 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_361
timestamp 1698431365
transform 1 0 41776 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_382
timestamp 1698431365
transform 1 0 44128 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_384
timestamp 1698431365
transform 1 0 44352 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_387
timestamp 1698431365
transform 1 0 44688 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_389
timestamp 1698431365
transform 1 0 44912 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_437
timestamp 1698431365
transform 1 0 50288 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_439
timestamp 1698431365
transform 1 0 50512 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_448
timestamp 1698431365
transform 1 0 51520 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_452
timestamp 1698431365
transform 1 0 51968 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_454
timestamp 1698431365
transform 1 0 52192 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_457
timestamp 1698431365
transform 1 0 52528 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_461
timestamp 1698431365
transform 1 0 52976 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_527
timestamp 1698431365
transform 1 0 60368 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_591
timestamp 1698431365
transform 1 0 67536 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_597
timestamp 1698431365
transform 1 0 68208 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_646
timestamp 1698431365
transform 1 0 73696 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_648
timestamp 1698431365
transform 1 0 73920 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_664
timestamp 1698431365
transform 1 0 75712 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_685
timestamp 1698431365
transform 1 0 78064 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_687
timestamp 1698431365
transform 1 0 78288 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_8
timestamp 1698431365
transform 1 0 2240 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_12
timestamp 1698431365
transform 1 0 2688 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_44
timestamp 1698431365
transform 1 0 6272 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_60
timestamp 1698431365
transform 1 0 8064 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_68
timestamp 1698431365
transform 1 0 8960 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_72
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_136
timestamp 1698431365
transform 1 0 16576 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_150
timestamp 1698431365
transform 1 0 18144 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_154
timestamp 1698431365
transform 1 0 18592 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_158
timestamp 1698431365
transform 1 0 19040 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_170
timestamp 1698431365
transform 1 0 20384 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_174
timestamp 1698431365
transform 1 0 20832 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_176
timestamp 1698431365
transform 1 0 21056 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_185
timestamp 1698431365
transform 1 0 22064 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_193
timestamp 1698431365
transform 1 0 22960 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_197
timestamp 1698431365
transform 1 0 23408 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_200
timestamp 1698431365
transform 1 0 23744 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698431365
transform 1 0 24752 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_223
timestamp 1698431365
transform 1 0 26320 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_231
timestamp 1698431365
transform 1 0 27216 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_273
timestamp 1698431365
transform 1 0 31920 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_277
timestamp 1698431365
transform 1 0 32368 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_279
timestamp 1698431365
transform 1 0 32592 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_282
timestamp 1698431365
transform 1 0 32928 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_393
timestamp 1698431365
transform 1 0 45360 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_395
timestamp 1698431365
transform 1 0 45584 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_419
timestamp 1698431365
transform 1 0 48272 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_422
timestamp 1698431365
transform 1 0 48608 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_426
timestamp 1698431365
transform 1 0 49056 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_430
timestamp 1698431365
transform 1 0 49504 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_434
timestamp 1698431365
transform 1 0 49952 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_436
timestamp 1698431365
transform 1 0 50176 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_439
timestamp 1698431365
transform 1 0 50512 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_443
timestamp 1698431365
transform 1 0 50960 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_475
timestamp 1698431365
transform 1 0 54544 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_483
timestamp 1698431365
transform 1 0 55440 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_487
timestamp 1698431365
transform 1 0 55888 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_489
timestamp 1698431365
transform 1 0 56112 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_492
timestamp 1698431365
transform 1 0 56448 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_556
timestamp 1698431365
transform 1 0 63616 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_562
timestamp 1698431365
transform 1 0 64288 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_626
timestamp 1698431365
transform 1 0 71456 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_668
timestamp 1698431365
transform 1 0 76160 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_678
timestamp 1698431365
transform 1 0 77280 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_685
timestamp 1698431365
transform 1 0 78064 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_687
timestamp 1698431365
transform 1 0 78288 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_8
timestamp 1698431365
transform 1 0 2240 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_12
timestamp 1698431365
transform 1 0 2688 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_28
timestamp 1698431365
transform 1 0 4480 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_32
timestamp 1698431365
transform 1 0 4928 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698431365
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698431365
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698431365
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_107
timestamp 1698431365
transform 1 0 13328 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_123
timestamp 1698431365
transform 1 0 15120 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_131
timestamp 1698431365
transform 1 0 16016 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_135
timestamp 1698431365
transform 1 0 16464 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_171
timestamp 1698431365
transform 1 0 20496 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_185
timestamp 1698431365
transform 1 0 22064 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_189
timestamp 1698431365
transform 1 0 22512 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_193
timestamp 1698431365
transform 1 0 22960 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_230
timestamp 1698431365
transform 1 0 27104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_240
timestamp 1698431365
transform 1 0 28224 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_244
timestamp 1698431365
transform 1 0 28672 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_247
timestamp 1698431365
transform 1 0 29008 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_279
timestamp 1698431365
transform 1 0 32592 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_287
timestamp 1698431365
transform 1 0 33488 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_293
timestamp 1698431365
transform 1 0 34160 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_297
timestamp 1698431365
transform 1 0 34608 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_301
timestamp 1698431365
transform 1 0 35056 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_317
timestamp 1698431365
transform 1 0 36848 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_368
timestamp 1698431365
transform 1 0 42560 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_372
timestamp 1698431365
transform 1 0 43008 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_376
timestamp 1698431365
transform 1 0 43456 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_380
timestamp 1698431365
transform 1 0 43904 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_384
timestamp 1698431365
transform 1 0 44352 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_387
timestamp 1698431365
transform 1 0 44688 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_391
timestamp 1698431365
transform 1 0 45136 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_395
timestamp 1698431365
transform 1 0 45584 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_415
timestamp 1698431365
transform 1 0 47824 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_419
timestamp 1698431365
transform 1 0 48272 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_423
timestamp 1698431365
transform 1 0 48720 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_427
timestamp 1698431365
transform 1 0 49168 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_431
timestamp 1698431365
transform 1 0 49616 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_447
timestamp 1698431365
transform 1 0 51408 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_457
timestamp 1698431365
transform 1 0 52528 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_521
timestamp 1698431365
transform 1 0 59696 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_527
timestamp 1698431365
transform 1 0 60368 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_543
timestamp 1698431365
transform 1 0 62160 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_547
timestamp 1698431365
transform 1 0 62608 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_558
timestamp 1698431365
transform 1 0 63840 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_562
timestamp 1698431365
transform 1 0 64288 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_594
timestamp 1698431365
transform 1 0 67872 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_597
timestamp 1698431365
transform 1 0 68208 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_629
timestamp 1698431365
transform 1 0 71792 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_631
timestamp 1698431365
transform 1 0 72016 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_634
timestamp 1698431365
transform 1 0 72352 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_638
timestamp 1698431365
transform 1 0 72800 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_657
timestamp 1698431365
transform 1 0 74928 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_685
timestamp 1698431365
transform 1 0 78064 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_687
timestamp 1698431365
transform 1 0 78288 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698431365
transform 1 0 1568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698431365
transform 1 0 8736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_72
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_136
timestamp 1698431365
transform 1 0 16576 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_147
timestamp 1698431365
transform 1 0 17808 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_151
timestamp 1698431365
transform 1 0 18256 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_159
timestamp 1698431365
transform 1 0 19152 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_202
timestamp 1698431365
transform 1 0 23968 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_220
timestamp 1698431365
transform 1 0 25984 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_261
timestamp 1698431365
transform 1 0 30576 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_277
timestamp 1698431365
transform 1 0 32368 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_279
timestamp 1698431365
transform 1 0 32592 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_282
timestamp 1698431365
transform 1 0 32928 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_298
timestamp 1698431365
transform 1 0 34720 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_358
timestamp 1698431365
transform 1 0 41440 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_368
timestamp 1698431365
transform 1 0 42560 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_370
timestamp 1698431365
transform 1 0 42784 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_384
timestamp 1698431365
transform 1 0 44352 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_388
timestamp 1698431365
transform 1 0 44800 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_402
timestamp 1698431365
transform 1 0 46368 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_406
timestamp 1698431365
transform 1 0 46816 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_410
timestamp 1698431365
transform 1 0 47264 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_418
timestamp 1698431365
transform 1 0 48160 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_422
timestamp 1698431365
transform 1 0 48608 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_486
timestamp 1698431365
transform 1 0 55776 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_492
timestamp 1698431365
transform 1 0 56448 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_524
timestamp 1698431365
transform 1 0 60032 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_540
timestamp 1698431365
transform 1 0 61824 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_548
timestamp 1698431365
transform 1 0 62720 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_557
timestamp 1698431365
transform 1 0 63728 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_559
timestamp 1698431365
transform 1 0 63952 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_562
timestamp 1698431365
transform 1 0 64288 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_566
timestamp 1698431365
transform 1 0 64736 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_598
timestamp 1698431365
transform 1 0 68320 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_614
timestamp 1698431365
transform 1 0 70112 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_622
timestamp 1698431365
transform 1 0 71008 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_626
timestamp 1698431365
transform 1 0 71456 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_668
timestamp 1698431365
transform 1 0 76160 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_672
timestamp 1698431365
transform 1 0 76608 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_685
timestamp 1698431365
transform 1 0 78064 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_687
timestamp 1698431365
transform 1 0 78288 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_8
timestamp 1698431365
transform 1 0 2240 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_12
timestamp 1698431365
transform 1 0 2688 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_28
timestamp 1698431365
transform 1 0 4480 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_32
timestamp 1698431365
transform 1 0 4928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698431365
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698431365
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698431365
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_107
timestamp 1698431365
transform 1 0 13328 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_171
timestamp 1698431365
transform 1 0 20496 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_177
timestamp 1698431365
transform 1 0 21168 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_241
timestamp 1698431365
transform 1 0 28336 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_247
timestamp 1698431365
transform 1 0 29008 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_279
timestamp 1698431365
transform 1 0 32592 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_295
timestamp 1698431365
transform 1 0 34384 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_312
timestamp 1698431365
transform 1 0 36288 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_314
timestamp 1698431365
transform 1 0 36512 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_317
timestamp 1698431365
transform 1 0 36848 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_340
timestamp 1698431365
transform 1 0 39424 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_344
timestamp 1698431365
transform 1 0 39872 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_410
timestamp 1698431365
transform 1 0 47264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_414
timestamp 1698431365
transform 1 0 47712 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_446
timestamp 1698431365
transform 1 0 51296 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_454
timestamp 1698431365
transform 1 0 52192 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_457
timestamp 1698431365
transform 1 0 52528 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_521
timestamp 1698431365
transform 1 0 59696 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_527
timestamp 1698431365
transform 1 0 60368 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_591
timestamp 1698431365
transform 1 0 67536 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_597
timestamp 1698431365
transform 1 0 68208 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_613
timestamp 1698431365
transform 1 0 70000 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_615
timestamp 1698431365
transform 1 0 70224 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_618
timestamp 1698431365
transform 1 0 70560 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_652
timestamp 1698431365
transform 1 0 74368 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_656
timestamp 1698431365
transform 1 0 74816 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_658
timestamp 1698431365
transform 1 0 75040 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_673
timestamp 1698431365
transform 1 0 76720 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_681
timestamp 1698431365
transform 1 0 77616 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_8
timestamp 1698431365
transform 1 0 2240 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_12
timestamp 1698431365
transform 1 0 2688 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_44
timestamp 1698431365
transform 1 0 6272 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_60
timestamp 1698431365
transform 1 0 8064 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_68
timestamp 1698431365
transform 1 0 8960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_72
timestamp 1698431365
transform 1 0 9408 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_136
timestamp 1698431365
transform 1 0 16576 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_142
timestamp 1698431365
transform 1 0 17248 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_206
timestamp 1698431365
transform 1 0 24416 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_212
timestamp 1698431365
transform 1 0 25088 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_276
timestamp 1698431365
transform 1 0 32256 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_282
timestamp 1698431365
transform 1 0 32928 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_286
timestamp 1698431365
transform 1 0 33376 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_349
timestamp 1698431365
transform 1 0 40432 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_373
timestamp 1698431365
transform 1 0 43120 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_392
timestamp 1698431365
transform 1 0 45248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_418
timestamp 1698431365
transform 1 0 48160 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_432
timestamp 1698431365
transform 1 0 49728 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_436
timestamp 1698431365
transform 1 0 50176 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_440
timestamp 1698431365
transform 1 0 50624 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_472
timestamp 1698431365
transform 1 0 54208 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_488
timestamp 1698431365
transform 1 0 56000 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_492
timestamp 1698431365
transform 1 0 56448 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_556
timestamp 1698431365
transform 1 0 63616 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_562
timestamp 1698431365
transform 1 0 64288 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_594
timestamp 1698431365
transform 1 0 67872 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_610
timestamp 1698431365
transform 1 0 69664 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_618
timestamp 1698431365
transform 1 0 70560 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_622
timestamp 1698431365
transform 1 0 71008 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_626
timestamp 1698431365
transform 1 0 71456 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_632
timestamp 1698431365
transform 1 0 72128 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_634
timestamp 1698431365
transform 1 0 72352 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_637
timestamp 1698431365
transform 1 0 72688 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_664
timestamp 1698431365
transform 1 0 75712 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_666
timestamp 1698431365
transform 1 0 75936 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_675
timestamp 1698431365
transform 1 0 76944 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_685
timestamp 1698431365
transform 1 0 78064 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_687
timestamp 1698431365
transform 1 0 78288 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_8
timestamp 1698431365
transform 1 0 2240 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_12
timestamp 1698431365
transform 1 0 2688 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_28
timestamp 1698431365
transform 1 0 4480 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_32
timestamp 1698431365
transform 1 0 4928 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698431365
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698431365
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698431365
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_107
timestamp 1698431365
transform 1 0 13328 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_171
timestamp 1698431365
transform 1 0 20496 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_177
timestamp 1698431365
transform 1 0 21168 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_241
timestamp 1698431365
transform 1 0 28336 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_247
timestamp 1698431365
transform 1 0 29008 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_279
timestamp 1698431365
transform 1 0 32592 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_287
timestamp 1698431365
transform 1 0 33488 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_338
timestamp 1698431365
transform 1 0 39200 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_366
timestamp 1698431365
transform 1 0 42336 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_370
timestamp 1698431365
transform 1 0 42784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_374
timestamp 1698431365
transform 1 0 43232 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_382
timestamp 1698431365
transform 1 0 44128 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_384
timestamp 1698431365
transform 1 0 44352 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_391
timestamp 1698431365
transform 1 0 45136 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_395
timestamp 1698431365
transform 1 0 45584 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_399
timestamp 1698431365
transform 1 0 46032 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_401
timestamp 1698431365
transform 1 0 46256 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_418
timestamp 1698431365
transform 1 0 48160 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_422
timestamp 1698431365
transform 1 0 48608 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_434
timestamp 1698431365
transform 1 0 49952 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_438
timestamp 1698431365
transform 1 0 50400 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_442
timestamp 1698431365
transform 1 0 50848 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_450
timestamp 1698431365
transform 1 0 51744 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_454
timestamp 1698431365
transform 1 0 52192 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_457
timestamp 1698431365
transform 1 0 52528 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_521
timestamp 1698431365
transform 1 0 59696 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_527
timestamp 1698431365
transform 1 0 60368 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_591
timestamp 1698431365
transform 1 0 67536 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_597
timestamp 1698431365
transform 1 0 68208 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_613
timestamp 1698431365
transform 1 0 70000 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_615
timestamp 1698431365
transform 1 0 70224 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_624
timestamp 1698431365
transform 1 0 71232 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_630
timestamp 1698431365
transform 1 0 71904 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_634
timestamp 1698431365
transform 1 0 72352 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_646
timestamp 1698431365
transform 1 0 73696 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_650
timestamp 1698431365
transform 1 0 74144 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_652
timestamp 1698431365
transform 1 0 74368 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_685
timestamp 1698431365
transform 1 0 78064 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_687
timestamp 1698431365
transform 1 0 78288 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698431365
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1698431365
transform 1 0 9408 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698431365
transform 1 0 16576 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_142
timestamp 1698431365
transform 1 0 17248 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_206
timestamp 1698431365
transform 1 0 24416 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698431365
transform 1 0 25088 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698431365
transform 1 0 32256 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_282
timestamp 1698431365
transform 1 0 32928 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_298
timestamp 1698431365
transform 1 0 34720 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_300
timestamp 1698431365
transform 1 0 34944 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_316
timestamp 1698431365
transform 1 0 36736 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_320
timestamp 1698431365
transform 1 0 37184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_337
timestamp 1698431365
transform 1 0 39088 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_341
timestamp 1698431365
transform 1 0 39536 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_345
timestamp 1698431365
transform 1 0 39984 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_347
timestamp 1698431365
transform 1 0 40208 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_365
timestamp 1698431365
transform 1 0 42224 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_369
timestamp 1698431365
transform 1 0 42672 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_385
timestamp 1698431365
transform 1 0 44464 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_393
timestamp 1698431365
transform 1 0 45360 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_409
timestamp 1698431365
transform 1 0 47152 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_417
timestamp 1698431365
transform 1 0 48048 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_419
timestamp 1698431365
transform 1 0 48272 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_422
timestamp 1698431365
transform 1 0 48608 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_486
timestamp 1698431365
transform 1 0 55776 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_492
timestamp 1698431365
transform 1 0 56448 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_556
timestamp 1698431365
transform 1 0 63616 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_562
timestamp 1698431365
transform 1 0 64288 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_594
timestamp 1698431365
transform 1 0 67872 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_610
timestamp 1698431365
transform 1 0 69664 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_612
timestamp 1698431365
transform 1 0 69888 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_623
timestamp 1698431365
transform 1 0 71120 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_625
timestamp 1698431365
transform 1 0 71344 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_628
timestamp 1698431365
transform 1 0 71680 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_632
timestamp 1698431365
transform 1 0 72128 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_634
timestamp 1698431365
transform 1 0 72352 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_667
timestamp 1698431365
transform 1 0 76048 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_685
timestamp 1698431365
transform 1 0 78064 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_687
timestamp 1698431365
transform 1 0 78288 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_8
timestamp 1698431365
transform 1 0 2240 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_12
timestamp 1698431365
transform 1 0 2688 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_28
timestamp 1698431365
transform 1 0 4480 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_32
timestamp 1698431365
transform 1 0 4928 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698431365
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698431365
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698431365
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698431365
transform 1 0 13328 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698431365
transform 1 0 20496 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698431365
transform 1 0 21168 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698431365
transform 1 0 28336 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698431365
transform 1 0 29008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698431365
transform 1 0 36176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_317
timestamp 1698431365
transform 1 0 36848 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_321
timestamp 1698431365
transform 1 0 37296 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_387
timestamp 1698431365
transform 1 0 44688 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_451
timestamp 1698431365
transform 1 0 51856 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_457
timestamp 1698431365
transform 1 0 52528 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_521
timestamp 1698431365
transform 1 0 59696 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_527
timestamp 1698431365
transform 1 0 60368 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_591
timestamp 1698431365
transform 1 0 67536 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_597
timestamp 1698431365
transform 1 0 68208 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_605
timestamp 1698431365
transform 1 0 69104 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_609
timestamp 1698431365
transform 1 0 69552 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_611
timestamp 1698431365
transform 1 0 69776 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_627
timestamp 1698431365
transform 1 0 71568 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_640
timestamp 1698431365
transform 1 0 73024 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_642
timestamp 1698431365
transform 1 0 73248 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_663
timestamp 1698431365
transform 1 0 75600 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_683
timestamp 1698431365
transform 1 0 77840 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_687
timestamp 1698431365
transform 1 0 78288 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_8
timestamp 1698431365
transform 1 0 2240 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_12
timestamp 1698431365
transform 1 0 2688 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_44
timestamp 1698431365
transform 1 0 6272 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_60
timestamp 1698431365
transform 1 0 8064 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_68
timestamp 1698431365
transform 1 0 8960 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698431365
transform 1 0 9408 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698431365
transform 1 0 16576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698431365
transform 1 0 17248 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698431365
transform 1 0 24416 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698431365
transform 1 0 25088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698431365
transform 1 0 32256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698431365
transform 1 0 32928 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_346
timestamp 1698431365
transform 1 0 40096 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_352
timestamp 1698431365
transform 1 0 40768 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_384
timestamp 1698431365
transform 1 0 44352 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_391
timestamp 1698431365
transform 1 0 45136 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_407
timestamp 1698431365
transform 1 0 46928 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_415
timestamp 1698431365
transform 1 0 47824 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_419
timestamp 1698431365
transform 1 0 48272 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_422
timestamp 1698431365
transform 1 0 48608 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_486
timestamp 1698431365
transform 1 0 55776 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_492
timestamp 1698431365
transform 1 0 56448 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_556
timestamp 1698431365
transform 1 0 63616 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_562
timestamp 1698431365
transform 1 0 64288 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_594
timestamp 1698431365
transform 1 0 67872 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_610
timestamp 1698431365
transform 1 0 69664 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_618
timestamp 1698431365
transform 1 0 70560 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_622
timestamp 1698431365
transform 1 0 71008 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_626
timestamp 1698431365
transform 1 0 71456 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_632
timestamp 1698431365
transform 1 0 72128 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_634
timestamp 1698431365
transform 1 0 72352 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_643
timestamp 1698431365
transform 1 0 73360 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_659
timestamp 1698431365
transform 1 0 75152 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_669
timestamp 1698431365
transform 1 0 76272 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_685
timestamp 1698431365
transform 1 0 78064 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_687
timestamp 1698431365
transform 1 0 78288 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698431365
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698431365
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698431365
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698431365
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698431365
transform 1 0 13328 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698431365
transform 1 0 20496 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698431365
transform 1 0 21168 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698431365
transform 1 0 28336 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698431365
transform 1 0 29008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698431365
transform 1 0 36176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_317
timestamp 1698431365
transform 1 0 36848 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_381
timestamp 1698431365
transform 1 0 44016 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_387
timestamp 1698431365
transform 1 0 44688 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_395
timestamp 1698431365
transform 1 0 45584 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_412
timestamp 1698431365
transform 1 0 47488 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_428
timestamp 1698431365
transform 1 0 49280 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_436
timestamp 1698431365
transform 1 0 50176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_440
timestamp 1698431365
transform 1 0 50624 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_450
timestamp 1698431365
transform 1 0 51744 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_454
timestamp 1698431365
transform 1 0 52192 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_457
timestamp 1698431365
transform 1 0 52528 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_461
timestamp 1698431365
transform 1 0 52976 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_527
timestamp 1698431365
transform 1 0 60368 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_591
timestamp 1698431365
transform 1 0 67536 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_597
timestamp 1698431365
transform 1 0 68208 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_613
timestamp 1698431365
transform 1 0 70000 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_621
timestamp 1698431365
transform 1 0 70896 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_651
timestamp 1698431365
transform 1 0 74256 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_655
timestamp 1698431365
transform 1 0 74704 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_681
timestamp 1698431365
transform 1 0 77616 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_8
timestamp 1698431365
transform 1 0 2240 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_12
timestamp 1698431365
transform 1 0 2688 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_44
timestamp 1698431365
transform 1 0 6272 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_60
timestamp 1698431365
transform 1 0 8064 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_68
timestamp 1698431365
transform 1 0 8960 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698431365
transform 1 0 9408 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698431365
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698431365
transform 1 0 17248 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698431365
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698431365
transform 1 0 25088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698431365
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698431365
transform 1 0 32928 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_346
timestamp 1698431365
transform 1 0 40096 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_352
timestamp 1698431365
transform 1 0 40768 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_368
timestamp 1698431365
transform 1 0 42560 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_376
timestamp 1698431365
transform 1 0 43456 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_380
timestamp 1698431365
transform 1 0 43904 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_387
timestamp 1698431365
transform 1 0 44688 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_389
timestamp 1698431365
transform 1 0 44912 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_410
timestamp 1698431365
transform 1 0 47264 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_418
timestamp 1698431365
transform 1 0 48160 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_422
timestamp 1698431365
transform 1 0 48608 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_438
timestamp 1698431365
transform 1 0 50400 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_464
timestamp 1698431365
transform 1 0 53312 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_468
timestamp 1698431365
transform 1 0 53760 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_484
timestamp 1698431365
transform 1 0 55552 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_488
timestamp 1698431365
transform 1 0 56000 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_492
timestamp 1698431365
transform 1 0 56448 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_556
timestamp 1698431365
transform 1 0 63616 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_562
timestamp 1698431365
transform 1 0 64288 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_626
timestamp 1698431365
transform 1 0 71456 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_640
timestamp 1698431365
transform 1 0 73024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_644
timestamp 1698431365
transform 1 0 73472 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_653
timestamp 1698431365
transform 1 0 74480 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_657
timestamp 1698431365
transform 1 0 74928 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_675
timestamp 1698431365
transform 1 0 76944 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_685
timestamp 1698431365
transform 1 0 78064 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_687
timestamp 1698431365
transform 1 0 78288 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_8
timestamp 1698431365
transform 1 0 2240 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_12
timestamp 1698431365
transform 1 0 2688 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_28
timestamp 1698431365
transform 1 0 4480 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_32
timestamp 1698431365
transform 1 0 4928 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698431365
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698431365
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698431365
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698431365
transform 1 0 13328 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698431365
transform 1 0 20496 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698431365
transform 1 0 21168 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698431365
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698431365
transform 1 0 29008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698431365
transform 1 0 36176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_317
timestamp 1698431365
transform 1 0 36848 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_381
timestamp 1698431365
transform 1 0 44016 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_395
timestamp 1698431365
transform 1 0 45584 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_404
timestamp 1698431365
transform 1 0 46592 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_436
timestamp 1698431365
transform 1 0 50176 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_444
timestamp 1698431365
transform 1 0 51072 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_457
timestamp 1698431365
transform 1 0 52528 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_461
timestamp 1698431365
transform 1 0 52976 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_527
timestamp 1698431365
transform 1 0 60368 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_591
timestamp 1698431365
transform 1 0 67536 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_597
timestamp 1698431365
transform 1 0 68208 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_629
timestamp 1698431365
transform 1 0 71792 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_632
timestamp 1698431365
transform 1 0 72128 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_638
timestamp 1698431365
transform 1 0 72800 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_650
timestamp 1698431365
transform 1 0 74144 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_654
timestamp 1698431365
transform 1 0 74592 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_663
timestamp 1698431365
transform 1 0 75600 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_675
timestamp 1698431365
transform 1 0 76944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_685
timestamp 1698431365
transform 1 0 78064 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_687
timestamp 1698431365
transform 1 0 78288 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698431365
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698431365
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698431365
transform 1 0 9408 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698431365
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698431365
transform 1 0 17248 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698431365
transform 1 0 24416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698431365
transform 1 0 25088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698431365
transform 1 0 32256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698431365
transform 1 0 32928 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_346
timestamp 1698431365
transform 1 0 40096 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_352
timestamp 1698431365
transform 1 0 40768 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_384
timestamp 1698431365
transform 1 0 44352 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_388
timestamp 1698431365
transform 1 0 44800 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_391
timestamp 1698431365
transform 1 0 45136 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_407
timestamp 1698431365
transform 1 0 46928 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_415
timestamp 1698431365
transform 1 0 47824 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_419
timestamp 1698431365
transform 1 0 48272 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_422
timestamp 1698431365
transform 1 0 48608 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_486
timestamp 1698431365
transform 1 0 55776 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_492
timestamp 1698431365
transform 1 0 56448 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_556
timestamp 1698431365
transform 1 0 63616 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_562
timestamp 1698431365
transform 1 0 64288 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_594
timestamp 1698431365
transform 1 0 67872 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_610
timestamp 1698431365
transform 1 0 69664 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_618
timestamp 1698431365
transform 1 0 70560 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_646
timestamp 1698431365
transform 1 0 73696 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_665
timestamp 1698431365
transform 1 0 75824 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_669
timestamp 1698431365
transform 1 0 76272 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_678
timestamp 1698431365
transform 1 0 77280 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_8
timestamp 1698431365
transform 1 0 2240 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_12
timestamp 1698431365
transform 1 0 2688 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_28
timestamp 1698431365
transform 1 0 4480 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_32
timestamp 1698431365
transform 1 0 4928 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698431365
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698431365
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698431365
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698431365
transform 1 0 13328 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698431365
transform 1 0 20496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698431365
transform 1 0 21168 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698431365
transform 1 0 28336 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698431365
transform 1 0 29008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698431365
transform 1 0 36176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_317
timestamp 1698431365
transform 1 0 36848 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_381
timestamp 1698431365
transform 1 0 44016 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_387
timestamp 1698431365
transform 1 0 44688 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_391
timestamp 1698431365
transform 1 0 45136 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_407
timestamp 1698431365
transform 1 0 46928 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_439
timestamp 1698431365
transform 1 0 50512 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_457
timestamp 1698431365
transform 1 0 52528 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_465
timestamp 1698431365
transform 1 0 53424 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_471
timestamp 1698431365
transform 1 0 54096 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_503
timestamp 1698431365
transform 1 0 57680 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_519
timestamp 1698431365
transform 1 0 59472 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_523
timestamp 1698431365
transform 1 0 59920 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_527
timestamp 1698431365
transform 1 0 60368 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_591
timestamp 1698431365
transform 1 0 67536 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_597
timestamp 1698431365
transform 1 0 68208 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_613
timestamp 1698431365
transform 1 0 70000 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_621
timestamp 1698431365
transform 1 0 70896 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_625
timestamp 1698431365
transform 1 0 71344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_635
timestamp 1698431365
transform 1 0 72464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_639
timestamp 1698431365
transform 1 0 72912 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_641
timestamp 1698431365
transform 1 0 73136 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_667
timestamp 1698431365
transform 1 0 76048 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_669
timestamp 1698431365
transform 1 0 76272 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_684
timestamp 1698431365
transform 1 0 77952 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_8
timestamp 1698431365
transform 1 0 2240 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_12
timestamp 1698431365
transform 1 0 2688 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_44
timestamp 1698431365
transform 1 0 6272 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_60
timestamp 1698431365
transform 1 0 8064 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_68
timestamp 1698431365
transform 1 0 8960 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698431365
transform 1 0 9408 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698431365
transform 1 0 16576 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698431365
transform 1 0 17248 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698431365
transform 1 0 24416 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698431365
transform 1 0 25088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698431365
transform 1 0 32256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698431365
transform 1 0 32928 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_346
timestamp 1698431365
transform 1 0 40096 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_352
timestamp 1698431365
transform 1 0 40768 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_368
timestamp 1698431365
transform 1 0 42560 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_376
timestamp 1698431365
transform 1 0 43456 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_380
timestamp 1698431365
transform 1 0 43904 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_387
timestamp 1698431365
transform 1 0 44688 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_419
timestamp 1698431365
transform 1 0 48272 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_422
timestamp 1698431365
transform 1 0 48608 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_454
timestamp 1698431365
transform 1 0 52192 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_458
timestamp 1698431365
transform 1 0 52640 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_469
timestamp 1698431365
transform 1 0 53872 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_480
timestamp 1698431365
transform 1 0 55104 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_484
timestamp 1698431365
transform 1 0 55552 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_488
timestamp 1698431365
transform 1 0 56000 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_492
timestamp 1698431365
transform 1 0 56448 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_556
timestamp 1698431365
transform 1 0 63616 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_562
timestamp 1698431365
transform 1 0 64288 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_594
timestamp 1698431365
transform 1 0 67872 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_610
timestamp 1698431365
transform 1 0 69664 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_618
timestamp 1698431365
transform 1 0 70560 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_622
timestamp 1698431365
transform 1 0 71008 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_626
timestamp 1698431365
transform 1 0 71456 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_632
timestamp 1698431365
transform 1 0 72128 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_640
timestamp 1698431365
transform 1 0 73024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_644
timestamp 1698431365
transform 1 0 73472 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_663
timestamp 1698431365
transform 1 0 75600 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_667
timestamp 1698431365
transform 1 0 76048 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_684
timestamp 1698431365
transform 1 0 77952 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_8
timestamp 1698431365
transform 1 0 2240 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_12
timestamp 1698431365
transform 1 0 2688 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_28
timestamp 1698431365
transform 1 0 4480 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_32
timestamp 1698431365
transform 1 0 4928 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698431365
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698431365
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698431365
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698431365
transform 1 0 13328 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698431365
transform 1 0 20496 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698431365
transform 1 0 21168 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698431365
transform 1 0 28336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698431365
transform 1 0 29008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698431365
transform 1 0 36176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_317
timestamp 1698431365
transform 1 0 36848 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_381
timestamp 1698431365
transform 1 0 44016 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_391
timestamp 1698431365
transform 1 0 45136 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_401
timestamp 1698431365
transform 1 0 46256 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_433
timestamp 1698431365
transform 1 0 49840 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_449
timestamp 1698431365
transform 1 0 51632 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_453
timestamp 1698431365
transform 1 0 52080 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_457
timestamp 1698431365
transform 1 0 52528 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_461
timestamp 1698431365
transform 1 0 52976 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_463
timestamp 1698431365
transform 1 0 53200 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_482
timestamp 1698431365
transform 1 0 55328 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_486
timestamp 1698431365
transform 1 0 55776 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_518
timestamp 1698431365
transform 1 0 59360 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_522
timestamp 1698431365
transform 1 0 59808 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_524
timestamp 1698431365
transform 1 0 60032 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_527
timestamp 1698431365
transform 1 0 60368 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_591
timestamp 1698431365
transform 1 0 67536 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_597
timestamp 1698431365
transform 1 0 68208 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_613
timestamp 1698431365
transform 1 0 70000 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_617
timestamp 1698431365
transform 1 0 70448 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_619
timestamp 1698431365
transform 1 0 70672 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_652
timestamp 1698431365
transform 1 0 74368 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698431365
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698431365
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698431365
transform 1 0 9408 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698431365
transform 1 0 16576 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698431365
transform 1 0 17248 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698431365
transform 1 0 24416 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698431365
transform 1 0 25088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698431365
transform 1 0 32256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698431365
transform 1 0 32928 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_346
timestamp 1698431365
transform 1 0 40096 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_352
timestamp 1698431365
transform 1 0 40768 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_368
timestamp 1698431365
transform 1 0 42560 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_376
timestamp 1698431365
transform 1 0 43456 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_380
timestamp 1698431365
transform 1 0 43904 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_382
timestamp 1698431365
transform 1 0 44128 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_389
timestamp 1698431365
transform 1 0 44912 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_409
timestamp 1698431365
transform 1 0 47152 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_417
timestamp 1698431365
transform 1 0 48048 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_419
timestamp 1698431365
transform 1 0 48272 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_422
timestamp 1698431365
transform 1 0 48608 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_454
timestamp 1698431365
transform 1 0 52192 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_470
timestamp 1698431365
transform 1 0 53984 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_472
timestamp 1698431365
transform 1 0 54208 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_475
timestamp 1698431365
transform 1 0 54544 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_483
timestamp 1698431365
transform 1 0 55440 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_487
timestamp 1698431365
transform 1 0 55888 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_489
timestamp 1698431365
transform 1 0 56112 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_492
timestamp 1698431365
transform 1 0 56448 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_556
timestamp 1698431365
transform 1 0 63616 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_562
timestamp 1698431365
transform 1 0 64288 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_626
timestamp 1698431365
transform 1 0 71456 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_632
timestamp 1698431365
transform 1 0 72128 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_634
timestamp 1698431365
transform 1 0 72352 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_669
timestamp 1698431365
transform 1 0 76272 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_678
timestamp 1698431365
transform 1 0 77280 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_8
timestamp 1698431365
transform 1 0 2240 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_12
timestamp 1698431365
transform 1 0 2688 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_28
timestamp 1698431365
transform 1 0 4480 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_32
timestamp 1698431365
transform 1 0 4928 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698431365
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698431365
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698431365
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698431365
transform 1 0 13328 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698431365
transform 1 0 20496 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698431365
transform 1 0 21168 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698431365
transform 1 0 28336 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698431365
transform 1 0 29008 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698431365
transform 1 0 36176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_317
timestamp 1698431365
transform 1 0 36848 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_381
timestamp 1698431365
transform 1 0 44016 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_391
timestamp 1698431365
transform 1 0 45136 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_395
timestamp 1698431365
transform 1 0 45584 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_427
timestamp 1698431365
transform 1 0 49168 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_443
timestamp 1698431365
transform 1 0 50960 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_451
timestamp 1698431365
transform 1 0 51856 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_457
timestamp 1698431365
transform 1 0 52528 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_521
timestamp 1698431365
transform 1 0 59696 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_527
timestamp 1698431365
transform 1 0 60368 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_591
timestamp 1698431365
transform 1 0 67536 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_597
timestamp 1698431365
transform 1 0 68208 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_601
timestamp 1698431365
transform 1 0 68656 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_603
timestamp 1698431365
transform 1 0 68880 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_606
timestamp 1698431365
transform 1 0 69216 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_622
timestamp 1698431365
transform 1 0 71008 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_625
timestamp 1698431365
transform 1 0 71344 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_631
timestamp 1698431365
transform 1 0 72016 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_633
timestamp 1698431365
transform 1 0 72240 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_636
timestamp 1698431365
transform 1 0 72576 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_640
timestamp 1698431365
transform 1 0 73024 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_644
timestamp 1698431365
transform 1 0 73472 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_646
timestamp 1698431365
transform 1 0 73696 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_649
timestamp 1698431365
transform 1 0 74032 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_8
timestamp 1698431365
transform 1 0 2240 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_12
timestamp 1698431365
transform 1 0 2688 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_44
timestamp 1698431365
transform 1 0 6272 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_60
timestamp 1698431365
transform 1 0 8064 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_68
timestamp 1698431365
transform 1 0 8960 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698431365
transform 1 0 9408 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698431365
transform 1 0 16576 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_142
timestamp 1698431365
transform 1 0 17248 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_206
timestamp 1698431365
transform 1 0 24416 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_212
timestamp 1698431365
transform 1 0 25088 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_276
timestamp 1698431365
transform 1 0 32256 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698431365
transform 1 0 32928 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_346
timestamp 1698431365
transform 1 0 40096 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_352
timestamp 1698431365
transform 1 0 40768 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_416
timestamp 1698431365
transform 1 0 47936 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_422
timestamp 1698431365
transform 1 0 48608 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_486
timestamp 1698431365
transform 1 0 55776 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_492
timestamp 1698431365
transform 1 0 56448 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_556
timestamp 1698431365
transform 1 0 63616 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_562
timestamp 1698431365
transform 1 0 64288 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_594
timestamp 1698431365
transform 1 0 67872 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_597
timestamp 1698431365
transform 1 0 68208 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_599
timestamp 1698431365
transform 1 0 68432 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_612
timestamp 1698431365
transform 1 0 69888 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_616
timestamp 1698431365
transform 1 0 70336 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_629
timestamp 1698431365
transform 1 0 71792 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_648
timestamp 1698431365
transform 1 0 73920 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_663
timestamp 1698431365
transform 1 0 75600 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_2
timestamp 1698431365
transform 1 0 1568 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_12
timestamp 1698431365
transform 1 0 2688 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_16
timestamp 1698431365
transform 1 0 3136 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_32
timestamp 1698431365
transform 1 0 4928 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_34
timestamp 1698431365
transform 1 0 5152 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_37
timestamp 1698431365
transform 1 0 5488 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_101
timestamp 1698431365
transform 1 0 12656 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_107
timestamp 1698431365
transform 1 0 13328 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_171
timestamp 1698431365
transform 1 0 20496 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_177
timestamp 1698431365
transform 1 0 21168 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_241
timestamp 1698431365
transform 1 0 28336 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_247
timestamp 1698431365
transform 1 0 29008 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_311
timestamp 1698431365
transform 1 0 36176 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_317
timestamp 1698431365
transform 1 0 36848 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_381
timestamp 1698431365
transform 1 0 44016 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_387
timestamp 1698431365
transform 1 0 44688 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_451
timestamp 1698431365
transform 1 0 51856 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_457
timestamp 1698431365
transform 1 0 52528 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_521
timestamp 1698431365
transform 1 0 59696 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_527
timestamp 1698431365
transform 1 0 60368 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_559
timestamp 1698431365
transform 1 0 63952 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_575
timestamp 1698431365
transform 1 0 65744 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_583
timestamp 1698431365
transform 1 0 66640 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_616
timestamp 1698431365
transform 1 0 70336 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_620
timestamp 1698431365
transform 1 0 70784 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_629
timestamp 1698431365
transform 1 0 71792 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_661
timestamp 1698431365
transform 1 0 75376 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_683
timestamp 1698431365
transform 1 0 77840 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_687
timestamp 1698431365
transform 1 0 78288 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_28
timestamp 1698431365
transform 1 0 4480 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_60
timestamp 1698431365
transform 1 0 8064 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_68
timestamp 1698431365
transform 1 0 8960 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_72
timestamp 1698431365
transform 1 0 9408 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_136
timestamp 1698431365
transform 1 0 16576 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_142
timestamp 1698431365
transform 1 0 17248 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_206
timestamp 1698431365
transform 1 0 24416 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_212
timestamp 1698431365
transform 1 0 25088 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_276
timestamp 1698431365
transform 1 0 32256 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_282
timestamp 1698431365
transform 1 0 32928 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_346
timestamp 1698431365
transform 1 0 40096 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_352
timestamp 1698431365
transform 1 0 40768 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_375
timestamp 1698431365
transform 1 0 43344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_379
timestamp 1698431365
transform 1 0 43792 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_383
timestamp 1698431365
transform 1 0 44240 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_415
timestamp 1698431365
transform 1 0 47824 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_419
timestamp 1698431365
transform 1 0 48272 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_422
timestamp 1698431365
transform 1 0 48608 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_486
timestamp 1698431365
transform 1 0 55776 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_492
timestamp 1698431365
transform 1 0 56448 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_524
timestamp 1698431365
transform 1 0 60032 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_548
timestamp 1698431365
transform 1 0 62720 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_556
timestamp 1698431365
transform 1 0 63616 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_562
timestamp 1698431365
transform 1 0 64288 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_604
timestamp 1698431365
transform 1 0 68992 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_608
timestamp 1698431365
transform 1 0 69440 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_612
timestamp 1698431365
transform 1 0 69888 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_614
timestamp 1698431365
transform 1 0 70112 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_623
timestamp 1698431365
transform 1 0 71120 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_627
timestamp 1698431365
transform 1 0 71568 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_629
timestamp 1698431365
transform 1 0 71792 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_632
timestamp 1698431365
transform 1 0 72128 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_647
timestamp 1698431365
transform 1 0 73808 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_654
timestamp 1698431365
transform 1 0 74592 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_661
timestamp 1698431365
transform 1 0 75376 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_28
timestamp 1698431365
transform 1 0 4480 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_32
timestamp 1698431365
transform 1 0 4928 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_34
timestamp 1698431365
transform 1 0 5152 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_37
timestamp 1698431365
transform 1 0 5488 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_101
timestamp 1698431365
transform 1 0 12656 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_107
timestamp 1698431365
transform 1 0 13328 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_171
timestamp 1698431365
transform 1 0 20496 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_177
timestamp 1698431365
transform 1 0 21168 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_241
timestamp 1698431365
transform 1 0 28336 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_247
timestamp 1698431365
transform 1 0 29008 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_311
timestamp 1698431365
transform 1 0 36176 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_317
timestamp 1698431365
transform 1 0 36848 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_381
timestamp 1698431365
transform 1 0 44016 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_387
timestamp 1698431365
transform 1 0 44688 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_451
timestamp 1698431365
transform 1 0 51856 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_457
timestamp 1698431365
transform 1 0 52528 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_521
timestamp 1698431365
transform 1 0 59696 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_527
timestamp 1698431365
transform 1 0 60368 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_531
timestamp 1698431365
transform 1 0 60816 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_533
timestamp 1698431365
transform 1 0 61040 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_536
timestamp 1698431365
transform 1 0 61376 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_542
timestamp 1698431365
transform 1 0 62048 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_550
timestamp 1698431365
transform 1 0 62944 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_556
timestamp 1698431365
transform 1 0 63616 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_585
timestamp 1698431365
transform 1 0 66864 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_589
timestamp 1698431365
transform 1 0 67312 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_593
timestamp 1698431365
transform 1 0 67760 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_610
timestamp 1698431365
transform 1 0 69664 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_628
timestamp 1698431365
transform 1 0 71680 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_632
timestamp 1698431365
transform 1 0 72128 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_636
timestamp 1698431365
transform 1 0 72576 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_652
timestamp 1698431365
transform 1 0 74368 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_656
timestamp 1698431365
transform 1 0 74816 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_26
timestamp 1698431365
transform 1 0 4256 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_30
timestamp 1698431365
transform 1 0 4704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_34
timestamp 1698431365
transform 1 0 5152 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_47_38
timestamp 1698431365
transform 1 0 5600 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_72
timestamp 1698431365
transform 1 0 9408 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_136
timestamp 1698431365
transform 1 0 16576 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_142
timestamp 1698431365
transform 1 0 17248 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_206
timestamp 1698431365
transform 1 0 24416 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_212
timestamp 1698431365
transform 1 0 25088 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_276
timestamp 1698431365
transform 1 0 32256 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_282
timestamp 1698431365
transform 1 0 32928 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_346
timestamp 1698431365
transform 1 0 40096 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_352
timestamp 1698431365
transform 1 0 40768 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_416
timestamp 1698431365
transform 1 0 47936 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_422
timestamp 1698431365
transform 1 0 48608 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_486
timestamp 1698431365
transform 1 0 55776 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_492
timestamp 1698431365
transform 1 0 56448 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_508
timestamp 1698431365
transform 1 0 58240 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_516
timestamp 1698431365
transform 1 0 59136 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_520
timestamp 1698431365
transform 1 0 59584 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_534
timestamp 1698431365
transform 1 0 61152 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_588
timestamp 1698431365
transform 1 0 67200 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_592
timestamp 1698431365
transform 1 0 67648 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_612
timestamp 1698431365
transform 1 0 69888 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_616
timestamp 1698431365
transform 1 0 70336 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_623
timestamp 1698431365
transform 1 0 71120 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_627
timestamp 1698431365
transform 1 0 71568 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_629
timestamp 1698431365
transform 1 0 71792 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_632
timestamp 1698431365
transform 1 0 72128 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_636
timestamp 1698431365
transform 1 0 72576 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_640
timestamp 1698431365
transform 1 0 73024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_28
timestamp 1698431365
transform 1 0 4480 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_32
timestamp 1698431365
transform 1 0 4928 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_34
timestamp 1698431365
transform 1 0 5152 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_37
timestamp 1698431365
transform 1 0 5488 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_101
timestamp 1698431365
transform 1 0 12656 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_107
timestamp 1698431365
transform 1 0 13328 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_171
timestamp 1698431365
transform 1 0 20496 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_177
timestamp 1698431365
transform 1 0 21168 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_241
timestamp 1698431365
transform 1 0 28336 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_247
timestamp 1698431365
transform 1 0 29008 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_311
timestamp 1698431365
transform 1 0 36176 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_317
timestamp 1698431365
transform 1 0 36848 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_381
timestamp 1698431365
transform 1 0 44016 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_387
timestamp 1698431365
transform 1 0 44688 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_451
timestamp 1698431365
transform 1 0 51856 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_457
timestamp 1698431365
transform 1 0 52528 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_473
timestamp 1698431365
transform 1 0 54320 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_477
timestamp 1698431365
transform 1 0 54768 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_489
timestamp 1698431365
transform 1 0 56112 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_493
timestamp 1698431365
transform 1 0 56560 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_497
timestamp 1698431365
transform 1 0 57008 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_500
timestamp 1698431365
transform 1 0 57344 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_504
timestamp 1698431365
transform 1 0 57792 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_566
timestamp 1698431365
transform 1 0 64736 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_570
timestamp 1698431365
transform 1 0 65184 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_572
timestamp 1698431365
transform 1 0 65408 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_586
timestamp 1698431365
transform 1 0 66976 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_594
timestamp 1698431365
transform 1 0 67872 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_597
timestamp 1698431365
transform 1 0 68208 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_601
timestamp 1698431365
transform 1 0 68656 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_611
timestamp 1698431365
transform 1 0 69776 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_630
timestamp 1698431365
transform 1 0 71904 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_638
timestamp 1698431365
transform 1 0 72800 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_640
timestamp 1698431365
transform 1 0 73024 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_683
timestamp 1698431365
transform 1 0 77840 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_687
timestamp 1698431365
transform 1 0 78288 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_28
timestamp 1698431365
transform 1 0 4480 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_32
timestamp 1698431365
transform 1 0 4928 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_64
timestamp 1698431365
transform 1 0 8512 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_68
timestamp 1698431365
transform 1 0 8960 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_72
timestamp 1698431365
transform 1 0 9408 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_136
timestamp 1698431365
transform 1 0 16576 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_142
timestamp 1698431365
transform 1 0 17248 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_206
timestamp 1698431365
transform 1 0 24416 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_212
timestamp 1698431365
transform 1 0 25088 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_276
timestamp 1698431365
transform 1 0 32256 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_282
timestamp 1698431365
transform 1 0 32928 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_346
timestamp 1698431365
transform 1 0 40096 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_352
timestamp 1698431365
transform 1 0 40768 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_416
timestamp 1698431365
transform 1 0 47936 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_422
timestamp 1698431365
transform 1 0 48608 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_454
timestamp 1698431365
transform 1 0 52192 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_470
timestamp 1698431365
transform 1 0 53984 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_474
timestamp 1698431365
transform 1 0 54432 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_476
timestamp 1698431365
transform 1 0 54656 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_487
timestamp 1698431365
transform 1 0 55888 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_489
timestamp 1698431365
transform 1 0 56112 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_508
timestamp 1698431365
transform 1 0 58240 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_516
timestamp 1698431365
transform 1 0 59136 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_520
timestamp 1698431365
transform 1 0 59584 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_522
timestamp 1698431365
transform 1 0 59808 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_531
timestamp 1698431365
transform 1 0 60816 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_535
timestamp 1698431365
transform 1 0 61264 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_544
timestamp 1698431365
transform 1 0 62272 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_554
timestamp 1698431365
transform 1 0 63392 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_558
timestamp 1698431365
transform 1 0 63840 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_570
timestamp 1698431365
transform 1 0 65184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_574
timestamp 1698431365
transform 1 0 65632 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_578
timestamp 1698431365
transform 1 0 66080 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_612
timestamp 1698431365
transform 1 0 69888 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_616
timestamp 1698431365
transform 1 0 70336 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_620
timestamp 1698431365
transform 1 0 70784 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_624
timestamp 1698431365
transform 1 0 71232 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_628
timestamp 1698431365
transform 1 0 71680 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_632
timestamp 1698431365
transform 1 0 72128 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_648
timestamp 1698431365
transform 1 0 73920 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_651
timestamp 1698431365
transform 1 0 74256 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_653
timestamp 1698431365
transform 1 0 74480 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_28
timestamp 1698431365
transform 1 0 4480 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_32
timestamp 1698431365
transform 1 0 4928 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_34
timestamp 1698431365
transform 1 0 5152 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_37
timestamp 1698431365
transform 1 0 5488 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_101
timestamp 1698431365
transform 1 0 12656 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_107
timestamp 1698431365
transform 1 0 13328 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_171
timestamp 1698431365
transform 1 0 20496 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_177
timestamp 1698431365
transform 1 0 21168 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_241
timestamp 1698431365
transform 1 0 28336 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_247
timestamp 1698431365
transform 1 0 29008 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_311
timestamp 1698431365
transform 1 0 36176 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_317
timestamp 1698431365
transform 1 0 36848 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_381
timestamp 1698431365
transform 1 0 44016 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_387
timestamp 1698431365
transform 1 0 44688 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_451
timestamp 1698431365
transform 1 0 51856 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_457
timestamp 1698431365
transform 1 0 52528 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_473
timestamp 1698431365
transform 1 0 54320 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_481
timestamp 1698431365
transform 1 0 55216 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_490
timestamp 1698431365
transform 1 0 56224 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_492
timestamp 1698431365
transform 1 0 56448 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_509
timestamp 1698431365
transform 1 0 58352 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_527
timestamp 1698431365
transform 1 0 60368 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_543
timestamp 1698431365
transform 1 0 62160 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_546
timestamp 1698431365
transform 1 0 62496 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_578
timestamp 1698431365
transform 1 0 66080 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_594
timestamp 1698431365
transform 1 0 67872 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_597
timestamp 1698431365
transform 1 0 68208 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_661
timestamp 1698431365
transform 1 0 75376 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_667
timestamp 1698431365
transform 1 0 76048 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_2
timestamp 1698431365
transform 1 0 1568 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_4
timestamp 1698431365
transform 1 0 1792 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_51_17
timestamp 1698431365
transform 1 0 3248 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_49
timestamp 1698431365
transform 1 0 6832 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_65
timestamp 1698431365
transform 1 0 8624 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_69
timestamp 1698431365
transform 1 0 9072 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_72
timestamp 1698431365
transform 1 0 9408 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_136
timestamp 1698431365
transform 1 0 16576 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_142
timestamp 1698431365
transform 1 0 17248 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_206
timestamp 1698431365
transform 1 0 24416 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_212
timestamp 1698431365
transform 1 0 25088 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_276
timestamp 1698431365
transform 1 0 32256 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_282
timestamp 1698431365
transform 1 0 32928 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_346
timestamp 1698431365
transform 1 0 40096 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_352
timestamp 1698431365
transform 1 0 40768 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_416
timestamp 1698431365
transform 1 0 47936 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_422
timestamp 1698431365
transform 1 0 48608 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_486
timestamp 1698431365
transform 1 0 55776 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_51_500
timestamp 1698431365
transform 1 0 57344 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_532
timestamp 1698431365
transform 1 0 60928 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_548
timestamp 1698431365
transform 1 0 62720 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_556
timestamp 1698431365
transform 1 0 63616 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_562
timestamp 1698431365
transform 1 0 64288 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_626
timestamp 1698431365
transform 1 0 71456 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_51_632
timestamp 1698431365
transform 1 0 72128 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_664
timestamp 1698431365
transform 1 0 75712 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_672
timestamp 1698431365
transform 1 0 76608 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_684
timestamp 1698431365
transform 1 0 77952 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_28
timestamp 1698431365
transform 1 0 4480 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_32
timestamp 1698431365
transform 1 0 4928 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_34
timestamp 1698431365
transform 1 0 5152 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_37
timestamp 1698431365
transform 1 0 5488 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_101
timestamp 1698431365
transform 1 0 12656 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_107
timestamp 1698431365
transform 1 0 13328 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_171
timestamp 1698431365
transform 1 0 20496 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_177
timestamp 1698431365
transform 1 0 21168 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_241
timestamp 1698431365
transform 1 0 28336 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_247
timestamp 1698431365
transform 1 0 29008 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_311
timestamp 1698431365
transform 1 0 36176 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_317
timestamp 1698431365
transform 1 0 36848 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_381
timestamp 1698431365
transform 1 0 44016 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_387
timestamp 1698431365
transform 1 0 44688 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_451
timestamp 1698431365
transform 1 0 51856 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_457
timestamp 1698431365
transform 1 0 52528 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_521
timestamp 1698431365
transform 1 0 59696 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_527
timestamp 1698431365
transform 1 0 60368 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_591
timestamp 1698431365
transform 1 0 67536 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_597
timestamp 1698431365
transform 1 0 68208 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_661
timestamp 1698431365
transform 1 0 75376 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_667
timestamp 1698431365
transform 1 0 76048 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_683
timestamp 1698431365
transform 1 0 77840 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_685
timestamp 1698431365
transform 1 0 78064 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_53_28
timestamp 1698431365
transform 1 0 4480 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_60
timestamp 1698431365
transform 1 0 8064 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_68
timestamp 1698431365
transform 1 0 8960 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_72
timestamp 1698431365
transform 1 0 9408 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_136
timestamp 1698431365
transform 1 0 16576 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_142
timestamp 1698431365
transform 1 0 17248 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_206
timestamp 1698431365
transform 1 0 24416 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_212
timestamp 1698431365
transform 1 0 25088 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_276
timestamp 1698431365
transform 1 0 32256 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_282
timestamp 1698431365
transform 1 0 32928 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_346
timestamp 1698431365
transform 1 0 40096 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_352
timestamp 1698431365
transform 1 0 40768 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_416
timestamp 1698431365
transform 1 0 47936 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_422
timestamp 1698431365
transform 1 0 48608 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_486
timestamp 1698431365
transform 1 0 55776 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_492
timestamp 1698431365
transform 1 0 56448 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_556
timestamp 1698431365
transform 1 0 63616 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_562
timestamp 1698431365
transform 1 0 64288 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_626
timestamp 1698431365
transform 1 0 71456 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_53_632
timestamp 1698431365
transform 1 0 72128 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_664
timestamp 1698431365
transform 1 0 75712 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_2
timestamp 1698431365
transform 1 0 1568 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_4
timestamp 1698431365
transform 1 0 1792 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_23
timestamp 1698431365
transform 1 0 3920 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_27
timestamp 1698431365
transform 1 0 4368 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_37
timestamp 1698431365
transform 1 0 5488 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_101
timestamp 1698431365
transform 1 0 12656 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_107
timestamp 1698431365
transform 1 0 13328 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_171
timestamp 1698431365
transform 1 0 20496 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_177
timestamp 1698431365
transform 1 0 21168 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_241
timestamp 1698431365
transform 1 0 28336 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_247
timestamp 1698431365
transform 1 0 29008 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_311
timestamp 1698431365
transform 1 0 36176 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_317
timestamp 1698431365
transform 1 0 36848 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_381
timestamp 1698431365
transform 1 0 44016 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_387
timestamp 1698431365
transform 1 0 44688 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_451
timestamp 1698431365
transform 1 0 51856 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_457
timestamp 1698431365
transform 1 0 52528 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_521
timestamp 1698431365
transform 1 0 59696 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_527
timestamp 1698431365
transform 1 0 60368 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_591
timestamp 1698431365
transform 1 0 67536 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_597
timestamp 1698431365
transform 1 0 68208 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_661
timestamp 1698431365
transform 1 0 75376 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_667
timestamp 1698431365
transform 1 0 76048 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_675
timestamp 1698431365
transform 1 0 76944 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_679
timestamp 1698431365
transform 1 0 77392 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_55_28
timestamp 1698431365
transform 1 0 4480 0 -1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_60
timestamp 1698431365
transform 1 0 8064 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_68
timestamp 1698431365
transform 1 0 8960 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_72
timestamp 1698431365
transform 1 0 9408 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_136
timestamp 1698431365
transform 1 0 16576 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_142
timestamp 1698431365
transform 1 0 17248 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_206
timestamp 1698431365
transform 1 0 24416 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_212
timestamp 1698431365
transform 1 0 25088 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_276
timestamp 1698431365
transform 1 0 32256 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_282
timestamp 1698431365
transform 1 0 32928 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_346
timestamp 1698431365
transform 1 0 40096 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_352
timestamp 1698431365
transform 1 0 40768 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_416
timestamp 1698431365
transform 1 0 47936 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_422
timestamp 1698431365
transform 1 0 48608 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_486
timestamp 1698431365
transform 1 0 55776 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_492
timestamp 1698431365
transform 1 0 56448 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_556
timestamp 1698431365
transform 1 0 63616 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_562
timestamp 1698431365
transform 1 0 64288 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_626
timestamp 1698431365
transform 1 0 71456 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_55_632
timestamp 1698431365
transform 1 0 72128 0 -1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_664
timestamp 1698431365
transform 1 0 75712 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_680
timestamp 1698431365
transform 1 0 77504 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_28
timestamp 1698431365
transform 1 0 4480 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_32
timestamp 1698431365
transform 1 0 4928 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_34
timestamp 1698431365
transform 1 0 5152 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_37
timestamp 1698431365
transform 1 0 5488 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_101
timestamp 1698431365
transform 1 0 12656 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_107
timestamp 1698431365
transform 1 0 13328 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_171
timestamp 1698431365
transform 1 0 20496 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_177
timestamp 1698431365
transform 1 0 21168 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_241
timestamp 1698431365
transform 1 0 28336 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_247
timestamp 1698431365
transform 1 0 29008 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_311
timestamp 1698431365
transform 1 0 36176 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_317
timestamp 1698431365
transform 1 0 36848 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_381
timestamp 1698431365
transform 1 0 44016 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_387
timestamp 1698431365
transform 1 0 44688 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_451
timestamp 1698431365
transform 1 0 51856 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_457
timestamp 1698431365
transform 1 0 52528 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_521
timestamp 1698431365
transform 1 0 59696 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_527
timestamp 1698431365
transform 1 0 60368 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_591
timestamp 1698431365
transform 1 0 67536 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_597
timestamp 1698431365
transform 1 0 68208 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_661
timestamp 1698431365
transform 1 0 75376 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_667
timestamp 1698431365
transform 1 0 76048 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_675
timestamp 1698431365
transform 1 0 76944 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_679
timestamp 1698431365
transform 1 0 77392 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_2
timestamp 1698431365
transform 1 0 1568 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_4
timestamp 1698431365
transform 1 0 1792 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_57_23
timestamp 1698431365
transform 1 0 3920 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_55
timestamp 1698431365
transform 1 0 7504 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_63
timestamp 1698431365
transform 1 0 8400 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_67
timestamp 1698431365
transform 1 0 8848 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_69
timestamp 1698431365
transform 1 0 9072 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_72
timestamp 1698431365
transform 1 0 9408 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_136
timestamp 1698431365
transform 1 0 16576 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_142
timestamp 1698431365
transform 1 0 17248 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_206
timestamp 1698431365
transform 1 0 24416 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_212
timestamp 1698431365
transform 1 0 25088 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_276
timestamp 1698431365
transform 1 0 32256 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_282
timestamp 1698431365
transform 1 0 32928 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_346
timestamp 1698431365
transform 1 0 40096 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_352
timestamp 1698431365
transform 1 0 40768 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_416
timestamp 1698431365
transform 1 0 47936 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_422
timestamp 1698431365
transform 1 0 48608 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_486
timestamp 1698431365
transform 1 0 55776 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_492
timestamp 1698431365
transform 1 0 56448 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_556
timestamp 1698431365
transform 1 0 63616 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_562
timestamp 1698431365
transform 1 0 64288 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_626
timestamp 1698431365
transform 1 0 71456 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_57_632
timestamp 1698431365
transform 1 0 72128 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_664
timestamp 1698431365
transform 1 0 75712 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_28
timestamp 1698431365
transform 1 0 4480 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_32
timestamp 1698431365
transform 1 0 4928 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_34
timestamp 1698431365
transform 1 0 5152 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_37
timestamp 1698431365
transform 1 0 5488 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_101
timestamp 1698431365
transform 1 0 12656 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_107
timestamp 1698431365
transform 1 0 13328 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_171
timestamp 1698431365
transform 1 0 20496 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_177
timestamp 1698431365
transform 1 0 21168 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_241
timestamp 1698431365
transform 1 0 28336 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_247
timestamp 1698431365
transform 1 0 29008 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_311
timestamp 1698431365
transform 1 0 36176 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_317
timestamp 1698431365
transform 1 0 36848 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_381
timestamp 1698431365
transform 1 0 44016 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_387
timestamp 1698431365
transform 1 0 44688 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_451
timestamp 1698431365
transform 1 0 51856 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_457
timestamp 1698431365
transform 1 0 52528 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_521
timestamp 1698431365
transform 1 0 59696 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_527
timestamp 1698431365
transform 1 0 60368 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_591
timestamp 1698431365
transform 1 0 67536 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_597
timestamp 1698431365
transform 1 0 68208 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_661
timestamp 1698431365
transform 1 0 75376 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_667
timestamp 1698431365
transform 1 0 76048 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_675
timestamp 1698431365
transform 1 0 76944 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_679
timestamp 1698431365
transform 1 0 77392 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_59_28
timestamp 1698431365
transform 1 0 4480 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_60
timestamp 1698431365
transform 1 0 8064 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_68
timestamp 1698431365
transform 1 0 8960 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_72
timestamp 1698431365
transform 1 0 9408 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_136
timestamp 1698431365
transform 1 0 16576 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_142
timestamp 1698431365
transform 1 0 17248 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_206
timestamp 1698431365
transform 1 0 24416 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_212
timestamp 1698431365
transform 1 0 25088 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_276
timestamp 1698431365
transform 1 0 32256 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_282
timestamp 1698431365
transform 1 0 32928 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_346
timestamp 1698431365
transform 1 0 40096 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_352
timestamp 1698431365
transform 1 0 40768 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_416
timestamp 1698431365
transform 1 0 47936 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_422
timestamp 1698431365
transform 1 0 48608 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_486
timestamp 1698431365
transform 1 0 55776 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_492
timestamp 1698431365
transform 1 0 56448 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_556
timestamp 1698431365
transform 1 0 63616 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_562
timestamp 1698431365
transform 1 0 64288 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_626
timestamp 1698431365
transform 1 0 71456 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_59_632
timestamp 1698431365
transform 1 0 72128 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_664
timestamp 1698431365
transform 1 0 75712 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_680
timestamp 1698431365
transform 1 0 77504 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_28
timestamp 1698431365
transform 1 0 4480 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_32
timestamp 1698431365
transform 1 0 4928 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_34
timestamp 1698431365
transform 1 0 5152 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_37
timestamp 1698431365
transform 1 0 5488 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_101
timestamp 1698431365
transform 1 0 12656 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_107
timestamp 1698431365
transform 1 0 13328 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_171
timestamp 1698431365
transform 1 0 20496 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_177
timestamp 1698431365
transform 1 0 21168 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_241
timestamp 1698431365
transform 1 0 28336 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_247
timestamp 1698431365
transform 1 0 29008 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_311
timestamp 1698431365
transform 1 0 36176 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_317
timestamp 1698431365
transform 1 0 36848 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_381
timestamp 1698431365
transform 1 0 44016 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_387
timestamp 1698431365
transform 1 0 44688 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_451
timestamp 1698431365
transform 1 0 51856 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_457
timestamp 1698431365
transform 1 0 52528 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_521
timestamp 1698431365
transform 1 0 59696 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_527
timestamp 1698431365
transform 1 0 60368 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_591
timestamp 1698431365
transform 1 0 67536 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_597
timestamp 1698431365
transform 1 0 68208 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_661
timestamp 1698431365
transform 1 0 75376 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_667
timestamp 1698431365
transform 1 0 76048 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_675
timestamp 1698431365
transform 1 0 76944 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_679
timestamp 1698431365
transform 1 0 77392 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_2
timestamp 1698431365
transform 1 0 1568 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_24
timestamp 1698431365
transform 1 0 4032 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_56
timestamp 1698431365
transform 1 0 7616 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_64
timestamp 1698431365
transform 1 0 8512 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_68
timestamp 1698431365
transform 1 0 8960 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_72
timestamp 1698431365
transform 1 0 9408 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_136
timestamp 1698431365
transform 1 0 16576 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_142
timestamp 1698431365
transform 1 0 17248 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_206
timestamp 1698431365
transform 1 0 24416 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_212
timestamp 1698431365
transform 1 0 25088 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_276
timestamp 1698431365
transform 1 0 32256 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_282
timestamp 1698431365
transform 1 0 32928 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_346
timestamp 1698431365
transform 1 0 40096 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_352
timestamp 1698431365
transform 1 0 40768 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_416
timestamp 1698431365
transform 1 0 47936 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_422
timestamp 1698431365
transform 1 0 48608 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_486
timestamp 1698431365
transform 1 0 55776 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_492
timestamp 1698431365
transform 1 0 56448 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_556
timestamp 1698431365
transform 1 0 63616 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_562
timestamp 1698431365
transform 1 0 64288 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_626
timestamp 1698431365
transform 1 0 71456 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_632
timestamp 1698431365
transform 1 0 72128 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_664
timestamp 1698431365
transform 1 0 75712 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_28
timestamp 1698431365
transform 1 0 4480 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_32
timestamp 1698431365
transform 1 0 4928 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_34
timestamp 1698431365
transform 1 0 5152 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_37
timestamp 1698431365
transform 1 0 5488 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_101
timestamp 1698431365
transform 1 0 12656 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_107
timestamp 1698431365
transform 1 0 13328 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_171
timestamp 1698431365
transform 1 0 20496 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_177
timestamp 1698431365
transform 1 0 21168 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_241
timestamp 1698431365
transform 1 0 28336 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_247
timestamp 1698431365
transform 1 0 29008 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_311
timestamp 1698431365
transform 1 0 36176 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_317
timestamp 1698431365
transform 1 0 36848 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_381
timestamp 1698431365
transform 1 0 44016 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_387
timestamp 1698431365
transform 1 0 44688 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_451
timestamp 1698431365
transform 1 0 51856 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_457
timestamp 1698431365
transform 1 0 52528 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_521
timestamp 1698431365
transform 1 0 59696 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_527
timestamp 1698431365
transform 1 0 60368 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_591
timestamp 1698431365
transform 1 0 67536 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_597
timestamp 1698431365
transform 1 0 68208 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_661
timestamp 1698431365
transform 1 0 75376 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_667
timestamp 1698431365
transform 1 0 76048 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_683
timestamp 1698431365
transform 1 0 77840 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_687
timestamp 1698431365
transform 1 0 78288 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_63_28
timestamp 1698431365
transform 1 0 4480 0 -1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_60
timestamp 1698431365
transform 1 0 8064 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_68
timestamp 1698431365
transform 1 0 8960 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_72
timestamp 1698431365
transform 1 0 9408 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_136
timestamp 1698431365
transform 1 0 16576 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_142
timestamp 1698431365
transform 1 0 17248 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_206
timestamp 1698431365
transform 1 0 24416 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_212
timestamp 1698431365
transform 1 0 25088 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_276
timestamp 1698431365
transform 1 0 32256 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_282
timestamp 1698431365
transform 1 0 32928 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_346
timestamp 1698431365
transform 1 0 40096 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_352
timestamp 1698431365
transform 1 0 40768 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_416
timestamp 1698431365
transform 1 0 47936 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_422
timestamp 1698431365
transform 1 0 48608 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_486
timestamp 1698431365
transform 1 0 55776 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_492
timestamp 1698431365
transform 1 0 56448 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_556
timestamp 1698431365
transform 1 0 63616 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_562
timestamp 1698431365
transform 1 0 64288 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_626
timestamp 1698431365
transform 1 0 71456 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_63_632
timestamp 1698431365
transform 1 0 72128 0 -1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_664
timestamp 1698431365
transform 1 0 75712 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_2
timestamp 1698431365
transform 1 0 1568 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_24
timestamp 1698431365
transform 1 0 4032 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_32
timestamp 1698431365
transform 1 0 4928 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_34
timestamp 1698431365
transform 1 0 5152 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_37
timestamp 1698431365
transform 1 0 5488 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_101
timestamp 1698431365
transform 1 0 12656 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_107
timestamp 1698431365
transform 1 0 13328 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_171
timestamp 1698431365
transform 1 0 20496 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_177
timestamp 1698431365
transform 1 0 21168 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_241
timestamp 1698431365
transform 1 0 28336 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_247
timestamp 1698431365
transform 1 0 29008 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_311
timestamp 1698431365
transform 1 0 36176 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_317
timestamp 1698431365
transform 1 0 36848 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_381
timestamp 1698431365
transform 1 0 44016 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_387
timestamp 1698431365
transform 1 0 44688 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_451
timestamp 1698431365
transform 1 0 51856 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_457
timestamp 1698431365
transform 1 0 52528 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_521
timestamp 1698431365
transform 1 0 59696 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_527
timestamp 1698431365
transform 1 0 60368 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_591
timestamp 1698431365
transform 1 0 67536 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_597
timestamp 1698431365
transform 1 0 68208 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_661
timestamp 1698431365
transform 1 0 75376 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_667
timestamp 1698431365
transform 1 0 76048 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_675
timestamp 1698431365
transform 1 0 76944 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_679
timestamp 1698431365
transform 1 0 77392 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_65_28
timestamp 1698431365
transform 1 0 4480 0 -1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_60
timestamp 1698431365
transform 1 0 8064 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_68
timestamp 1698431365
transform 1 0 8960 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_72
timestamp 1698431365
transform 1 0 9408 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_136
timestamp 1698431365
transform 1 0 16576 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_142
timestamp 1698431365
transform 1 0 17248 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_206
timestamp 1698431365
transform 1 0 24416 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_212
timestamp 1698431365
transform 1 0 25088 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_276
timestamp 1698431365
transform 1 0 32256 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_282
timestamp 1698431365
transform 1 0 32928 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_346
timestamp 1698431365
transform 1 0 40096 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_352
timestamp 1698431365
transform 1 0 40768 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_416
timestamp 1698431365
transform 1 0 47936 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_422
timestamp 1698431365
transform 1 0 48608 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_486
timestamp 1698431365
transform 1 0 55776 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_492
timestamp 1698431365
transform 1 0 56448 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_556
timestamp 1698431365
transform 1 0 63616 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_562
timestamp 1698431365
transform 1 0 64288 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_626
timestamp 1698431365
transform 1 0 71456 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_65_632
timestamp 1698431365
transform 1 0 72128 0 -1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_664
timestamp 1698431365
transform 1 0 75712 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_680
timestamp 1698431365
transform 1 0 77504 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_28
timestamp 1698431365
transform 1 0 4480 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_32
timestamp 1698431365
transform 1 0 4928 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_34
timestamp 1698431365
transform 1 0 5152 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_37
timestamp 1698431365
transform 1 0 5488 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_101
timestamp 1698431365
transform 1 0 12656 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_107
timestamp 1698431365
transform 1 0 13328 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_171
timestamp 1698431365
transform 1 0 20496 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_177
timestamp 1698431365
transform 1 0 21168 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_241
timestamp 1698431365
transform 1 0 28336 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_247
timestamp 1698431365
transform 1 0 29008 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_311
timestamp 1698431365
transform 1 0 36176 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_317
timestamp 1698431365
transform 1 0 36848 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_381
timestamp 1698431365
transform 1 0 44016 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_387
timestamp 1698431365
transform 1 0 44688 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_451
timestamp 1698431365
transform 1 0 51856 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_457
timestamp 1698431365
transform 1 0 52528 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_521
timestamp 1698431365
transform 1 0 59696 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_527
timestamp 1698431365
transform 1 0 60368 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_591
timestamp 1698431365
transform 1 0 67536 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_597
timestamp 1698431365
transform 1 0 68208 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_661
timestamp 1698431365
transform 1 0 75376 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_667
timestamp 1698431365
transform 1 0 76048 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_675
timestamp 1698431365
transform 1 0 76944 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_679
timestamp 1698431365
transform 1 0 77392 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_2
timestamp 1698431365
transform 1 0 1568 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_4
timestamp 1698431365
transform 1 0 1792 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_23
timestamp 1698431365
transform 1 0 3920 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_55
timestamp 1698431365
transform 1 0 7504 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_63
timestamp 1698431365
transform 1 0 8400 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_67
timestamp 1698431365
transform 1 0 8848 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_69
timestamp 1698431365
transform 1 0 9072 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_67_72
timestamp 1698431365
transform 1 0 9408 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_136
timestamp 1698431365
transform 1 0 16576 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_67_142
timestamp 1698431365
transform 1 0 17248 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_206
timestamp 1698431365
transform 1 0 24416 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_67_212
timestamp 1698431365
transform 1 0 25088 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_276
timestamp 1698431365
transform 1 0 32256 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_67_282
timestamp 1698431365
transform 1 0 32928 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_346
timestamp 1698431365
transform 1 0 40096 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_67_352
timestamp 1698431365
transform 1 0 40768 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_416
timestamp 1698431365
transform 1 0 47936 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_67_422
timestamp 1698431365
transform 1 0 48608 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_486
timestamp 1698431365
transform 1 0 55776 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_67_492
timestamp 1698431365
transform 1 0 56448 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_556
timestamp 1698431365
transform 1 0 63616 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_67_562
timestamp 1698431365
transform 1 0 64288 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_626
timestamp 1698431365
transform 1 0 71456 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_632
timestamp 1698431365
transform 1 0 72128 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_664
timestamp 1698431365
transform 1 0 75712 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_672
timestamp 1698431365
transform 1 0 76608 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_676
timestamp 1698431365
transform 1 0 77056 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_34
timestamp 1698431365
transform 1 0 5152 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_68_37
timestamp 1698431365
transform 1 0 5488 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_101
timestamp 1698431365
transform 1 0 12656 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_68_107
timestamp 1698431365
transform 1 0 13328 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_171
timestamp 1698431365
transform 1 0 20496 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_68_177
timestamp 1698431365
transform 1 0 21168 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_241
timestamp 1698431365
transform 1 0 28336 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_68_247
timestamp 1698431365
transform 1 0 29008 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_311
timestamp 1698431365
transform 1 0 36176 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_68_317
timestamp 1698431365
transform 1 0 36848 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_381
timestamp 1698431365
transform 1 0 44016 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_68_387
timestamp 1698431365
transform 1 0 44688 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_451
timestamp 1698431365
transform 1 0 51856 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_68_457
timestamp 1698431365
transform 1 0 52528 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_521
timestamp 1698431365
transform 1 0 59696 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_68_527
timestamp 1698431365
transform 1 0 60368 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_591
timestamp 1698431365
transform 1 0 67536 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_68_597
timestamp 1698431365
transform 1 0 68208 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_661
timestamp 1698431365
transform 1 0 75376 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_68_667
timestamp 1698431365
transform 1 0 76048 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_675
timestamp 1698431365
transform 1 0 76944 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_679
timestamp 1698431365
transform 1 0 77392 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_69_28
timestamp 1698431365
transform 1 0 4480 0 -1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_69_60
timestamp 1698431365
transform 1 0 8064 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_68
timestamp 1698431365
transform 1 0 8960 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_69_72
timestamp 1698431365
transform 1 0 9408 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_136
timestamp 1698431365
transform 1 0 16576 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_69_142
timestamp 1698431365
transform 1 0 17248 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_206
timestamp 1698431365
transform 1 0 24416 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_69_212
timestamp 1698431365
transform 1 0 25088 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_276
timestamp 1698431365
transform 1 0 32256 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_69_282
timestamp 1698431365
transform 1 0 32928 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_346
timestamp 1698431365
transform 1 0 40096 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_69_352
timestamp 1698431365
transform 1 0 40768 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_416
timestamp 1698431365
transform 1 0 47936 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_69_422
timestamp 1698431365
transform 1 0 48608 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_486
timestamp 1698431365
transform 1 0 55776 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_69_492
timestamp 1698431365
transform 1 0 56448 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_556
timestamp 1698431365
transform 1 0 63616 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_69_562
timestamp 1698431365
transform 1 0 64288 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_626
timestamp 1698431365
transform 1 0 71456 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_69_632
timestamp 1698431365
transform 1 0 72128 0 -1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_69_664
timestamp 1698431365
transform 1 0 75712 0 -1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_69_680
timestamp 1698431365
transform 1 0 77504 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_28
timestamp 1698431365
transform 1 0 4480 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_32
timestamp 1698431365
transform 1 0 4928 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_34
timestamp 1698431365
transform 1 0 5152 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_70_37
timestamp 1698431365
transform 1 0 5488 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_101
timestamp 1698431365
transform 1 0 12656 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_70_107
timestamp 1698431365
transform 1 0 13328 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_171
timestamp 1698431365
transform 1 0 20496 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_70_177
timestamp 1698431365
transform 1 0 21168 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_241
timestamp 1698431365
transform 1 0 28336 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_70_247
timestamp 1698431365
transform 1 0 29008 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_311
timestamp 1698431365
transform 1 0 36176 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_70_317
timestamp 1698431365
transform 1 0 36848 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_381
timestamp 1698431365
transform 1 0 44016 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_70_387
timestamp 1698431365
transform 1 0 44688 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_451
timestamp 1698431365
transform 1 0 51856 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_70_457
timestamp 1698431365
transform 1 0 52528 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_521
timestamp 1698431365
transform 1 0 59696 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_70_527
timestamp 1698431365
transform 1 0 60368 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_591
timestamp 1698431365
transform 1 0 67536 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_70_597
timestamp 1698431365
transform 1 0 68208 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_661
timestamp 1698431365
transform 1 0 75376 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_70_667
timestamp 1698431365
transform 1 0 76048 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_675
timestamp 1698431365
transform 1 0 76944 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_679
timestamp 1698431365
transform 1 0 77392 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_2
timestamp 1698431365
transform 1 0 1568 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_4
timestamp 1698431365
transform 1 0 1792 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_17
timestamp 1698431365
transform 1 0 3248 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_71_21
timestamp 1698431365
transform 1 0 3696 0 -1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_71_53
timestamp 1698431365
transform 1 0 7280 0 -1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_69
timestamp 1698431365
transform 1 0 9072 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_71_72
timestamp 1698431365
transform 1 0 9408 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_136
timestamp 1698431365
transform 1 0 16576 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_71_142
timestamp 1698431365
transform 1 0 17248 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_206
timestamp 1698431365
transform 1 0 24416 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_71_212
timestamp 1698431365
transform 1 0 25088 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_276
timestamp 1698431365
transform 1 0 32256 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_71_282
timestamp 1698431365
transform 1 0 32928 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_346
timestamp 1698431365
transform 1 0 40096 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_71_352
timestamp 1698431365
transform 1 0 40768 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_416
timestamp 1698431365
transform 1 0 47936 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_71_422
timestamp 1698431365
transform 1 0 48608 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_486
timestamp 1698431365
transform 1 0 55776 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_71_492
timestamp 1698431365
transform 1 0 56448 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_556
timestamp 1698431365
transform 1 0 63616 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_71_562
timestamp 1698431365
transform 1 0 64288 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_626
timestamp 1698431365
transform 1 0 71456 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_71_632
timestamp 1698431365
transform 1 0 72128 0 -1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_71_664
timestamp 1698431365
transform 1 0 75712 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_672
timestamp 1698431365
transform 1 0 76608 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_676
timestamp 1698431365
transform 1 0 77056 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_28
timestamp 1698431365
transform 1 0 4480 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_32
timestamp 1698431365
transform 1 0 4928 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_34
timestamp 1698431365
transform 1 0 5152 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_72_37
timestamp 1698431365
transform 1 0 5488 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_101
timestamp 1698431365
transform 1 0 12656 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_72_107
timestamp 1698431365
transform 1 0 13328 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_171
timestamp 1698431365
transform 1 0 20496 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_72_177
timestamp 1698431365
transform 1 0 21168 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_241
timestamp 1698431365
transform 1 0 28336 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_72_247
timestamp 1698431365
transform 1 0 29008 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_311
timestamp 1698431365
transform 1 0 36176 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_72_317
timestamp 1698431365
transform 1 0 36848 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_381
timestamp 1698431365
transform 1 0 44016 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_72_387
timestamp 1698431365
transform 1 0 44688 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_451
timestamp 1698431365
transform 1 0 51856 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_72_457
timestamp 1698431365
transform 1 0 52528 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_521
timestamp 1698431365
transform 1 0 59696 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_72_527
timestamp 1698431365
transform 1 0 60368 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_591
timestamp 1698431365
transform 1 0 67536 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_72_597
timestamp 1698431365
transform 1 0 68208 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_661
timestamp 1698431365
transform 1 0 75376 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_72_667
timestamp 1698431365
transform 1 0 76048 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_683
timestamp 1698431365
transform 1 0 77840 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_687
timestamp 1698431365
transform 1 0 78288 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_73_28
timestamp 1698431365
transform 1 0 4480 0 -1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_73_60
timestamp 1698431365
transform 1 0 8064 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_68
timestamp 1698431365
transform 1 0 8960 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_73_72
timestamp 1698431365
transform 1 0 9408 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_136
timestamp 1698431365
transform 1 0 16576 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_73_142
timestamp 1698431365
transform 1 0 17248 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_206
timestamp 1698431365
transform 1 0 24416 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_73_212
timestamp 1698431365
transform 1 0 25088 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_276
timestamp 1698431365
transform 1 0 32256 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_73_282
timestamp 1698431365
transform 1 0 32928 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_346
timestamp 1698431365
transform 1 0 40096 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_73_352
timestamp 1698431365
transform 1 0 40768 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_416
timestamp 1698431365
transform 1 0 47936 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_73_422
timestamp 1698431365
transform 1 0 48608 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_486
timestamp 1698431365
transform 1 0 55776 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_73_492
timestamp 1698431365
transform 1 0 56448 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_556
timestamp 1698431365
transform 1 0 63616 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_73_562
timestamp 1698431365
transform 1 0 64288 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_626
timestamp 1698431365
transform 1 0 71456 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_73_632
timestamp 1698431365
transform 1 0 72128 0 -1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_73_664
timestamp 1698431365
transform 1 0 75712 0 -1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_2
timestamp 1698431365
transform 1 0 1568 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_4
timestamp 1698431365
transform 1 0 1792 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_23
timestamp 1698431365
transform 1 0 3920 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_74_27
timestamp 1698431365
transform 1 0 4368 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_74_37
timestamp 1698431365
transform 1 0 5488 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_101
timestamp 1698431365
transform 1 0 12656 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_74_107
timestamp 1698431365
transform 1 0 13328 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_171
timestamp 1698431365
transform 1 0 20496 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_74_177
timestamp 1698431365
transform 1 0 21168 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_241
timestamp 1698431365
transform 1 0 28336 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_74_247
timestamp 1698431365
transform 1 0 29008 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_311
timestamp 1698431365
transform 1 0 36176 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_74_317
timestamp 1698431365
transform 1 0 36848 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_381
timestamp 1698431365
transform 1 0 44016 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_74_387
timestamp 1698431365
transform 1 0 44688 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_451
timestamp 1698431365
transform 1 0 51856 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_74_457
timestamp 1698431365
transform 1 0 52528 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_521
timestamp 1698431365
transform 1 0 59696 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_74_527
timestamp 1698431365
transform 1 0 60368 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_591
timestamp 1698431365
transform 1 0 67536 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_74_597
timestamp 1698431365
transform 1 0 68208 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_661
timestamp 1698431365
transform 1 0 75376 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_74_667
timestamp 1698431365
transform 1 0 76048 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_675
timestamp 1698431365
transform 1 0 76944 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_679
timestamp 1698431365
transform 1 0 77392 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_75_28
timestamp 1698431365
transform 1 0 4480 0 -1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_75_60
timestamp 1698431365
transform 1 0 8064 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_68
timestamp 1698431365
transform 1 0 8960 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_75_72
timestamp 1698431365
transform 1 0 9408 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_136
timestamp 1698431365
transform 1 0 16576 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_75_142
timestamp 1698431365
transform 1 0 17248 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_206
timestamp 1698431365
transform 1 0 24416 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_75_212
timestamp 1698431365
transform 1 0 25088 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_276
timestamp 1698431365
transform 1 0 32256 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_75_282
timestamp 1698431365
transform 1 0 32928 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_346
timestamp 1698431365
transform 1 0 40096 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_75_352
timestamp 1698431365
transform 1 0 40768 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_416
timestamp 1698431365
transform 1 0 47936 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_75_422
timestamp 1698431365
transform 1 0 48608 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_486
timestamp 1698431365
transform 1 0 55776 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_75_492
timestamp 1698431365
transform 1 0 56448 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_556
timestamp 1698431365
transform 1 0 63616 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_75_562
timestamp 1698431365
transform 1 0 64288 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_626
timestamp 1698431365
transform 1 0 71456 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_75_632
timestamp 1698431365
transform 1 0 72128 0 -1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_75_664
timestamp 1698431365
transform 1 0 75712 0 -1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_75_680
timestamp 1698431365
transform 1 0 77504 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_28
timestamp 1698431365
transform 1 0 4480 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_32
timestamp 1698431365
transform 1 0 4928 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_34
timestamp 1698431365
transform 1 0 5152 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_76_37
timestamp 1698431365
transform 1 0 5488 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_101
timestamp 1698431365
transform 1 0 12656 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_76_107
timestamp 1698431365
transform 1 0 13328 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_171
timestamp 1698431365
transform 1 0 20496 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_76_177
timestamp 1698431365
transform 1 0 21168 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_241
timestamp 1698431365
transform 1 0 28336 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_76_247
timestamp 1698431365
transform 1 0 29008 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_311
timestamp 1698431365
transform 1 0 36176 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_76_317
timestamp 1698431365
transform 1 0 36848 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_381
timestamp 1698431365
transform 1 0 44016 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_76_387
timestamp 1698431365
transform 1 0 44688 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_451
timestamp 1698431365
transform 1 0 51856 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_76_457
timestamp 1698431365
transform 1 0 52528 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_521
timestamp 1698431365
transform 1 0 59696 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_76_527
timestamp 1698431365
transform 1 0 60368 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_591
timestamp 1698431365
transform 1 0 67536 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_76_597
timestamp 1698431365
transform 1 0 68208 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_661
timestamp 1698431365
transform 1 0 75376 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_76_667
timestamp 1698431365
transform 1 0 76048 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_675
timestamp 1698431365
transform 1 0 76944 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_677
timestamp 1698431365
transform 1 0 77168 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_2
timestamp 1698431365
transform 1 0 1568 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_77_24
timestamp 1698431365
transform 1 0 4032 0 -1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_77_56
timestamp 1698431365
transform 1 0 7616 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_64
timestamp 1698431365
transform 1 0 8512 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_68
timestamp 1698431365
transform 1 0 8960 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_77_72
timestamp 1698431365
transform 1 0 9408 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_136
timestamp 1698431365
transform 1 0 16576 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_77_142
timestamp 1698431365
transform 1 0 17248 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_206
timestamp 1698431365
transform 1 0 24416 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_77_212
timestamp 1698431365
transform 1 0 25088 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_276
timestamp 1698431365
transform 1 0 32256 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_77_282
timestamp 1698431365
transform 1 0 32928 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_346
timestamp 1698431365
transform 1 0 40096 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_77_352
timestamp 1698431365
transform 1 0 40768 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_416
timestamp 1698431365
transform 1 0 47936 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_77_422
timestamp 1698431365
transform 1 0 48608 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_486
timestamp 1698431365
transform 1 0 55776 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_77_492
timestamp 1698431365
transform 1 0 56448 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_556
timestamp 1698431365
transform 1 0 63616 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_77_562
timestamp 1698431365
transform 1 0 64288 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_626
timestamp 1698431365
transform 1 0 71456 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_77_632
timestamp 1698431365
transform 1 0 72128 0 -1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_77_664
timestamp 1698431365
transform 1 0 75712 0 -1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_28
timestamp 1698431365
transform 1 0 4480 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_32
timestamp 1698431365
transform 1 0 4928 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_34
timestamp 1698431365
transform 1 0 5152 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_78_37
timestamp 1698431365
transform 1 0 5488 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_101
timestamp 1698431365
transform 1 0 12656 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_78_107
timestamp 1698431365
transform 1 0 13328 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_171
timestamp 1698431365
transform 1 0 20496 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_78_177
timestamp 1698431365
transform 1 0 21168 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_241
timestamp 1698431365
transform 1 0 28336 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_78_247
timestamp 1698431365
transform 1 0 29008 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_311
timestamp 1698431365
transform 1 0 36176 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_78_317
timestamp 1698431365
transform 1 0 36848 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_381
timestamp 1698431365
transform 1 0 44016 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_78_387
timestamp 1698431365
transform 1 0 44688 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_451
timestamp 1698431365
transform 1 0 51856 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_78_457
timestamp 1698431365
transform 1 0 52528 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_521
timestamp 1698431365
transform 1 0 59696 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_78_527
timestamp 1698431365
transform 1 0 60368 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_591
timestamp 1698431365
transform 1 0 67536 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_78_597
timestamp 1698431365
transform 1 0 68208 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_661
timestamp 1698431365
transform 1 0 75376 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_78_667
timestamp 1698431365
transform 1 0 76048 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_675
timestamp 1698431365
transform 1 0 76944 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_677
timestamp 1698431365
transform 1 0 77168 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_79_28
timestamp 1698431365
transform 1 0 4480 0 -1 65856
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_79_60
timestamp 1698431365
transform 1 0 8064 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_68
timestamp 1698431365
transform 1 0 8960 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_79_72
timestamp 1698431365
transform 1 0 9408 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_136
timestamp 1698431365
transform 1 0 16576 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_79_142
timestamp 1698431365
transform 1 0 17248 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_206
timestamp 1698431365
transform 1 0 24416 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_79_212
timestamp 1698431365
transform 1 0 25088 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_276
timestamp 1698431365
transform 1 0 32256 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_79_282
timestamp 1698431365
transform 1 0 32928 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_346
timestamp 1698431365
transform 1 0 40096 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_79_352
timestamp 1698431365
transform 1 0 40768 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_416
timestamp 1698431365
transform 1 0 47936 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_79_422
timestamp 1698431365
transform 1 0 48608 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_486
timestamp 1698431365
transform 1 0 55776 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_79_492
timestamp 1698431365
transform 1 0 56448 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_556
timestamp 1698431365
transform 1 0 63616 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_79_562
timestamp 1698431365
transform 1 0 64288 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_626
timestamp 1698431365
transform 1 0 71456 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_79_632
timestamp 1698431365
transform 1 0 72128 0 -1 65856
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_79_664
timestamp 1698431365
transform 1 0 75712 0 -1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_79_680
timestamp 1698431365
transform 1 0 77504 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_28
timestamp 1698431365
transform 1 0 4480 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_32
timestamp 1698431365
transform 1 0 4928 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_34
timestamp 1698431365
transform 1 0 5152 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_80_37
timestamp 1698431365
transform 1 0 5488 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_101
timestamp 1698431365
transform 1 0 12656 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_80_107
timestamp 1698431365
transform 1 0 13328 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_171
timestamp 1698431365
transform 1 0 20496 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_80_177
timestamp 1698431365
transform 1 0 21168 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_241
timestamp 1698431365
transform 1 0 28336 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_80_247
timestamp 1698431365
transform 1 0 29008 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_311
timestamp 1698431365
transform 1 0 36176 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_80_317
timestamp 1698431365
transform 1 0 36848 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_381
timestamp 1698431365
transform 1 0 44016 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_80_387
timestamp 1698431365
transform 1 0 44688 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_451
timestamp 1698431365
transform 1 0 51856 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_80_457
timestamp 1698431365
transform 1 0 52528 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_521
timestamp 1698431365
transform 1 0 59696 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_80_527
timestamp 1698431365
transform 1 0 60368 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_591
timestamp 1698431365
transform 1 0 67536 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_80_597
timestamp 1698431365
transform 1 0 68208 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_661
timestamp 1698431365
transform 1 0 75376 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_80_667
timestamp 1698431365
transform 1 0 76048 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_675
timestamp 1698431365
transform 1 0 76944 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_677
timestamp 1698431365
transform 1 0 77168 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_2
timestamp 1698431365
transform 1 0 1568 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_4
timestamp 1698431365
transform 1 0 1792 0 -1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_81_29
timestamp 1698431365
transform 1 0 4592 0 -1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_81_61
timestamp 1698431365
transform 1 0 8176 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_69
timestamp 1698431365
transform 1 0 9072 0 -1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_81_72
timestamp 1698431365
transform 1 0 9408 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_136
timestamp 1698431365
transform 1 0 16576 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_81_142
timestamp 1698431365
transform 1 0 17248 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_206
timestamp 1698431365
transform 1 0 24416 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_81_212
timestamp 1698431365
transform 1 0 25088 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_276
timestamp 1698431365
transform 1 0 32256 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_81_282
timestamp 1698431365
transform 1 0 32928 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_346
timestamp 1698431365
transform 1 0 40096 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_81_352
timestamp 1698431365
transform 1 0 40768 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_416
timestamp 1698431365
transform 1 0 47936 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_81_422
timestamp 1698431365
transform 1 0 48608 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_486
timestamp 1698431365
transform 1 0 55776 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_81_492
timestamp 1698431365
transform 1 0 56448 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_556
timestamp 1698431365
transform 1 0 63616 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_81_562
timestamp 1698431365
transform 1 0 64288 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_626
timestamp 1698431365
transform 1 0 71456 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_81_632
timestamp 1698431365
transform 1 0 72128 0 -1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_81_664
timestamp 1698431365
transform 1 0 75712 0 -1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_28
timestamp 1698431365
transform 1 0 4480 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_32
timestamp 1698431365
transform 1 0 4928 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_34
timestamp 1698431365
transform 1 0 5152 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_82_37
timestamp 1698431365
transform 1 0 5488 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_101
timestamp 1698431365
transform 1 0 12656 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_82_107
timestamp 1698431365
transform 1 0 13328 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_171
timestamp 1698431365
transform 1 0 20496 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_82_177
timestamp 1698431365
transform 1 0 21168 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_241
timestamp 1698431365
transform 1 0 28336 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_82_247
timestamp 1698431365
transform 1 0 29008 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_311
timestamp 1698431365
transform 1 0 36176 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_82_317
timestamp 1698431365
transform 1 0 36848 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_381
timestamp 1698431365
transform 1 0 44016 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_82_387
timestamp 1698431365
transform 1 0 44688 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_451
timestamp 1698431365
transform 1 0 51856 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_82_457
timestamp 1698431365
transform 1 0 52528 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_521
timestamp 1698431365
transform 1 0 59696 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_82_527
timestamp 1698431365
transform 1 0 60368 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_591
timestamp 1698431365
transform 1 0 67536 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_82_597
timestamp 1698431365
transform 1 0 68208 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_661
timestamp 1698431365
transform 1 0 75376 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_82_667
timestamp 1698431365
transform 1 0 76048 0 1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_683
timestamp 1698431365
transform 1 0 77840 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_687
timestamp 1698431365
transform 1 0 78288 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_83_28
timestamp 1698431365
transform 1 0 4480 0 -1 68992
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_83_60
timestamp 1698431365
transform 1 0 8064 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_68
timestamp 1698431365
transform 1 0 8960 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_83_72
timestamp 1698431365
transform 1 0 9408 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_136
timestamp 1698431365
transform 1 0 16576 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_83_142
timestamp 1698431365
transform 1 0 17248 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_206
timestamp 1698431365
transform 1 0 24416 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_83_212
timestamp 1698431365
transform 1 0 25088 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_276
timestamp 1698431365
transform 1 0 32256 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_83_282
timestamp 1698431365
transform 1 0 32928 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_346
timestamp 1698431365
transform 1 0 40096 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_83_352
timestamp 1698431365
transform 1 0 40768 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_416
timestamp 1698431365
transform 1 0 47936 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_83_422
timestamp 1698431365
transform 1 0 48608 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_486
timestamp 1698431365
transform 1 0 55776 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_83_492
timestamp 1698431365
transform 1 0 56448 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_556
timestamp 1698431365
transform 1 0 63616 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_83_562
timestamp 1698431365
transform 1 0 64288 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_626
timestamp 1698431365
transform 1 0 71456 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_83_632
timestamp 1698431365
transform 1 0 72128 0 -1 68992
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_83_664
timestamp 1698431365
transform 1 0 75712 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_672
timestamp 1698431365
transform 1 0 76608 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_676
timestamp 1698431365
transform 1 0 77056 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_2
timestamp 1698431365
transform 1 0 1568 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_4
timestamp 1698431365
transform 1 0 1792 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_84_17
timestamp 1698431365
transform 1 0 3248 0 1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_33
timestamp 1698431365
transform 1 0 5040 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_84_37
timestamp 1698431365
transform 1 0 5488 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_101
timestamp 1698431365
transform 1 0 12656 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_84_107
timestamp 1698431365
transform 1 0 13328 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_171
timestamp 1698431365
transform 1 0 20496 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_84_177
timestamp 1698431365
transform 1 0 21168 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_241
timestamp 1698431365
transform 1 0 28336 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_84_247
timestamp 1698431365
transform 1 0 29008 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_311
timestamp 1698431365
transform 1 0 36176 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_84_317
timestamp 1698431365
transform 1 0 36848 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_381
timestamp 1698431365
transform 1 0 44016 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_84_387
timestamp 1698431365
transform 1 0 44688 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_451
timestamp 1698431365
transform 1 0 51856 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_84_457
timestamp 1698431365
transform 1 0 52528 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_521
timestamp 1698431365
transform 1 0 59696 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_84_527
timestamp 1698431365
transform 1 0 60368 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_591
timestamp 1698431365
transform 1 0 67536 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_84_597
timestamp 1698431365
transform 1 0 68208 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_661
timestamp 1698431365
transform 1 0 75376 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_84_667
timestamp 1698431365
transform 1 0 76048 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_675
timestamp 1698431365
transform 1 0 76944 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_679
timestamp 1698431365
transform 1 0 77392 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_85_28
timestamp 1698431365
transform 1 0 4480 0 -1 70560
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_85_60
timestamp 1698431365
transform 1 0 8064 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_68
timestamp 1698431365
transform 1 0 8960 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_85_72
timestamp 1698431365
transform 1 0 9408 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_136
timestamp 1698431365
transform 1 0 16576 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_85_142
timestamp 1698431365
transform 1 0 17248 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_206
timestamp 1698431365
transform 1 0 24416 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_85_212
timestamp 1698431365
transform 1 0 25088 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_276
timestamp 1698431365
transform 1 0 32256 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_85_282
timestamp 1698431365
transform 1 0 32928 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_346
timestamp 1698431365
transform 1 0 40096 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_85_352
timestamp 1698431365
transform 1 0 40768 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_416
timestamp 1698431365
transform 1 0 47936 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_85_422
timestamp 1698431365
transform 1 0 48608 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_486
timestamp 1698431365
transform 1 0 55776 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_85_492
timestamp 1698431365
transform 1 0 56448 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_556
timestamp 1698431365
transform 1 0 63616 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_85_562
timestamp 1698431365
transform 1 0 64288 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_626
timestamp 1698431365
transform 1 0 71456 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_85_632
timestamp 1698431365
transform 1 0 72128 0 -1 70560
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_85_664
timestamp 1698431365
transform 1 0 75712 0 -1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_85_680
timestamp 1698431365
transform 1 0 77504 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_28
timestamp 1698431365
transform 1 0 4480 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_32
timestamp 1698431365
transform 1 0 4928 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_86_34
timestamp 1698431365
transform 1 0 5152 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_86_37
timestamp 1698431365
transform 1 0 5488 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_101
timestamp 1698431365
transform 1 0 12656 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_86_107
timestamp 1698431365
transform 1 0 13328 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_171
timestamp 1698431365
transform 1 0 20496 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_86_177
timestamp 1698431365
transform 1 0 21168 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_241
timestamp 1698431365
transform 1 0 28336 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_86_247
timestamp 1698431365
transform 1 0 29008 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_311
timestamp 1698431365
transform 1 0 36176 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_86_317
timestamp 1698431365
transform 1 0 36848 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_381
timestamp 1698431365
transform 1 0 44016 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_86_387
timestamp 1698431365
transform 1 0 44688 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_451
timestamp 1698431365
transform 1 0 51856 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_86_457
timestamp 1698431365
transform 1 0 52528 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_521
timestamp 1698431365
transform 1 0 59696 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_86_527
timestamp 1698431365
transform 1 0 60368 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_591
timestamp 1698431365
transform 1 0 67536 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_86_597
timestamp 1698431365
transform 1 0 68208 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_661
timestamp 1698431365
transform 1 0 75376 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_86_667
timestamp 1698431365
transform 1 0 76048 0 1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_675
timestamp 1698431365
transform 1 0 76944 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_86_677
timestamp 1698431365
transform 1 0 77168 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_2
timestamp 1698431365
transform 1 0 1568 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_87_24
timestamp 1698431365
transform 1 0 4032 0 -1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_87_56
timestamp 1698431365
transform 1 0 7616 0 -1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_64
timestamp 1698431365
transform 1 0 8512 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_68
timestamp 1698431365
transform 1 0 8960 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_72
timestamp 1698431365
transform 1 0 9408 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_136
timestamp 1698431365
transform 1 0 16576 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_142
timestamp 1698431365
transform 1 0 17248 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_206
timestamp 1698431365
transform 1 0 24416 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_212
timestamp 1698431365
transform 1 0 25088 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_276
timestamp 1698431365
transform 1 0 32256 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_282
timestamp 1698431365
transform 1 0 32928 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_346
timestamp 1698431365
transform 1 0 40096 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_352
timestamp 1698431365
transform 1 0 40768 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_416
timestamp 1698431365
transform 1 0 47936 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_422
timestamp 1698431365
transform 1 0 48608 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_486
timestamp 1698431365
transform 1 0 55776 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_492
timestamp 1698431365
transform 1 0 56448 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_556
timestamp 1698431365
transform 1 0 63616 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_562
timestamp 1698431365
transform 1 0 64288 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_626
timestamp 1698431365
transform 1 0 71456 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_87_632
timestamp 1698431365
transform 1 0 72128 0 -1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_87_664
timestamp 1698431365
transform 1 0 75712 0 -1 72128
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_88_34
timestamp 1698431365
transform 1 0 5152 0 1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_88_37
timestamp 1698431365
transform 1 0 5488 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_101
timestamp 1698431365
transform 1 0 12656 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_107
timestamp 1698431365
transform 1 0 13328 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_111
timestamp 1698431365
transform 1 0 13776 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_88_113
timestamp 1698431365
transform 1 0 14000 0 1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_88_116
timestamp 1698431365
transform 1 0 14336 0 1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_88_148
timestamp 1698431365
transform 1 0 17920 0 1 72128
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_88_164
timestamp 1698431365
transform 1 0 19712 0 1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_172
timestamp 1698431365
transform 1 0 20608 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_88_174
timestamp 1698431365
transform 1 0 20832 0 1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_88_177
timestamp 1698431365
transform 1 0 21168 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_241
timestamp 1698431365
transform 1 0 28336 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_88_247
timestamp 1698431365
transform 1 0 29008 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_311
timestamp 1698431365
transform 1 0 36176 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_88_317
timestamp 1698431365
transform 1 0 36848 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_381
timestamp 1698431365
transform 1 0 44016 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_88_387
timestamp 1698431365
transform 1 0 44688 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_451
timestamp 1698431365
transform 1 0 51856 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_88_457
timestamp 1698431365
transform 1 0 52528 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_521
timestamp 1698431365
transform 1 0 59696 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_88_527
timestamp 1698431365
transform 1 0 60368 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_591
timestamp 1698431365
transform 1 0 67536 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_88_597
timestamp 1698431365
transform 1 0 68208 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_661
timestamp 1698431365
transform 1 0 75376 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_88_667
timestamp 1698431365
transform 1 0 76048 0 1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_88_675
timestamp 1698431365
transform 1 0 76944 0 1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_678
timestamp 1698431365
transform 1 0 77280 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_89_34
timestamp 1698431365
transform 1 0 5152 0 -1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_66
timestamp 1698431365
transform 1 0 8736 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_89_72
timestamp 1698431365
transform 1 0 9408 0 -1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_142
timestamp 1698431365
transform 1 0 17248 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_146
timestamp 1698431365
transform 1 0 17696 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_89_148
timestamp 1698431365
transform 1 0 17920 0 -1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_89_151
timestamp 1698431365
transform 1 0 18256 0 -1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_89_183
timestamp 1698431365
transform 1 0 21840 0 -1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_89_199
timestamp 1698431365
transform 1 0 23632 0 -1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_207
timestamp 1698431365
transform 1 0 24528 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_89_209
timestamp 1698431365
transform 1 0 24752 0 -1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_89_212
timestamp 1698431365
transform 1 0 25088 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_276
timestamp 1698431365
transform 1 0 32256 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_89_282
timestamp 1698431365
transform 1 0 32928 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_346
timestamp 1698431365
transform 1 0 40096 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_89_352
timestamp 1698431365
transform 1 0 40768 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_416
timestamp 1698431365
transform 1 0 47936 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_89_422
timestamp 1698431365
transform 1 0 48608 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_486
timestamp 1698431365
transform 1 0 55776 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_89_492
timestamp 1698431365
transform 1 0 56448 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_556
timestamp 1698431365
transform 1 0 63616 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_89_562
timestamp 1698431365
transform 1 0 64288 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_626
timestamp 1698431365
transform 1 0 71456 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_89_632
timestamp 1698431365
transform 1 0 72128 0 -1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_664
timestamp 1698431365
transform 1 0 75712 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_668
timestamp 1698431365
transform 1 0 76160 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_672
timestamp 1698431365
transform 1 0 76608 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_676
timestamp 1698431365
transform 1 0 77056 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_34
timestamp 1698431365
transform 1 0 5152 0 1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_90_37
timestamp 1698431365
transform 1 0 5488 0 1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_90_69
timestamp 1698431365
transform 1 0 9072 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_77
timestamp 1698431365
transform 1 0 9968 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_107
timestamp 1698431365
transform 1 0 13328 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_111
timestamp 1698431365
transform 1 0 13776 0 1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_114
timestamp 1698431365
transform 1 0 14112 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_118
timestamp 1698431365
transform 1 0 14560 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_122
timestamp 1698431365
transform 1 0 15008 0 1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_90_177
timestamp 1698431365
transform 1 0 21168 0 1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_90_195
timestamp 1698431365
transform 1 0 23184 0 1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_90_227
timestamp 1698431365
transform 1 0 26768 0 1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_243
timestamp 1698431365
transform 1 0 28560 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_90_247
timestamp 1698431365
transform 1 0 29008 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_311
timestamp 1698431365
transform 1 0 36176 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_90_317
timestamp 1698431365
transform 1 0 36848 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_381
timestamp 1698431365
transform 1 0 44016 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_90_387
timestamp 1698431365
transform 1 0 44688 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_451
timestamp 1698431365
transform 1 0 51856 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_90_457
timestamp 1698431365
transform 1 0 52528 0 1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_90_489
timestamp 1698431365
transform 1 0 56112 0 1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_505
timestamp 1698431365
transform 1 0 57904 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_509
timestamp 1698431365
transform 1 0 58352 0 1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_512
timestamp 1698431365
transform 1 0 58688 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_514
timestamp 1698431365
transform 1 0 58912 0 1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_517
timestamp 1698431365
transform 1 0 59248 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_521
timestamp 1698431365
transform 1 0 59696 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_90_527
timestamp 1698431365
transform 1 0 60368 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_591
timestamp 1698431365
transform 1 0 67536 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_90_597
timestamp 1698431365
transform 1 0 68208 0 1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_90_629
timestamp 1698431365
transform 1 0 71792 0 1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_90_645
timestamp 1698431365
transform 1 0 73584 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_653
timestamp 1698431365
transform 1 0 74480 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_657
timestamp 1698431365
transform 1 0 74928 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_661
timestamp 1698431365
transform 1 0 75376 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_667
timestamp 1698431365
transform 1 0 76048 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_671
timestamp 1698431365
transform 1 0 76496 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_673
timestamp 1698431365
transform 1 0 76720 0 1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_682
timestamp 1698431365
transform 1 0 77728 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_686
timestamp 1698431365
transform 1 0 78176 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_91_34
timestamp 1698431365
transform 1 0 5152 0 -1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_66
timestamp 1698431365
transform 1 0 8736 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_91_72
timestamp 1698431365
transform 1 0 9408 0 -1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_142
timestamp 1698431365
transform 1 0 17248 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_146
timestamp 1698431365
transform 1 0 17696 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_149
timestamp 1698431365
transform 1 0 18032 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_91_153
timestamp 1698431365
transform 1 0 18480 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_163
timestamp 1698431365
transform 1 0 19600 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_91_201
timestamp 1698431365
transform 1 0 23856 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_209
timestamp 1698431365
transform 1 0 24752 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_91_212
timestamp 1698431365
transform 1 0 25088 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_276
timestamp 1698431365
transform 1 0 32256 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_91_282
timestamp 1698431365
transform 1 0 32928 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_290
timestamp 1698431365
transform 1 0 33824 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_294
timestamp 1698431365
transform 1 0 34272 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_296
timestamp 1698431365
transform 1 0 34496 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_305
timestamp 1698431365
transform 1 0 35504 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_91_309
timestamp 1698431365
transform 1 0 35952 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_317
timestamp 1698431365
transform 1 0 36848 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_91_323
timestamp 1698431365
transform 1 0 37520 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_331
timestamp 1698431365
transform 1 0 38416 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_91_337
timestamp 1698431365
transform 1 0 39088 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_345
timestamp 1698431365
transform 1 0 39984 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_349
timestamp 1698431365
transform 1 0 40432 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_91_352
timestamp 1698431365
transform 1 0 40768 0 -1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_91_384
timestamp 1698431365
transform 1 0 44352 0 -1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_400
timestamp 1698431365
transform 1 0 46144 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_404
timestamp 1698431365
transform 1 0 46592 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_91_407
timestamp 1698431365
transform 1 0 46928 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_415
timestamp 1698431365
transform 1 0 47824 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_419
timestamp 1698431365
transform 1 0 48272 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_91_422
timestamp 1698431365
transform 1 0 48608 0 -1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_454
timestamp 1698431365
transform 1 0 52192 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_460
timestamp 1698431365
transform 1 0 52864 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_464
timestamp 1698431365
transform 1 0 53312 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_467
timestamp 1698431365
transform 1 0 53648 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_471
timestamp 1698431365
transform 1 0 54096 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_475
timestamp 1698431365
transform 1 0 54544 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_479
timestamp 1698431365
transform 1 0 54992 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_483
timestamp 1698431365
transform 1 0 55440 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_487
timestamp 1698431365
transform 1 0 55888 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_489
timestamp 1698431365
transform 1 0 56112 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_91_492
timestamp 1698431365
transform 1 0 56448 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_500
timestamp 1698431365
transform 1 0 57344 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_529
timestamp 1698431365
transform 1 0 60592 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_533
timestamp 1698431365
transform 1 0 61040 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_537
timestamp 1698431365
transform 1 0 61488 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_541
timestamp 1698431365
transform 1 0 61936 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_91_545
timestamp 1698431365
transform 1 0 62384 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_553
timestamp 1698431365
transform 1 0 63280 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_557
timestamp 1698431365
transform 1 0 63728 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_559
timestamp 1698431365
transform 1 0 63952 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_91_562
timestamp 1698431365
transform 1 0 64288 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_626
timestamp 1698431365
transform 1 0 71456 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_91_632
timestamp 1698431365
transform 1 0 72128 0 -1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_650
timestamp 1698431365
transform 1 0 74144 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_654
timestamp 1698431365
transform 1 0 74592 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_658
timestamp 1698431365
transform 1 0 75040 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_34
timestamp 1698431365
transform 1 0 5152 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_92_37
timestamp 1698431365
transform 1 0 5488 0 1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_92_69
timestamp 1698431365
transform 1 0 9072 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_77
timestamp 1698431365
transform 1 0 9968 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_107
timestamp 1698431365
transform 1 0 13328 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_111
timestamp 1698431365
transform 1 0 13776 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_113
timestamp 1698431365
transform 1 0 14000 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_116
timestamp 1698431365
transform 1 0 14336 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_120
timestamp 1698431365
transform 1 0 14784 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_122
timestamp 1698431365
transform 1 0 15008 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_207
timestamp 1698431365
transform 1 0 24528 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_211
timestamp 1698431365
transform 1 0 24976 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_92_215
timestamp 1698431365
transform 1 0 25424 0 1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_92_231
timestamp 1698431365
transform 1 0 27216 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_239
timestamp 1698431365
transform 1 0 28112 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_243
timestamp 1698431365
transform 1 0 28560 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_92_247
timestamp 1698431365
transform 1 0 29008 0 1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_289
timestamp 1698431365
transform 1 0 33712 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_301
timestamp 1698431365
transform 1 0 35056 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_311
timestamp 1698431365
transform 1 0 36176 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_317
timestamp 1698431365
transform 1 0 36848 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_323
timestamp 1698431365
transform 1 0 37520 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_343
timestamp 1698431365
transform 1 0 39760 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_347
timestamp 1698431365
transform 1 0 40208 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_351
timestamp 1698431365
transform 1 0 40656 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_355
timestamp 1698431365
transform 1 0 41104 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_365
timestamp 1698431365
transform 1 0 42224 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_369
timestamp 1698431365
transform 1 0 42672 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_373
timestamp 1698431365
transform 1 0 43120 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_376
timestamp 1698431365
transform 1 0 43456 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_378
timestamp 1698431365
transform 1 0 43680 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_381
timestamp 1698431365
transform 1 0 44016 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_387
timestamp 1698431365
transform 1 0 44688 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_397
timestamp 1698431365
transform 1 0 45808 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_401
timestamp 1698431365
transform 1 0 46256 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_405
timestamp 1698431365
transform 1 0 46704 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_415
timestamp 1698431365
transform 1 0 47824 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_419
timestamp 1698431365
transform 1 0 48272 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_423
timestamp 1698431365
transform 1 0 48720 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_427
timestamp 1698431365
transform 1 0 49168 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_439
timestamp 1698431365
transform 1 0 50512 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_443
timestamp 1698431365
transform 1 0 50960 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_447
timestamp 1698431365
transform 1 0 51408 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_451
timestamp 1698431365
transform 1 0 51856 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_465
timestamp 1698431365
transform 1 0 53424 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_523
timestamp 1698431365
transform 1 0 59920 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_545
timestamp 1698431365
transform 1 0 62384 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_549
timestamp 1698431365
transform 1 0 62832 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_553
timestamp 1698431365
transform 1 0 63280 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_557
timestamp 1698431365
transform 1 0 63728 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_561
timestamp 1698431365
transform 1 0 64176 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_565
timestamp 1698431365
transform 1 0 64624 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_575
timestamp 1698431365
transform 1 0 65744 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_579
timestamp 1698431365
transform 1 0 66192 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_583
timestamp 1698431365
transform 1 0 66640 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_587
timestamp 1698431365
transform 1 0 67088 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_589
timestamp 1698431365
transform 1 0 67312 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_592
timestamp 1698431365
transform 1 0 67648 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_594
timestamp 1698431365
transform 1 0 67872 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_597
timestamp 1698431365
transform 1 0 68208 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_601
timestamp 1698431365
transform 1 0 68656 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_605
timestamp 1698431365
transform 1 0 69104 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_609
timestamp 1698431365
transform 1 0 69552 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_611
timestamp 1698431365
transform 1 0 69776 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_614
timestamp 1698431365
transform 1 0 70112 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_620
timestamp 1698431365
transform 1 0 70784 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_626
timestamp 1698431365
transform 1 0 71456 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_628
timestamp 1698431365
transform 1 0 71680 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_631
timestamp 1698431365
transform 1 0 72016 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_641
timestamp 1698431365
transform 1 0 73136 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_645
timestamp 1698431365
transform 1 0 73584 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_649
timestamp 1698431365
transform 1 0 74032 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_651
timestamp 1698431365
transform 1 0 74256 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_654
timestamp 1698431365
transform 1 0 74592 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_656
timestamp 1698431365
transform 1 0 74816 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_679
timestamp 1698431365
transform 1 0 77392 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_681
timestamp 1698431365
transform 1 0 77616 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_93_42
timestamp 1698431365
transform 1 0 6048 0 -1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_93_58
timestamp 1698431365
transform 1 0 7840 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_66
timestamp 1698431365
transform 1 0 8736 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_70
timestamp 1698431365
transform 1 0 9184 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_74
timestamp 1698431365
transform 1 0 9632 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_104
timestamp 1698431365
transform 1 0 12992 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_108
timestamp 1698431365
transform 1 0 13440 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_138
timestamp 1698431365
transform 1 0 16800 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_142
timestamp 1698431365
transform 1 0 17248 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_172
timestamp 1698431365
transform 1 0 20608 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_206
timestamp 1698431365
transform 1 0 24416 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_208
timestamp 1698431365
transform 1 0 24640 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_213
timestamp 1698431365
transform 1 0 25200 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_219
timestamp 1698431365
transform 1 0 25872 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_225
timestamp 1698431365
transform 1 0 26544 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_231
timestamp 1698431365
transform 1 0 27216 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_237
timestamp 1698431365
transform 1 0 27888 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_244
timestamp 1698431365
transform 1 0 28672 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_249
timestamp 1698431365
transform 1 0 29232 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_255
timestamp 1698431365
transform 1 0 29904 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_261
timestamp 1698431365
transform 1 0 30576 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_267
timestamp 1698431365
transform 1 0 31248 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_274
timestamp 1698431365
transform 1 0 32032 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_279
timestamp 1698431365
transform 1 0 32592 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_308
timestamp 1698431365
transform 1 0 35840 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_331
timestamp 1698431365
transform 1 0 38416 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_342
timestamp 1698431365
transform 1 0 39648 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_344
timestamp 1698431365
transform 1 0 39872 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_361
timestamp 1698431365
transform 1 0 41776 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_373
timestamp 1698431365
transform 1 0 43120 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_478
timestamp 1698431365
transform 1 0 54880 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_482
timestamp 1698431365
transform 1 0 55328 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_576
timestamp 1698431365
transform 1 0 65856 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_610
timestamp 1698431365
transform 1 0 69664 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_644
timestamp 1698431365
transform 1 0 73472 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1698431365
transform 1 0 24192 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698431365
transform 1 0 29792 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input3
timestamp 1698431365
transform 1 0 31136 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1698431365
transform 1 0 27328 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input5
timestamp 1698431365
transform 1 0 28448 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1698431365
transform 1 0 29120 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1698431365
transform 1 0 29792 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1698431365
transform 1 0 30464 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input9
timestamp 1698431365
transform 1 0 31136 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input10
timestamp 1698431365
transform 1 0 32256 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input11
timestamp 1698431365
transform 1 0 32928 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input12
timestamp 1698431365
transform 1 0 22176 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input13
timestamp 1698431365
transform 1 0 33600 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input14
timestamp 1698431365
transform 1 0 34272 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input15
timestamp 1698431365
transform 1 0 34944 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input16
timestamp 1698431365
transform -1 0 49056 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input17
timestamp 1698431365
transform -1 0 49728 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input18
timestamp 1698431365
transform -1 0 42336 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input19
timestamp 1698431365
transform -1 0 49280 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input20
timestamp 1698431365
transform -1 0 50400 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input21
timestamp 1698431365
transform 1 0 47488 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input22
timestamp 1698431365
transform -1 0 49504 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input23
timestamp 1698431365
transform 1 0 20832 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input24
timestamp 1698431365
transform -1 0 49280 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input25
timestamp 1698431365
transform -1 0 50176 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input26
timestamp 1698431365
transform 1 0 22848 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input27
timestamp 1698431365
transform 1 0 22176 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input28
timestamp 1698431365
transform 1 0 23520 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input29
timestamp 1698431365
transform 1 0 30576 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input30
timestamp 1698431365
transform 1 0 25312 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input31
timestamp 1698431365
transform 1 0 25984 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input32
timestamp 1698431365
transform 1 0 26656 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input33
timestamp 1698431365
transform -1 0 50848 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input34
timestamp 1698431365
transform 1 0 3808 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input35
timestamp 1698431365
transform 1 0 7168 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input36
timestamp 1698431365
transform 1 0 6944 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input37
timestamp 1698431365
transform 1 0 7616 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input38
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input39
timestamp 1698431365
transform 1 0 8512 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input40
timestamp 1698431365
transform 1 0 8288 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input41
timestamp 1698431365
transform 1 0 9408 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input42
timestamp 1698431365
transform 1 0 10080 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input43
timestamp 1698431365
transform 1 0 11424 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input44
timestamp 1698431365
transform 1 0 12096 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input45
timestamp 1698431365
transform 1 0 3136 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input46
timestamp 1698431365
transform 1 0 13216 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input47
timestamp 1698431365
transform 1 0 13888 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input48
timestamp 1698431365
transform 1 0 14560 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input49
timestamp 1698431365
transform 1 0 18144 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input50
timestamp 1698431365
transform 1 0 15904 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input51
timestamp 1698431365
transform 1 0 17696 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input52
timestamp 1698431365
transform 1 0 18368 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input53
timestamp 1698431365
transform 1 0 19040 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input54
timestamp 1698431365
transform 1 0 22176 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input55
timestamp 1698431365
transform 1 0 23520 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input56
timestamp 1698431365
transform 1 0 4480 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input57
timestamp 1698431365
transform 1 0 24192 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input58
timestamp 1698431365
transform 1 0 19712 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input59
timestamp 1698431365
transform 1 0 5152 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input60
timestamp 1698431365
transform 1 0 3808 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input61
timestamp 1698431365
transform -1 0 8512 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input62
timestamp 1698431365
transform 1 0 6272 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input63
timestamp 1698431365
transform 1 0 4480 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input64
timestamp 1698431365
transform 1 0 5600 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input65
timestamp 1698431365
transform 1 0 6272 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input66
timestamp 1698431365
transform 1 0 51072 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input67
timestamp 1698431365
transform -1 0 52640 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input68
timestamp 1698431365
transform -1 0 53312 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input69
timestamp 1698431365
transform -1 0 53984 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input70
timestamp 1698431365
transform 1 0 2240 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input71
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input72
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input73
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input74
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input75
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input76
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input77
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input78
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input79
timestamp 1698431365
transform 1 0 1568 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input80
timestamp 1698431365
transform 1 0 1568 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input81
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input82
timestamp 1698431365
transform 1 0 1568 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input83
timestamp 1698431365
transform 1 0 1568 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input84
timestamp 1698431365
transform 1 0 1568 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input85
timestamp 1698431365
transform 1 0 1568 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input86
timestamp 1698431365
transform 1 0 1568 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input87
timestamp 1698431365
transform 1 0 1568 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input88
timestamp 1698431365
transform 1 0 1568 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input89
timestamp 1698431365
transform 1 0 1568 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input90
timestamp 1698431365
transform 1 0 1568 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input91
timestamp 1698431365
transform 1 0 1568 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input92
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input93
timestamp 1698431365
transform 1 0 1568 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input94
timestamp 1698431365
transform 1 0 1568 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input95
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input96
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input97
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input98
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input99
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input100
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input101
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input102
timestamp 1698431365
transform 1 0 74928 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input103
timestamp 1698431365
transform -1 0 78400 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input104
timestamp 1698431365
transform -1 0 78400 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input105
timestamp 1698431365
transform -1 0 78400 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input106
timestamp 1698431365
transform -1 0 78400 0 1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input107
timestamp 1698431365
transform -1 0 78400 0 1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input108
timestamp 1698431365
transform -1 0 78400 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input109
timestamp 1698431365
transform -1 0 78400 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input110
timestamp 1698431365
transform -1 0 78400 0 1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input111
timestamp 1698431365
transform -1 0 78400 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input112
timestamp 1698431365
transform -1 0 78400 0 -1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input113
timestamp 1698431365
transform -1 0 78400 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input114
timestamp 1698431365
transform -1 0 78400 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input115
timestamp 1698431365
transform -1 0 78400 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input116
timestamp 1698431365
transform -1 0 78400 0 -1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input117
timestamp 1698431365
transform -1 0 78400 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input118
timestamp 1698431365
transform -1 0 78400 0 1 68992
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input119
timestamp 1698431365
transform -1 0 78400 0 1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input120
timestamp 1698431365
transform -1 0 78400 0 -1 72128
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input121
timestamp 1698431365
transform -1 0 78400 0 1 72128
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input122
timestamp 1698431365
transform -1 0 78400 0 -1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input123
timestamp 1698431365
transform -1 0 78400 0 -1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input124
timestamp 1698431365
transform -1 0 78400 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input125
timestamp 1698431365
transform -1 0 78400 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input126
timestamp 1698431365
transform -1 0 77056 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input127
timestamp 1698431365
transform -1 0 77728 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input128
timestamp 1698431365
transform -1 0 78400 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input129
timestamp 1698431365
transform -1 0 78400 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input130
timestamp 1698431365
transform -1 0 78400 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input131
timestamp 1698431365
transform -1 0 78400 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input132
timestamp 1698431365
transform -1 0 78400 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input133
timestamp 1698431365
transform -1 0 78400 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input134
timestamp 1698431365
transform -1 0 78400 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input135
timestamp 1698431365
transform -1 0 77504 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input136
timestamp 1698431365
transform -1 0 78400 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input137
timestamp 1698431365
transform -1 0 78400 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input138
timestamp 1698431365
transform -1 0 77728 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input139
timestamp 1698431365
transform -1 0 78400 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input140
timestamp 1698431365
transform 1 0 74592 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input141
timestamp 1698431365
transform -1 0 77728 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input142
timestamp 1698431365
transform -1 0 78400 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input143
timestamp 1698431365
transform -1 0 78400 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input144
timestamp 1698431365
transform 1 0 76048 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input145
timestamp 1698431365
transform 1 0 75152 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input146
timestamp 1698431365
transform 1 0 74480 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input147
timestamp 1698431365
transform -1 0 77056 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input148
timestamp 1698431365
transform -1 0 78400 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input149
timestamp 1698431365
transform 1 0 73584 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input150
timestamp 1698431365
transform 1 0 75376 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input151
timestamp 1698431365
transform 1 0 75152 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input152
timestamp 1698431365
transform 1 0 73808 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input153
timestamp 1698431365
transform -1 0 78400 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input154
timestamp 1698431365
transform 1 0 74480 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input155
timestamp 1698431365
transform -1 0 78400 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input156
timestamp 1698431365
transform 1 0 74032 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input157
timestamp 1698431365
transform 1 0 75152 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input158
timestamp 1698431365
transform -1 0 77728 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input159
timestamp 1698431365
transform 1 0 77728 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input160
timestamp 1698431365
transform -1 0 76832 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input161
timestamp 1698431365
transform -1 0 78400 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input162
timestamp 1698431365
transform -1 0 78400 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input163
timestamp 1698431365
transform -1 0 78400 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input164
timestamp 1698431365
transform -1 0 78400 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input165
timestamp 1698431365
transform -1 0 78400 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input166
timestamp 1698431365
transform -1 0 78400 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input167
timestamp 1698431365
transform -1 0 78400 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input168
timestamp 1698431365
transform 1 0 34160 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input169
timestamp 1698431365
transform 1 0 40880 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input170
timestamp 1698431365
transform 1 0 41552 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input171
timestamp 1698431365
transform 1 0 42224 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input172
timestamp 1698431365
transform 1 0 43456 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input173
timestamp 1698431365
transform 1 0 44352 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input174
timestamp 1698431365
transform 1 0 45248 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input175
timestamp 1698431365
transform 1 0 44912 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input176
timestamp 1698431365
transform 1 0 46144 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input177
timestamp 1698431365
transform 1 0 47264 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input178
timestamp 1698431365
transform 1 0 46928 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input179
timestamp 1698431365
transform -1 0 35504 0 -1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input180
timestamp 1698431365
transform 1 0 48160 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input181
timestamp 1698431365
transform 1 0 49056 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input182
timestamp 1698431365
transform 1 0 49952 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input183
timestamp 1698431365
transform 1 0 49616 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input184
timestamp 1698431365
transform 1 0 51072 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input185
timestamp 1698431365
transform 1 0 51968 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input186
timestamp 1698431365
transform 1 0 52864 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input187
timestamp 1698431365
transform 1 0 52528 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input188
timestamp 1698431365
transform 1 0 53760 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input189
timestamp 1698431365
transform 1 0 53648 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input190
timestamp 1698431365
transform 1 0 35504 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input191
timestamp 1698431365
transform 1 0 54544 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input192
timestamp 1698431365
transform 1 0 55440 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input193
timestamp 1698431365
transform -1 0 36624 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input194
timestamp 1698431365
transform 1 0 36624 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input195
timestamp 1698431365
transform 1 0 37520 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input196
timestamp 1698431365
transform 1 0 37968 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input197
timestamp 1698431365
transform 1 0 38864 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input198
timestamp 1698431365
transform -1 0 39424 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input199
timestamp 1698431365
transform 1 0 39984 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input200
timestamp 1698431365
transform 1 0 32816 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input201
timestamp 1698431365
transform 1 0 59248 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input202
timestamp 1698431365
transform 1 0 65072 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input203
timestamp 1698431365
transform 1 0 66304 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input204
timestamp 1698431365
transform 1 0 66976 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input205
timestamp 1698431365
transform 1 0 67648 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input206
timestamp 1698431365
transform 1 0 68320 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input207
timestamp 1698431365
transform 1 0 68992 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input208
timestamp 1698431365
transform 1 0 70112 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input209
timestamp 1698431365
transform 1 0 70784 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input210
timestamp 1698431365
transform -1 0 72128 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input211
timestamp 1698431365
transform -1 0 72800 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input212
timestamp 1698431365
transform 1 0 60368 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input213
timestamp 1698431365
transform -1 0 73472 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input214
timestamp 1698431365
transform 1 0 72464 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input215
timestamp 1698431365
transform 1 0 73920 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input216
timestamp 1698431365
transform -1 0 75264 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input217
timestamp 1698431365
transform -1 0 75936 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input218
timestamp 1698431365
transform -1 0 76608 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input219
timestamp 1698431365
transform 1 0 76048 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input220
timestamp 1698431365
transform 1 0 76720 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input221
timestamp 1698431365
transform 1 0 77728 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input222
timestamp 1698431365
transform 1 0 77056 0 -1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input223
timestamp 1698431365
transform -1 0 62272 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input224
timestamp 1698431365
transform 1 0 75152 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input225
timestamp 1698431365
transform -1 0 76160 0 -1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input226
timestamp 1698431365
transform 1 0 61040 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input227
timestamp 1698431365
transform 1 0 61712 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input228
timestamp 1698431365
transform 1 0 62496 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input229
timestamp 1698431365
transform 1 0 63168 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input230
timestamp 1698431365
transform 1 0 63840 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input231
timestamp 1698431365
transform 1 0 64512 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input232
timestamp 1698431365
transform 1 0 65184 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output233 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 13104 0 1 73696
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output234
timestamp 1698431365
transform 1 0 18032 0 1 73696
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output235
timestamp 1698431365
transform -1 0 20944 0 1 75264
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output236
timestamp 1698431365
transform -1 0 20384 0 -1 76832
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output237
timestamp 1698431365
transform -1 0 22960 0 -1 75264
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output238
timestamp 1698431365
transform -1 0 24080 0 1 75264
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output239
timestamp 1698431365
transform -1 0 24192 0 -1 76832
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output240
timestamp 1698431365
transform -1 0 14112 0 -1 73696
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output241
timestamp 1698431365
transform -1 0 13104 0 1 75264
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output242
timestamp 1698431365
transform -1 0 14112 0 -1 75264
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output243
timestamp 1698431365
transform -1 0 12768 0 -1 76832
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output244
timestamp 1698431365
transform -1 0 17024 0 -1 73696
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output245
timestamp 1698431365
transform 1 0 14112 0 -1 75264
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output246
timestamp 1698431365
transform -1 0 18032 0 1 73696
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output247
timestamp 1698431365
transform -1 0 16576 0 -1 76832
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output248
timestamp 1698431365
transform -1 0 18032 0 1 75264
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output249
timestamp 1698431365
transform 1 0 52752 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output250
timestamp 1698431365
transform 1 0 59696 0 -1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output251
timestamp 1698431365
transform 1 0 60368 0 1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output252
timestamp 1698431365
transform 1 0 63280 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output253
timestamp 1698431365
transform 1 0 64288 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output254
timestamp 1698431365
transform 1 0 66304 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output255
timestamp 1698431365
transform 1 0 63280 0 1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output256
timestamp 1698431365
transform 1 0 64288 0 -1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output257
timestamp 1698431365
transform 1 0 67200 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output258
timestamp 1698431365
transform 1 0 70112 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output259
timestamp 1698431365
transform 1 0 67200 0 -1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output260
timestamp 1698431365
transform 1 0 54880 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output261
timestamp 1698431365
transform 1 0 68208 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output262
timestamp 1698431365
transform 1 0 66864 0 -1 7840
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output263
timestamp 1698431365
transform 1 0 68208 0 1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output264
timestamp 1698431365
transform 1 0 71120 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output265
timestamp 1698431365
transform 1 0 72128 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output266
timestamp 1698431365
transform 1 0 73920 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output267
timestamp 1698431365
transform 1 0 71120 0 1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output268
timestamp 1698431365
transform 1 0 72128 0 -1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output269
timestamp 1698431365
transform 1 0 75040 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output270
timestamp 1698431365
transform 1 0 72240 0 -1 7840
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output271
timestamp 1698431365
transform 1 0 54096 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output272
timestamp 1698431365
transform -1 0 77952 0 -1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output273
timestamp 1698431365
transform 1 0 75152 0 -1 7840
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output274
timestamp 1698431365
transform 1 0 56448 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output275
timestamp 1698431365
transform -1 0 61600 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output276
timestamp 1698431365
transform 1 0 57008 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output277
timestamp 1698431365
transform 1 0 56784 0 -1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output278
timestamp 1698431365
transform -1 0 62272 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output279
timestamp 1698431365
transform 1 0 62496 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output280
timestamp 1698431365
transform 1 0 60368 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output281
timestamp 1698431365
transform 1 0 49392 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output282
timestamp 1698431365
transform 1 0 1568 0 -1 39200
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output283
timestamp 1698431365
transform -1 0 4480 0 1 39200
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output284
timestamp 1698431365
transform -1 0 4480 0 1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output285
timestamp 1698431365
transform -1 0 4480 0 -1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output286
timestamp 1698431365
transform -1 0 4480 0 1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output287
timestamp 1698431365
transform -1 0 4480 0 -1 54880
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output288
timestamp 1698431365
transform 1 0 1568 0 1 54880
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output289
timestamp 1698431365
transform -1 0 4480 0 1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output290
timestamp 1698431365
transform -1 0 4480 0 -1 58016
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output291
timestamp 1698431365
transform 1 0 1568 0 1 58016
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output292
timestamp 1698431365
transform -1 0 4480 0 1 59584
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output293
timestamp 1698431365
transform 1 0 1568 0 -1 61152
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output294
timestamp 1698431365
transform -1 0 4480 0 -1 62720
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output295
timestamp 1698431365
transform -1 0 4480 0 1 62720
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output296
timestamp 1698431365
transform -1 0 4480 0 1 64288
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output297
timestamp 1698431365
transform 1 0 1568 0 1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output298
timestamp 1698431365
transform 1 0 1568 0 -1 65856
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output299
timestamp 1698431365
transform -1 0 4480 0 1 65856
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output300
timestamp 1698431365
transform -1 0 4480 0 1 67424
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output301
timestamp 1698431365
transform 1 0 1568 0 -1 68992
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output302
timestamp 1698431365
transform -1 0 4480 0 -1 70560
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output303
timestamp 1698431365
transform -1 0 4480 0 1 70560
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output304
timestamp 1698431365
transform -1 0 4480 0 1 72128
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output305
timestamp 1698431365
transform -1 0 4480 0 -1 73696
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output306
timestamp 1698431365
transform -1 0 4480 0 1 73696
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output307
timestamp 1698431365
transform -1 0 4480 0 1 75264
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output308
timestamp 1698431365
transform 1 0 1568 0 -1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output309
timestamp 1698431365
transform -1 0 4480 0 -1 76832
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output310
timestamp 1698431365
transform -1 0 4480 0 -1 75264
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output311
timestamp 1698431365
transform -1 0 4480 0 -1 47040
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output312
timestamp 1698431365
transform 1 0 1568 0 1 47040
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output313
timestamp 1698431365
transform -1 0 4480 0 1 48608
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output314
timestamp 1698431365
transform -1 0 4480 0 -1 50176
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output315
timestamp 1698431365
transform -1 0 4480 0 1 50176
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output316
timestamp 1698431365
transform -1 0 4480 0 1 51744
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output317
timestamp 1698431365
transform -1 0 4480 0 -1 53312
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output318
timestamp 1698431365
transform 1 0 75488 0 -1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output319
timestamp 1698431365
transform -1 0 78400 0 -1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output320
timestamp 1698431365
transform -1 0 75824 0 1 7840
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output321
timestamp 1698431365
transform -1 0 78400 0 -1 10976
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output322
timestamp 1698431365
transform -1 0 75488 0 -1 9408
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output323
timestamp 1698431365
transform 1 0 75488 0 -1 9408
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output324
timestamp 1698431365
transform -1 0 35616 0 -1 76832
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output325
timestamp 1698431365
transform -1 0 58464 0 -1 76832
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output326
timestamp 1698431365
transform -1 0 59248 0 1 75264
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output327
timestamp 1698431365
transform 1 0 58688 0 -1 76832
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output328
timestamp 1698431365
transform -1 0 60592 0 -1 75264
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_94 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 78624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_95
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 78624 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_96
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 78624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_97
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 78624 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_98
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 78624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_99
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 78624 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_100
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 78624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_101
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 78624 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_102
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 78624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_103
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 78624 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_104
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 78624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_105
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 78624 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_106
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 78624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_107
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 78624 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_108
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 78624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_109
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 78624 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_110
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 78624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_111
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 78624 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_112
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 78624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_113
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 78624 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_114
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 78624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_115
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 78624 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_116
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 78624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_117
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 78624 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_118
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 78624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_119
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 78624 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_120
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 78624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_121
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 78624 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_122
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 78624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_123
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 78624 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_124
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 78624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_125
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 78624 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_126
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 78624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_127
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 78624 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_128
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 78624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_129
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 78624 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_130
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 78624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_131
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 78624 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_132
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 78624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_133
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 78624 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_134
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 78624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_135
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 78624 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_136
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 78624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_137
timestamp 1698431365
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698431365
transform -1 0 78624 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_138
timestamp 1698431365
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698431365
transform -1 0 78624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_139
timestamp 1698431365
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698431365
transform -1 0 78624 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_140
timestamp 1698431365
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698431365
transform -1 0 78624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_141
timestamp 1698431365
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698431365
transform -1 0 78624 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_142
timestamp 1698431365
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698431365
transform -1 0 78624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_143
timestamp 1698431365
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698431365
transform -1 0 78624 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Left_144
timestamp 1698431365
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1698431365
transform -1 0 78624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Left_145
timestamp 1698431365
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1698431365
transform -1 0 78624 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Left_146
timestamp 1698431365
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Right_52
timestamp 1698431365
transform -1 0 78624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Left_147
timestamp 1698431365
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Right_53
timestamp 1698431365
transform -1 0 78624 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Left_148
timestamp 1698431365
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Right_54
timestamp 1698431365
transform -1 0 78624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Left_149
timestamp 1698431365
transform 1 0 1344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Right_55
timestamp 1698431365
transform -1 0 78624 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Left_150
timestamp 1698431365
transform 1 0 1344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Right_56
timestamp 1698431365
transform -1 0 78624 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Left_151
timestamp 1698431365
transform 1 0 1344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Right_57
timestamp 1698431365
transform -1 0 78624 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Left_152
timestamp 1698431365
transform 1 0 1344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Right_58
timestamp 1698431365
transform -1 0 78624 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Left_153
timestamp 1698431365
transform 1 0 1344 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Right_59
timestamp 1698431365
transform -1 0 78624 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Left_154
timestamp 1698431365
transform 1 0 1344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Right_60
timestamp 1698431365
transform -1 0 78624 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Left_155
timestamp 1698431365
transform 1 0 1344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Right_61
timestamp 1698431365
transform -1 0 78624 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Left_156
timestamp 1698431365
transform 1 0 1344 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Right_62
timestamp 1698431365
transform -1 0 78624 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Left_157
timestamp 1698431365
transform 1 0 1344 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Right_63
timestamp 1698431365
transform -1 0 78624 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Left_158
timestamp 1698431365
transform 1 0 1344 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Right_64
timestamp 1698431365
transform -1 0 78624 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Left_159
timestamp 1698431365
transform 1 0 1344 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Right_65
timestamp 1698431365
transform -1 0 78624 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Left_160
timestamp 1698431365
transform 1 0 1344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Right_66
timestamp 1698431365
transform -1 0 78624 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Left_161
timestamp 1698431365
transform 1 0 1344 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Right_67
timestamp 1698431365
transform -1 0 78624 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_68_Left_162
timestamp 1698431365
transform 1 0 1344 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_68_Right_68
timestamp 1698431365
transform -1 0 78624 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_69_Left_163
timestamp 1698431365
transform 1 0 1344 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_69_Right_69
timestamp 1698431365
transform -1 0 78624 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_70_Left_164
timestamp 1698431365
transform 1 0 1344 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_70_Right_70
timestamp 1698431365
transform -1 0 78624 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_71_Left_165
timestamp 1698431365
transform 1 0 1344 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_71_Right_71
timestamp 1698431365
transform -1 0 78624 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_72_Left_166
timestamp 1698431365
transform 1 0 1344 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_72_Right_72
timestamp 1698431365
transform -1 0 78624 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_73_Left_167
timestamp 1698431365
transform 1 0 1344 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_73_Right_73
timestamp 1698431365
transform -1 0 78624 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_74_Left_168
timestamp 1698431365
transform 1 0 1344 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_74_Right_74
timestamp 1698431365
transform -1 0 78624 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_75_Left_169
timestamp 1698431365
transform 1 0 1344 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_75_Right_75
timestamp 1698431365
transform -1 0 78624 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_76_Left_170
timestamp 1698431365
transform 1 0 1344 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_76_Right_76
timestamp 1698431365
transform -1 0 78624 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_77_Left_171
timestamp 1698431365
transform 1 0 1344 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_77_Right_77
timestamp 1698431365
transform -1 0 78624 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_78_Left_172
timestamp 1698431365
transform 1 0 1344 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_78_Right_78
timestamp 1698431365
transform -1 0 78624 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_79_Left_173
timestamp 1698431365
transform 1 0 1344 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_79_Right_79
timestamp 1698431365
transform -1 0 78624 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_80_Left_174
timestamp 1698431365
transform 1 0 1344 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_80_Right_80
timestamp 1698431365
transform -1 0 78624 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_81_Left_175
timestamp 1698431365
transform 1 0 1344 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_81_Right_81
timestamp 1698431365
transform -1 0 78624 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_82_Left_176
timestamp 1698431365
transform 1 0 1344 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_82_Right_82
timestamp 1698431365
transform -1 0 78624 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_83_Left_177
timestamp 1698431365
transform 1 0 1344 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_83_Right_83
timestamp 1698431365
transform -1 0 78624 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_84_Left_178
timestamp 1698431365
transform 1 0 1344 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_84_Right_84
timestamp 1698431365
transform -1 0 78624 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_85_Left_179
timestamp 1698431365
transform 1 0 1344 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_85_Right_85
timestamp 1698431365
transform -1 0 78624 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_86_Left_180
timestamp 1698431365
transform 1 0 1344 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_86_Right_86
timestamp 1698431365
transform -1 0 78624 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_87_Left_181
timestamp 1698431365
transform 1 0 1344 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_87_Right_87
timestamp 1698431365
transform -1 0 78624 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_88_Left_182
timestamp 1698431365
transform 1 0 1344 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_88_Right_88
timestamp 1698431365
transform -1 0 78624 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_89_Left_183
timestamp 1698431365
transform 1 0 1344 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_89_Right_89
timestamp 1698431365
transform -1 0 78624 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_90_Left_184
timestamp 1698431365
transform 1 0 1344 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_90_Right_90
timestamp 1698431365
transform -1 0 78624 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_91_Left_185
timestamp 1698431365
transform 1 0 1344 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_91_Right_91
timestamp 1698431365
transform -1 0 78624 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_92_Left_186
timestamp 1698431365
transform 1 0 1344 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_92_Right_92
timestamp 1698431365
transform -1 0 78624 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_93_Left_187
timestamp 1698431365
transform 1 0 1344 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_93_Right_93
timestamp 1698431365
transform -1 0 78624 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  simple_interconnect_343 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 20832 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  simple_interconnect_344
timestamp 1698431365
transform -1 0 23408 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  simple_interconnect_345
timestamp 1698431365
transform -1 0 23856 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  simple_interconnect_346
timestamp 1698431365
transform -1 0 24528 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  simple_interconnect_347
timestamp 1698431365
transform -1 0 25200 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  simple_interconnect_348
timestamp 1698431365
transform -1 0 25872 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  simple_interconnect_349
timestamp 1698431365
transform -1 0 26544 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  simple_interconnect_350
timestamp 1698431365
transform -1 0 27216 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  simple_interconnect_351
timestamp 1698431365
transform -1 0 27888 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  simple_interconnect_352
timestamp 1698431365
transform -1 0 28672 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  simple_interconnect_353
timestamp 1698431365
transform -1 0 29232 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  simple_interconnect_354
timestamp 1698431365
transform -1 0 29904 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  simple_interconnect_355
timestamp 1698431365
transform -1 0 30576 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  simple_interconnect_356
timestamp 1698431365
transform -1 0 31248 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  simple_interconnect_357
timestamp 1698431365
transform -1 0 31808 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  simple_interconnect_358
timestamp 1698431365
transform -1 0 32592 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_188 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_189
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_190
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_191
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_192
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_193
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_194
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_195
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_196
timestamp 1698431365
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_197
timestamp 1698431365
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_198
timestamp 1698431365
transform 1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_199
timestamp 1698431365
transform 1 0 47040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_200
timestamp 1698431365
transform 1 0 50848 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_201
timestamp 1698431365
transform 1 0 54656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_202
timestamp 1698431365
transform 1 0 58464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_203
timestamp 1698431365
transform 1 0 62272 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_204
timestamp 1698431365
transform 1 0 66080 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_205
timestamp 1698431365
transform 1 0 69888 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_206
timestamp 1698431365
transform 1 0 73696 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_207
timestamp 1698431365
transform 1 0 77504 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_208
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_209
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_210
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_211
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_212
timestamp 1698431365
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_213
timestamp 1698431365
transform 1 0 48384 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_214
timestamp 1698431365
transform 1 0 56224 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_215
timestamp 1698431365
transform 1 0 64064 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_216
timestamp 1698431365
transform 1 0 71904 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_217
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_218
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_219
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_220
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_221
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_222
timestamp 1698431365
transform 1 0 44464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_223
timestamp 1698431365
transform 1 0 52304 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_224
timestamp 1698431365
transform 1 0 60144 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_225
timestamp 1698431365
transform 1 0 67984 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_226
timestamp 1698431365
transform 1 0 75824 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_227
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_228
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_229
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_230
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_231
timestamp 1698431365
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_232
timestamp 1698431365
transform 1 0 48384 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_233
timestamp 1698431365
transform 1 0 56224 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_234
timestamp 1698431365
transform 1 0 64064 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_235
timestamp 1698431365
transform 1 0 71904 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_236
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_237
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_238
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_239
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_240
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_241
timestamp 1698431365
transform 1 0 44464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_242
timestamp 1698431365
transform 1 0 52304 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_243
timestamp 1698431365
transform 1 0 60144 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_244
timestamp 1698431365
transform 1 0 67984 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_245
timestamp 1698431365
transform 1 0 75824 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_246
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_247
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_248
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_249
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_250
timestamp 1698431365
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_251
timestamp 1698431365
transform 1 0 48384 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_252
timestamp 1698431365
transform 1 0 56224 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_253
timestamp 1698431365
transform 1 0 64064 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_254
timestamp 1698431365
transform 1 0 71904 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_255
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_256
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_257
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_258
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_259
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_260
timestamp 1698431365
transform 1 0 44464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_261
timestamp 1698431365
transform 1 0 52304 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_262
timestamp 1698431365
transform 1 0 60144 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_263
timestamp 1698431365
transform 1 0 67984 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_264
timestamp 1698431365
transform 1 0 75824 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_265
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_266
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_267
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_268
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_269
timestamp 1698431365
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_270
timestamp 1698431365
transform 1 0 48384 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_271
timestamp 1698431365
transform 1 0 56224 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_272
timestamp 1698431365
transform 1 0 64064 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_273
timestamp 1698431365
transform 1 0 71904 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_274
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_275
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_276
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_277
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_278
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_279
timestamp 1698431365
transform 1 0 44464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_280
timestamp 1698431365
transform 1 0 52304 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_281
timestamp 1698431365
transform 1 0 60144 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_282
timestamp 1698431365
transform 1 0 67984 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_283
timestamp 1698431365
transform 1 0 75824 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_284
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_285
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_286
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_287
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_288
timestamp 1698431365
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_289
timestamp 1698431365
transform 1 0 48384 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_290
timestamp 1698431365
transform 1 0 56224 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_291
timestamp 1698431365
transform 1 0 64064 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_292
timestamp 1698431365
transform 1 0 71904 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_293
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_294
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_295
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_296
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_297
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_298
timestamp 1698431365
transform 1 0 44464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_299
timestamp 1698431365
transform 1 0 52304 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_300
timestamp 1698431365
transform 1 0 60144 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_301
timestamp 1698431365
transform 1 0 67984 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_302
timestamp 1698431365
transform 1 0 75824 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_303
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_304
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_305
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_306
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_307
timestamp 1698431365
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_308
timestamp 1698431365
transform 1 0 48384 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_309
timestamp 1698431365
transform 1 0 56224 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_310
timestamp 1698431365
transform 1 0 64064 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_311
timestamp 1698431365
transform 1 0 71904 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_312
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_313
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_314
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_315
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_316
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_317
timestamp 1698431365
transform 1 0 44464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_318
timestamp 1698431365
transform 1 0 52304 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_319
timestamp 1698431365
transform 1 0 60144 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_320
timestamp 1698431365
transform 1 0 67984 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_321
timestamp 1698431365
transform 1 0 75824 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_322
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_323
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_324
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_325
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_326
timestamp 1698431365
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_327
timestamp 1698431365
transform 1 0 48384 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_328
timestamp 1698431365
transform 1 0 56224 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_329
timestamp 1698431365
transform 1 0 64064 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_330
timestamp 1698431365
transform 1 0 71904 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_331
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_332
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_333
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_334
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_335
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_336
timestamp 1698431365
transform 1 0 44464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_337
timestamp 1698431365
transform 1 0 52304 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_338
timestamp 1698431365
transform 1 0 60144 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_339
timestamp 1698431365
transform 1 0 67984 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_340
timestamp 1698431365
transform 1 0 75824 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_341
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_342
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_343
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_344
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_345
timestamp 1698431365
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_346
timestamp 1698431365
transform 1 0 48384 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_347
timestamp 1698431365
transform 1 0 56224 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_348
timestamp 1698431365
transform 1 0 64064 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_349
timestamp 1698431365
transform 1 0 71904 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_350
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_351
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_352
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_353
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_354
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_355
timestamp 1698431365
transform 1 0 44464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_356
timestamp 1698431365
transform 1 0 52304 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_357
timestamp 1698431365
transform 1 0 60144 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_358
timestamp 1698431365
transform 1 0 67984 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_359
timestamp 1698431365
transform 1 0 75824 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_360
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_361
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_362
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_363
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_364
timestamp 1698431365
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_365
timestamp 1698431365
transform 1 0 48384 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_366
timestamp 1698431365
transform 1 0 56224 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_367
timestamp 1698431365
transform 1 0 64064 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_368
timestamp 1698431365
transform 1 0 71904 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_369
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_370
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_371
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_372
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_373
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_374
timestamp 1698431365
transform 1 0 44464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_375
timestamp 1698431365
transform 1 0 52304 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_376
timestamp 1698431365
transform 1 0 60144 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_377
timestamp 1698431365
transform 1 0 67984 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_378
timestamp 1698431365
transform 1 0 75824 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_379
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_380
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_381
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_382
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_383
timestamp 1698431365
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_384
timestamp 1698431365
transform 1 0 48384 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_385
timestamp 1698431365
transform 1 0 56224 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_386
timestamp 1698431365
transform 1 0 64064 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_387
timestamp 1698431365
transform 1 0 71904 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_388
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_389
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_390
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_391
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_392
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_393
timestamp 1698431365
transform 1 0 44464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_394
timestamp 1698431365
transform 1 0 52304 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_395
timestamp 1698431365
transform 1 0 60144 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_396
timestamp 1698431365
transform 1 0 67984 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_397
timestamp 1698431365
transform 1 0 75824 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_398
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_399
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_400
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_401
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_402
timestamp 1698431365
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_403
timestamp 1698431365
transform 1 0 48384 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_404
timestamp 1698431365
transform 1 0 56224 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_405
timestamp 1698431365
transform 1 0 64064 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_406
timestamp 1698431365
transform 1 0 71904 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_407
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_408
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_409
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_410
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_411
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_412
timestamp 1698431365
transform 1 0 44464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_413
timestamp 1698431365
transform 1 0 52304 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_414
timestamp 1698431365
transform 1 0 60144 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_415
timestamp 1698431365
transform 1 0 67984 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_416
timestamp 1698431365
transform 1 0 75824 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_417
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_418
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_419
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_420
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_421
timestamp 1698431365
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_422
timestamp 1698431365
transform 1 0 48384 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_423
timestamp 1698431365
transform 1 0 56224 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_424
timestamp 1698431365
transform 1 0 64064 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_425
timestamp 1698431365
transform 1 0 71904 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_426
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_427
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_428
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_429
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_430
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_431
timestamp 1698431365
transform 1 0 44464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_432
timestamp 1698431365
transform 1 0 52304 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_433
timestamp 1698431365
transform 1 0 60144 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_434
timestamp 1698431365
transform 1 0 67984 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_435
timestamp 1698431365
transform 1 0 75824 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_436
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_437
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_438
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_439
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_440
timestamp 1698431365
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_441
timestamp 1698431365
transform 1 0 48384 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_442
timestamp 1698431365
transform 1 0 56224 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_443
timestamp 1698431365
transform 1 0 64064 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_444
timestamp 1698431365
transform 1 0 71904 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_445
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_446
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_447
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_448
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_449
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_450
timestamp 1698431365
transform 1 0 44464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_451
timestamp 1698431365
transform 1 0 52304 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_452
timestamp 1698431365
transform 1 0 60144 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_453
timestamp 1698431365
transform 1 0 67984 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_454
timestamp 1698431365
transform 1 0 75824 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_455
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_456
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_457
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_458
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_459
timestamp 1698431365
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_460
timestamp 1698431365
transform 1 0 48384 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_461
timestamp 1698431365
transform 1 0 56224 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_462
timestamp 1698431365
transform 1 0 64064 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_463
timestamp 1698431365
transform 1 0 71904 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_464
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_465
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_466
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_467
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_468
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_469
timestamp 1698431365
transform 1 0 44464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_470
timestamp 1698431365
transform 1 0 52304 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_471
timestamp 1698431365
transform 1 0 60144 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_472
timestamp 1698431365
transform 1 0 67984 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_473
timestamp 1698431365
transform 1 0 75824 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_474
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_475
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_476
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_477
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_478
timestamp 1698431365
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_479
timestamp 1698431365
transform 1 0 48384 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_480
timestamp 1698431365
transform 1 0 56224 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_481
timestamp 1698431365
transform 1 0 64064 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_482
timestamp 1698431365
transform 1 0 71904 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_483
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_484
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_485
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_486
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_487
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_488
timestamp 1698431365
transform 1 0 44464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_489
timestamp 1698431365
transform 1 0 52304 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_490
timestamp 1698431365
transform 1 0 60144 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_491
timestamp 1698431365
transform 1 0 67984 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_492
timestamp 1698431365
transform 1 0 75824 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_493
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_494
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_495
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_496
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_497
timestamp 1698431365
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_498
timestamp 1698431365
transform 1 0 48384 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_499
timestamp 1698431365
transform 1 0 56224 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_500
timestamp 1698431365
transform 1 0 64064 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_501
timestamp 1698431365
transform 1 0 71904 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_502
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_503
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_504
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_505
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_506
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_507
timestamp 1698431365
transform 1 0 44464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_508
timestamp 1698431365
transform 1 0 52304 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_509
timestamp 1698431365
transform 1 0 60144 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_510
timestamp 1698431365
transform 1 0 67984 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_511
timestamp 1698431365
transform 1 0 75824 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_512
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_513
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_514
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_515
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_516
timestamp 1698431365
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_517
timestamp 1698431365
transform 1 0 48384 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_518
timestamp 1698431365
transform 1 0 56224 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_519
timestamp 1698431365
transform 1 0 64064 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_520
timestamp 1698431365
transform 1 0 71904 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_521
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_522
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_523
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_524
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_525
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_526
timestamp 1698431365
transform 1 0 44464 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_527
timestamp 1698431365
transform 1 0 52304 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_528
timestamp 1698431365
transform 1 0 60144 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_529
timestamp 1698431365
transform 1 0 67984 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_530
timestamp 1698431365
transform 1 0 75824 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_531
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_532
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_533
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_534
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_535
timestamp 1698431365
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_536
timestamp 1698431365
transform 1 0 48384 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_537
timestamp 1698431365
transform 1 0 56224 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_538
timestamp 1698431365
transform 1 0 64064 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_539
timestamp 1698431365
transform 1 0 71904 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_540
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_541
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_542
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_543
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_544
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_545
timestamp 1698431365
transform 1 0 44464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_546
timestamp 1698431365
transform 1 0 52304 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_547
timestamp 1698431365
transform 1 0 60144 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_548
timestamp 1698431365
transform 1 0 67984 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_549
timestamp 1698431365
transform 1 0 75824 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_550
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_551
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_552
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_553
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_554
timestamp 1698431365
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_555
timestamp 1698431365
transform 1 0 48384 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_556
timestamp 1698431365
transform 1 0 56224 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_557
timestamp 1698431365
transform 1 0 64064 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_558
timestamp 1698431365
transform 1 0 71904 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_559
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_560
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_561
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_562
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_563
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_564
timestamp 1698431365
transform 1 0 44464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_565
timestamp 1698431365
transform 1 0 52304 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_566
timestamp 1698431365
transform 1 0 60144 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_567
timestamp 1698431365
transform 1 0 67984 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_568
timestamp 1698431365
transform 1 0 75824 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_569
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_570
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_571
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_572
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_573
timestamp 1698431365
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_574
timestamp 1698431365
transform 1 0 48384 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_575
timestamp 1698431365
transform 1 0 56224 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_576
timestamp 1698431365
transform 1 0 64064 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_577
timestamp 1698431365
transform 1 0 71904 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_578
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_579
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_580
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_581
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_582
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_583
timestamp 1698431365
transform 1 0 44464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_584
timestamp 1698431365
transform 1 0 52304 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_585
timestamp 1698431365
transform 1 0 60144 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_586
timestamp 1698431365
transform 1 0 67984 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_587
timestamp 1698431365
transform 1 0 75824 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_588
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_589
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_590
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_591
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_592
timestamp 1698431365
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_593
timestamp 1698431365
transform 1 0 48384 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_594
timestamp 1698431365
transform 1 0 56224 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_595
timestamp 1698431365
transform 1 0 64064 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_596
timestamp 1698431365
transform 1 0 71904 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_597
timestamp 1698431365
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_598
timestamp 1698431365
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_599
timestamp 1698431365
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_600
timestamp 1698431365
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_601
timestamp 1698431365
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_602
timestamp 1698431365
transform 1 0 44464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_603
timestamp 1698431365
transform 1 0 52304 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_604
timestamp 1698431365
transform 1 0 60144 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_605
timestamp 1698431365
transform 1 0 67984 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_606
timestamp 1698431365
transform 1 0 75824 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_607
timestamp 1698431365
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_608
timestamp 1698431365
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_609
timestamp 1698431365
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_610
timestamp 1698431365
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_611
timestamp 1698431365
transform 1 0 40544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_612
timestamp 1698431365
transform 1 0 48384 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_613
timestamp 1698431365
transform 1 0 56224 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_614
timestamp 1698431365
transform 1 0 64064 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_615
timestamp 1698431365
transform 1 0 71904 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_616
timestamp 1698431365
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_617
timestamp 1698431365
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_618
timestamp 1698431365
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_619
timestamp 1698431365
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_620
timestamp 1698431365
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_621
timestamp 1698431365
transform 1 0 44464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_622
timestamp 1698431365
transform 1 0 52304 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_623
timestamp 1698431365
transform 1 0 60144 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_624
timestamp 1698431365
transform 1 0 67984 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_625
timestamp 1698431365
transform 1 0 75824 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_626
timestamp 1698431365
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_627
timestamp 1698431365
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_628
timestamp 1698431365
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_629
timestamp 1698431365
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_630
timestamp 1698431365
transform 1 0 40544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_631
timestamp 1698431365
transform 1 0 48384 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_632
timestamp 1698431365
transform 1 0 56224 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_633
timestamp 1698431365
transform 1 0 64064 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_634
timestamp 1698431365
transform 1 0 71904 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_635
timestamp 1698431365
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_636
timestamp 1698431365
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_637
timestamp 1698431365
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_638
timestamp 1698431365
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_639
timestamp 1698431365
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_640
timestamp 1698431365
transform 1 0 44464 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_641
timestamp 1698431365
transform 1 0 52304 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_642
timestamp 1698431365
transform 1 0 60144 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_643
timestamp 1698431365
transform 1 0 67984 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_644
timestamp 1698431365
transform 1 0 75824 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_645
timestamp 1698431365
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_646
timestamp 1698431365
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_647
timestamp 1698431365
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_648
timestamp 1698431365
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_649
timestamp 1698431365
transform 1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_650
timestamp 1698431365
transform 1 0 48384 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_651
timestamp 1698431365
transform 1 0 56224 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_652
timestamp 1698431365
transform 1 0 64064 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_653
timestamp 1698431365
transform 1 0 71904 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_654
timestamp 1698431365
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_655
timestamp 1698431365
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_656
timestamp 1698431365
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_657
timestamp 1698431365
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_658
timestamp 1698431365
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_659
timestamp 1698431365
transform 1 0 44464 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_660
timestamp 1698431365
transform 1 0 52304 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_661
timestamp 1698431365
transform 1 0 60144 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_662
timestamp 1698431365
transform 1 0 67984 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_663
timestamp 1698431365
transform 1 0 75824 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_664
timestamp 1698431365
transform 1 0 9184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_665
timestamp 1698431365
transform 1 0 17024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_666
timestamp 1698431365
transform 1 0 24864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_667
timestamp 1698431365
transform 1 0 32704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_668
timestamp 1698431365
transform 1 0 40544 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_669
timestamp 1698431365
transform 1 0 48384 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_670
timestamp 1698431365
transform 1 0 56224 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_671
timestamp 1698431365
transform 1 0 64064 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_672
timestamp 1698431365
transform 1 0 71904 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_673
timestamp 1698431365
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_674
timestamp 1698431365
transform 1 0 13104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_675
timestamp 1698431365
transform 1 0 20944 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_676
timestamp 1698431365
transform 1 0 28784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_677
timestamp 1698431365
transform 1 0 36624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_678
timestamp 1698431365
transform 1 0 44464 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_679
timestamp 1698431365
transform 1 0 52304 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_680
timestamp 1698431365
transform 1 0 60144 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_681
timestamp 1698431365
transform 1 0 67984 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_682
timestamp 1698431365
transform 1 0 75824 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_683
timestamp 1698431365
transform 1 0 9184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_684
timestamp 1698431365
transform 1 0 17024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_685
timestamp 1698431365
transform 1 0 24864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_686
timestamp 1698431365
transform 1 0 32704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_687
timestamp 1698431365
transform 1 0 40544 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_688
timestamp 1698431365
transform 1 0 48384 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_689
timestamp 1698431365
transform 1 0 56224 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_690
timestamp 1698431365
transform 1 0 64064 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_691
timestamp 1698431365
transform 1 0 71904 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_692
timestamp 1698431365
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_693
timestamp 1698431365
transform 1 0 13104 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_694
timestamp 1698431365
transform 1 0 20944 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_695
timestamp 1698431365
transform 1 0 28784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_696
timestamp 1698431365
transform 1 0 36624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_697
timestamp 1698431365
transform 1 0 44464 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_698
timestamp 1698431365
transform 1 0 52304 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_699
timestamp 1698431365
transform 1 0 60144 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_700
timestamp 1698431365
transform 1 0 67984 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_701
timestamp 1698431365
transform 1 0 75824 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_702
timestamp 1698431365
transform 1 0 9184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_703
timestamp 1698431365
transform 1 0 17024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_704
timestamp 1698431365
transform 1 0 24864 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_705
timestamp 1698431365
transform 1 0 32704 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_706
timestamp 1698431365
transform 1 0 40544 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_707
timestamp 1698431365
transform 1 0 48384 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_708
timestamp 1698431365
transform 1 0 56224 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_709
timestamp 1698431365
transform 1 0 64064 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_710
timestamp 1698431365
transform 1 0 71904 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_711
timestamp 1698431365
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_712
timestamp 1698431365
transform 1 0 13104 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_713
timestamp 1698431365
transform 1 0 20944 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_714
timestamp 1698431365
transform 1 0 28784 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_715
timestamp 1698431365
transform 1 0 36624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_716
timestamp 1698431365
transform 1 0 44464 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_717
timestamp 1698431365
transform 1 0 52304 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_718
timestamp 1698431365
transform 1 0 60144 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_719
timestamp 1698431365
transform 1 0 67984 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_720
timestamp 1698431365
transform 1 0 75824 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_721
timestamp 1698431365
transform 1 0 9184 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_722
timestamp 1698431365
transform 1 0 17024 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_723
timestamp 1698431365
transform 1 0 24864 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_724
timestamp 1698431365
transform 1 0 32704 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_725
timestamp 1698431365
transform 1 0 40544 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_726
timestamp 1698431365
transform 1 0 48384 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_727
timestamp 1698431365
transform 1 0 56224 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_728
timestamp 1698431365
transform 1 0 64064 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_729
timestamp 1698431365
transform 1 0 71904 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_730
timestamp 1698431365
transform 1 0 5264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_731
timestamp 1698431365
transform 1 0 13104 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_732
timestamp 1698431365
transform 1 0 20944 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_733
timestamp 1698431365
transform 1 0 28784 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_734
timestamp 1698431365
transform 1 0 36624 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_735
timestamp 1698431365
transform 1 0 44464 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_736
timestamp 1698431365
transform 1 0 52304 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_737
timestamp 1698431365
transform 1 0 60144 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_738
timestamp 1698431365
transform 1 0 67984 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_739
timestamp 1698431365
transform 1 0 75824 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_740
timestamp 1698431365
transform 1 0 9184 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_741
timestamp 1698431365
transform 1 0 17024 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_742
timestamp 1698431365
transform 1 0 24864 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_743
timestamp 1698431365
transform 1 0 32704 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_744
timestamp 1698431365
transform 1 0 40544 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_745
timestamp 1698431365
transform 1 0 48384 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_746
timestamp 1698431365
transform 1 0 56224 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_747
timestamp 1698431365
transform 1 0 64064 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_748
timestamp 1698431365
transform 1 0 71904 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_749
timestamp 1698431365
transform 1 0 5264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_750
timestamp 1698431365
transform 1 0 13104 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_751
timestamp 1698431365
transform 1 0 20944 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_752
timestamp 1698431365
transform 1 0 28784 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_753
timestamp 1698431365
transform 1 0 36624 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_754
timestamp 1698431365
transform 1 0 44464 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_755
timestamp 1698431365
transform 1 0 52304 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_756
timestamp 1698431365
transform 1 0 60144 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_757
timestamp 1698431365
transform 1 0 67984 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_758
timestamp 1698431365
transform 1 0 75824 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_759
timestamp 1698431365
transform 1 0 9184 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_760
timestamp 1698431365
transform 1 0 17024 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_761
timestamp 1698431365
transform 1 0 24864 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_762
timestamp 1698431365
transform 1 0 32704 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_763
timestamp 1698431365
transform 1 0 40544 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_764
timestamp 1698431365
transform 1 0 48384 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_765
timestamp 1698431365
transform 1 0 56224 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_766
timestamp 1698431365
transform 1 0 64064 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_767
timestamp 1698431365
transform 1 0 71904 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_768
timestamp 1698431365
transform 1 0 5264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_769
timestamp 1698431365
transform 1 0 13104 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_770
timestamp 1698431365
transform 1 0 20944 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_771
timestamp 1698431365
transform 1 0 28784 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_772
timestamp 1698431365
transform 1 0 36624 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_773
timestamp 1698431365
transform 1 0 44464 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_774
timestamp 1698431365
transform 1 0 52304 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_775
timestamp 1698431365
transform 1 0 60144 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_776
timestamp 1698431365
transform 1 0 67984 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_777
timestamp 1698431365
transform 1 0 75824 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_778
timestamp 1698431365
transform 1 0 9184 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_779
timestamp 1698431365
transform 1 0 17024 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_780
timestamp 1698431365
transform 1 0 24864 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_781
timestamp 1698431365
transform 1 0 32704 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_782
timestamp 1698431365
transform 1 0 40544 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_783
timestamp 1698431365
transform 1 0 48384 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_784
timestamp 1698431365
transform 1 0 56224 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_785
timestamp 1698431365
transform 1 0 64064 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_786
timestamp 1698431365
transform 1 0 71904 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_787
timestamp 1698431365
transform 1 0 5264 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_788
timestamp 1698431365
transform 1 0 13104 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_789
timestamp 1698431365
transform 1 0 20944 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_790
timestamp 1698431365
transform 1 0 28784 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_791
timestamp 1698431365
transform 1 0 36624 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_792
timestamp 1698431365
transform 1 0 44464 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_793
timestamp 1698431365
transform 1 0 52304 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_794
timestamp 1698431365
transform 1 0 60144 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_795
timestamp 1698431365
transform 1 0 67984 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_796
timestamp 1698431365
transform 1 0 75824 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_797
timestamp 1698431365
transform 1 0 9184 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_798
timestamp 1698431365
transform 1 0 17024 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_799
timestamp 1698431365
transform 1 0 24864 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_800
timestamp 1698431365
transform 1 0 32704 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_801
timestamp 1698431365
transform 1 0 40544 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_802
timestamp 1698431365
transform 1 0 48384 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_803
timestamp 1698431365
transform 1 0 56224 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_804
timestamp 1698431365
transform 1 0 64064 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_805
timestamp 1698431365
transform 1 0 71904 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_806
timestamp 1698431365
transform 1 0 5264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_807
timestamp 1698431365
transform 1 0 13104 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_808
timestamp 1698431365
transform 1 0 20944 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_809
timestamp 1698431365
transform 1 0 28784 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_810
timestamp 1698431365
transform 1 0 36624 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_811
timestamp 1698431365
transform 1 0 44464 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_812
timestamp 1698431365
transform 1 0 52304 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_813
timestamp 1698431365
transform 1 0 60144 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_814
timestamp 1698431365
transform 1 0 67984 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_815
timestamp 1698431365
transform 1 0 75824 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_816
timestamp 1698431365
transform 1 0 9184 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_817
timestamp 1698431365
transform 1 0 17024 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_818
timestamp 1698431365
transform 1 0 24864 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_819
timestamp 1698431365
transform 1 0 32704 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_820
timestamp 1698431365
transform 1 0 40544 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_821
timestamp 1698431365
transform 1 0 48384 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_822
timestamp 1698431365
transform 1 0 56224 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_823
timestamp 1698431365
transform 1 0 64064 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_824
timestamp 1698431365
transform 1 0 71904 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_825
timestamp 1698431365
transform 1 0 5264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_826
timestamp 1698431365
transform 1 0 13104 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_827
timestamp 1698431365
transform 1 0 20944 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_828
timestamp 1698431365
transform 1 0 28784 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_829
timestamp 1698431365
transform 1 0 36624 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_830
timestamp 1698431365
transform 1 0 44464 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_831
timestamp 1698431365
transform 1 0 52304 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_832
timestamp 1698431365
transform 1 0 60144 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_833
timestamp 1698431365
transform 1 0 67984 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_834
timestamp 1698431365
transform 1 0 75824 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_835
timestamp 1698431365
transform 1 0 9184 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_836
timestamp 1698431365
transform 1 0 17024 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_837
timestamp 1698431365
transform 1 0 24864 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_838
timestamp 1698431365
transform 1 0 32704 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_839
timestamp 1698431365
transform 1 0 40544 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_840
timestamp 1698431365
transform 1 0 48384 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_841
timestamp 1698431365
transform 1 0 56224 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_842
timestamp 1698431365
transform 1 0 64064 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_843
timestamp 1698431365
transform 1 0 71904 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_844
timestamp 1698431365
transform 1 0 5264 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_845
timestamp 1698431365
transform 1 0 13104 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_846
timestamp 1698431365
transform 1 0 20944 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_847
timestamp 1698431365
transform 1 0 28784 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_848
timestamp 1698431365
transform 1 0 36624 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_849
timestamp 1698431365
transform 1 0 44464 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_850
timestamp 1698431365
transform 1 0 52304 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_851
timestamp 1698431365
transform 1 0 60144 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_852
timestamp 1698431365
transform 1 0 67984 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_853
timestamp 1698431365
transform 1 0 75824 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_854
timestamp 1698431365
transform 1 0 9184 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_855
timestamp 1698431365
transform 1 0 17024 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_856
timestamp 1698431365
transform 1 0 24864 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_857
timestamp 1698431365
transform 1 0 32704 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_858
timestamp 1698431365
transform 1 0 40544 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_859
timestamp 1698431365
transform 1 0 48384 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_860
timestamp 1698431365
transform 1 0 56224 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_861
timestamp 1698431365
transform 1 0 64064 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_862
timestamp 1698431365
transform 1 0 71904 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_863
timestamp 1698431365
transform 1 0 5264 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_864
timestamp 1698431365
transform 1 0 13104 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_865
timestamp 1698431365
transform 1 0 20944 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_866
timestamp 1698431365
transform 1 0 28784 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_867
timestamp 1698431365
transform 1 0 36624 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_868
timestamp 1698431365
transform 1 0 44464 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_869
timestamp 1698431365
transform 1 0 52304 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_870
timestamp 1698431365
transform 1 0 60144 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_871
timestamp 1698431365
transform 1 0 67984 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_872
timestamp 1698431365
transform 1 0 75824 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_873
timestamp 1698431365
transform 1 0 9184 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_874
timestamp 1698431365
transform 1 0 17024 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_875
timestamp 1698431365
transform 1 0 24864 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_876
timestamp 1698431365
transform 1 0 32704 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_877
timestamp 1698431365
transform 1 0 40544 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_878
timestamp 1698431365
transform 1 0 48384 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_879
timestamp 1698431365
transform 1 0 56224 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_880
timestamp 1698431365
transform 1 0 64064 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_881
timestamp 1698431365
transform 1 0 71904 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_882
timestamp 1698431365
transform 1 0 5264 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_883
timestamp 1698431365
transform 1 0 13104 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_884
timestamp 1698431365
transform 1 0 20944 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_885
timestamp 1698431365
transform 1 0 28784 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_886
timestamp 1698431365
transform 1 0 36624 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_887
timestamp 1698431365
transform 1 0 44464 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_888
timestamp 1698431365
transform 1 0 52304 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_889
timestamp 1698431365
transform 1 0 60144 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_890
timestamp 1698431365
transform 1 0 67984 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_891
timestamp 1698431365
transform 1 0 75824 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_892
timestamp 1698431365
transform 1 0 9184 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_893
timestamp 1698431365
transform 1 0 17024 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_894
timestamp 1698431365
transform 1 0 24864 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_895
timestamp 1698431365
transform 1 0 32704 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_896
timestamp 1698431365
transform 1 0 40544 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_897
timestamp 1698431365
transform 1 0 48384 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_898
timestamp 1698431365
transform 1 0 56224 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_899
timestamp 1698431365
transform 1 0 64064 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_900
timestamp 1698431365
transform 1 0 71904 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_901
timestamp 1698431365
transform 1 0 5264 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_902
timestamp 1698431365
transform 1 0 13104 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_903
timestamp 1698431365
transform 1 0 20944 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_904
timestamp 1698431365
transform 1 0 28784 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_905
timestamp 1698431365
transform 1 0 36624 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_906
timestamp 1698431365
transform 1 0 44464 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_907
timestamp 1698431365
transform 1 0 52304 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_908
timestamp 1698431365
transform 1 0 60144 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_909
timestamp 1698431365
transform 1 0 67984 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_910
timestamp 1698431365
transform 1 0 75824 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_911
timestamp 1698431365
transform 1 0 9184 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_912
timestamp 1698431365
transform 1 0 17024 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_913
timestamp 1698431365
transform 1 0 24864 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_914
timestamp 1698431365
transform 1 0 32704 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_915
timestamp 1698431365
transform 1 0 40544 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_916
timestamp 1698431365
transform 1 0 48384 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_917
timestamp 1698431365
transform 1 0 56224 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_918
timestamp 1698431365
transform 1 0 64064 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_919
timestamp 1698431365
transform 1 0 71904 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_920
timestamp 1698431365
transform 1 0 5264 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_921
timestamp 1698431365
transform 1 0 13104 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_922
timestamp 1698431365
transform 1 0 20944 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_923
timestamp 1698431365
transform 1 0 28784 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_924
timestamp 1698431365
transform 1 0 36624 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_925
timestamp 1698431365
transform 1 0 44464 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_926
timestamp 1698431365
transform 1 0 52304 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_927
timestamp 1698431365
transform 1 0 60144 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_928
timestamp 1698431365
transform 1 0 67984 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_929
timestamp 1698431365
transform 1 0 75824 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_930
timestamp 1698431365
transform 1 0 9184 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_931
timestamp 1698431365
transform 1 0 17024 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_932
timestamp 1698431365
transform 1 0 24864 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_933
timestamp 1698431365
transform 1 0 32704 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_934
timestamp 1698431365
transform 1 0 40544 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_935
timestamp 1698431365
transform 1 0 48384 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_936
timestamp 1698431365
transform 1 0 56224 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_937
timestamp 1698431365
transform 1 0 64064 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_938
timestamp 1698431365
transform 1 0 71904 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_939
timestamp 1698431365
transform 1 0 5264 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_940
timestamp 1698431365
transform 1 0 13104 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_941
timestamp 1698431365
transform 1 0 20944 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_942
timestamp 1698431365
transform 1 0 28784 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_943
timestamp 1698431365
transform 1 0 36624 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_944
timestamp 1698431365
transform 1 0 44464 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_945
timestamp 1698431365
transform 1 0 52304 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_946
timestamp 1698431365
transform 1 0 60144 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_947
timestamp 1698431365
transform 1 0 67984 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_948
timestamp 1698431365
transform 1 0 75824 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_949
timestamp 1698431365
transform 1 0 9184 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_950
timestamp 1698431365
transform 1 0 17024 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_951
timestamp 1698431365
transform 1 0 24864 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_952
timestamp 1698431365
transform 1 0 32704 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_953
timestamp 1698431365
transform 1 0 40544 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_954
timestamp 1698431365
transform 1 0 48384 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_955
timestamp 1698431365
transform 1 0 56224 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_956
timestamp 1698431365
transform 1 0 64064 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_957
timestamp 1698431365
transform 1 0 71904 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_958
timestamp 1698431365
transform 1 0 5264 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_959
timestamp 1698431365
transform 1 0 13104 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_960
timestamp 1698431365
transform 1 0 20944 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_961
timestamp 1698431365
transform 1 0 28784 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_962
timestamp 1698431365
transform 1 0 36624 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_963
timestamp 1698431365
transform 1 0 44464 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_964
timestamp 1698431365
transform 1 0 52304 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_965
timestamp 1698431365
transform 1 0 60144 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_966
timestamp 1698431365
transform 1 0 67984 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_967
timestamp 1698431365
transform 1 0 75824 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_968
timestamp 1698431365
transform 1 0 9184 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_969
timestamp 1698431365
transform 1 0 17024 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_970
timestamp 1698431365
transform 1 0 24864 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_971
timestamp 1698431365
transform 1 0 32704 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_972
timestamp 1698431365
transform 1 0 40544 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_973
timestamp 1698431365
transform 1 0 48384 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_974
timestamp 1698431365
transform 1 0 56224 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_975
timestamp 1698431365
transform 1 0 64064 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_976
timestamp 1698431365
transform 1 0 71904 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_977
timestamp 1698431365
transform 1 0 5264 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_978
timestamp 1698431365
transform 1 0 13104 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_979
timestamp 1698431365
transform 1 0 20944 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_980
timestamp 1698431365
transform 1 0 28784 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_981
timestamp 1698431365
transform 1 0 36624 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_982
timestamp 1698431365
transform 1 0 44464 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_983
timestamp 1698431365
transform 1 0 52304 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_984
timestamp 1698431365
transform 1 0 60144 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_985
timestamp 1698431365
transform 1 0 67984 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_986
timestamp 1698431365
transform 1 0 75824 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_987
timestamp 1698431365
transform 1 0 9184 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_988
timestamp 1698431365
transform 1 0 17024 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_989
timestamp 1698431365
transform 1 0 24864 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_990
timestamp 1698431365
transform 1 0 32704 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_991
timestamp 1698431365
transform 1 0 40544 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_992
timestamp 1698431365
transform 1 0 48384 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_993
timestamp 1698431365
transform 1 0 56224 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_994
timestamp 1698431365
transform 1 0 64064 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_995
timestamp 1698431365
transform 1 0 71904 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_996
timestamp 1698431365
transform 1 0 5264 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_997
timestamp 1698431365
transform 1 0 13104 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_998
timestamp 1698431365
transform 1 0 20944 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_999
timestamp 1698431365
transform 1 0 28784 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_1000
timestamp 1698431365
transform 1 0 36624 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_1001
timestamp 1698431365
transform 1 0 44464 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_1002
timestamp 1698431365
transform 1 0 52304 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_1003
timestamp 1698431365
transform 1 0 60144 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_1004
timestamp 1698431365
transform 1 0 67984 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_1005
timestamp 1698431365
transform 1 0 75824 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_1006
timestamp 1698431365
transform 1 0 9184 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_1007
timestamp 1698431365
transform 1 0 17024 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_1008
timestamp 1698431365
transform 1 0 24864 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_1009
timestamp 1698431365
transform 1 0 32704 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_1010
timestamp 1698431365
transform 1 0 40544 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_1011
timestamp 1698431365
transform 1 0 48384 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_1012
timestamp 1698431365
transform 1 0 56224 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_1013
timestamp 1698431365
transform 1 0 64064 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_1014
timestamp 1698431365
transform 1 0 71904 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_1015
timestamp 1698431365
transform 1 0 5264 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_1016
timestamp 1698431365
transform 1 0 13104 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_1017
timestamp 1698431365
transform 1 0 20944 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_1018
timestamp 1698431365
transform 1 0 28784 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_1019
timestamp 1698431365
transform 1 0 36624 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_1020
timestamp 1698431365
transform 1 0 44464 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_1021
timestamp 1698431365
transform 1 0 52304 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_1022
timestamp 1698431365
transform 1 0 60144 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_1023
timestamp 1698431365
transform 1 0 67984 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_1024
timestamp 1698431365
transform 1 0 75824 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_1025
timestamp 1698431365
transform 1 0 9184 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_1026
timestamp 1698431365
transform 1 0 17024 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_1027
timestamp 1698431365
transform 1 0 24864 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_1028
timestamp 1698431365
transform 1 0 32704 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_1029
timestamp 1698431365
transform 1 0 40544 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_1030
timestamp 1698431365
transform 1 0 48384 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_1031
timestamp 1698431365
transform 1 0 56224 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_1032
timestamp 1698431365
transform 1 0 64064 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_1033
timestamp 1698431365
transform 1 0 71904 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_1034
timestamp 1698431365
transform 1 0 5264 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_1035
timestamp 1698431365
transform 1 0 13104 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_1036
timestamp 1698431365
transform 1 0 20944 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_1037
timestamp 1698431365
transform 1 0 28784 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_1038
timestamp 1698431365
transform 1 0 36624 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_1039
timestamp 1698431365
transform 1 0 44464 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_1040
timestamp 1698431365
transform 1 0 52304 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_1041
timestamp 1698431365
transform 1 0 60144 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_1042
timestamp 1698431365
transform 1 0 67984 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_1043
timestamp 1698431365
transform 1 0 75824 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_1044
timestamp 1698431365
transform 1 0 9184 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_1045
timestamp 1698431365
transform 1 0 17024 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_1046
timestamp 1698431365
transform 1 0 24864 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_1047
timestamp 1698431365
transform 1 0 32704 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_1048
timestamp 1698431365
transform 1 0 40544 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_1049
timestamp 1698431365
transform 1 0 48384 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_1050
timestamp 1698431365
transform 1 0 56224 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_1051
timestamp 1698431365
transform 1 0 64064 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_1052
timestamp 1698431365
transform 1 0 71904 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_1053
timestamp 1698431365
transform 1 0 5264 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_1054
timestamp 1698431365
transform 1 0 13104 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_1055
timestamp 1698431365
transform 1 0 20944 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_1056
timestamp 1698431365
transform 1 0 28784 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_1057
timestamp 1698431365
transform 1 0 36624 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_1058
timestamp 1698431365
transform 1 0 44464 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_1059
timestamp 1698431365
transform 1 0 52304 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_1060
timestamp 1698431365
transform 1 0 60144 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_1061
timestamp 1698431365
transform 1 0 67984 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_1062
timestamp 1698431365
transform 1 0 75824 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_1063
timestamp 1698431365
transform 1 0 9184 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_1064
timestamp 1698431365
transform 1 0 17024 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_1065
timestamp 1698431365
transform 1 0 24864 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_1066
timestamp 1698431365
transform 1 0 32704 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_1067
timestamp 1698431365
transform 1 0 40544 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_1068
timestamp 1698431365
transform 1 0 48384 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_1069
timestamp 1698431365
transform 1 0 56224 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_1070
timestamp 1698431365
transform 1 0 64064 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_1071
timestamp 1698431365
transform 1 0 71904 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_1072
timestamp 1698431365
transform 1 0 5264 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_1073
timestamp 1698431365
transform 1 0 13104 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_1074
timestamp 1698431365
transform 1 0 20944 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_1075
timestamp 1698431365
transform 1 0 28784 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_1076
timestamp 1698431365
transform 1 0 36624 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_1077
timestamp 1698431365
transform 1 0 44464 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_1078
timestamp 1698431365
transform 1 0 52304 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_1079
timestamp 1698431365
transform 1 0 60144 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_1080
timestamp 1698431365
transform 1 0 67984 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_1081
timestamp 1698431365
transform 1 0 75824 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1082
timestamp 1698431365
transform 1 0 5152 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1083
timestamp 1698431365
transform 1 0 8960 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1084
timestamp 1698431365
transform 1 0 12768 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1085
timestamp 1698431365
transform 1 0 16576 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1086
timestamp 1698431365
transform 1 0 20384 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1087
timestamp 1698431365
transform 1 0 24192 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1088
timestamp 1698431365
transform 1 0 28000 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1089
timestamp 1698431365
transform 1 0 31808 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1090
timestamp 1698431365
transform 1 0 35616 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1091
timestamp 1698431365
transform 1 0 39424 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1092
timestamp 1698431365
transform 1 0 43232 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1093
timestamp 1698431365
transform 1 0 47040 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1094
timestamp 1698431365
transform 1 0 50848 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1095
timestamp 1698431365
transform 1 0 54656 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1096
timestamp 1698431365
transform 1 0 58464 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1097
timestamp 1698431365
transform 1 0 62272 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1098
timestamp 1698431365
transform 1 0 66080 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1099
timestamp 1698431365
transform 1 0 69888 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1100
timestamp 1698431365
transform 1 0 73696 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1101
timestamp 1698431365
transform 1 0 77504 0 -1 76832
box -86 -86 310 870
<< labels >>
flabel metal2 s 74144 0 74256 800 0 FreeSans 448 90 0 0 clk
port 0 nsew signal input
flabel metal2 s 448 79200 560 80000 0 FreeSans 448 90 0 0 gpio_in[0]
port 1 nsew signal input
flabel metal2 s 7168 79200 7280 80000 0 FreeSans 448 90 0 0 gpio_in[10]
port 2 nsew signal input
flabel metal2 s 7840 79200 7952 80000 0 FreeSans 448 90 0 0 gpio_in[11]
port 3 nsew signal input
flabel metal2 s 8512 79200 8624 80000 0 FreeSans 448 90 0 0 gpio_in[12]
port 4 nsew signal input
flabel metal2 s 9184 79200 9296 80000 0 FreeSans 448 90 0 0 gpio_in[13]
port 5 nsew signal input
flabel metal2 s 9856 79200 9968 80000 0 FreeSans 448 90 0 0 gpio_in[14]
port 6 nsew signal input
flabel metal2 s 10528 79200 10640 80000 0 FreeSans 448 90 0 0 gpio_in[15]
port 7 nsew signal input
flabel metal2 s 1120 79200 1232 80000 0 FreeSans 448 90 0 0 gpio_in[1]
port 8 nsew signal input
flabel metal2 s 1792 79200 1904 80000 0 FreeSans 448 90 0 0 gpio_in[2]
port 9 nsew signal input
flabel metal2 s 2464 79200 2576 80000 0 FreeSans 448 90 0 0 gpio_in[3]
port 10 nsew signal input
flabel metal2 s 3136 79200 3248 80000 0 FreeSans 448 90 0 0 gpio_in[4]
port 11 nsew signal input
flabel metal2 s 3808 79200 3920 80000 0 FreeSans 448 90 0 0 gpio_in[5]
port 12 nsew signal input
flabel metal2 s 4480 79200 4592 80000 0 FreeSans 448 90 0 0 gpio_in[6]
port 13 nsew signal input
flabel metal2 s 5152 79200 5264 80000 0 FreeSans 448 90 0 0 gpio_in[7]
port 14 nsew signal input
flabel metal2 s 5824 79200 5936 80000 0 FreeSans 448 90 0 0 gpio_in[8]
port 15 nsew signal input
flabel metal2 s 6496 79200 6608 80000 0 FreeSans 448 90 0 0 gpio_in[9]
port 16 nsew signal input
flabel metal2 s 21952 79200 22064 80000 0 FreeSans 448 90 0 0 gpio_oeb[0]
port 17 nsew signal tristate
flabel metal2 s 28672 79200 28784 80000 0 FreeSans 448 90 0 0 gpio_oeb[10]
port 18 nsew signal tristate
flabel metal2 s 29344 79200 29456 80000 0 FreeSans 448 90 0 0 gpio_oeb[11]
port 19 nsew signal tristate
flabel metal2 s 30016 79200 30128 80000 0 FreeSans 448 90 0 0 gpio_oeb[12]
port 20 nsew signal tristate
flabel metal2 s 30688 79200 30800 80000 0 FreeSans 448 90 0 0 gpio_oeb[13]
port 21 nsew signal tristate
flabel metal2 s 31360 79200 31472 80000 0 FreeSans 448 90 0 0 gpio_oeb[14]
port 22 nsew signal tristate
flabel metal2 s 32032 79200 32144 80000 0 FreeSans 448 90 0 0 gpio_oeb[15]
port 23 nsew signal tristate
flabel metal2 s 22624 79200 22736 80000 0 FreeSans 448 90 0 0 gpio_oeb[1]
port 24 nsew signal tristate
flabel metal2 s 23296 79200 23408 80000 0 FreeSans 448 90 0 0 gpio_oeb[2]
port 25 nsew signal tristate
flabel metal2 s 23968 79200 24080 80000 0 FreeSans 448 90 0 0 gpio_oeb[3]
port 26 nsew signal tristate
flabel metal2 s 24640 79200 24752 80000 0 FreeSans 448 90 0 0 gpio_oeb[4]
port 27 nsew signal tristate
flabel metal2 s 25312 79200 25424 80000 0 FreeSans 448 90 0 0 gpio_oeb[5]
port 28 nsew signal tristate
flabel metal2 s 25984 79200 26096 80000 0 FreeSans 448 90 0 0 gpio_oeb[6]
port 29 nsew signal tristate
flabel metal2 s 26656 79200 26768 80000 0 FreeSans 448 90 0 0 gpio_oeb[7]
port 30 nsew signal tristate
flabel metal2 s 27328 79200 27440 80000 0 FreeSans 448 90 0 0 gpio_oeb[8]
port 31 nsew signal tristate
flabel metal2 s 28000 79200 28112 80000 0 FreeSans 448 90 0 0 gpio_oeb[9]
port 32 nsew signal tristate
flabel metal2 s 11200 79200 11312 80000 0 FreeSans 448 90 0 0 gpio_out[0]
port 33 nsew signal tristate
flabel metal2 s 17920 79200 18032 80000 0 FreeSans 448 90 0 0 gpio_out[10]
port 34 nsew signal tristate
flabel metal2 s 18592 79200 18704 80000 0 FreeSans 448 90 0 0 gpio_out[11]
port 35 nsew signal tristate
flabel metal2 s 19264 79200 19376 80000 0 FreeSans 448 90 0 0 gpio_out[12]
port 36 nsew signal tristate
flabel metal2 s 19936 79200 20048 80000 0 FreeSans 448 90 0 0 gpio_out[13]
port 37 nsew signal tristate
flabel metal2 s 20608 79200 20720 80000 0 FreeSans 448 90 0 0 gpio_out[14]
port 38 nsew signal tristate
flabel metal2 s 21280 79200 21392 80000 0 FreeSans 448 90 0 0 gpio_out[15]
port 39 nsew signal tristate
flabel metal2 s 11872 79200 11984 80000 0 FreeSans 448 90 0 0 gpio_out[1]
port 40 nsew signal tristate
flabel metal2 s 12544 79200 12656 80000 0 FreeSans 448 90 0 0 gpio_out[2]
port 41 nsew signal tristate
flabel metal2 s 13216 79200 13328 80000 0 FreeSans 448 90 0 0 gpio_out[3]
port 42 nsew signal tristate
flabel metal2 s 13888 79200 14000 80000 0 FreeSans 448 90 0 0 gpio_out[4]
port 43 nsew signal tristate
flabel metal2 s 14560 79200 14672 80000 0 FreeSans 448 90 0 0 gpio_out[5]
port 44 nsew signal tristate
flabel metal2 s 15232 79200 15344 80000 0 FreeSans 448 90 0 0 gpio_out[6]
port 45 nsew signal tristate
flabel metal2 s 15904 79200 16016 80000 0 FreeSans 448 90 0 0 gpio_out[7]
port 46 nsew signal tristate
flabel metal2 s 16576 79200 16688 80000 0 FreeSans 448 90 0 0 gpio_out[8]
port 47 nsew signal tristate
flabel metal2 s 17248 79200 17360 80000 0 FreeSans 448 90 0 0 gpio_out[9]
port 48 nsew signal tristate
flabel metal2 s 26432 0 26544 800 0 FreeSans 448 90 0 0 mem_addr[0]
port 49 nsew signal input
flabel metal2 s 33152 0 33264 800 0 FreeSans 448 90 0 0 mem_addr[10]
port 50 nsew signal input
flabel metal2 s 33824 0 33936 800 0 FreeSans 448 90 0 0 mem_addr[11]
port 51 nsew signal input
flabel metal2 s 34496 0 34608 800 0 FreeSans 448 90 0 0 mem_addr[12]
port 52 nsew signal input
flabel metal2 s 35168 0 35280 800 0 FreeSans 448 90 0 0 mem_addr[13]
port 53 nsew signal input
flabel metal2 s 35840 0 35952 800 0 FreeSans 448 90 0 0 mem_addr[14]
port 54 nsew signal input
flabel metal2 s 36512 0 36624 800 0 FreeSans 448 90 0 0 mem_addr[15]
port 55 nsew signal input
flabel metal2 s 37184 0 37296 800 0 FreeSans 448 90 0 0 mem_addr[16]
port 56 nsew signal input
flabel metal2 s 37856 0 37968 800 0 FreeSans 448 90 0 0 mem_addr[17]
port 57 nsew signal input
flabel metal2 s 38528 0 38640 800 0 FreeSans 448 90 0 0 mem_addr[18]
port 58 nsew signal input
flabel metal2 s 39200 0 39312 800 0 FreeSans 448 90 0 0 mem_addr[19]
port 59 nsew signal input
flabel metal2 s 27104 0 27216 800 0 FreeSans 448 90 0 0 mem_addr[1]
port 60 nsew signal input
flabel metal2 s 39872 0 39984 800 0 FreeSans 448 90 0 0 mem_addr[20]
port 61 nsew signal input
flabel metal2 s 40544 0 40656 800 0 FreeSans 448 90 0 0 mem_addr[21]
port 62 nsew signal input
flabel metal2 s 41216 0 41328 800 0 FreeSans 448 90 0 0 mem_addr[22]
port 63 nsew signal input
flabel metal2 s 41888 0 42000 800 0 FreeSans 448 90 0 0 mem_addr[23]
port 64 nsew signal input
flabel metal2 s 42560 0 42672 800 0 FreeSans 448 90 0 0 mem_addr[24]
port 65 nsew signal input
flabel metal2 s 43232 0 43344 800 0 FreeSans 448 90 0 0 mem_addr[25]
port 66 nsew signal input
flabel metal2 s 43904 0 44016 800 0 FreeSans 448 90 0 0 mem_addr[26]
port 67 nsew signal input
flabel metal2 s 44576 0 44688 800 0 FreeSans 448 90 0 0 mem_addr[27]
port 68 nsew signal input
flabel metal2 s 45248 0 45360 800 0 FreeSans 448 90 0 0 mem_addr[28]
port 69 nsew signal input
flabel metal2 s 45920 0 46032 800 0 FreeSans 448 90 0 0 mem_addr[29]
port 70 nsew signal input
flabel metal2 s 27776 0 27888 800 0 FreeSans 448 90 0 0 mem_addr[2]
port 71 nsew signal input
flabel metal2 s 46592 0 46704 800 0 FreeSans 448 90 0 0 mem_addr[30]
port 72 nsew signal input
flabel metal2 s 47264 0 47376 800 0 FreeSans 448 90 0 0 mem_addr[31]
port 73 nsew signal input
flabel metal2 s 28448 0 28560 800 0 FreeSans 448 90 0 0 mem_addr[3]
port 74 nsew signal input
flabel metal2 s 29120 0 29232 800 0 FreeSans 448 90 0 0 mem_addr[4]
port 75 nsew signal input
flabel metal2 s 29792 0 29904 800 0 FreeSans 448 90 0 0 mem_addr[5]
port 76 nsew signal input
flabel metal2 s 30464 0 30576 800 0 FreeSans 448 90 0 0 mem_addr[6]
port 77 nsew signal input
flabel metal2 s 31136 0 31248 800 0 FreeSans 448 90 0 0 mem_addr[7]
port 78 nsew signal input
flabel metal2 s 31808 0 31920 800 0 FreeSans 448 90 0 0 mem_addr[8]
port 79 nsew signal input
flabel metal2 s 32480 0 32592 800 0 FreeSans 448 90 0 0 mem_addr[9]
port 80 nsew signal input
flabel metal2 s 48608 0 48720 800 0 FreeSans 448 90 0 0 mem_instr
port 81 nsew signal input
flabel metal2 s 52640 0 52752 800 0 FreeSans 448 90 0 0 mem_rdata[0]
port 82 nsew signal tristate
flabel metal2 s 59360 0 59472 800 0 FreeSans 448 90 0 0 mem_rdata[10]
port 83 nsew signal tristate
flabel metal2 s 60032 0 60144 800 0 FreeSans 448 90 0 0 mem_rdata[11]
port 84 nsew signal tristate
flabel metal2 s 60704 0 60816 800 0 FreeSans 448 90 0 0 mem_rdata[12]
port 85 nsew signal tristate
flabel metal2 s 61376 0 61488 800 0 FreeSans 448 90 0 0 mem_rdata[13]
port 86 nsew signal tristate
flabel metal2 s 62048 0 62160 800 0 FreeSans 448 90 0 0 mem_rdata[14]
port 87 nsew signal tristate
flabel metal2 s 62720 0 62832 800 0 FreeSans 448 90 0 0 mem_rdata[15]
port 88 nsew signal tristate
flabel metal2 s 63392 0 63504 800 0 FreeSans 448 90 0 0 mem_rdata[16]
port 89 nsew signal tristate
flabel metal2 s 64064 0 64176 800 0 FreeSans 448 90 0 0 mem_rdata[17]
port 90 nsew signal tristate
flabel metal2 s 64736 0 64848 800 0 FreeSans 448 90 0 0 mem_rdata[18]
port 91 nsew signal tristate
flabel metal2 s 65408 0 65520 800 0 FreeSans 448 90 0 0 mem_rdata[19]
port 92 nsew signal tristate
flabel metal2 s 53312 0 53424 800 0 FreeSans 448 90 0 0 mem_rdata[1]
port 93 nsew signal tristate
flabel metal2 s 66080 0 66192 800 0 FreeSans 448 90 0 0 mem_rdata[20]
port 94 nsew signal tristate
flabel metal2 s 66752 0 66864 800 0 FreeSans 448 90 0 0 mem_rdata[21]
port 95 nsew signal tristate
flabel metal2 s 67424 0 67536 800 0 FreeSans 448 90 0 0 mem_rdata[22]
port 96 nsew signal tristate
flabel metal2 s 68096 0 68208 800 0 FreeSans 448 90 0 0 mem_rdata[23]
port 97 nsew signal tristate
flabel metal2 s 68768 0 68880 800 0 FreeSans 448 90 0 0 mem_rdata[24]
port 98 nsew signal tristate
flabel metal2 s 69440 0 69552 800 0 FreeSans 448 90 0 0 mem_rdata[25]
port 99 nsew signal tristate
flabel metal2 s 70112 0 70224 800 0 FreeSans 448 90 0 0 mem_rdata[26]
port 100 nsew signal tristate
flabel metal2 s 70784 0 70896 800 0 FreeSans 448 90 0 0 mem_rdata[27]
port 101 nsew signal tristate
flabel metal2 s 71456 0 71568 800 0 FreeSans 448 90 0 0 mem_rdata[28]
port 102 nsew signal tristate
flabel metal2 s 72128 0 72240 800 0 FreeSans 448 90 0 0 mem_rdata[29]
port 103 nsew signal tristate
flabel metal2 s 53984 0 54096 800 0 FreeSans 448 90 0 0 mem_rdata[2]
port 104 nsew signal tristate
flabel metal2 s 72800 0 72912 800 0 FreeSans 448 90 0 0 mem_rdata[30]
port 105 nsew signal tristate
flabel metal2 s 73472 0 73584 800 0 FreeSans 448 90 0 0 mem_rdata[31]
port 106 nsew signal tristate
flabel metal2 s 54656 0 54768 800 0 FreeSans 448 90 0 0 mem_rdata[3]
port 107 nsew signal tristate
flabel metal2 s 55328 0 55440 800 0 FreeSans 448 90 0 0 mem_rdata[4]
port 108 nsew signal tristate
flabel metal2 s 56000 0 56112 800 0 FreeSans 448 90 0 0 mem_rdata[5]
port 109 nsew signal tristate
flabel metal2 s 56672 0 56784 800 0 FreeSans 448 90 0 0 mem_rdata[6]
port 110 nsew signal tristate
flabel metal2 s 57344 0 57456 800 0 FreeSans 448 90 0 0 mem_rdata[7]
port 111 nsew signal tristate
flabel metal2 s 58016 0 58128 800 0 FreeSans 448 90 0 0 mem_rdata[8]
port 112 nsew signal tristate
flabel metal2 s 58688 0 58800 800 0 FreeSans 448 90 0 0 mem_rdata[9]
port 113 nsew signal tristate
flabel metal2 s 49280 0 49392 800 0 FreeSans 448 90 0 0 mem_ready
port 114 nsew signal tristate
flabel metal2 s 47936 0 48048 800 0 FreeSans 448 90 0 0 mem_valid
port 115 nsew signal input
flabel metal2 s 4928 0 5040 800 0 FreeSans 448 90 0 0 mem_wdata[0]
port 116 nsew signal input
flabel metal2 s 11648 0 11760 800 0 FreeSans 448 90 0 0 mem_wdata[10]
port 117 nsew signal input
flabel metal2 s 12320 0 12432 800 0 FreeSans 448 90 0 0 mem_wdata[11]
port 118 nsew signal input
flabel metal2 s 12992 0 13104 800 0 FreeSans 448 90 0 0 mem_wdata[12]
port 119 nsew signal input
flabel metal2 s 13664 0 13776 800 0 FreeSans 448 90 0 0 mem_wdata[13]
port 120 nsew signal input
flabel metal2 s 14336 0 14448 800 0 FreeSans 448 90 0 0 mem_wdata[14]
port 121 nsew signal input
flabel metal2 s 15008 0 15120 800 0 FreeSans 448 90 0 0 mem_wdata[15]
port 122 nsew signal input
flabel metal2 s 15680 0 15792 800 0 FreeSans 448 90 0 0 mem_wdata[16]
port 123 nsew signal input
flabel metal2 s 16352 0 16464 800 0 FreeSans 448 90 0 0 mem_wdata[17]
port 124 nsew signal input
flabel metal2 s 17024 0 17136 800 0 FreeSans 448 90 0 0 mem_wdata[18]
port 125 nsew signal input
flabel metal2 s 17696 0 17808 800 0 FreeSans 448 90 0 0 mem_wdata[19]
port 126 nsew signal input
flabel metal2 s 5600 0 5712 800 0 FreeSans 448 90 0 0 mem_wdata[1]
port 127 nsew signal input
flabel metal2 s 18368 0 18480 800 0 FreeSans 448 90 0 0 mem_wdata[20]
port 128 nsew signal input
flabel metal2 s 19040 0 19152 800 0 FreeSans 448 90 0 0 mem_wdata[21]
port 129 nsew signal input
flabel metal2 s 19712 0 19824 800 0 FreeSans 448 90 0 0 mem_wdata[22]
port 130 nsew signal input
flabel metal2 s 20384 0 20496 800 0 FreeSans 448 90 0 0 mem_wdata[23]
port 131 nsew signal input
flabel metal2 s 21056 0 21168 800 0 FreeSans 448 90 0 0 mem_wdata[24]
port 132 nsew signal input
flabel metal2 s 21728 0 21840 800 0 FreeSans 448 90 0 0 mem_wdata[25]
port 133 nsew signal input
flabel metal2 s 22400 0 22512 800 0 FreeSans 448 90 0 0 mem_wdata[26]
port 134 nsew signal input
flabel metal2 s 23072 0 23184 800 0 FreeSans 448 90 0 0 mem_wdata[27]
port 135 nsew signal input
flabel metal2 s 23744 0 23856 800 0 FreeSans 448 90 0 0 mem_wdata[28]
port 136 nsew signal input
flabel metal2 s 24416 0 24528 800 0 FreeSans 448 90 0 0 mem_wdata[29]
port 137 nsew signal input
flabel metal2 s 6272 0 6384 800 0 FreeSans 448 90 0 0 mem_wdata[2]
port 138 nsew signal input
flabel metal2 s 25088 0 25200 800 0 FreeSans 448 90 0 0 mem_wdata[30]
port 139 nsew signal input
flabel metal2 s 25760 0 25872 800 0 FreeSans 448 90 0 0 mem_wdata[31]
port 140 nsew signal input
flabel metal2 s 6944 0 7056 800 0 FreeSans 448 90 0 0 mem_wdata[3]
port 141 nsew signal input
flabel metal2 s 7616 0 7728 800 0 FreeSans 448 90 0 0 mem_wdata[4]
port 142 nsew signal input
flabel metal2 s 8288 0 8400 800 0 FreeSans 448 90 0 0 mem_wdata[5]
port 143 nsew signal input
flabel metal2 s 8960 0 9072 800 0 FreeSans 448 90 0 0 mem_wdata[6]
port 144 nsew signal input
flabel metal2 s 9632 0 9744 800 0 FreeSans 448 90 0 0 mem_wdata[7]
port 145 nsew signal input
flabel metal2 s 10304 0 10416 800 0 FreeSans 448 90 0 0 mem_wdata[8]
port 146 nsew signal input
flabel metal2 s 10976 0 11088 800 0 FreeSans 448 90 0 0 mem_wdata[9]
port 147 nsew signal input
flabel metal2 s 49952 0 50064 800 0 FreeSans 448 90 0 0 mem_wstrb[0]
port 148 nsew signal input
flabel metal2 s 50624 0 50736 800 0 FreeSans 448 90 0 0 mem_wstrb[1]
port 149 nsew signal input
flabel metal2 s 51296 0 51408 800 0 FreeSans 448 90 0 0 mem_wstrb[2]
port 150 nsew signal input
flabel metal2 s 51968 0 52080 800 0 FreeSans 448 90 0 0 mem_wstrb[3]
port 151 nsew signal input
flabel metal3 s 0 38080 800 38192 0 FreeSans 448 0 0 0 ram_gwenb[0]
port 152 nsew signal tristate
flabel metal3 s 0 39200 800 39312 0 FreeSans 448 0 0 0 ram_gwenb[1]
port 153 nsew signal tristate
flabel metal3 s 0 40320 800 40432 0 FreeSans 448 0 0 0 ram_gwenb[2]
port 154 nsew signal tristate
flabel metal3 s 0 41440 800 41552 0 FreeSans 448 0 0 0 ram_gwenb[3]
port 155 nsew signal tristate
flabel metal3 s 0 2240 800 2352 0 FreeSans 448 0 0 0 ram_rdata[0]
port 156 nsew signal input
flabel metal3 s 0 13440 800 13552 0 FreeSans 448 0 0 0 ram_rdata[10]
port 157 nsew signal input
flabel metal3 s 0 14560 800 14672 0 FreeSans 448 0 0 0 ram_rdata[11]
port 158 nsew signal input
flabel metal3 s 0 15680 800 15792 0 FreeSans 448 0 0 0 ram_rdata[12]
port 159 nsew signal input
flabel metal3 s 0 16800 800 16912 0 FreeSans 448 0 0 0 ram_rdata[13]
port 160 nsew signal input
flabel metal3 s 0 17920 800 18032 0 FreeSans 448 0 0 0 ram_rdata[14]
port 161 nsew signal input
flabel metal3 s 0 19040 800 19152 0 FreeSans 448 0 0 0 ram_rdata[15]
port 162 nsew signal input
flabel metal3 s 0 20160 800 20272 0 FreeSans 448 0 0 0 ram_rdata[16]
port 163 nsew signal input
flabel metal3 s 0 21280 800 21392 0 FreeSans 448 0 0 0 ram_rdata[17]
port 164 nsew signal input
flabel metal3 s 0 22400 800 22512 0 FreeSans 448 0 0 0 ram_rdata[18]
port 165 nsew signal input
flabel metal3 s 0 23520 800 23632 0 FreeSans 448 0 0 0 ram_rdata[19]
port 166 nsew signal input
flabel metal3 s 0 3360 800 3472 0 FreeSans 448 0 0 0 ram_rdata[1]
port 167 nsew signal input
flabel metal3 s 0 24640 800 24752 0 FreeSans 448 0 0 0 ram_rdata[20]
port 168 nsew signal input
flabel metal3 s 0 25760 800 25872 0 FreeSans 448 0 0 0 ram_rdata[21]
port 169 nsew signal input
flabel metal3 s 0 26880 800 26992 0 FreeSans 448 0 0 0 ram_rdata[22]
port 170 nsew signal input
flabel metal3 s 0 28000 800 28112 0 FreeSans 448 0 0 0 ram_rdata[23]
port 171 nsew signal input
flabel metal3 s 0 29120 800 29232 0 FreeSans 448 0 0 0 ram_rdata[24]
port 172 nsew signal input
flabel metal3 s 0 30240 800 30352 0 FreeSans 448 0 0 0 ram_rdata[25]
port 173 nsew signal input
flabel metal3 s 0 31360 800 31472 0 FreeSans 448 0 0 0 ram_rdata[26]
port 174 nsew signal input
flabel metal3 s 0 32480 800 32592 0 FreeSans 448 0 0 0 ram_rdata[27]
port 175 nsew signal input
flabel metal3 s 0 33600 800 33712 0 FreeSans 448 0 0 0 ram_rdata[28]
port 176 nsew signal input
flabel metal3 s 0 34720 800 34832 0 FreeSans 448 0 0 0 ram_rdata[29]
port 177 nsew signal input
flabel metal3 s 0 4480 800 4592 0 FreeSans 448 0 0 0 ram_rdata[2]
port 178 nsew signal input
flabel metal3 s 0 35840 800 35952 0 FreeSans 448 0 0 0 ram_rdata[30]
port 179 nsew signal input
flabel metal3 s 0 36960 800 37072 0 FreeSans 448 0 0 0 ram_rdata[31]
port 180 nsew signal input
flabel metal3 s 0 5600 800 5712 0 FreeSans 448 0 0 0 ram_rdata[3]
port 181 nsew signal input
flabel metal3 s 0 6720 800 6832 0 FreeSans 448 0 0 0 ram_rdata[4]
port 182 nsew signal input
flabel metal3 s 0 7840 800 7952 0 FreeSans 448 0 0 0 ram_rdata[5]
port 183 nsew signal input
flabel metal3 s 0 8960 800 9072 0 FreeSans 448 0 0 0 ram_rdata[6]
port 184 nsew signal input
flabel metal3 s 0 10080 800 10192 0 FreeSans 448 0 0 0 ram_rdata[7]
port 185 nsew signal input
flabel metal3 s 0 11200 800 11312 0 FreeSans 448 0 0 0 ram_rdata[8]
port 186 nsew signal input
flabel metal3 s 0 12320 800 12432 0 FreeSans 448 0 0 0 ram_rdata[9]
port 187 nsew signal input
flabel metal3 s 0 42560 800 42672 0 FreeSans 448 0 0 0 ram_wenb[0]
port 188 nsew signal tristate
flabel metal3 s 0 53760 800 53872 0 FreeSans 448 0 0 0 ram_wenb[10]
port 189 nsew signal tristate
flabel metal3 s 0 54880 800 54992 0 FreeSans 448 0 0 0 ram_wenb[11]
port 190 nsew signal tristate
flabel metal3 s 0 56000 800 56112 0 FreeSans 448 0 0 0 ram_wenb[12]
port 191 nsew signal tristate
flabel metal3 s 0 57120 800 57232 0 FreeSans 448 0 0 0 ram_wenb[13]
port 192 nsew signal tristate
flabel metal3 s 0 58240 800 58352 0 FreeSans 448 0 0 0 ram_wenb[14]
port 193 nsew signal tristate
flabel metal3 s 0 59360 800 59472 0 FreeSans 448 0 0 0 ram_wenb[15]
port 194 nsew signal tristate
flabel metal3 s 0 60480 800 60592 0 FreeSans 448 0 0 0 ram_wenb[16]
port 195 nsew signal tristate
flabel metal3 s 0 61600 800 61712 0 FreeSans 448 0 0 0 ram_wenb[17]
port 196 nsew signal tristate
flabel metal3 s 0 62720 800 62832 0 FreeSans 448 0 0 0 ram_wenb[18]
port 197 nsew signal tristate
flabel metal3 s 0 63840 800 63952 0 FreeSans 448 0 0 0 ram_wenb[19]
port 198 nsew signal tristate
flabel metal3 s 0 43680 800 43792 0 FreeSans 448 0 0 0 ram_wenb[1]
port 199 nsew signal tristate
flabel metal3 s 0 64960 800 65072 0 FreeSans 448 0 0 0 ram_wenb[20]
port 200 nsew signal tristate
flabel metal3 s 0 66080 800 66192 0 FreeSans 448 0 0 0 ram_wenb[21]
port 201 nsew signal tristate
flabel metal3 s 0 67200 800 67312 0 FreeSans 448 0 0 0 ram_wenb[22]
port 202 nsew signal tristate
flabel metal3 s 0 68320 800 68432 0 FreeSans 448 0 0 0 ram_wenb[23]
port 203 nsew signal tristate
flabel metal3 s 0 69440 800 69552 0 FreeSans 448 0 0 0 ram_wenb[24]
port 204 nsew signal tristate
flabel metal3 s 0 70560 800 70672 0 FreeSans 448 0 0 0 ram_wenb[25]
port 205 nsew signal tristate
flabel metal3 s 0 71680 800 71792 0 FreeSans 448 0 0 0 ram_wenb[26]
port 206 nsew signal tristate
flabel metal3 s 0 72800 800 72912 0 FreeSans 448 0 0 0 ram_wenb[27]
port 207 nsew signal tristate
flabel metal3 s 0 73920 800 74032 0 FreeSans 448 0 0 0 ram_wenb[28]
port 208 nsew signal tristate
flabel metal3 s 0 75040 800 75152 0 FreeSans 448 0 0 0 ram_wenb[29]
port 209 nsew signal tristate
flabel metal3 s 0 44800 800 44912 0 FreeSans 448 0 0 0 ram_wenb[2]
port 210 nsew signal tristate
flabel metal3 s 0 76160 800 76272 0 FreeSans 448 0 0 0 ram_wenb[30]
port 211 nsew signal tristate
flabel metal3 s 0 77280 800 77392 0 FreeSans 448 0 0 0 ram_wenb[31]
port 212 nsew signal tristate
flabel metal3 s 0 45920 800 46032 0 FreeSans 448 0 0 0 ram_wenb[3]
port 213 nsew signal tristate
flabel metal3 s 0 47040 800 47152 0 FreeSans 448 0 0 0 ram_wenb[4]
port 214 nsew signal tristate
flabel metal3 s 0 48160 800 48272 0 FreeSans 448 0 0 0 ram_wenb[5]
port 215 nsew signal tristate
flabel metal3 s 0 49280 800 49392 0 FreeSans 448 0 0 0 ram_wenb[6]
port 216 nsew signal tristate
flabel metal3 s 0 50400 800 50512 0 FreeSans 448 0 0 0 ram_wenb[7]
port 217 nsew signal tristate
flabel metal3 s 0 51520 800 51632 0 FreeSans 448 0 0 0 ram_wenb[8]
port 218 nsew signal tristate
flabel metal3 s 0 52640 800 52752 0 FreeSans 448 0 0 0 ram_wenb[9]
port 219 nsew signal tristate
flabel metal2 s 74816 0 74928 800 0 FreeSans 448 90 0 0 resetn
port 220 nsew signal input
flabel metal3 s 79200 42112 80000 42224 0 FreeSans 448 0 0 0 simpleuart_dat_re
port 221 nsew signal tristate
flabel metal3 s 79200 40992 80000 41104 0 FreeSans 448 0 0 0 simpleuart_dat_we
port 222 nsew signal tristate
flabel metal3 s 79200 672 80000 784 0 FreeSans 448 0 0 0 simpleuart_div_we[0]
port 223 nsew signal tristate
flabel metal3 s 79200 1792 80000 1904 0 FreeSans 448 0 0 0 simpleuart_div_we[1]
port 224 nsew signal tristate
flabel metal3 s 79200 2912 80000 3024 0 FreeSans 448 0 0 0 simpleuart_div_we[2]
port 225 nsew signal tristate
flabel metal3 s 79200 4032 80000 4144 0 FreeSans 448 0 0 0 simpleuart_div_we[3]
port 226 nsew signal tristate
flabel metal3 s 79200 43232 80000 43344 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[0]
port 227 nsew signal input
flabel metal3 s 79200 54432 80000 54544 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[10]
port 228 nsew signal input
flabel metal3 s 79200 55552 80000 55664 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[11]
port 229 nsew signal input
flabel metal3 s 79200 56672 80000 56784 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[12]
port 230 nsew signal input
flabel metal3 s 79200 57792 80000 57904 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[13]
port 231 nsew signal input
flabel metal3 s 79200 58912 80000 59024 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[14]
port 232 nsew signal input
flabel metal3 s 79200 60032 80000 60144 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[15]
port 233 nsew signal input
flabel metal3 s 79200 61152 80000 61264 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[16]
port 234 nsew signal input
flabel metal3 s 79200 62272 80000 62384 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[17]
port 235 nsew signal input
flabel metal3 s 79200 63392 80000 63504 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[18]
port 236 nsew signal input
flabel metal3 s 79200 64512 80000 64624 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[19]
port 237 nsew signal input
flabel metal3 s 79200 44352 80000 44464 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[1]
port 238 nsew signal input
flabel metal3 s 79200 65632 80000 65744 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[20]
port 239 nsew signal input
flabel metal3 s 79200 66752 80000 66864 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[21]
port 240 nsew signal input
flabel metal3 s 79200 67872 80000 67984 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[22]
port 241 nsew signal input
flabel metal3 s 79200 68992 80000 69104 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[23]
port 242 nsew signal input
flabel metal3 s 79200 70112 80000 70224 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[24]
port 243 nsew signal input
flabel metal3 s 79200 71232 80000 71344 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[25]
port 244 nsew signal input
flabel metal3 s 79200 72352 80000 72464 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[26]
port 245 nsew signal input
flabel metal3 s 79200 73472 80000 73584 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[27]
port 246 nsew signal input
flabel metal3 s 79200 74592 80000 74704 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[28]
port 247 nsew signal input
flabel metal3 s 79200 75712 80000 75824 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[29]
port 248 nsew signal input
flabel metal3 s 79200 45472 80000 45584 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[2]
port 249 nsew signal input
flabel metal3 s 79200 76832 80000 76944 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[30]
port 250 nsew signal input
flabel metal3 s 79200 77952 80000 78064 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[31]
port 251 nsew signal input
flabel metal3 s 79200 46592 80000 46704 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[3]
port 252 nsew signal input
flabel metal3 s 79200 47712 80000 47824 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[4]
port 253 nsew signal input
flabel metal3 s 79200 48832 80000 48944 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[5]
port 254 nsew signal input
flabel metal3 s 79200 49952 80000 50064 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[6]
port 255 nsew signal input
flabel metal3 s 79200 51072 80000 51184 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[7]
port 256 nsew signal input
flabel metal3 s 79200 52192 80000 52304 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[8]
port 257 nsew signal input
flabel metal3 s 79200 53312 80000 53424 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[9]
port 258 nsew signal input
flabel metal3 s 79200 79072 80000 79184 0 FreeSans 448 0 0 0 simpleuart_reg_dat_wait
port 259 nsew signal input
flabel metal3 s 79200 5152 80000 5264 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[0]
port 260 nsew signal input
flabel metal3 s 79200 16352 80000 16464 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[10]
port 261 nsew signal input
flabel metal3 s 79200 17472 80000 17584 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[11]
port 262 nsew signal input
flabel metal3 s 79200 18592 80000 18704 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[12]
port 263 nsew signal input
flabel metal3 s 79200 19712 80000 19824 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[13]
port 264 nsew signal input
flabel metal3 s 79200 20832 80000 20944 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[14]
port 265 nsew signal input
flabel metal3 s 79200 21952 80000 22064 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[15]
port 266 nsew signal input
flabel metal3 s 79200 23072 80000 23184 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[16]
port 267 nsew signal input
flabel metal3 s 79200 24192 80000 24304 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[17]
port 268 nsew signal input
flabel metal3 s 79200 25312 80000 25424 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[18]
port 269 nsew signal input
flabel metal3 s 79200 26432 80000 26544 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[19]
port 270 nsew signal input
flabel metal3 s 79200 6272 80000 6384 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[1]
port 271 nsew signal input
flabel metal3 s 79200 27552 80000 27664 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[20]
port 272 nsew signal input
flabel metal3 s 79200 28672 80000 28784 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[21]
port 273 nsew signal input
flabel metal3 s 79200 29792 80000 29904 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[22]
port 274 nsew signal input
flabel metal3 s 79200 30912 80000 31024 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[23]
port 275 nsew signal input
flabel metal3 s 79200 32032 80000 32144 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[24]
port 276 nsew signal input
flabel metal3 s 79200 33152 80000 33264 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[25]
port 277 nsew signal input
flabel metal3 s 79200 34272 80000 34384 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[26]
port 278 nsew signal input
flabel metal3 s 79200 35392 80000 35504 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[27]
port 279 nsew signal input
flabel metal3 s 79200 36512 80000 36624 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[28]
port 280 nsew signal input
flabel metal3 s 79200 37632 80000 37744 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[29]
port 281 nsew signal input
flabel metal3 s 79200 7392 80000 7504 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[2]
port 282 nsew signal input
flabel metal3 s 79200 38752 80000 38864 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[30]
port 283 nsew signal input
flabel metal3 s 79200 39872 80000 39984 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[31]
port 284 nsew signal input
flabel metal3 s 79200 8512 80000 8624 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[3]
port 285 nsew signal input
flabel metal3 s 79200 9632 80000 9744 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[4]
port 286 nsew signal input
flabel metal3 s 79200 10752 80000 10864 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[5]
port 287 nsew signal input
flabel metal3 s 79200 11872 80000 11984 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[6]
port 288 nsew signal input
flabel metal3 s 79200 12992 80000 13104 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[7]
port 289 nsew signal input
flabel metal3 s 79200 14112 80000 14224 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[8]
port 290 nsew signal input
flabel metal3 s 79200 15232 80000 15344 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[9]
port 291 nsew signal input
flabel metal2 s 34048 79200 34160 80000 0 FreeSans 448 90 0 0 spimem_rdata[0]
port 292 nsew signal input
flabel metal2 s 40768 79200 40880 80000 0 FreeSans 448 90 0 0 spimem_rdata[10]
port 293 nsew signal input
flabel metal2 s 41440 79200 41552 80000 0 FreeSans 448 90 0 0 spimem_rdata[11]
port 294 nsew signal input
flabel metal2 s 42112 79200 42224 80000 0 FreeSans 448 90 0 0 spimem_rdata[12]
port 295 nsew signal input
flabel metal2 s 42784 79200 42896 80000 0 FreeSans 448 90 0 0 spimem_rdata[13]
port 296 nsew signal input
flabel metal2 s 43456 79200 43568 80000 0 FreeSans 448 90 0 0 spimem_rdata[14]
port 297 nsew signal input
flabel metal2 s 44128 79200 44240 80000 0 FreeSans 448 90 0 0 spimem_rdata[15]
port 298 nsew signal input
flabel metal2 s 44800 79200 44912 80000 0 FreeSans 448 90 0 0 spimem_rdata[16]
port 299 nsew signal input
flabel metal2 s 45472 79200 45584 80000 0 FreeSans 448 90 0 0 spimem_rdata[17]
port 300 nsew signal input
flabel metal2 s 46144 79200 46256 80000 0 FreeSans 448 90 0 0 spimem_rdata[18]
port 301 nsew signal input
flabel metal2 s 46816 79200 46928 80000 0 FreeSans 448 90 0 0 spimem_rdata[19]
port 302 nsew signal input
flabel metal2 s 34720 79200 34832 80000 0 FreeSans 448 90 0 0 spimem_rdata[1]
port 303 nsew signal input
flabel metal2 s 47488 79200 47600 80000 0 FreeSans 448 90 0 0 spimem_rdata[20]
port 304 nsew signal input
flabel metal2 s 48160 79200 48272 80000 0 FreeSans 448 90 0 0 spimem_rdata[21]
port 305 nsew signal input
flabel metal2 s 48832 79200 48944 80000 0 FreeSans 448 90 0 0 spimem_rdata[22]
port 306 nsew signal input
flabel metal2 s 49504 79200 49616 80000 0 FreeSans 448 90 0 0 spimem_rdata[23]
port 307 nsew signal input
flabel metal2 s 50176 79200 50288 80000 0 FreeSans 448 90 0 0 spimem_rdata[24]
port 308 nsew signal input
flabel metal2 s 50848 79200 50960 80000 0 FreeSans 448 90 0 0 spimem_rdata[25]
port 309 nsew signal input
flabel metal2 s 51520 79200 51632 80000 0 FreeSans 448 90 0 0 spimem_rdata[26]
port 310 nsew signal input
flabel metal2 s 52192 79200 52304 80000 0 FreeSans 448 90 0 0 spimem_rdata[27]
port 311 nsew signal input
flabel metal2 s 52864 79200 52976 80000 0 FreeSans 448 90 0 0 spimem_rdata[28]
port 312 nsew signal input
flabel metal2 s 53536 79200 53648 80000 0 FreeSans 448 90 0 0 spimem_rdata[29]
port 313 nsew signal input
flabel metal2 s 35392 79200 35504 80000 0 FreeSans 448 90 0 0 spimem_rdata[2]
port 314 nsew signal input
flabel metal2 s 54208 79200 54320 80000 0 FreeSans 448 90 0 0 spimem_rdata[30]
port 315 nsew signal input
flabel metal2 s 54880 79200 54992 80000 0 FreeSans 448 90 0 0 spimem_rdata[31]
port 316 nsew signal input
flabel metal2 s 36064 79200 36176 80000 0 FreeSans 448 90 0 0 spimem_rdata[3]
port 317 nsew signal input
flabel metal2 s 36736 79200 36848 80000 0 FreeSans 448 90 0 0 spimem_rdata[4]
port 318 nsew signal input
flabel metal2 s 37408 79200 37520 80000 0 FreeSans 448 90 0 0 spimem_rdata[5]
port 319 nsew signal input
flabel metal2 s 38080 79200 38192 80000 0 FreeSans 448 90 0 0 spimem_rdata[6]
port 320 nsew signal input
flabel metal2 s 38752 79200 38864 80000 0 FreeSans 448 90 0 0 spimem_rdata[7]
port 321 nsew signal input
flabel metal2 s 39424 79200 39536 80000 0 FreeSans 448 90 0 0 spimem_rdata[8]
port 322 nsew signal input
flabel metal2 s 40096 79200 40208 80000 0 FreeSans 448 90 0 0 spimem_rdata[9]
port 323 nsew signal input
flabel metal2 s 32704 79200 32816 80000 0 FreeSans 448 90 0 0 spimem_ready
port 324 nsew signal input
flabel metal2 s 33376 79200 33488 80000 0 FreeSans 448 90 0 0 spimem_valid
port 325 nsew signal tristate
flabel metal2 s 58240 79200 58352 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[0]
port 326 nsew signal input
flabel metal2 s 64960 79200 65072 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[10]
port 327 nsew signal input
flabel metal2 s 65632 79200 65744 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[11]
port 328 nsew signal input
flabel metal2 s 66304 79200 66416 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[12]
port 329 nsew signal input
flabel metal2 s 66976 79200 67088 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[13]
port 330 nsew signal input
flabel metal2 s 67648 79200 67760 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[14]
port 331 nsew signal input
flabel metal2 s 68320 79200 68432 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[15]
port 332 nsew signal input
flabel metal2 s 68992 79200 69104 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[16]
port 333 nsew signal input
flabel metal2 s 69664 79200 69776 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[17]
port 334 nsew signal input
flabel metal2 s 70336 79200 70448 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[18]
port 335 nsew signal input
flabel metal2 s 71008 79200 71120 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[19]
port 336 nsew signal input
flabel metal2 s 58912 79200 59024 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[1]
port 337 nsew signal input
flabel metal2 s 71680 79200 71792 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[20]
port 338 nsew signal input
flabel metal2 s 72352 79200 72464 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[21]
port 339 nsew signal input
flabel metal2 s 73024 79200 73136 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[22]
port 340 nsew signal input
flabel metal2 s 73696 79200 73808 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[23]
port 341 nsew signal input
flabel metal2 s 74368 79200 74480 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[24]
port 342 nsew signal input
flabel metal2 s 75040 79200 75152 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[25]
port 343 nsew signal input
flabel metal2 s 75712 79200 75824 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[26]
port 344 nsew signal input
flabel metal2 s 76384 79200 76496 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[27]
port 345 nsew signal input
flabel metal2 s 77056 79200 77168 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[28]
port 346 nsew signal input
flabel metal2 s 77728 79200 77840 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[29]
port 347 nsew signal input
flabel metal2 s 59584 79200 59696 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[2]
port 348 nsew signal input
flabel metal2 s 78400 79200 78512 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[30]
port 349 nsew signal input
flabel metal2 s 79072 79200 79184 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[31]
port 350 nsew signal input
flabel metal2 s 60256 79200 60368 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[3]
port 351 nsew signal input
flabel metal2 s 60928 79200 61040 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[4]
port 352 nsew signal input
flabel metal2 s 61600 79200 61712 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[5]
port 353 nsew signal input
flabel metal2 s 62272 79200 62384 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[6]
port 354 nsew signal input
flabel metal2 s 62944 79200 63056 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[7]
port 355 nsew signal input
flabel metal2 s 63616 79200 63728 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[8]
port 356 nsew signal input
flabel metal2 s 64288 79200 64400 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[9]
port 357 nsew signal input
flabel metal2 s 55552 79200 55664 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_we[0]
port 358 nsew signal tristate
flabel metal2 s 56224 79200 56336 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_we[1]
port 359 nsew signal tristate
flabel metal2 s 56896 79200 57008 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_we[2]
port 360 nsew signal tristate
flabel metal2 s 57568 79200 57680 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_we[3]
port 361 nsew signal tristate
flabel metal4 s 4448 3076 4768 76892 0 FreeSans 1280 90 0 0 vdd
port 362 nsew power bidirectional
flabel metal4 s 35168 3076 35488 76892 0 FreeSans 1280 90 0 0 vdd
port 362 nsew power bidirectional
flabel metal4 s 65888 3076 66208 76892 0 FreeSans 1280 90 0 0 vdd
port 362 nsew power bidirectional
flabel metal4 s 19808 3076 20128 76892 0 FreeSans 1280 90 0 0 vss
port 363 nsew ground bidirectional
flabel metal4 s 50528 3076 50848 76892 0 FreeSans 1280 90 0 0 vss
port 363 nsew ground bidirectional
rlabel metal1 39984 76048 39984 76048 0 vdd
rlabel metal1 39984 76832 39984 76832 0 vss
rlabel metal3 41720 38808 41720 38808 0 _0000_
rlabel metal2 16184 10248 16184 10248 0 _0001_
rlabel metal2 15400 8624 15400 8624 0 _0002_
rlabel metal2 15736 7056 15736 7056 0 _0003_
rlabel metal3 17080 5208 17080 5208 0 _0004_
rlabel metal2 17640 12432 17640 12432 0 _0005_
rlabel metal2 20496 12040 20496 12040 0 _0006_
rlabel metal3 18928 10472 18928 10472 0 _0007_
rlabel metal2 19152 8344 19152 8344 0 _0008_
rlabel metal3 23912 4200 23912 4200 0 _0009_
rlabel metal2 23688 5320 23688 5320 0 _0010_
rlabel metal2 23464 6944 23464 6944 0 _0011_
rlabel metal2 27608 8624 27608 8624 0 _0012_
rlabel metal2 22400 8344 22400 8344 0 _0013_
rlabel metal3 25536 11256 25536 11256 0 _0014_
rlabel metal2 22344 11760 22344 11760 0 _0015_
rlabel metal2 23688 13328 23688 13328 0 _0016_
rlabel metal2 30184 8624 30184 8624 0 _0017_
rlabel metal2 33208 10416 33208 10416 0 _0018_
rlabel metal2 29960 11760 29960 11760 0 _0019_
rlabel metal2 29176 10248 29176 10248 0 _0020_
rlabel metal3 34160 8904 34160 8904 0 _0021_
rlabel metal2 30856 5544 30856 5544 0 _0022_
rlabel metal2 30408 6104 30408 6104 0 _0023_
rlabel metal2 35168 7560 35168 7560 0 _0024_
rlabel metal3 28560 23016 28560 23016 0 _0025_
rlabel metal2 24808 24304 24808 24304 0 _0026_
rlabel metal2 27888 24024 27888 24024 0 _0027_
rlabel metal2 26488 22008 26488 22008 0 _0028_
rlabel metal2 17528 23576 17528 23576 0 _0029_
rlabel metal2 21448 24472 21448 24472 0 _0030_
rlabel metal2 17864 22008 17864 22008 0 _0031_
rlabel metal2 21952 22456 21952 22456 0 _0032_
rlabel metal2 19544 21168 19544 21168 0 _0033_
rlabel metal2 19320 17024 19320 17024 0 _0034_
rlabel metal2 22568 17472 22568 17472 0 _0035_
rlabel metal2 22680 19600 22680 19600 0 _0036_
rlabel metal2 27496 19600 27496 19600 0 _0037_
rlabel metal2 29960 18536 29960 18536 0 _0038_
rlabel metal2 30408 19600 30408 19600 0 _0039_
rlabel metal2 29848 21168 29848 21168 0 _0040_
rlabel metal2 36008 14896 36008 14896 0 _0041_
rlabel metal2 35896 13328 35896 13328 0 _0042_
rlabel metal2 33544 14168 33544 14168 0 _0043_
rlabel metal2 33544 15568 33544 15568 0 _0044_
rlabel metal2 26712 17696 26712 17696 0 _0045_
rlabel metal2 29288 16464 29288 16464 0 _0046_
rlabel metal2 25816 15540 25816 15540 0 _0047_
rlabel metal2 29232 13832 29232 13832 0 _0048_
rlabel metal2 39928 13104 39928 13104 0 _0049_
rlabel metal2 42896 13048 42896 13048 0 _0050_
rlabel metal2 42504 15148 42504 15148 0 _0051_
rlabel metal2 40264 15148 40264 15148 0 _0052_
rlabel metal2 39704 11088 39704 11088 0 _0053_
rlabel metal2 42504 10192 42504 10192 0 _0054_
rlabel metal2 38248 8456 38248 8456 0 _0055_
rlabel metal2 42616 9240 42616 9240 0 _0056_
rlabel metal2 37968 6776 37968 6776 0 _0057_
rlabel metal3 9632 8904 9632 8904 0 _0058_
rlabel metal3 8736 9688 8736 9688 0 _0059_
rlabel metal2 9464 11760 9464 11760 0 _0060_
rlabel metal2 13384 11088 13384 11088 0 _0061_
rlabel metal2 10920 7728 10920 7728 0 _0062_
rlabel metal2 10696 5488 10696 5488 0 _0063_
rlabel metal3 9632 4200 9632 4200 0 _0064_
rlabel metal3 13216 4200 13216 4200 0 _0065_
rlabel metal3 32312 6776 32312 6776 0 _0066_
rlabel metal2 31864 7560 31864 7560 0 _0067_
rlabel metal3 34496 7672 34496 7672 0 _0068_
rlabel metal2 25928 17976 25928 17976 0 _0069_
rlabel metal2 21784 19656 21784 19656 0 _0070_
rlabel metal2 26152 24024 26152 24024 0 _0071_
rlabel metal2 19320 21168 19320 21168 0 _0072_
rlabel metal2 24360 23296 24360 23296 0 _0073_
rlabel metal3 26488 23128 26488 23128 0 _0074_
rlabel metal2 24696 23576 24696 23576 0 _0075_
rlabel metal3 25480 23688 25480 23688 0 _0076_
rlabel metal2 25760 21560 25760 21560 0 _0077_
rlabel metal2 17976 22288 17976 22288 0 _0078_
rlabel metal2 17416 24136 17416 24136 0 _0079_
rlabel metal2 17808 23352 17808 23352 0 _0080_
rlabel metal2 21896 24192 21896 24192 0 _0081_
rlabel metal3 16688 21784 16688 21784 0 _0082_
rlabel metal2 20384 23128 20384 23128 0 _0083_
rlabel metal2 19992 18144 19992 18144 0 _0084_
rlabel metal3 19264 19992 19264 19992 0 _0085_
rlabel metal2 20048 20216 20048 20216 0 _0086_
rlabel metal2 19544 17472 19544 17472 0 _0087_
rlabel metal2 19208 17920 19208 17920 0 _0088_
rlabel metal2 22120 19488 22120 19488 0 _0089_
rlabel metal2 27608 19880 27608 19880 0 _0090_
rlabel metal3 25368 19096 25368 19096 0 _0091_
rlabel metal2 26152 19880 26152 19880 0 _0092_
rlabel metal3 28056 18984 28056 18984 0 _0093_
rlabel metal3 24136 18928 24136 18928 0 _0094_
rlabel metal3 27552 20552 27552 20552 0 _0095_
rlabel metal2 29512 13552 29512 13552 0 _0096_
rlabel metal3 34216 13832 34216 13832 0 _0097_
rlabel metal2 28280 12600 28280 12600 0 _0098_
rlabel metal2 32928 12936 32928 12936 0 _0099_
rlabel metal2 33992 13832 33992 13832 0 _0100_
rlabel metal3 35112 12936 35112 12936 0 _0101_
rlabel metal2 33096 13440 33096 13440 0 _0102_
rlabel metal2 32984 15204 32984 15204 0 _0103_
rlabel metal2 26712 15288 26712 15288 0 _0104_
rlabel metal2 26432 13720 26432 13720 0 _0105_
rlabel metal2 27048 15456 27048 15456 0 _0106_
rlabel metal3 28896 15848 28896 15848 0 _0107_
rlabel metal2 25928 14224 25928 14224 0 _0108_
rlabel metal2 29624 13888 29624 13888 0 _0109_
rlabel metal2 42504 14112 42504 14112 0 _0110_
rlabel metal2 37632 11256 37632 11256 0 _0111_
rlabel metal2 39592 13104 39592 13104 0 _0112_
rlabel metal2 36232 12656 36232 12656 0 _0113_
rlabel metal2 37240 13384 37240 13384 0 _0114_
rlabel metal2 39704 14616 39704 14616 0 _0115_
rlabel metal2 39816 11200 39816 11200 0 _0116_
rlabel metal2 38696 10192 38696 10192 0 _0117_
rlabel metal2 39032 10640 39032 10640 0 _0118_
rlabel metal3 40096 9576 40096 9576 0 _0119_
rlabel metal2 39144 8848 39144 8848 0 _0120_
rlabel metal2 43400 9520 43400 9520 0 _0121_
rlabel metal2 38136 7952 38136 7952 0 _0122_
rlabel metal2 9016 6216 9016 6216 0 _0123_
rlabel metal3 8792 6888 8792 6888 0 _0124_
rlabel metal2 9352 7952 9352 7952 0 _0125_
rlabel metal3 21112 9520 21112 9520 0 _0126_
rlabel metal3 13832 9576 13832 9576 0 _0127_
rlabel metal2 11928 10864 11928 10864 0 _0128_
rlabel metal3 10584 8792 10584 8792 0 _0129_
rlabel metal2 8008 8176 8008 8176 0 _0130_
rlabel metal2 8232 10248 8232 10248 0 _0131_
rlabel metal2 8792 7784 8792 7784 0 _0132_
rlabel metal3 10584 11256 10584 11256 0 _0133_
rlabel metal2 8512 7672 8512 7672 0 _0134_
rlabel metal2 13664 9912 13664 9912 0 _0135_
rlabel metal3 6664 4088 6664 4088 0 _0136_
rlabel metal2 6776 4480 6776 4480 0 _0137_
rlabel metal2 13496 6664 13496 6664 0 _0138_
rlabel metal3 13440 6440 13440 6440 0 _0139_
rlabel metal3 12376 7336 12376 7336 0 _0140_
rlabel metal2 6272 4536 6272 4536 0 _0141_
rlabel metal2 10808 6048 10808 6048 0 _0142_
rlabel metal2 8008 4480 8008 4480 0 _0143_
rlabel metal2 8344 4816 8344 4816 0 _0144_
rlabel metal3 10304 5096 10304 5096 0 _0145_
rlabel metal2 12040 5544 12040 5544 0 _0146_
rlabel metal2 47320 5040 47320 5040 0 _0147_
rlabel metal2 47096 6160 47096 6160 0 _0148_
rlabel metal3 43736 5992 43736 5992 0 _0149_
rlabel metal2 40936 5544 40936 5544 0 _0150_
rlabel metal2 43064 3472 43064 3472 0 _0151_
rlabel metal2 42280 3472 42280 3472 0 _0152_
rlabel metal2 46424 5488 46424 5488 0 _0153_
rlabel metal2 43736 4032 43736 4032 0 _0154_
rlabel metal2 33992 4592 33992 4592 0 _0155_
rlabel metal2 34216 4480 34216 4480 0 _0156_
rlabel metal2 42504 3276 42504 3276 0 _0157_
rlabel metal2 39648 5992 39648 5992 0 _0158_
rlabel metal2 36792 4536 36792 4536 0 _0159_
rlabel metal2 39368 3808 39368 3808 0 _0160_
rlabel metal2 44968 16968 44968 16968 0 _0161_
rlabel metal3 44352 18312 44352 18312 0 _0162_
rlabel metal2 40936 7616 40936 7616 0 _0163_
rlabel metal2 39536 5096 39536 5096 0 _0164_
rlabel metal2 41608 5264 41608 5264 0 _0165_
rlabel metal2 44016 18536 44016 18536 0 _0166_
rlabel metal2 42616 4648 42616 4648 0 _0167_
rlabel metal2 46760 17304 46760 17304 0 _0168_
rlabel metal2 43680 8120 43680 8120 0 _0169_
rlabel metal2 42504 8008 42504 8008 0 _0170_
rlabel metal3 43904 8232 43904 8232 0 _0171_
rlabel metal2 43120 8008 43120 8008 0 _0172_
rlabel metal2 44296 17752 44296 17752 0 _0173_
rlabel metal2 41608 7392 41608 7392 0 _0174_
rlabel metal2 39760 8008 39760 8008 0 _0175_
rlabel metal2 43064 7168 43064 7168 0 _0176_
rlabel metal2 42504 23688 42504 23688 0 _0177_
rlabel metal2 71232 18648 71232 18648 0 _0178_
rlabel metal3 73752 38864 73752 38864 0 _0179_
rlabel metal3 74760 41272 74760 41272 0 _0180_
rlabel metal2 74984 6608 74984 6608 0 _0181_
rlabel metal2 77056 6664 77056 6664 0 _0182_
rlabel metal2 76216 7448 76216 7448 0 _0183_
rlabel metal2 71736 41440 71736 41440 0 _0184_
rlabel metal2 74816 41384 74816 41384 0 _0185_
rlabel metal2 41720 8512 41720 8512 0 _0186_
rlabel metal2 55048 41832 55048 41832 0 _0187_
rlabel metal2 60648 41888 60648 41888 0 _0188_
rlabel metal2 60536 40768 60536 40768 0 _0189_
rlabel metal2 55384 41552 55384 41552 0 _0190_
rlabel metal2 55720 42448 55720 42448 0 _0191_
rlabel metal2 55944 41776 55944 41776 0 _0192_
rlabel metal2 56672 42168 56672 42168 0 _0193_
rlabel metal2 57568 42168 57568 42168 0 _0194_
rlabel metal3 72800 38808 72800 38808 0 _0195_
rlabel metal2 72912 38920 72912 38920 0 _0196_
rlabel metal2 75376 26264 75376 26264 0 _0197_
rlabel metal2 77448 6664 77448 6664 0 _0198_
rlabel metal3 75992 11368 75992 11368 0 _0199_
rlabel metal2 77896 5768 77896 5768 0 _0200_
rlabel metal2 77448 5768 77448 5768 0 _0201_
rlabel metal2 76552 5768 76552 5768 0 _0202_
rlabel metal3 29792 23128 29792 23128 0 _0203_
rlabel metal2 43400 23240 43400 23240 0 _0204_
rlabel metal2 41384 21224 41384 21224 0 _0205_
rlabel metal2 37352 21896 37352 21896 0 _0206_
rlabel metal2 74144 26264 74144 26264 0 _0207_
rlabel metal2 76888 23240 76888 23240 0 _0208_
rlabel metal2 75656 23520 75656 23520 0 _0209_
rlabel metal2 74760 26208 74760 26208 0 _0210_
rlabel metal3 54208 38920 54208 38920 0 _0211_
rlabel metal2 64680 39200 64680 39200 0 _0212_
rlabel metal2 61712 40376 61712 40376 0 _0213_
rlabel metal2 58856 36456 58856 36456 0 _0214_
rlabel metal2 36344 25312 36344 25312 0 _0215_
rlabel metal2 34664 19768 34664 19768 0 _0216_
rlabel metal3 35728 21560 35728 21560 0 _0217_
rlabel metal2 33992 19544 33992 19544 0 _0218_
rlabel metal2 40376 24472 40376 24472 0 _0219_
rlabel metal3 40320 20552 40320 20552 0 _0220_
rlabel metal2 35672 21168 35672 21168 0 _0221_
rlabel metal2 35056 20104 35056 20104 0 _0222_
rlabel metal2 36568 23408 36568 23408 0 _0223_
rlabel metal2 41384 25984 41384 25984 0 _0224_
rlabel metal2 36456 27440 36456 27440 0 _0225_
rlabel metal2 40488 25536 40488 25536 0 _0226_
rlabel metal2 35560 27440 35560 27440 0 _0227_
rlabel metal2 36008 25424 36008 25424 0 _0228_
rlabel metal2 26600 25312 26600 25312 0 _0229_
rlabel metal2 74480 35560 74480 35560 0 _0230_
rlabel metal3 74928 24024 74928 24024 0 _0231_
rlabel metal2 60648 38808 60648 38808 0 _0232_
rlabel metal2 35784 23968 35784 23968 0 _0233_
rlabel metal2 33432 20888 33432 20888 0 _0234_
rlabel metal2 35168 21672 35168 21672 0 _0235_
rlabel metal2 36064 23912 36064 23912 0 _0236_
rlabel metal2 34888 26600 34888 26600 0 _0237_
rlabel metal3 34160 24584 34160 24584 0 _0238_
rlabel metal2 73304 35336 73304 35336 0 _0239_
rlabel metal2 73752 33488 73752 33488 0 _0240_
rlabel metal2 75768 23688 75768 23688 0 _0241_
rlabel metal2 60088 31920 60088 31920 0 _0242_
rlabel metal2 35336 24752 35336 24752 0 _0243_
rlabel metal2 34328 20440 34328 20440 0 _0244_
rlabel metal2 34552 21560 34552 21560 0 _0245_
rlabel metal3 35784 24808 35784 24808 0 _0246_
rlabel metal2 36120 27300 36120 27300 0 _0247_
rlabel metal2 26712 20832 26712 20832 0 _0248_
rlabel metal3 71680 34776 71680 34776 0 _0249_
rlabel metal3 72296 25256 72296 25256 0 _0250_
rlabel metal2 73528 24640 73528 24640 0 _0251_
rlabel metal2 62552 41104 62552 41104 0 _0252_
rlabel metal2 71736 25032 71736 25032 0 _0253_
rlabel metal2 68936 23016 68936 23016 0 _0254_
rlabel metal2 33880 20552 33880 20552 0 _0255_
rlabel metal2 35336 20944 35336 20944 0 _0256_
rlabel metal2 35000 21952 35000 21952 0 _0257_
rlabel metal2 35952 23464 35952 23464 0 _0258_
rlabel metal2 20328 23632 20328 23632 0 _0259_
rlabel metal3 40096 23240 40096 23240 0 _0260_
rlabel metal2 63448 23968 63448 23968 0 _0261_
rlabel metal2 77336 23240 77336 23240 0 _0262_
rlabel metal2 63672 22736 63672 22736 0 _0263_
rlabel metal2 63560 40656 63560 40656 0 _0264_
rlabel metal2 62608 40152 62608 40152 0 _0265_
rlabel metal2 63560 24136 63560 24136 0 _0266_
rlabel metal3 35336 19208 35336 19208 0 _0267_
rlabel metal2 33880 17304 33880 17304 0 _0268_
rlabel metal3 36512 19096 36512 19096 0 _0269_
rlabel metal2 35672 17416 35672 17416 0 _0270_
rlabel metal3 37912 22344 37912 22344 0 _0271_
rlabel metal2 38248 27440 38248 27440 0 _0272_
rlabel metal3 39424 26264 39424 26264 0 _0273_
rlabel metal2 38472 22876 38472 22876 0 _0274_
rlabel metal2 23800 24080 23800 24080 0 _0275_
rlabel metal2 63336 24976 63336 24976 0 _0276_
rlabel metal2 63784 23856 63784 23856 0 _0277_
rlabel metal2 62776 37772 62776 37772 0 _0278_
rlabel metal2 37800 24136 37800 24136 0 _0279_
rlabel metal2 34328 18088 34328 18088 0 _0280_
rlabel metal2 35448 19376 35448 19376 0 _0281_
rlabel metal2 38024 23856 38024 23856 0 _0282_
rlabel metal2 38584 25480 38584 25480 0 _0283_
rlabel metal2 20104 22624 20104 22624 0 _0284_
rlabel metal2 72184 29232 72184 29232 0 _0285_
rlabel metal3 71848 30968 71848 30968 0 _0286_
rlabel metal2 71792 25928 71792 25928 0 _0287_
rlabel metal2 72072 24360 72072 24360 0 _0288_
rlabel metal3 67704 25480 67704 25480 0 _0289_
rlabel metal3 36512 22120 36512 22120 0 _0290_
rlabel metal3 35896 16856 35896 16856 0 _0291_
rlabel metal2 37072 17752 37072 17752 0 _0292_
rlabel metal2 35784 22848 35784 22848 0 _0293_
rlabel metal2 37576 24248 37576 24248 0 _0294_
rlabel metal2 24696 22400 24696 22400 0 _0295_
rlabel metal2 72744 30184 72744 30184 0 _0296_
rlabel metal2 72520 25928 72520 25928 0 _0297_
rlabel metal2 73752 25200 73752 25200 0 _0298_
rlabel metal2 65576 39984 65576 39984 0 _0299_
rlabel metal3 68376 26488 68376 26488 0 _0300_
rlabel metal3 39816 23072 39816 23072 0 _0301_
rlabel metal3 35336 15736 35336 15736 0 _0302_
rlabel metal2 36008 18256 36008 18256 0 _0303_
rlabel metal2 36568 21840 36568 21840 0 _0304_
rlabel metal2 39872 21672 39872 21672 0 _0305_
rlabel metal2 20552 20216 20552 20216 0 _0306_
rlabel metal2 42952 18368 42952 18368 0 _0307_
rlabel metal3 72072 23800 72072 23800 0 _0308_
rlabel metal2 76552 18816 76552 18816 0 _0309_
rlabel metal2 72744 20440 72744 20440 0 _0310_
rlabel metal2 66808 40768 66808 40768 0 _0311_
rlabel metal3 68936 20888 68936 20888 0 _0312_
rlabel metal2 40040 18928 40040 18928 0 _0313_
rlabel metal2 39816 18032 39816 18032 0 _0314_
rlabel metal2 39704 15960 39704 15960 0 _0315_
rlabel metal3 39424 16856 39424 16856 0 _0316_
rlabel metal2 39032 17808 39032 17808 0 _0317_
rlabel metal2 40264 19600 40264 19600 0 _0318_
rlabel metal2 42056 26320 42056 26320 0 _0319_
rlabel metal2 40936 25928 40936 25928 0 _0320_
rlabel metal2 40824 28056 40824 28056 0 _0321_
rlabel metal2 21672 17360 21672 17360 0 _0322_
rlabel metal2 72800 21560 72800 21560 0 _0323_
rlabel metal2 73528 21504 73528 21504 0 _0324_
rlabel metal3 69104 21672 69104 21672 0 _0325_
rlabel metal2 41496 16912 41496 16912 0 _0326_
rlabel metal2 38528 16296 38528 16296 0 _0327_
rlabel metal2 41384 17192 41384 17192 0 _0328_
rlabel metal2 41720 18144 41720 18144 0 _0329_
rlabel metal3 40320 19208 40320 19208 0 _0330_
rlabel metal2 25144 18536 25144 18536 0 _0331_
rlabel metal2 72912 28504 72912 28504 0 _0332_
rlabel metal3 73584 26488 73584 26488 0 _0333_
rlabel metal3 77784 18144 77784 18144 0 _0334_
rlabel metal2 66976 40600 66976 40600 0 _0335_
rlabel metal2 41384 18872 41384 18872 0 _0336_
rlabel metal3 38696 16296 38696 16296 0 _0337_
rlabel metal2 39704 17920 39704 17920 0 _0338_
rlabel metal2 41384 17920 41384 17920 0 _0339_
rlabel metal2 41496 21840 41496 21840 0 _0340_
rlabel metal2 24808 20552 24808 20552 0 _0341_
rlabel metal2 76832 30968 76832 30968 0 _0342_
rlabel metal2 73528 27440 73528 27440 0 _0343_
rlabel metal2 73136 26824 73136 26824 0 _0344_
rlabel metal2 76664 18928 76664 18928 0 _0345_
rlabel metal2 68712 37632 68712 37632 0 _0346_
rlabel metal2 68320 39592 68320 39592 0 _0347_
rlabel metal2 73080 23296 73080 23296 0 _0348_
rlabel metal2 40600 19376 40600 19376 0 _0349_
rlabel metal2 39032 15624 39032 15624 0 _0350_
rlabel metal2 39816 16912 39816 16912 0 _0351_
rlabel metal2 40824 19320 40824 19320 0 _0352_
rlabel metal2 41160 23744 41160 23744 0 _0353_
rlabel via2 46760 19320 46760 19320 0 _0354_
rlabel metal3 43792 21672 43792 21672 0 _0355_
rlabel metal2 72912 24472 72912 24472 0 _0356_
rlabel metal2 76888 21336 76888 21336 0 _0357_
rlabel metal2 73304 22008 73304 22008 0 _0358_
rlabel metal2 68600 38976 68600 38976 0 _0359_
rlabel metal3 69776 23352 69776 23352 0 _0360_
rlabel metal2 41944 19656 41944 19656 0 _0361_
rlabel metal3 38892 19208 38892 19208 0 _0362_
rlabel metal2 38920 18144 38920 18144 0 _0363_
rlabel metal2 38696 18368 38696 18368 0 _0364_
rlabel metal2 41832 18760 41832 18760 0 _0365_
rlabel metal3 43344 18200 43344 18200 0 _0366_
rlabel metal2 43064 25256 43064 25256 0 _0367_
rlabel metal2 44296 25928 44296 25928 0 _0368_
rlabel metal3 44016 20104 44016 20104 0 _0369_
rlabel metal2 44744 15960 44744 15960 0 _0370_
rlabel metal2 72856 23352 72856 23352 0 _0371_
rlabel metal2 73416 22120 73416 22120 0 _0372_
rlabel metal3 70616 22456 70616 22456 0 _0373_
rlabel metal2 43512 16072 43512 16072 0 _0374_
rlabel metal2 38024 17360 38024 17360 0 _0375_
rlabel metal2 43400 16352 43400 16352 0 _0376_
rlabel metal2 43680 16072 43680 16072 0 _0377_
rlabel metal2 44072 24416 44072 24416 0 _0378_
rlabel metal2 47208 19488 47208 19488 0 _0379_
rlabel metal2 76944 28616 76944 28616 0 _0380_
rlabel metal2 75040 23128 75040 23128 0 _0381_
rlabel metal2 77000 20048 77000 20048 0 _0382_
rlabel metal2 70560 39032 70560 39032 0 _0383_
rlabel metal3 44968 15848 44968 15848 0 _0384_
rlabel metal2 40040 19712 40040 19712 0 _0385_
rlabel metal2 43960 17024 43960 17024 0 _0386_
rlabel metal2 44072 17080 44072 17080 0 _0387_
rlabel metal2 44520 24584 44520 24584 0 _0388_
rlabel metal2 44184 20888 44184 20888 0 _0389_
rlabel metal2 77112 27776 77112 27776 0 _0390_
rlabel metal2 74872 22960 74872 22960 0 _0391_
rlabel metal3 75992 21000 75992 21000 0 _0392_
rlabel metal3 69720 38808 69720 38808 0 _0393_
rlabel metal2 69496 31304 69496 31304 0 _0394_
rlabel metal2 43848 22512 43848 22512 0 _0395_
rlabel metal3 37240 19208 37240 19208 0 _0396_
rlabel metal3 43736 22120 43736 22120 0 _0397_
rlabel metal2 44072 21840 44072 21840 0 _0398_
rlabel metal2 45304 23688 45304 23688 0 _0399_
rlabel metal3 36680 14504 36680 14504 0 _0400_
rlabel metal3 52024 14504 52024 14504 0 _0401_
rlabel metal2 47768 16352 47768 16352 0 _0402_
rlabel metal3 70728 27888 70728 27888 0 _0403_
rlabel metal2 77896 31416 77896 31416 0 _0404_
rlabel metal2 77112 25200 77112 25200 0 _0405_
rlabel metal3 72184 26264 72184 26264 0 _0406_
rlabel metal3 72184 40488 72184 40488 0 _0407_
rlabel metal2 71008 38920 71008 38920 0 _0408_
rlabel metal2 70280 33600 70280 33600 0 _0409_
rlabel metal3 48720 23240 48720 23240 0 _0410_
rlabel metal2 46032 26264 46032 26264 0 _0411_
rlabel metal2 46200 22008 46200 22008 0 _0412_
rlabel metal2 48048 20216 48048 20216 0 _0413_
rlabel metal2 45584 24920 45584 24920 0 _0414_
rlabel metal2 45976 22736 45976 22736 0 _0415_
rlabel metal4 47656 22288 47656 22288 0 _0416_
rlabel metal2 47544 18200 47544 18200 0 _0417_
rlabel metal2 45528 21448 45528 21448 0 _0418_
rlabel metal2 48552 20272 48552 20272 0 _0419_
rlabel metal2 47768 20552 47768 20552 0 _0420_
rlabel metal2 46984 21392 46984 21392 0 _0421_
rlabel metal2 46872 17472 46872 17472 0 _0422_
rlabel metal2 45528 14784 45528 14784 0 _0423_
rlabel metal2 70728 27272 70728 27272 0 _0424_
rlabel metal2 70448 26824 70448 26824 0 _0425_
rlabel metal2 71064 31024 71064 31024 0 _0426_
rlabel metal2 47376 23352 47376 23352 0 _0427_
rlabel metal2 48104 21952 48104 21952 0 _0428_
rlabel metal2 46312 22792 46312 22792 0 _0429_
rlabel metal2 47208 15904 47208 15904 0 _0430_
rlabel metal2 47712 15400 47712 15400 0 _0431_
rlabel metal2 48328 14504 48328 14504 0 _0432_
rlabel metal3 75432 28616 75432 28616 0 _0433_
rlabel metal2 70728 29456 70728 29456 0 _0434_
rlabel metal3 70672 25032 70672 25032 0 _0435_
rlabel metal2 70504 38668 70504 38668 0 _0436_
rlabel metal2 49056 23352 49056 23352 0 _0437_
rlabel metal2 46648 22568 46648 22568 0 _0438_
rlabel metal2 46760 23296 46760 23296 0 _0439_
rlabel metal4 46872 19096 46872 19096 0 _0440_
rlabel metal2 48104 16968 48104 16968 0 _0441_
rlabel metal2 47320 15736 47320 15736 0 _0442_
rlabel metal2 76664 30016 76664 30016 0 _0443_
rlabel metal2 74424 29680 74424 29680 0 _0444_
rlabel metal2 75432 27272 75432 27272 0 _0445_
rlabel metal3 71288 37912 71288 37912 0 _0446_
rlabel metal3 71904 35224 71904 35224 0 _0447_
rlabel metal2 47544 23912 47544 23912 0 _0448_
rlabel metal2 45192 23632 45192 23632 0 _0449_
rlabel metal2 47432 23744 47432 23744 0 _0450_
rlabel metal2 47768 23576 47768 23576 0 _0451_
rlabel metal2 49560 17920 49560 17920 0 _0452_
rlabel metal2 26824 17192 26824 17192 0 _0453_
rlabel metal2 51128 18816 51128 18816 0 _0454_
rlabel metal2 72072 30520 72072 30520 0 _0455_
rlabel metal2 77560 28560 77560 28560 0 _0456_
rlabel metal4 71960 27552 71960 27552 0 _0457_
rlabel metal2 72744 37520 72744 37520 0 _0458_
rlabel metal2 72352 37128 72352 37128 0 _0459_
rlabel metal2 50512 30744 50512 30744 0 _0460_
rlabel metal3 47320 26376 47320 26376 0 _0461_
rlabel metal2 47152 25704 47152 25704 0 _0462_
rlabel metal2 46984 26208 46984 26208 0 _0463_
rlabel metal2 49336 26152 49336 26152 0 _0464_
rlabel metal2 50064 18424 50064 18424 0 _0465_
rlabel metal2 49952 21672 49952 21672 0 _0466_
rlabel metal3 49672 20776 49672 20776 0 _0467_
rlabel metal2 48888 18872 48888 18872 0 _0468_
rlabel metal3 33432 16968 33432 16968 0 _0469_
rlabel metal2 73752 29792 73752 29792 0 _0470_
rlabel metal4 73864 26572 73864 26572 0 _0471_
rlabel metal2 72968 31920 72968 31920 0 _0472_
rlabel metal3 65828 30408 65828 30408 0 _0473_
rlabel metal3 45752 26264 45752 26264 0 _0474_
rlabel metal3 47712 26264 47712 26264 0 _0475_
rlabel metal2 48832 26040 48832 26040 0 _0476_
rlabel metal2 49392 16968 49392 16968 0 _0477_
rlabel metal2 46312 17248 46312 17248 0 _0478_
rlabel metal3 76720 34216 76720 34216 0 _0479_
rlabel metal3 73836 31528 73836 31528 0 _0480_
rlabel metal2 77672 28224 77672 28224 0 _0481_
rlabel metal2 72912 36792 72912 36792 0 _0482_
rlabel metal3 50176 26936 50176 26936 0 _0483_
rlabel metal2 47320 26992 47320 26992 0 _0484_
rlabel metal3 48552 27048 48552 27048 0 _0485_
rlabel metal2 49728 22792 49728 22792 0 _0486_
rlabel metal2 49336 19152 49336 19152 0 _0487_
rlabel metal2 49448 14056 49448 14056 0 _0488_
rlabel metal2 77000 32256 77000 32256 0 _0489_
rlabel metal3 75432 31192 75432 31192 0 _0490_
rlabel metal2 77672 30016 77672 30016 0 _0491_
rlabel metal2 71680 37464 71680 37464 0 _0492_
rlabel metal2 73640 31528 73640 31528 0 _0493_
rlabel metal2 60424 29064 60424 29064 0 _0494_
rlabel metal2 46424 27160 46424 27160 0 _0495_
rlabel metal2 49000 27160 49000 27160 0 _0496_
rlabel metal2 49336 26656 49336 26656 0 _0497_
rlabel metal2 49224 18592 49224 18592 0 _0498_
rlabel metal2 41608 13888 41608 13888 0 _0499_
rlabel metal2 52024 14056 52024 14056 0 _0500_
rlabel metal2 75320 33656 75320 33656 0 _0501_
rlabel metal3 75096 32648 75096 32648 0 _0502_
rlabel metal2 74872 33096 74872 33096 0 _0503_
rlabel metal3 75712 40600 75712 40600 0 _0504_
rlabel metal2 74648 33936 74648 33936 0 _0505_
rlabel metal3 51632 30072 51632 30072 0 _0506_
rlabel metal2 46200 31360 46200 31360 0 _0507_
rlabel metal2 44968 29848 44968 29848 0 _0508_
rlabel metal2 46312 31024 46312 31024 0 _0509_
rlabel metal3 49056 30184 49056 30184 0 _0510_
rlabel metal3 52024 22680 52024 22680 0 _0511_
rlabel metal3 53368 20104 53368 20104 0 _0512_
rlabel metal3 52360 19208 52360 19208 0 _0513_
rlabel metal2 51520 20216 51520 20216 0 _0514_
rlabel metal2 42784 12824 42784 12824 0 _0515_
rlabel metal3 75600 34104 75600 34104 0 _0516_
rlabel metal2 77896 32088 77896 32088 0 _0517_
rlabel metal2 75096 35784 75096 35784 0 _0518_
rlabel metal3 53144 31976 53144 31976 0 _0519_
rlabel metal3 45136 30184 45136 30184 0 _0520_
rlabel metal2 52472 30688 52472 30688 0 _0521_
rlabel metal2 53424 30856 53424 30856 0 _0522_
rlabel metal2 53816 16744 53816 16744 0 _0523_
rlabel metal2 42728 14616 42728 14616 0 _0524_
rlabel metal2 76664 37296 76664 37296 0 _0525_
rlabel metal2 76664 35392 76664 35392 0 _0526_
rlabel metal2 76776 34272 76776 34272 0 _0527_
rlabel metal2 76048 34888 76048 34888 0 _0528_
rlabel metal2 51800 30688 51800 30688 0 _0529_
rlabel metal2 45752 31248 45752 31248 0 _0530_
rlabel metal2 51464 30912 51464 30912 0 _0531_
rlabel metal2 52080 30296 52080 30296 0 _0532_
rlabel metal2 52360 17808 52360 17808 0 _0533_
rlabel metal3 42448 15848 42448 15848 0 _0534_
rlabel metal3 76608 38696 76608 38696 0 _0535_
rlabel metal2 76888 37016 76888 37016 0 _0536_
rlabel metal2 75432 35224 75432 35224 0 _0537_
rlabel metal2 69608 41216 69608 41216 0 _0538_
rlabel metal2 76328 39788 76328 39788 0 _0539_
rlabel metal3 52192 31640 52192 31640 0 _0540_
rlabel metal3 45360 31752 45360 31752 0 _0541_
rlabel metal3 48720 31752 48720 31752 0 _0542_
rlabel metal2 51856 31528 51856 31528 0 _0543_
rlabel metal2 52024 20608 52024 20608 0 _0544_
rlabel metal2 41720 12432 41720 12432 0 _0545_
rlabel metal2 55160 17416 55160 17416 0 _0546_
rlabel metal3 76832 38584 76832 38584 0 _0547_
rlabel metal2 74816 39480 74816 39480 0 _0548_
rlabel metal2 74872 36624 74872 36624 0 _0549_
rlabel metal2 77616 42728 77616 42728 0 _0550_
rlabel metal2 77840 39256 77840 39256 0 _0551_
rlabel metal3 53592 34216 53592 34216 0 _0552_
rlabel metal3 46256 35784 46256 35784 0 _0553_
rlabel metal3 44968 33320 44968 33320 0 _0554_
rlabel metal2 46088 32984 46088 32984 0 _0555_
rlabel metal2 45752 33600 45752 33600 0 _0556_
rlabel metal2 53200 17640 53200 17640 0 _0557_
rlabel metal2 54376 21616 54376 21616 0 _0558_
rlabel metal2 53592 20384 53592 20384 0 _0559_
rlabel metal2 53480 17584 53480 17584 0 _0560_
rlabel metal2 45192 11200 45192 11200 0 _0561_
rlabel metal2 77560 38472 77560 38472 0 _0562_
rlabel metal2 78120 36904 78120 36904 0 _0563_
rlabel metal2 77112 40768 77112 40768 0 _0564_
rlabel metal2 54376 37464 54376 37464 0 _0565_
rlabel metal2 45192 34888 45192 34888 0 _0566_
rlabel metal3 49616 34888 49616 34888 0 _0567_
rlabel metal3 53312 33768 53312 33768 0 _0568_
rlabel metal3 53704 18536 53704 18536 0 _0569_
rlabel metal2 40936 9632 40936 9632 0 _0570_
rlabel metal2 75320 39480 75320 39480 0 _0571_
rlabel metal2 78008 37352 78008 37352 0 _0572_
rlabel metal2 77224 41832 77224 41832 0 _0573_
rlabel metal2 54600 34272 54600 34272 0 _0574_
rlabel metal3 45080 35672 45080 35672 0 _0575_
rlabel metal2 54264 34720 54264 34720 0 _0576_
rlabel metal2 54600 26600 54600 26600 0 _0577_
rlabel metal2 54824 20048 54824 20048 0 _0578_
rlabel metal2 43960 9240 43960 9240 0 _0579_
rlabel metal2 73584 39032 73584 39032 0 _0580_
rlabel metal2 74088 39872 74088 39872 0 _0581_
rlabel metal2 73192 40096 73192 40096 0 _0582_
rlabel metal2 54824 34832 54824 34832 0 _0583_
rlabel metal2 46984 36008 46984 36008 0 _0584_
rlabel metal2 54488 35224 54488 35224 0 _0585_
rlabel metal2 55160 31920 55160 31920 0 _0586_
rlabel metal2 55384 20664 55384 20664 0 _0587_
rlabel metal2 78120 39872 78120 39872 0 _0588_
rlabel metal2 30072 6552 30072 6552 0 _0589_
rlabel metal2 33320 4368 33320 4368 0 _0590_
rlabel metal2 16856 7280 16856 7280 0 _0591_
rlabel metal2 11256 4704 11256 4704 0 _0592_
rlabel metal2 14168 5264 14168 5264 0 _0593_
rlabel metal2 28280 6272 28280 6272 0 _0594_
rlabel metal2 19712 7448 19712 7448 0 _0595_
rlabel metal2 18088 6832 18088 6832 0 _0596_
rlabel metal2 23128 8176 23128 8176 0 _0597_
rlabel metal2 18760 8624 18760 8624 0 _0598_
rlabel metal3 17248 8904 17248 8904 0 _0599_
rlabel metal2 15568 6104 15568 6104 0 _0600_
rlabel metal3 16912 8344 16912 8344 0 _0601_
rlabel metal3 15372 7560 15372 7560 0 _0602_
rlabel metal3 17192 7336 17192 7336 0 _0603_
rlabel metal2 14728 5544 14728 5544 0 _0604_
rlabel metal2 17976 5880 17976 5880 0 _0605_
rlabel metal2 17976 4704 17976 4704 0 _0606_
rlabel metal2 17304 6384 17304 6384 0 _0607_
rlabel metal2 19208 12824 19208 12824 0 _0608_
rlabel metal2 19880 12208 19880 12208 0 _0609_
rlabel metal3 18648 12040 18648 12040 0 _0610_
rlabel metal2 15624 4088 15624 4088 0 _0611_
rlabel metal2 20160 12264 20160 12264 0 _0612_
rlabel metal2 19544 5544 19544 5544 0 _0613_
rlabel metal2 18480 10696 18480 10696 0 _0614_
rlabel metal2 17864 5096 17864 5096 0 _0615_
rlabel metal2 19880 8400 19880 8400 0 _0616_
rlabel metal2 20328 5208 20328 5208 0 _0617_
rlabel metal2 23016 4480 23016 4480 0 _0618_
rlabel metal3 22456 4424 22456 4424 0 _0619_
rlabel metal2 26712 8288 26712 8288 0 _0620_
rlabel metal2 25704 7616 25704 7616 0 _0621_
rlabel metal2 26376 7840 26376 7840 0 _0622_
rlabel metal2 22008 5096 22008 5096 0 _0623_
rlabel metal2 21224 4872 21224 4872 0 _0624_
rlabel metal2 23352 6384 23352 6384 0 _0625_
rlabel metal2 22456 6216 22456 6216 0 _0626_
rlabel metal3 24808 7336 24808 7336 0 _0627_
rlabel metal2 21672 5432 21672 5432 0 _0628_
rlabel metal3 27160 8344 27160 8344 0 _0629_
rlabel metal2 21504 5320 21504 5320 0 _0630_
rlabel metal2 20664 6832 20664 6832 0 _0631_
rlabel metal2 25256 11928 25256 11928 0 _0632_
rlabel metal2 24696 9632 24696 9632 0 _0633_
rlabel metal2 26096 12152 26096 12152 0 _0634_
rlabel metal3 23408 10472 23408 10472 0 _0635_
rlabel metal2 21784 5432 21784 5432 0 _0636_
rlabel metal3 25424 10808 25424 10808 0 _0637_
rlabel metal2 19096 5488 19096 5488 0 _0638_
rlabel metal2 22512 11592 22512 11592 0 _0639_
rlabel metal2 21560 6160 21560 6160 0 _0640_
rlabel metal3 25200 13048 25200 13048 0 _0641_
rlabel metal3 29680 5880 29680 5880 0 _0642_
rlabel metal3 25480 5656 25480 5656 0 _0643_
rlabel metal2 26488 5768 26488 5768 0 _0644_
rlabel metal2 32200 7168 32200 7168 0 _0645_
rlabel metal2 31584 9576 31584 9576 0 _0646_
rlabel metal2 32312 9744 32312 9744 0 _0647_
rlabel metal2 30296 9240 30296 9240 0 _0648_
rlabel metal2 25480 6664 25480 6664 0 _0649_
rlabel metal2 32984 10024 32984 10024 0 _0650_
rlabel metal2 27832 5768 27832 5768 0 _0651_
rlabel metal3 30744 11256 30744 11256 0 _0652_
rlabel metal2 25032 6328 25032 6328 0 _0653_
rlabel metal2 29512 10248 29512 10248 0 _0654_
rlabel metal2 28952 6552 28952 6552 0 _0655_
rlabel metal2 28392 6104 28392 6104 0 _0656_
rlabel metal2 34104 7224 34104 7224 0 _0657_
rlabel metal2 33320 6720 33320 6720 0 _0658_
rlabel metal2 34216 8568 34216 8568 0 _0659_
rlabel metal3 30072 5096 30072 5096 0 _0660_
rlabel metal2 30968 5544 30968 5544 0 _0661_
rlabel metal2 27832 5264 27832 5264 0 _0662_
rlabel metal2 74200 2478 74200 2478 0 clk
rlabel metal2 23800 16464 23800 16464 0 clknet_0_clk
rlabel metal2 15400 10640 15400 10640 0 clknet_3_0__leaf_clk
rlabel metal3 19208 9016 19208 9016 0 clknet_3_1__leaf_clk
rlabel metal2 16744 22344 16744 22344 0 clknet_3_2__leaf_clk
rlabel metal2 21336 22848 21336 22848 0 clknet_3_3__leaf_clk
rlabel metal2 33264 11368 33264 11368 0 clknet_3_4__leaf_clk
rlabel metal3 40656 15176 40656 15176 0 clknet_3_5__leaf_clk
rlabel metal2 26488 19376 26488 19376 0 clknet_3_6__leaf_clk
rlabel metal2 41048 21224 41048 21224 0 clknet_3_7__leaf_clk
rlabel metal2 27160 7616 27160 7616 0 gpio\[16\]
rlabel metal2 26432 6664 26432 6664 0 gpio\[17\]
rlabel metal2 25928 8232 25928 8232 0 gpio\[18\]
rlabel metal2 26824 8344 26824 8344 0 gpio\[19\]
rlabel metal2 24360 11312 24360 11312 0 gpio\[20\]
rlabel metal2 25928 11144 25928 11144 0 gpio\[21\]
rlabel metal2 25480 12824 25480 12824 0 gpio\[22\]
rlabel metal2 26488 13104 26488 13104 0 gpio\[23\]
rlabel metal2 31864 9912 31864 9912 0 gpio\[24\]
rlabel metal2 36008 11424 36008 11424 0 gpio\[25\]
rlabel metal2 32088 12152 32088 12152 0 gpio\[26\]
rlabel metal2 31696 11928 31696 11928 0 gpio\[27\]
rlabel metal2 38808 10360 38808 10360 0 gpio\[28\]
rlabel metal2 36456 7112 36456 7112 0 gpio\[29\]
rlabel metal2 38920 8904 38920 8904 0 gpio\[30\]
rlabel metal2 37352 7784 37352 7784 0 gpio\[31\]
rlabel metal2 11256 76706 11256 76706 0 gpio_out[0]
rlabel metal2 19208 74928 19208 74928 0 gpio_out[10]
rlabel metal2 18648 77490 18648 77490 0 gpio_out[11]
rlabel metal2 19264 76664 19264 76664 0 gpio_out[12]
rlabel metal2 20216 75152 20216 75152 0 gpio_out[13]
rlabel metal3 21112 75880 21112 75880 0 gpio_out[14]
rlabel metal2 21336 77770 21336 77770 0 gpio_out[15]
rlabel metal2 11928 78554 11928 78554 0 gpio_out[1]
rlabel metal2 12600 77546 12600 77546 0 gpio_out[2]
rlabel metal2 12936 75600 12936 75600 0 gpio_out[3]
rlabel metal2 11592 75880 11592 75880 0 gpio_out[4]
rlabel metal2 14616 76202 14616 76202 0 gpio_out[5]
rlabel metal2 15288 77154 15288 77154 0 gpio_out[6]
rlabel metal2 16072 75432 16072 75432 0 gpio_out[7]
rlabel metal3 16016 76664 16016 76664 0 gpio_out[8]
rlabel metal2 17304 78218 17304 78218 0 gpio_out[9]
rlabel metal2 31304 23072 31304 23072 0 iomem_rdata\[0\]
rlabel metal2 24752 16744 24752 16744 0 iomem_rdata\[10\]
rlabel metal2 24528 19880 24528 19880 0 iomem_rdata\[11\]
rlabel metal2 28840 19320 28840 19320 0 iomem_rdata\[12\]
rlabel metal2 32200 18872 32200 18872 0 iomem_rdata\[13\]
rlabel metal2 32536 20440 32536 20440 0 iomem_rdata\[14\]
rlabel metal2 32088 21504 32088 21504 0 iomem_rdata\[15\]
rlabel metal2 37968 15176 37968 15176 0 iomem_rdata\[16\]
rlabel metal2 38024 13664 38024 13664 0 iomem_rdata\[17\]
rlabel metal2 34384 14616 34384 14616 0 iomem_rdata\[18\]
rlabel metal2 35336 16128 35336 16128 0 iomem_rdata\[19\]
rlabel metal2 26936 24360 26936 24360 0 iomem_rdata\[1\]
rlabel metal2 28616 18032 28616 18032 0 iomem_rdata\[20\]
rlabel metal2 31584 16744 31584 16744 0 iomem_rdata\[21\]
rlabel metal2 28112 16184 28112 16184 0 iomem_rdata\[22\]
rlabel metal2 31248 13608 31248 13608 0 iomem_rdata\[23\]
rlabel metal2 42000 13048 42000 13048 0 iomem_rdata\[24\]
rlabel metal2 44968 13664 44968 13664 0 iomem_rdata\[25\]
rlabel metal2 44632 15148 44632 15148 0 iomem_rdata\[26\]
rlabel metal2 42168 15288 42168 15288 0 iomem_rdata\[27\]
rlabel metal2 40376 12096 40376 12096 0 iomem_rdata\[28\]
rlabel metal2 44296 10864 44296 10864 0 iomem_rdata\[29\]
rlabel metal2 29960 24640 29960 24640 0 iomem_rdata\[2\]
rlabel metal2 40376 9296 40376 9296 0 iomem_rdata\[30\]
rlabel metal2 44912 8904 44912 8904 0 iomem_rdata\[31\]
rlabel metal3 28784 22456 28784 22456 0 iomem_rdata\[3\]
rlabel metal2 19824 24024 19824 24024 0 iomem_rdata\[4\]
rlabel metal2 23296 24584 23296 24584 0 iomem_rdata\[5\]
rlabel metal2 19600 22456 19600 22456 0 iomem_rdata\[6\]
rlabel metal2 24416 22456 24416 22456 0 iomem_rdata\[7\]
rlabel metal2 21336 20776 21336 20776 0 iomem_rdata\[8\]
rlabel metal2 21392 16744 21392 16744 0 iomem_rdata\[9\]
rlabel metal2 44296 6888 44296 6888 0 iomem_ready
rlabel metal2 26488 1246 26488 1246 0 mem_addr[0]
rlabel metal3 29400 4984 29400 4984 0 mem_addr[10]
rlabel metal2 31416 5152 31416 5152 0 mem_addr[11]
rlabel metal3 31080 2296 31080 2296 0 mem_addr[12]
rlabel metal2 35224 854 35224 854 0 mem_addr[13]
rlabel metal2 35896 1302 35896 1302 0 mem_addr[14]
rlabel metal2 30128 3528 30128 3528 0 mem_addr[15]
rlabel metal2 24136 3192 24136 3192 0 mem_addr[16]
rlabel metal2 37912 1246 37912 1246 0 mem_addr[17]
rlabel metal2 38584 2086 38584 2086 0 mem_addr[18]
rlabel metal2 39256 1806 39256 1806 0 mem_addr[19]
rlabel metal2 22456 4144 22456 4144 0 mem_addr[1]
rlabel metal2 39928 2198 39928 2198 0 mem_addr[20]
rlabel metal2 40600 2142 40600 2142 0 mem_addr[21]
rlabel metal2 41272 2058 41272 2058 0 mem_addr[22]
rlabel metal2 51128 4480 51128 4480 0 mem_addr[23]
rlabel metal2 51576 4424 51576 4424 0 mem_addr[24]
rlabel metal2 42168 4872 42168 4872 0 mem_addr[25]
rlabel metal2 49112 4144 49112 4144 0 mem_addr[26]
rlabel metal2 53592 4536 53592 4536 0 mem_addr[27]
rlabel metal2 45248 3304 45248 3304 0 mem_addr[28]
rlabel metal2 49224 5208 49224 5208 0 mem_addr[29]
rlabel metal2 21112 3696 21112 3696 0 mem_addr[2]
rlabel metal2 49112 5320 49112 5320 0 mem_addr[30]
rlabel metal2 47320 2058 47320 2058 0 mem_addr[31]
rlabel metal2 23016 3808 23016 3808 0 mem_addr[3]
rlabel metal3 22848 3192 22848 3192 0 mem_addr[4]
rlabel metal2 23800 4984 23800 4984 0 mem_addr[5]
rlabel metal2 30520 2058 30520 2058 0 mem_addr[6]
rlabel metal2 25480 4536 25480 4536 0 mem_addr[7]
rlabel metal3 25760 3528 25760 3528 0 mem_addr[8]
rlabel metal2 23016 6776 23016 6776 0 mem_addr[9]
rlabel metal2 52696 2422 52696 2422 0 mem_rdata[0]
rlabel metal2 59416 3206 59416 3206 0 mem_rdata[10]
rlabel metal2 60088 3598 60088 3598 0 mem_rdata[11]
rlabel metal2 60760 2982 60760 2982 0 mem_rdata[12]
rlabel metal2 61432 1134 61432 1134 0 mem_rdata[13]
rlabel metal2 62104 2254 62104 2254 0 mem_rdata[14]
rlabel metal2 62776 3598 62776 3598 0 mem_rdata[15]
rlabel metal2 63448 854 63448 854 0 mem_rdata[16]
rlabel metal2 64120 2422 64120 2422 0 mem_rdata[17]
rlabel metal3 71288 3528 71288 3528 0 mem_rdata[18]
rlabel metal2 68936 4648 68936 4648 0 mem_rdata[19]
rlabel metal2 53368 2198 53368 2198 0 mem_rdata[1]
rlabel metal2 66136 1694 66136 1694 0 mem_rdata[20]
rlabel metal2 67816 6160 67816 6160 0 mem_rdata[21]
rlabel metal2 67480 1974 67480 1974 0 mem_rdata[22]
rlabel metal2 68152 2982 68152 2982 0 mem_rdata[23]
rlabel metal2 68824 2310 68824 2310 0 mem_rdata[24]
rlabel metal2 69496 2254 69496 2254 0 mem_rdata[25]
rlabel metal2 70168 1974 70168 1974 0 mem_rdata[26]
rlabel metal2 70840 3206 70840 3206 0 mem_rdata[27]
rlabel metal2 71512 2422 71512 2422 0 mem_rdata[28]
rlabel metal2 72184 2926 72184 2926 0 mem_rdata[29]
rlabel metal2 54040 2982 54040 2982 0 mem_rdata[2]
rlabel metal2 72856 3262 72856 3262 0 mem_rdata[30]
rlabel metal2 73528 2982 73528 2982 0 mem_rdata[31]
rlabel metal2 54712 2086 54712 2086 0 mem_rdata[3]
rlabel metal2 55384 2142 55384 2142 0 mem_rdata[4]
rlabel metal2 56056 1470 56056 1470 0 mem_rdata[5]
rlabel metal2 56728 3206 56728 3206 0 mem_rdata[6]
rlabel metal2 57400 2422 57400 2422 0 mem_rdata[7]
rlabel metal2 58072 2086 58072 2086 0 mem_rdata[8]
rlabel metal2 58744 2814 58744 2814 0 mem_rdata[9]
rlabel metal2 49336 2422 49336 2422 0 mem_ready
rlabel metal2 50568 5208 50568 5208 0 mem_valid
rlabel metal2 4368 728 4368 728 0 mem_wdata[0]
rlabel metal2 11704 2058 11704 2058 0 mem_wdata[10]
rlabel metal2 12376 1694 12376 1694 0 mem_wdata[11]
rlabel metal2 13048 1638 13048 1638 0 mem_wdata[12]
rlabel metal2 13664 3192 13664 3192 0 mem_wdata[13]
rlabel metal2 14336 3080 14336 3080 0 mem_wdata[14]
rlabel metal2 15008 3192 15008 3192 0 mem_wdata[15]
rlabel metal2 15736 1918 15736 1918 0 mem_wdata[16]
rlabel metal2 16408 1246 16408 1246 0 mem_wdata[17]
rlabel metal2 17080 2142 17080 2142 0 mem_wdata[18]
rlabel metal2 17752 2590 17752 2590 0 mem_wdata[19]
rlabel metal3 4536 3528 4536 3528 0 mem_wdata[1]
rlabel metal2 18424 2254 18424 2254 0 mem_wdata[20]
rlabel metal2 19096 2310 19096 2310 0 mem_wdata[21]
rlabel metal2 19768 854 19768 854 0 mem_wdata[22]
rlabel metal2 18312 4872 18312 4872 0 mem_wdata[23]
rlabel metal2 21112 2058 21112 2058 0 mem_wdata[24]
rlabel metal3 19824 3976 19824 3976 0 mem_wdata[25]
rlabel metal2 18648 3248 18648 3248 0 mem_wdata[26]
rlabel metal2 23128 2058 23128 2058 0 mem_wdata[27]
rlabel metal2 23800 2058 23800 2058 0 mem_wdata[28]
rlabel metal2 24472 1246 24472 1246 0 mem_wdata[29]
rlabel metal2 6328 2058 6328 2058 0 mem_wdata[2]
rlabel metal2 25144 854 25144 854 0 mem_wdata[30]
rlabel metal2 25816 1246 25816 1246 0 mem_wdata[31]
rlabel metal2 5432 4088 5432 4088 0 mem_wdata[3]
rlabel metal2 7616 3192 7616 3192 0 mem_wdata[4]
rlabel metal2 8232 5376 8232 5376 0 mem_wdata[5]
rlabel metal2 6552 4536 6552 4536 0 mem_wdata[6]
rlabel metal2 9688 2058 9688 2058 0 mem_wdata[7]
rlabel metal2 5880 3584 5880 3584 0 mem_wdata[8]
rlabel metal3 7392 3528 7392 3528 0 mem_wdata[9]
rlabel metal2 51688 4592 51688 4592 0 mem_wstrb[0]
rlabel metal3 51632 3528 51632 3528 0 mem_wstrb[1]
rlabel metal2 53032 3584 53032 3584 0 mem_wstrb[2]
rlabel metal2 53704 3640 53704 3640 0 mem_wstrb[3]
rlabel metal2 24696 3584 24696 3584 0 net1
rlabel metal2 32760 3920 32760 3920 0 net10
rlabel metal2 41048 12096 41048 12096 0 net100
rlabel metal2 38472 15512 38472 15512 0 net101
rlabel metal2 75544 5712 75544 5712 0 net102
rlabel metal2 75264 39144 75264 39144 0 net103
rlabel metal3 69160 55048 69160 55048 0 net104
rlabel metal3 71120 55944 71120 55944 0 net105
rlabel metal3 75992 56616 75992 56616 0 net106
rlabel metal3 73416 58184 73416 58184 0 net107
rlabel metal3 76776 59080 76776 59080 0 net108
rlabel metal2 78344 58408 78344 58408 0 net109
rlabel metal2 33432 3864 33432 3864 0 net11
rlabel metal3 77448 61320 77448 61320 0 net110
rlabel metal2 77336 63112 77336 63112 0 net111
rlabel metal3 77168 62216 77168 62216 0 net112
rlabel metal3 78288 64680 78288 64680 0 net113
rlabel metal2 78176 42392 78176 42392 0 net114
rlabel metal3 73864 66248 73864 66248 0 net115
rlabel metal3 76888 67144 76888 67144 0 net116
rlabel metal3 77000 67816 77000 67816 0 net117
rlabel metal2 77840 69160 77840 69160 0 net118
rlabel metal3 78344 71064 78344 71064 0 net119
rlabel metal2 22736 4424 22736 4424 0 net12
rlabel metal2 78680 71848 78680 71848 0 net120
rlabel metal2 78008 72296 78008 72296 0 net121
rlabel metal2 57008 41944 57008 41944 0 net122
rlabel metal3 77168 72520 77168 72520 0 net123
rlabel metal3 73640 75992 73640 75992 0 net124
rlabel metal2 73136 39368 73136 39368 0 net125
rlabel metal3 75264 74760 75264 74760 0 net126
rlabel metal3 75824 74088 75824 74088 0 net127
rlabel metal2 77896 46536 77896 46536 0 net128
rlabel metal2 73416 34496 73416 34496 0 net129
rlabel metal3 40488 5152 40488 5152 0 net13
rlabel metal3 78456 48776 78456 48776 0 net130
rlabel metal2 72072 33376 72072 33376 0 net131
rlabel metal2 77728 51464 77728 51464 0 net132
rlabel metal3 74368 53032 74368 53032 0 net133
rlabel metal2 77616 53032 77616 53032 0 net134
rlabel metal2 55608 37800 55608 37800 0 net135
rlabel metal2 77952 3416 77952 3416 0 net136
rlabel metal2 77952 17080 77952 17080 0 net137
rlabel metal2 77168 17528 77168 17528 0 net138
rlabel metal2 77896 18088 77896 18088 0 net139
rlabel metal2 40600 4536 40600 4536 0 net14
rlabel metal3 76384 20104 76384 20104 0 net140
rlabel metal2 77224 19544 77224 19544 0 net141
rlabel metal3 77336 18984 77336 18984 0 net142
rlabel metal2 77896 20944 77896 20944 0 net143
rlabel metal2 76608 22232 76608 22232 0 net144
rlabel metal2 77784 24360 77784 24360 0 net145
rlabel metal3 75152 27048 75152 27048 0 net146
rlabel metal2 76496 8008 76496 8008 0 net147
rlabel metal2 77000 26320 77000 26320 0 net148
rlabel metal2 74144 28392 74144 28392 0 net149
rlabel metal2 43176 4592 43176 4592 0 net15
rlabel metal3 76832 27944 76832 27944 0 net150
rlabel metal2 75656 29792 75656 29792 0 net151
rlabel metal2 74648 32592 74648 32592 0 net152
rlabel metal2 77896 30184 77896 30184 0 net153
rlabel metal2 76888 33544 76888 33544 0 net154
rlabel metal2 77896 33152 77896 33152 0 net155
rlabel metal2 74592 36456 74592 36456 0 net156
rlabel metal3 76944 34888 76944 34888 0 net157
rlabel metal2 77168 8120 77168 8120 0 net158
rlabel metal2 78232 36176 78232 36176 0 net159
rlabel metal2 42728 4704 42728 4704 0 net16
rlabel metal2 75208 41552 75208 41552 0 net160
rlabel metal2 77896 8176 77896 8176 0 net161
rlabel metal2 77896 10136 77896 10136 0 net162
rlabel metal2 77896 11704 77896 11704 0 net163
rlabel metal2 77896 12880 77896 12880 0 net164
rlabel metal2 77840 13944 77840 13944 0 net165
rlabel metal3 77616 14392 77616 14392 0 net166
rlabel metal2 77896 16296 77896 16296 0 net167
rlabel metal2 34720 27160 34720 27160 0 net168
rlabel metal2 41608 71764 41608 71764 0 net169
rlabel metal2 41272 4144 41272 4144 0 net17
rlabel metal2 42056 71316 42056 71316 0 net170
rlabel metal2 42616 55440 42616 55440 0 net171
rlabel metal2 44128 43680 44128 43680 0 net172
rlabel metal2 45024 76328 45024 76328 0 net173
rlabel metal2 46088 76328 46088 76328 0 net174
rlabel metal2 45640 71428 45640 71428 0 net175
rlabel metal3 47656 75880 47656 75880 0 net176
rlabel metal3 47488 76328 47488 76328 0 net177
rlabel metal2 47824 43680 47824 43680 0 net178
rlabel metal2 35000 27944 35000 27944 0 net179
rlabel metal2 44072 7840 44072 7840 0 net18
rlabel metal2 49560 20944 49560 20944 0 net180
rlabel metal2 49840 76328 49840 76328 0 net181
rlabel metal2 50960 27384 50960 27384 0 net182
rlabel metal2 50288 43680 50288 43680 0 net183
rlabel metal2 51408 55440 51408 55440 0 net184
rlabel metal2 53312 55440 53312 55440 0 net185
rlabel metal2 52920 23436 52920 23436 0 net186
rlabel metal2 53648 33544 53648 33544 0 net187
rlabel metal2 54208 31920 54208 31920 0 net188
rlabel metal2 53984 20776 53984 20776 0 net189
rlabel metal2 47152 6664 47152 6664 0 net19
rlabel metal3 36512 28056 36512 28056 0 net190
rlabel metal2 54880 37800 54880 37800 0 net191
rlabel metal2 55888 21784 55888 21784 0 net192
rlabel metal2 37128 28896 37128 28896 0 net193
rlabel metal2 37800 27944 37800 27944 0 net194
rlabel metal2 38080 76328 38080 76328 0 net195
rlabel metal2 33488 75880 33488 75880 0 net196
rlabel metal2 39760 75656 39760 75656 0 net197
rlabel metal2 31864 52024 31864 52024 0 net198
rlabel metal2 39816 27776 39816 27776 0 net199
rlabel metal3 32816 4984 32816 4984 0 net2
rlabel metal2 46648 5768 46648 5768 0 net20
rlabel metal2 30184 51856 30184 51856 0 net200
rlabel metal2 59192 42364 59192 42364 0 net201
rlabel metal2 66248 75432 66248 75432 0 net202
rlabel metal2 66808 71876 66808 71876 0 net203
rlabel metal1 68096 77112 68096 77112 0 net204
rlabel metal2 68488 37856 68488 37856 0 net205
rlabel metal2 67872 75992 67872 75992 0 net206
rlabel metal2 69384 76552 69384 76552 0 net207
rlabel metal2 71064 76776 71064 76776 0 net208
rlabel metal2 72408 39928 72408 39928 0 net209
rlabel metal2 46088 6328 46088 6328 0 net21
rlabel metal2 71624 71876 71624 71876 0 net210
rlabel metal2 72296 76384 72296 76384 0 net211
rlabel metal2 60984 40880 60984 40880 0 net212
rlabel metal2 72912 76552 72912 76552 0 net213
rlabel metal2 73136 75432 73136 75432 0 net214
rlabel metal2 74424 71876 74424 71876 0 net215
rlabel metal3 74256 73976 74256 73976 0 net216
rlabel metal2 75432 76720 75432 76720 0 net217
rlabel metal4 76048 55440 76048 55440 0 net218
rlabel metal3 75712 75768 75712 75768 0 net219
rlabel metal2 48216 4312 48216 4312 0 net22
rlabel metal3 74648 68824 74648 68824 0 net220
rlabel metal3 74368 76104 74368 76104 0 net221
rlabel metal3 70672 74984 70672 74984 0 net222
rlabel metal2 61320 40096 61320 40096 0 net223
rlabel metal3 74760 75656 74760 75656 0 net224
rlabel metal2 75376 61320 75376 61320 0 net225
rlabel metal2 61992 42364 61992 42364 0 net226
rlabel metal2 62384 75432 62384 75432 0 net227
rlabel metal2 63000 71876 63000 71876 0 net228
rlabel metal2 63616 55440 63616 55440 0 net229
rlabel metal2 21336 2464 21336 2464 0 net23
rlabel metal2 64792 71624 64792 71624 0 net230
rlabel metal2 65184 71848 65184 71848 0 net231
rlabel metal2 65688 71876 65688 71876 0 net232
rlabel metal2 12936 74032 12936 74032 0 net233
rlabel metal2 18200 74200 18200 74200 0 net234
rlabel metal2 19880 74312 19880 74312 0 net235
rlabel metal3 15568 74760 15568 74760 0 net236
rlabel metal2 22792 74424 22792 74424 0 net237
rlabel metal3 24248 75768 24248 75768 0 net238
rlabel metal2 23912 75824 23912 75824 0 net239
rlabel metal2 47992 4368 47992 4368 0 net24
rlabel metal3 14224 23464 14224 23464 0 net240
rlabel metal3 13160 75656 13160 75656 0 net241
rlabel metal3 11760 74872 11760 74872 0 net242
rlabel metal2 8344 50344 8344 50344 0 net243
rlabel metal3 15232 74088 15232 74088 0 net244
rlabel metal3 13832 22456 13832 22456 0 net245
rlabel metal2 17864 73640 17864 73640 0 net246
rlabel metal2 16408 76384 16408 76384 0 net247
rlabel metal2 17864 75320 17864 75320 0 net248
rlabel metal2 52640 5768 52640 5768 0 net249
rlabel metal2 48664 6328 48664 6328 0 net25
rlabel metal2 59864 6272 59864 6272 0 net250
rlabel metal2 60312 6664 60312 6664 0 net251
rlabel metal2 63224 4816 63224 4816 0 net252
rlabel metal2 65688 3976 65688 3976 0 net253
rlabel metal3 65576 5208 65576 5208 0 net254
rlabel metal2 63448 6328 63448 6328 0 net255
rlabel metal2 64456 5992 64456 5992 0 net256
rlabel metal2 67480 4760 67480 4760 0 net257
rlabel metal2 70280 3584 70280 3584 0 net258
rlabel metal3 52024 9296 52024 9296 0 net259
rlabel metal2 23464 3024 23464 3024 0 net26
rlabel metal2 55048 4256 55048 4256 0 net260
rlabel metal2 68488 5656 68488 5656 0 net261
rlabel metal2 67032 7504 67032 7504 0 net262
rlabel metal2 68152 6664 68152 6664 0 net263
rlabel metal2 71064 4816 71064 4816 0 net264
rlabel metal2 72296 4424 72296 4424 0 net265
rlabel metal2 70504 4088 70504 4088 0 net266
rlabel metal3 70504 6664 70504 6664 0 net267
rlabel metal3 72016 5880 72016 5880 0 net268
rlabel metal2 70504 5544 70504 5544 0 net269
rlabel metal2 28728 3864 28728 3864 0 net27
rlabel metal2 71736 7728 71736 7728 0 net270
rlabel metal2 54264 5600 54264 5600 0 net271
rlabel metal2 77336 5992 77336 5992 0 net272
rlabel metal2 75320 7560 75320 7560 0 net273
rlabel metal2 58072 3976 58072 3976 0 net274
rlabel metal2 61432 3584 61432 3584 0 net275
rlabel metal2 56840 5768 56840 5768 0 net276
rlabel metal2 56056 6272 56056 6272 0 net277
rlabel metal3 62104 4424 62104 4424 0 net278
rlabel metal2 63560 4144 63560 4144 0 net279
rlabel metal3 26432 4424 26432 4424 0 net28
rlabel metal2 60200 7168 60200 7168 0 net280
rlabel metal2 44128 18200 44128 18200 0 net281
rlabel metal3 3528 45864 3528 45864 0 net282
rlabel metal3 4088 40376 4088 40376 0 net283
rlabel metal3 4872 40488 4872 40488 0 net284
rlabel metal3 3864 40600 3864 40600 0 net285
rlabel metal2 2744 43176 2744 43176 0 net286
rlabel metal2 3528 54040 3528 54040 0 net287
rlabel metal2 2072 55720 2072 55720 0 net288
rlabel metal2 3752 56560 3752 56560 0 net289
rlabel metal2 31136 7560 31136 7560 0 net29
rlabel metal2 4480 56728 4480 56728 0 net290
rlabel metal2 2072 58856 2072 58856 0 net291
rlabel metal2 2744 59696 2744 59696 0 net292
rlabel metal2 2072 61040 2072 61040 0 net293
rlabel metal2 3416 61880 3416 61880 0 net294
rlabel metal2 3192 63560 3192 63560 0 net295
rlabel metal2 3528 64400 3528 64400 0 net296
rlabel metal2 2072 44016 2072 44016 0 net297
rlabel metal2 2072 66304 2072 66304 0 net298
rlabel metal2 3080 66696 3080 66696 0 net299
rlabel metal2 39592 7448 39592 7448 0 net3
rlabel metal2 25816 3864 25816 3864 0 net30
rlabel metal2 4088 67536 4088 67536 0 net300
rlabel metal2 2072 68880 2072 68880 0 net301
rlabel metal2 2744 69720 2744 69720 0 net302
rlabel metal3 3584 71960 3584 71960 0 net303
rlabel metal2 3528 72240 3528 72240 0 net304
rlabel metal2 4312 73360 4312 73360 0 net305
rlabel metal2 4648 74032 4648 74032 0 net306
rlabel metal2 4592 75096 4592 75096 0 net307
rlabel metal2 2072 45360 2072 45360 0 net308
rlabel metal2 4648 75712 4648 75712 0 net309
rlabel metal2 26712 4536 26712 4536 0 net31
rlabel metal2 4200 75768 4200 75768 0 net310
rlabel metal2 3416 46200 3416 46200 0 net311
rlabel metal2 2072 47880 2072 47880 0 net312
rlabel metal2 2744 48720 2744 48720 0 net313
rlabel metal2 3416 49112 3416 49112 0 net314
rlabel metal2 2856 51016 2856 51016 0 net315
rlabel metal2 3528 51856 3528 51856 0 net316
rlabel metal3 3584 53592 3584 53592 0 net317
rlabel metal2 75320 42000 75320 42000 0 net318
rlabel metal2 77896 39928 77896 39928 0 net319
rlabel metal2 27160 4144 27160 4144 0 net32
rlabel metal3 75768 9352 75768 9352 0 net320
rlabel metal2 78232 5264 78232 5264 0 net321
rlabel metal2 77224 5936 77224 5936 0 net322
rlabel metal2 76216 5544 76216 5544 0 net323
rlabel metal3 37800 74760 37800 74760 0 net324
rlabel metal3 57288 45304 57288 45304 0 net325
rlabel metal3 58296 43400 58296 43400 0 net326
rlabel metal2 57288 49140 57288 49140 0 net327
rlabel metal3 59080 42840 59080 42840 0 net328
rlabel metal2 2464 64120 2464 64120 0 net329
rlabel metal2 40040 5880 40040 5880 0 net33
rlabel metal2 2408 68236 2408 68236 0 net330
rlabel metal2 2296 65464 2296 65464 0 net331
rlabel metal2 4480 41272 4480 41272 0 net332
rlabel metal2 2408 57680 2408 57680 0 net333
rlabel metal2 3864 53144 3864 53144 0 net334
rlabel metal2 2352 53704 2352 53704 0 net335
rlabel metal3 2688 48216 2688 48216 0 net336
rlabel metal2 3192 50456 3192 50456 0 net337
rlabel metal2 2072 38472 2072 38472 0 net338
rlabel metal2 4648 72240 4648 72240 0 net339
rlabel metal2 4368 4536 4368 4536 0 net34
rlabel metal2 5264 76552 5264 76552 0 net340
rlabel metal3 5376 72520 5376 72520 0 net341
rlabel metal2 1904 71624 1904 71624 0 net342
rlabel metal3 21560 76664 21560 76664 0 net343
rlabel metal2 23128 76160 23128 76160 0 net344
rlabel metal2 23464 75096 23464 75096 0 net345
rlabel metal2 24136 75544 24136 75544 0 net346
rlabel metal2 24808 76664 24808 76664 0 net347
rlabel metal2 25480 76664 25480 76664 0 net348
rlabel metal2 26152 76664 26152 76664 0 net349
rlabel metal2 10920 3976 10920 3976 0 net35
rlabel metal2 26824 76664 26824 76664 0 net350
rlabel metal2 27496 76664 27496 76664 0 net351
rlabel metal2 28392 77280 28392 77280 0 net352
rlabel metal2 28840 76664 28840 76664 0 net353
rlabel metal2 29512 76664 29512 76664 0 net354
rlabel metal2 30184 76664 30184 76664 0 net355
rlabel metal2 30856 76664 30856 76664 0 net356
rlabel metal2 31472 76664 31472 76664 0 net357
rlabel metal2 32200 76664 32200 76664 0 net358
rlabel metal2 7448 3640 7448 3640 0 net36
rlabel metal2 8120 2800 8120 2800 0 net37
rlabel metal3 12712 3304 12712 3304 0 net38
rlabel metal2 19768 5544 19768 5544 0 net39
rlabel metal2 27832 3136 27832 3136 0 net4
rlabel metal3 13104 3192 13104 3192 0 net40
rlabel metal2 9912 3080 9912 3080 0 net41
rlabel metal2 10584 2856 10584 2856 0 net42
rlabel metal2 11928 3136 11928 3136 0 net43
rlabel metal2 21672 3472 21672 3472 0 net44
rlabel metal2 3640 4760 3640 4760 0 net45
rlabel metal2 20440 5264 20440 5264 0 net46
rlabel metal2 21896 5264 21896 5264 0 net47
rlabel metal2 15064 3864 15064 3864 0 net48
rlabel metal2 18648 5208 18648 5208 0 net49
rlabel metal2 28952 3192 28952 3192 0 net5
rlabel metal2 16408 3024 16408 3024 0 net50
rlabel metal2 18200 3808 18200 3808 0 net51
rlabel metal3 23128 3304 23128 3304 0 net52
rlabel metal3 22176 3528 22176 3528 0 net53
rlabel metal2 22680 5768 22680 5768 0 net54
rlabel metal2 29232 5096 29232 5096 0 net55
rlabel metal2 4984 5488 4984 5488 0 net56
rlabel metal3 24696 5264 24696 5264 0 net57
rlabel metal2 21000 8568 21000 8568 0 net58
rlabel metal2 5656 5208 5656 5208 0 net59
rlabel metal2 29680 3416 29680 3416 0 net6
rlabel metal2 4312 3752 4312 3752 0 net60
rlabel metal2 8008 5040 8008 5040 0 net61
rlabel metal2 7336 5040 7336 5040 0 net62
rlabel metal2 4928 3416 4928 3416 0 net63
rlabel metal2 6048 3416 6048 3416 0 net64
rlabel metal3 7588 3304 7588 3304 0 net65
rlabel metal2 51912 9408 51912 9408 0 net66
rlabel metal2 52304 3304 52304 3304 0 net67
rlabel metal2 51912 4928 51912 4928 0 net68
rlabel metal2 53480 5376 53480 5376 0 net69
rlabel metal2 30296 3808 30296 3808 0 net7
rlabel metal2 2744 4200 2744 4200 0 net70
rlabel metal3 36288 15960 36288 15960 0 net71
rlabel metal3 5236 15400 5236 15400 0 net72
rlabel metal2 2072 16128 2072 16128 0 net73
rlabel metal2 2072 17696 2072 17696 0 net74
rlabel metal2 2072 18424 2072 18424 0 net75
rlabel metal2 2072 19712 2072 19712 0 net76
rlabel metal2 2072 20776 2072 20776 0 net77
rlabel metal2 48216 21728 48216 21728 0 net78
rlabel metal2 2072 22904 2072 22904 0 net79
rlabel metal2 38696 3808 38696 3808 0 net8
rlabel metal2 2072 23856 2072 23856 0 net80
rlabel metal2 2072 4088 2072 4088 0 net81
rlabel metal2 2072 25480 2072 25480 0 net82
rlabel metal2 2072 26208 2072 26208 0 net83
rlabel metal2 2072 27104 2072 27104 0 net84
rlabel metal2 2072 28616 2072 28616 0 net85
rlabel metal2 44744 29512 44744 29512 0 net86
rlabel metal2 44296 31080 44296 31080 0 net87
rlabel metal2 2072 31696 2072 31696 0 net88
rlabel metal2 28504 32368 28504 32368 0 net89
rlabel metal2 39032 2436 39032 2436 0 net9
rlabel metal2 44296 34216 44296 34216 0 net90
rlabel metal2 44856 34720 44856 34720 0 net91
rlabel metal2 2072 5432 2072 5432 0 net92
rlabel metal2 44296 36064 44296 36064 0 net93
rlabel metal2 26936 36848 26936 36848 0 net94
rlabel metal2 2016 6104 2016 6104 0 net95
rlabel metal2 33824 16744 33824 16744 0 net96
rlabel metal2 2072 8260 2072 8260 0 net97
rlabel metal2 2072 10080 2072 10080 0 net98
rlabel metal3 32536 9912 32536 9912 0 net99
rlabel metal3 2086 38136 2086 38136 0 ram_gwenb[0]
rlabel metal3 1358 39256 1358 39256 0 ram_gwenb[1]
rlabel metal3 1358 40376 1358 40376 0 ram_gwenb[2]
rlabel metal3 1358 41496 1358 41496 0 ram_gwenb[3]
rlabel metal2 2408 2856 2408 2856 0 ram_rdata[0]
rlabel metal2 1736 13608 1736 13608 0 ram_rdata[10]
rlabel metal2 1736 14952 1736 14952 0 ram_rdata[11]
rlabel metal2 1736 15848 1736 15848 0 ram_rdata[12]
rlabel metal2 1736 17192 1736 17192 0 ram_rdata[13]
rlabel metal2 1736 18200 1736 18200 0 ram_rdata[14]
rlabel metal3 1246 19096 1246 19096 0 ram_rdata[15]
rlabel metal2 1736 20384 1736 20384 0 ram_rdata[16]
rlabel metal2 1736 21448 1736 21448 0 ram_rdata[17]
rlabel metal2 1736 22792 1736 22792 0 ram_rdata[18]
rlabel metal2 1736 23632 1736 23632 0 ram_rdata[19]
rlabel metal2 1848 3864 1848 3864 0 ram_rdata[1]
rlabel metal2 1736 24976 1736 24976 0 ram_rdata[20]
rlabel metal2 1736 26040 1736 26040 0 ram_rdata[21]
rlabel metal3 1246 26936 1246 26936 0 ram_rdata[22]
rlabel metal2 1736 28336 1736 28336 0 ram_rdata[23]
rlabel metal2 1736 29288 1736 29288 0 ram_rdata[24]
rlabel metal2 1736 30632 1736 30632 0 ram_rdata[25]
rlabel metal2 1736 31528 1736 31528 0 ram_rdata[26]
rlabel metal2 1736 32816 1736 32816 0 ram_rdata[27]
rlabel metal2 1736 33880 1736 33880 0 ram_rdata[28]
rlabel metal3 1246 34776 1246 34776 0 ram_rdata[29]
rlabel metal2 1736 4816 1736 4816 0 ram_rdata[2]
rlabel metal2 1736 36120 1736 36120 0 ram_rdata[30]
rlabel metal2 1736 37128 1736 37128 0 ram_rdata[31]
rlabel metal2 1736 5768 1736 5768 0 ram_rdata[3]
rlabel metal2 1736 7112 1736 7112 0 ram_rdata[4]
rlabel metal2 1736 8008 1736 8008 0 ram_rdata[5]
rlabel metal2 1736 9352 1736 9352 0 ram_rdata[6]
rlabel metal2 1736 10360 1736 10360 0 ram_rdata[7]
rlabel metal3 1246 11256 1246 11256 0 ram_rdata[8]
rlabel metal2 1736 12600 1736 12600 0 ram_rdata[9]
rlabel metal2 44296 22792 44296 22792 0 ram_ready
rlabel metal3 1358 42616 1358 42616 0 ram_wenb[0]
rlabel metal3 1358 53816 1358 53816 0 ram_wenb[10]
rlabel metal3 1750 54936 1750 54936 0 ram_wenb[11]
rlabel metal3 1358 56056 1358 56056 0 ram_wenb[12]
rlabel metal3 1358 57176 1358 57176 0 ram_wenb[13]
rlabel metal3 1750 58296 1750 58296 0 ram_wenb[14]
rlabel metal3 1358 59416 1358 59416 0 ram_wenb[15]
rlabel metal3 1750 60536 1750 60536 0 ram_wenb[16]
rlabel metal3 1358 61656 1358 61656 0 ram_wenb[17]
rlabel metal3 1358 62776 1358 62776 0 ram_wenb[18]
rlabel metal3 1358 63896 1358 63896 0 ram_wenb[19]
rlabel metal3 1750 43736 1750 43736 0 ram_wenb[1]
rlabel metal3 1750 65016 1750 65016 0 ram_wenb[20]
rlabel metal3 1358 66136 1358 66136 0 ram_wenb[21]
rlabel metal3 1358 67256 1358 67256 0 ram_wenb[22]
rlabel metal3 1750 68376 1750 68376 0 ram_wenb[23]
rlabel metal3 1358 69496 1358 69496 0 ram_wenb[24]
rlabel metal3 1358 70616 1358 70616 0 ram_wenb[25]
rlabel metal3 1358 71736 1358 71736 0 ram_wenb[26]
rlabel metal3 1358 72856 1358 72856 0 ram_wenb[27]
rlabel metal3 1358 73976 1358 73976 0 ram_wenb[28]
rlabel metal3 1358 75096 1358 75096 0 ram_wenb[29]
rlabel metal3 1750 44856 1750 44856 0 ram_wenb[2]
rlabel metal3 1358 76216 1358 76216 0 ram_wenb[30]
rlabel metal3 1470 77336 1470 77336 0 ram_wenb[31]
rlabel metal3 1358 45976 1358 45976 0 ram_wenb[3]
rlabel metal3 1750 47096 1750 47096 0 ram_wenb[4]
rlabel metal3 1358 48216 1358 48216 0 ram_wenb[5]
rlabel metal3 1358 49336 1358 49336 0 ram_wenb[6]
rlabel metal3 1358 50456 1358 50456 0 ram_wenb[7]
rlabel metal3 1358 51576 1358 51576 0 ram_wenb[8]
rlabel metal3 1358 52696 1358 52696 0 ram_wenb[9]
rlabel metal3 74256 3416 74256 3416 0 resetn
rlabel metal2 78008 42000 78008 42000 0 simpleuart_dat_re
rlabel metal2 76664 40768 76664 40768 0 simpleuart_dat_we
rlabel metal3 76930 728 76930 728 0 simpleuart_div_we[0]
rlabel metal2 75656 6776 75656 6776 0 simpleuart_div_we[1]
rlabel metal2 73920 4872 73920 4872 0 simpleuart_div_we[2]
rlabel metal3 78834 4088 78834 4088 0 simpleuart_div_we[3]
rlabel metal2 78120 43008 78120 43008 0 simpleuart_reg_dat_do[0]
rlabel metal2 78232 54824 78232 54824 0 simpleuart_reg_dat_do[10]
rlabel metal2 78232 55832 78232 55832 0 simpleuart_reg_dat_do[11]
rlabel metal3 78722 56728 78722 56728 0 simpleuart_reg_dat_do[12]
rlabel metal2 78232 58016 78232 58016 0 simpleuart_reg_dat_do[13]
rlabel metal2 78232 59080 78232 59080 0 simpleuart_reg_dat_do[14]
rlabel metal2 78232 60424 78232 60424 0 simpleuart_reg_dat_do[15]
rlabel metal2 78232 61264 78232 61264 0 simpleuart_reg_dat_do[16]
rlabel metal2 78232 62608 78232 62608 0 simpleuart_reg_dat_do[17]
rlabel metal2 78232 63672 78232 63672 0 simpleuart_reg_dat_do[18]
rlabel metal3 78722 64568 78722 64568 0 simpleuart_reg_dat_do[19]
rlabel metal2 78232 44744 78232 44744 0 simpleuart_reg_dat_do[1]
rlabel metal2 78232 65856 78232 65856 0 simpleuart_reg_dat_do[20]
rlabel metal2 78232 66920 78232 66920 0 simpleuart_reg_dat_do[21]
rlabel metal2 78232 68264 78232 68264 0 simpleuart_reg_dat_do[22]
rlabel metal2 78232 69104 78232 69104 0 simpleuart_reg_dat_do[23]
rlabel metal2 78232 70448 78232 70448 0 simpleuart_reg_dat_do[24]
rlabel metal2 78232 71512 78232 71512 0 simpleuart_reg_dat_do[25]
rlabel metal3 78722 72408 78722 72408 0 simpleuart_reg_dat_do[26]
rlabel metal3 78722 73528 78722 73528 0 simpleuart_reg_dat_do[27]
rlabel metal2 78120 74536 78120 74536 0 simpleuart_reg_dat_do[28]
rlabel metal2 78120 75544 78120 75544 0 simpleuart_reg_dat_do[29]
rlabel metal2 78232 45640 78232 45640 0 simpleuart_reg_dat_do[2]
rlabel metal2 76944 75096 76944 75096 0 simpleuart_reg_dat_do[30]
rlabel metal2 78008 76104 78008 76104 0 simpleuart_reg_dat_do[31]
rlabel metal2 78232 46984 78232 46984 0 simpleuart_reg_dat_do[3]
rlabel metal2 78232 47992 78232 47992 0 simpleuart_reg_dat_do[4]
rlabel metal3 78722 48888 78722 48888 0 simpleuart_reg_dat_do[5]
rlabel metal3 77952 50456 77952 50456 0 simpleuart_reg_dat_do[6]
rlabel metal2 78232 51240 78232 51240 0 simpleuart_reg_dat_do[7]
rlabel metal2 78232 52584 78232 52584 0 simpleuart_reg_dat_do[8]
rlabel metal2 78232 53480 78232 53480 0 simpleuart_reg_dat_do[9]
rlabel metal2 77224 77728 77224 77728 0 simpleuart_reg_dat_wait
rlabel metal3 78386 5208 78386 5208 0 simpleuart_reg_div_do[0]
rlabel metal3 78232 16856 78232 16856 0 simpleuart_reg_div_do[10]
rlabel metal3 78386 17528 78386 17528 0 simpleuart_reg_div_do[11]
rlabel metal2 78232 18144 78232 18144 0 simpleuart_reg_div_do[12]
rlabel metal2 74872 19880 74872 19880 0 simpleuart_reg_div_do[13]
rlabel metal3 77784 19096 77784 19096 0 simpleuart_reg_div_do[14]
rlabel metal3 78344 19208 78344 19208 0 simpleuart_reg_div_do[15]
rlabel metal2 78232 21952 78232 21952 0 simpleuart_reg_div_do[16]
rlabel metal2 76216 22904 76216 22904 0 simpleuart_reg_div_do[17]
rlabel metal2 71960 25816 71960 25816 0 simpleuart_reg_div_do[18]
rlabel metal3 75712 26600 75712 26600 0 simpleuart_reg_div_do[19]
rlabel metal2 76888 7336 76888 7336 0 simpleuart_reg_div_do[1]
rlabel metal2 78232 26544 78232 26544 0 simpleuart_reg_div_do[20]
rlabel metal3 73192 28616 73192 28616 0 simpleuart_reg_div_do[21]
rlabel metal2 75656 28168 75656 28168 0 simpleuart_reg_div_do[22]
rlabel metal2 75096 30576 75096 30576 0 simpleuart_reg_div_do[23]
rlabel metal2 74872 31640 74872 31640 0 simpleuart_reg_div_do[24]
rlabel metal2 70952 29176 70952 29176 0 simpleuart_reg_div_do[25]
rlabel metal2 74760 34832 74760 34832 0 simpleuart_reg_div_do[26]
rlabel metal3 78778 35448 78778 35448 0 simpleuart_reg_div_do[27]
rlabel metal2 77672 36456 77672 36456 0 simpleuart_reg_div_do[28]
rlabel metal2 75488 36456 75488 36456 0 simpleuart_reg_div_do[29]
rlabel metal2 77560 7784 77560 7784 0 simpleuart_reg_div_do[2]
rlabel metal3 78498 38808 78498 38808 0 simpleuart_reg_div_do[30]
rlabel metal2 76496 42728 76496 42728 0 simpleuart_reg_div_do[31]
rlabel metal2 78232 8316 78232 8316 0 simpleuart_reg_div_do[3]
rlabel metal3 78722 9688 78722 9688 0 simpleuart_reg_div_do[4]
rlabel metal2 78232 11032 78232 11032 0 simpleuart_reg_div_do[5]
rlabel metal2 78232 12040 78232 12040 0 simpleuart_reg_div_do[6]
rlabel metal2 78120 13608 78120 13608 0 simpleuart_reg_div_do[7]
rlabel metal2 78232 14280 78232 14280 0 simpleuart_reg_div_do[8]
rlabel metal2 78232 15624 78232 15624 0 simpleuart_reg_div_do[9]
rlabel metal2 34104 77490 34104 77490 0 spimem_rdata[0]
rlabel metal2 40936 76664 40936 76664 0 spimem_rdata[10]
rlabel metal2 41496 77490 41496 77490 0 spimem_rdata[11]
rlabel metal2 42280 76664 42280 76664 0 spimem_rdata[12]
rlabel metal2 43624 76832 43624 76832 0 spimem_rdata[13]
rlabel metal2 44520 76832 44520 76832 0 spimem_rdata[14]
rlabel metal3 44800 76664 44800 76664 0 spimem_rdata[15]
rlabel metal2 45192 76216 45192 76216 0 spimem_rdata[16]
rlabel metal2 46312 76832 46312 76832 0 spimem_rdata[17]
rlabel metal3 46816 76664 46816 76664 0 spimem_rdata[18]
rlabel metal2 47096 76104 47096 76104 0 spimem_rdata[19]
rlabel metal2 34776 77154 34776 77154 0 spimem_rdata[1]
rlabel metal2 48328 76832 48328 76832 0 spimem_rdata[20]
rlabel metal3 48720 76664 48720 76664 0 spimem_rdata[21]
rlabel metal2 50120 76832 50120 76832 0 spimem_rdata[22]
rlabel metal2 49560 77490 49560 77490 0 spimem_rdata[23]
rlabel metal2 50232 77938 50232 77938 0 spimem_rdata[24]
rlabel metal2 52136 76888 52136 76888 0 spimem_rdata[25]
rlabel metal2 53032 76832 53032 76832 0 spimem_rdata[26]
rlabel metal2 52248 77490 52248 77490 0 spimem_rdata[27]
rlabel metal3 53424 76664 53424 76664 0 spimem_rdata[28]
rlabel metal2 53816 76104 53816 76104 0 spimem_rdata[29]
rlabel metal2 35504 75768 35504 75768 0 spimem_rdata[2]
rlabel metal2 54712 76104 54712 76104 0 spimem_rdata[30]
rlabel metal2 55608 76048 55608 76048 0 spimem_rdata[31]
rlabel metal2 36344 76720 36344 76720 0 spimem_rdata[3]
rlabel metal2 36792 77938 36792 77938 0 spimem_rdata[4]
rlabel metal2 37576 76664 37576 76664 0 spimem_rdata[5]
rlabel metal2 38248 76104 38248 76104 0 spimem_rdata[6]
rlabel metal2 39032 76160 39032 76160 0 spimem_rdata[7]
rlabel metal2 39368 76664 39368 76664 0 spimem_rdata[8]
rlabel metal2 40152 77938 40152 77938 0 spimem_rdata[9]
rlabel metal2 32760 77490 32760 77490 0 spimem_ready
rlabel metal2 33432 77770 33432 77770 0 spimem_valid
rlabel metal3 58800 75544 58800 75544 0 spimemio_cfgreg_do[0]
rlabel metal2 65072 75768 65072 75768 0 spimemio_cfgreg_do[10]
rlabel metal2 66472 76832 66472 76832 0 spimemio_cfgreg_do[11]
rlabel metal2 67144 76888 67144 76888 0 spimemio_cfgreg_do[12]
rlabel metal2 67816 76832 67816 76832 0 spimemio_cfgreg_do[13]
rlabel metal2 68488 76832 68488 76832 0 spimemio_cfgreg_do[14]
rlabel metal3 68768 76664 68768 76664 0 spimemio_cfgreg_do[15]
rlabel metal2 70280 76888 70280 76888 0 spimemio_cfgreg_do[16]
rlabel metal3 70336 76552 70336 76552 0 spimemio_cfgreg_do[17]
rlabel metal2 71848 76720 71848 76720 0 spimemio_cfgreg_do[18]
rlabel metal2 72632 76832 72632 76832 0 spimemio_cfgreg_do[19]
rlabel metal3 59752 75432 59752 75432 0 spimemio_cfgreg_do[1]
rlabel metal2 73192 76496 73192 76496 0 spimemio_cfgreg_do[20]
rlabel metal2 72408 77490 72408 77490 0 spimemio_cfgreg_do[21]
rlabel metal3 73584 76664 73584 76664 0 spimemio_cfgreg_do[22]
rlabel metal2 74984 76496 74984 76496 0 spimemio_cfgreg_do[23]
rlabel metal2 75768 76776 75768 76776 0 spimemio_cfgreg_do[24]
rlabel metal2 76440 76944 76440 76944 0 spimemio_cfgreg_do[25]
rlabel metal2 76216 76552 76216 76552 0 spimemio_cfgreg_do[26]
rlabel metal2 76888 76552 76888 76552 0 spimemio_cfgreg_do[27]
rlabel metal2 77840 76440 77840 76440 0 spimemio_cfgreg_do[28]
rlabel metal2 77392 74872 77392 74872 0 spimemio_cfgreg_do[29]
rlabel metal2 62552 75656 62552 75656 0 spimemio_cfgreg_do[2]
rlabel metal2 75432 75768 75432 75768 0 spimemio_cfgreg_do[30]
rlabel metal2 75992 75096 75992 75096 0 spimemio_cfgreg_do[31]
rlabel metal3 60760 75544 60760 75544 0 spimemio_cfgreg_do[3]
rlabel metal2 62216 75152 62216 75152 0 spimemio_cfgreg_do[4]
rlabel metal2 62664 76776 62664 76776 0 spimemio_cfgreg_do[5]
rlabel metal2 63336 76832 63336 76832 0 spimemio_cfgreg_do[6]
rlabel metal2 64008 76888 64008 76888 0 spimemio_cfgreg_do[7]
rlabel metal2 64680 76832 64680 76832 0 spimemio_cfgreg_do[8]
rlabel metal2 65352 76832 65352 76832 0 spimemio_cfgreg_do[9]
rlabel metal2 55608 78498 55608 78498 0 spimemio_cfgreg_we[0]
rlabel metal2 56728 76608 56728 76608 0 spimemio_cfgreg_we[1]
rlabel metal2 56952 77938 56952 77938 0 spimemio_cfgreg_we[2]
rlabel metal2 57624 76986 57624 76986 0 spimemio_cfgreg_we[3]
<< properties >>
string FIXED_BBOX 0 0 80000 80000
<< end >>

magic
tech gf180mcuD
magscale 1 5
timestamp 1702205593
<< obsm1 >>
rect 672 1538 79791 138406
<< metal2 >>
rect 3584 139600 3640 140000
rect 10192 139600 10248 140000
rect 16800 139600 16856 140000
rect 23408 139600 23464 140000
rect 30016 139600 30072 140000
rect 36624 139600 36680 140000
rect 43232 139600 43288 140000
rect 49840 139600 49896 140000
rect 56448 139600 56504 140000
rect 63056 139600 63112 140000
rect 69664 139600 69720 140000
rect 76272 139600 76328 140000
<< obsm2 >>
rect 686 139570 3554 139600
rect 3670 139570 10162 139600
rect 10278 139570 16770 139600
rect 16886 139570 23378 139600
rect 23494 139570 29986 139600
rect 30102 139570 36594 139600
rect 36710 139570 43202 139600
rect 43318 139570 49810 139600
rect 49926 139570 56418 139600
rect 56534 139570 63026 139600
rect 63142 139570 69634 139600
rect 69750 139570 76242 139600
rect 76358 139570 79954 139600
rect 686 1353 79954 139570
<< metal3 >>
rect 0 138432 400 138488
rect 0 137088 400 137144
rect 79600 136528 80000 136584
rect 79600 135968 80000 136024
rect 0 135744 400 135800
rect 79600 135408 80000 135464
rect 79600 134848 80000 134904
rect 0 134400 400 134456
rect 79600 134288 80000 134344
rect 79600 133728 80000 133784
rect 79600 133168 80000 133224
rect 0 133056 400 133112
rect 79600 132608 80000 132664
rect 79600 132048 80000 132104
rect 0 131712 400 131768
rect 79600 131488 80000 131544
rect 79600 130928 80000 130984
rect 0 130368 400 130424
rect 79600 130368 80000 130424
rect 79600 129808 80000 129864
rect 79600 129248 80000 129304
rect 0 129024 400 129080
rect 79600 128688 80000 128744
rect 79600 128128 80000 128184
rect 0 127680 400 127736
rect 79600 127568 80000 127624
rect 79600 127008 80000 127064
rect 79600 126448 80000 126504
rect 0 126336 400 126392
rect 79600 125888 80000 125944
rect 79600 125328 80000 125384
rect 0 124992 400 125048
rect 79600 124768 80000 124824
rect 79600 124208 80000 124264
rect 0 123648 400 123704
rect 79600 123648 80000 123704
rect 79600 123088 80000 123144
rect 79600 122528 80000 122584
rect 0 122304 400 122360
rect 79600 121968 80000 122024
rect 79600 121408 80000 121464
rect 0 120960 400 121016
rect 79600 120848 80000 120904
rect 79600 120288 80000 120344
rect 79600 119728 80000 119784
rect 0 119616 400 119672
rect 79600 119168 80000 119224
rect 79600 118608 80000 118664
rect 0 118272 400 118328
rect 79600 118048 80000 118104
rect 79600 117488 80000 117544
rect 0 116928 400 116984
rect 79600 116928 80000 116984
rect 79600 116368 80000 116424
rect 79600 115808 80000 115864
rect 0 115584 400 115640
rect 79600 115248 80000 115304
rect 79600 114688 80000 114744
rect 0 114240 400 114296
rect 79600 114128 80000 114184
rect 79600 113568 80000 113624
rect 79600 113008 80000 113064
rect 0 112896 400 112952
rect 79600 112448 80000 112504
rect 79600 111888 80000 111944
rect 0 111552 400 111608
rect 79600 111328 80000 111384
rect 79600 110768 80000 110824
rect 0 110208 400 110264
rect 79600 110208 80000 110264
rect 79600 109648 80000 109704
rect 79600 109088 80000 109144
rect 0 108864 400 108920
rect 79600 108528 80000 108584
rect 79600 107968 80000 108024
rect 0 107520 400 107576
rect 79600 107408 80000 107464
rect 79600 106848 80000 106904
rect 79600 106288 80000 106344
rect 0 106176 400 106232
rect 79600 105728 80000 105784
rect 79600 105168 80000 105224
rect 0 104832 400 104888
rect 79600 104608 80000 104664
rect 79600 104048 80000 104104
rect 0 103488 400 103544
rect 79600 103488 80000 103544
rect 79600 102928 80000 102984
rect 79600 102368 80000 102424
rect 0 102144 400 102200
rect 79600 101808 80000 101864
rect 79600 101248 80000 101304
rect 0 100800 400 100856
rect 79600 100688 80000 100744
rect 79600 100128 80000 100184
rect 79600 99568 80000 99624
rect 0 99456 400 99512
rect 79600 99008 80000 99064
rect 79600 98448 80000 98504
rect 0 98112 400 98168
rect 79600 97888 80000 97944
rect 79600 97328 80000 97384
rect 0 96768 400 96824
rect 79600 96768 80000 96824
rect 79600 96208 80000 96264
rect 79600 95648 80000 95704
rect 0 95424 400 95480
rect 79600 95088 80000 95144
rect 79600 94528 80000 94584
rect 0 94080 400 94136
rect 79600 93968 80000 94024
rect 79600 93408 80000 93464
rect 79600 92848 80000 92904
rect 0 92736 400 92792
rect 79600 92288 80000 92344
rect 79600 91728 80000 91784
rect 0 91392 400 91448
rect 79600 91168 80000 91224
rect 79600 90608 80000 90664
rect 0 90048 400 90104
rect 79600 90048 80000 90104
rect 79600 89488 80000 89544
rect 79600 88928 80000 88984
rect 0 88704 400 88760
rect 79600 88368 80000 88424
rect 79600 87808 80000 87864
rect 0 87360 400 87416
rect 79600 87248 80000 87304
rect 79600 86688 80000 86744
rect 79600 86128 80000 86184
rect 0 86016 400 86072
rect 79600 85568 80000 85624
rect 79600 85008 80000 85064
rect 0 84672 400 84728
rect 79600 84448 80000 84504
rect 79600 83888 80000 83944
rect 0 83328 400 83384
rect 79600 83328 80000 83384
rect 79600 82768 80000 82824
rect 79600 82208 80000 82264
rect 0 81984 400 82040
rect 79600 81648 80000 81704
rect 79600 81088 80000 81144
rect 0 80640 400 80696
rect 79600 80528 80000 80584
rect 79600 79968 80000 80024
rect 79600 79408 80000 79464
rect 0 79296 400 79352
rect 79600 78848 80000 78904
rect 79600 78288 80000 78344
rect 0 77952 400 78008
rect 79600 77728 80000 77784
rect 79600 77168 80000 77224
rect 0 76608 400 76664
rect 79600 76608 80000 76664
rect 79600 76048 80000 76104
rect 79600 75488 80000 75544
rect 0 75264 400 75320
rect 79600 74928 80000 74984
rect 79600 74368 80000 74424
rect 0 73920 400 73976
rect 79600 73808 80000 73864
rect 79600 73248 80000 73304
rect 79600 72688 80000 72744
rect 0 72576 400 72632
rect 79600 72128 80000 72184
rect 79600 71568 80000 71624
rect 0 71232 400 71288
rect 79600 71008 80000 71064
rect 79600 70448 80000 70504
rect 0 69888 400 69944
rect 79600 69888 80000 69944
rect 79600 69328 80000 69384
rect 79600 68768 80000 68824
rect 0 68544 400 68600
rect 79600 68208 80000 68264
rect 79600 67648 80000 67704
rect 0 67200 400 67256
rect 79600 67088 80000 67144
rect 79600 66528 80000 66584
rect 79600 65968 80000 66024
rect 0 65856 400 65912
rect 79600 65408 80000 65464
rect 79600 64848 80000 64904
rect 0 64512 400 64568
rect 79600 64288 80000 64344
rect 79600 63728 80000 63784
rect 0 63168 400 63224
rect 79600 63168 80000 63224
rect 79600 62608 80000 62664
rect 79600 62048 80000 62104
rect 0 61824 400 61880
rect 79600 61488 80000 61544
rect 79600 60928 80000 60984
rect 0 60480 400 60536
rect 79600 60368 80000 60424
rect 79600 59808 80000 59864
rect 79600 59248 80000 59304
rect 0 59136 400 59192
rect 79600 58688 80000 58744
rect 79600 58128 80000 58184
rect 0 57792 400 57848
rect 79600 57568 80000 57624
rect 79600 57008 80000 57064
rect 0 56448 400 56504
rect 79600 56448 80000 56504
rect 79600 55888 80000 55944
rect 79600 55328 80000 55384
rect 0 55104 400 55160
rect 79600 54768 80000 54824
rect 79600 54208 80000 54264
rect 0 53760 400 53816
rect 79600 53648 80000 53704
rect 79600 53088 80000 53144
rect 79600 52528 80000 52584
rect 0 52416 400 52472
rect 79600 51968 80000 52024
rect 79600 51408 80000 51464
rect 0 51072 400 51128
rect 79600 50848 80000 50904
rect 79600 50288 80000 50344
rect 0 49728 400 49784
rect 79600 49728 80000 49784
rect 79600 49168 80000 49224
rect 79600 48608 80000 48664
rect 0 48384 400 48440
rect 79600 48048 80000 48104
rect 79600 47488 80000 47544
rect 0 47040 400 47096
rect 79600 46928 80000 46984
rect 79600 46368 80000 46424
rect 79600 45808 80000 45864
rect 0 45696 400 45752
rect 79600 45248 80000 45304
rect 79600 44688 80000 44744
rect 0 44352 400 44408
rect 79600 44128 80000 44184
rect 79600 43568 80000 43624
rect 0 43008 400 43064
rect 79600 43008 80000 43064
rect 79600 42448 80000 42504
rect 79600 41888 80000 41944
rect 0 41664 400 41720
rect 79600 41328 80000 41384
rect 79600 40768 80000 40824
rect 0 40320 400 40376
rect 79600 40208 80000 40264
rect 79600 39648 80000 39704
rect 79600 39088 80000 39144
rect 0 38976 400 39032
rect 79600 38528 80000 38584
rect 79600 37968 80000 38024
rect 0 37632 400 37688
rect 79600 37408 80000 37464
rect 79600 36848 80000 36904
rect 0 36288 400 36344
rect 79600 36288 80000 36344
rect 79600 35728 80000 35784
rect 79600 35168 80000 35224
rect 0 34944 400 35000
rect 79600 34608 80000 34664
rect 79600 34048 80000 34104
rect 0 33600 400 33656
rect 79600 33488 80000 33544
rect 79600 32928 80000 32984
rect 79600 32368 80000 32424
rect 0 32256 400 32312
rect 79600 31808 80000 31864
rect 79600 31248 80000 31304
rect 0 30912 400 30968
rect 79600 30688 80000 30744
rect 79600 30128 80000 30184
rect 0 29568 400 29624
rect 79600 29568 80000 29624
rect 79600 29008 80000 29064
rect 79600 28448 80000 28504
rect 0 28224 400 28280
rect 79600 27888 80000 27944
rect 79600 27328 80000 27384
rect 0 26880 400 26936
rect 79600 26768 80000 26824
rect 79600 26208 80000 26264
rect 79600 25648 80000 25704
rect 0 25536 400 25592
rect 79600 25088 80000 25144
rect 79600 24528 80000 24584
rect 0 24192 400 24248
rect 79600 23968 80000 24024
rect 79600 23408 80000 23464
rect 0 22848 400 22904
rect 79600 22848 80000 22904
rect 79600 22288 80000 22344
rect 79600 21728 80000 21784
rect 0 21504 400 21560
rect 79600 21168 80000 21224
rect 79600 20608 80000 20664
rect 0 20160 400 20216
rect 79600 20048 80000 20104
rect 79600 19488 80000 19544
rect 79600 18928 80000 18984
rect 0 18816 400 18872
rect 79600 18368 80000 18424
rect 79600 17808 80000 17864
rect 0 17472 400 17528
rect 79600 17248 80000 17304
rect 79600 16688 80000 16744
rect 0 16128 400 16184
rect 79600 16128 80000 16184
rect 79600 15568 80000 15624
rect 79600 15008 80000 15064
rect 0 14784 400 14840
rect 79600 14448 80000 14504
rect 79600 13888 80000 13944
rect 0 13440 400 13496
rect 79600 13328 80000 13384
rect 79600 12768 80000 12824
rect 79600 12208 80000 12264
rect 0 12096 400 12152
rect 79600 11648 80000 11704
rect 79600 11088 80000 11144
rect 0 10752 400 10808
rect 79600 10528 80000 10584
rect 79600 9968 80000 10024
rect 0 9408 400 9464
rect 79600 9408 80000 9464
rect 79600 8848 80000 8904
rect 79600 8288 80000 8344
rect 0 8064 400 8120
rect 79600 7728 80000 7784
rect 79600 7168 80000 7224
rect 0 6720 400 6776
rect 79600 6608 80000 6664
rect 79600 6048 80000 6104
rect 79600 5488 80000 5544
rect 0 5376 400 5432
rect 79600 4928 80000 4984
rect 79600 4368 80000 4424
rect 0 4032 400 4088
rect 79600 3808 80000 3864
rect 79600 3248 80000 3304
rect 0 2688 400 2744
rect 0 1344 400 1400
<< obsm3 >>
rect 430 138402 79959 138474
rect 400 137174 79959 138402
rect 430 137058 79959 137174
rect 400 136614 79959 137058
rect 400 136498 79570 136614
rect 400 136054 79959 136498
rect 400 135938 79570 136054
rect 400 135830 79959 135938
rect 430 135714 79959 135830
rect 400 135494 79959 135714
rect 400 135378 79570 135494
rect 400 134934 79959 135378
rect 400 134818 79570 134934
rect 400 134486 79959 134818
rect 430 134374 79959 134486
rect 430 134370 79570 134374
rect 400 134258 79570 134370
rect 400 133814 79959 134258
rect 400 133698 79570 133814
rect 400 133254 79959 133698
rect 400 133142 79570 133254
rect 430 133138 79570 133142
rect 430 133026 79959 133138
rect 400 132694 79959 133026
rect 400 132578 79570 132694
rect 400 132134 79959 132578
rect 400 132018 79570 132134
rect 400 131798 79959 132018
rect 430 131682 79959 131798
rect 400 131574 79959 131682
rect 400 131458 79570 131574
rect 400 131014 79959 131458
rect 400 130898 79570 131014
rect 400 130454 79959 130898
rect 430 130338 79570 130454
rect 400 129894 79959 130338
rect 400 129778 79570 129894
rect 400 129334 79959 129778
rect 400 129218 79570 129334
rect 400 129110 79959 129218
rect 430 128994 79959 129110
rect 400 128774 79959 128994
rect 400 128658 79570 128774
rect 400 128214 79959 128658
rect 400 128098 79570 128214
rect 400 127766 79959 128098
rect 430 127654 79959 127766
rect 430 127650 79570 127654
rect 400 127538 79570 127650
rect 400 127094 79959 127538
rect 400 126978 79570 127094
rect 400 126534 79959 126978
rect 400 126422 79570 126534
rect 430 126418 79570 126422
rect 430 126306 79959 126418
rect 400 125974 79959 126306
rect 400 125858 79570 125974
rect 400 125414 79959 125858
rect 400 125298 79570 125414
rect 400 125078 79959 125298
rect 430 124962 79959 125078
rect 400 124854 79959 124962
rect 400 124738 79570 124854
rect 400 124294 79959 124738
rect 400 124178 79570 124294
rect 400 123734 79959 124178
rect 430 123618 79570 123734
rect 400 123174 79959 123618
rect 400 123058 79570 123174
rect 400 122614 79959 123058
rect 400 122498 79570 122614
rect 400 122390 79959 122498
rect 430 122274 79959 122390
rect 400 122054 79959 122274
rect 400 121938 79570 122054
rect 400 121494 79959 121938
rect 400 121378 79570 121494
rect 400 121046 79959 121378
rect 430 120934 79959 121046
rect 430 120930 79570 120934
rect 400 120818 79570 120930
rect 400 120374 79959 120818
rect 400 120258 79570 120374
rect 400 119814 79959 120258
rect 400 119702 79570 119814
rect 430 119698 79570 119702
rect 430 119586 79959 119698
rect 400 119254 79959 119586
rect 400 119138 79570 119254
rect 400 118694 79959 119138
rect 400 118578 79570 118694
rect 400 118358 79959 118578
rect 430 118242 79959 118358
rect 400 118134 79959 118242
rect 400 118018 79570 118134
rect 400 117574 79959 118018
rect 400 117458 79570 117574
rect 400 117014 79959 117458
rect 430 116898 79570 117014
rect 400 116454 79959 116898
rect 400 116338 79570 116454
rect 400 115894 79959 116338
rect 400 115778 79570 115894
rect 400 115670 79959 115778
rect 430 115554 79959 115670
rect 400 115334 79959 115554
rect 400 115218 79570 115334
rect 400 114774 79959 115218
rect 400 114658 79570 114774
rect 400 114326 79959 114658
rect 430 114214 79959 114326
rect 430 114210 79570 114214
rect 400 114098 79570 114210
rect 400 113654 79959 114098
rect 400 113538 79570 113654
rect 400 113094 79959 113538
rect 400 112982 79570 113094
rect 430 112978 79570 112982
rect 430 112866 79959 112978
rect 400 112534 79959 112866
rect 400 112418 79570 112534
rect 400 111974 79959 112418
rect 400 111858 79570 111974
rect 400 111638 79959 111858
rect 430 111522 79959 111638
rect 400 111414 79959 111522
rect 400 111298 79570 111414
rect 400 110854 79959 111298
rect 400 110738 79570 110854
rect 400 110294 79959 110738
rect 430 110178 79570 110294
rect 400 109734 79959 110178
rect 400 109618 79570 109734
rect 400 109174 79959 109618
rect 400 109058 79570 109174
rect 400 108950 79959 109058
rect 430 108834 79959 108950
rect 400 108614 79959 108834
rect 400 108498 79570 108614
rect 400 108054 79959 108498
rect 400 107938 79570 108054
rect 400 107606 79959 107938
rect 430 107494 79959 107606
rect 430 107490 79570 107494
rect 400 107378 79570 107490
rect 400 106934 79959 107378
rect 400 106818 79570 106934
rect 400 106374 79959 106818
rect 400 106262 79570 106374
rect 430 106258 79570 106262
rect 430 106146 79959 106258
rect 400 105814 79959 106146
rect 400 105698 79570 105814
rect 400 105254 79959 105698
rect 400 105138 79570 105254
rect 400 104918 79959 105138
rect 430 104802 79959 104918
rect 400 104694 79959 104802
rect 400 104578 79570 104694
rect 400 104134 79959 104578
rect 400 104018 79570 104134
rect 400 103574 79959 104018
rect 430 103458 79570 103574
rect 400 103014 79959 103458
rect 400 102898 79570 103014
rect 400 102454 79959 102898
rect 400 102338 79570 102454
rect 400 102230 79959 102338
rect 430 102114 79959 102230
rect 400 101894 79959 102114
rect 400 101778 79570 101894
rect 400 101334 79959 101778
rect 400 101218 79570 101334
rect 400 100886 79959 101218
rect 430 100774 79959 100886
rect 430 100770 79570 100774
rect 400 100658 79570 100770
rect 400 100214 79959 100658
rect 400 100098 79570 100214
rect 400 99654 79959 100098
rect 400 99542 79570 99654
rect 430 99538 79570 99542
rect 430 99426 79959 99538
rect 400 99094 79959 99426
rect 400 98978 79570 99094
rect 400 98534 79959 98978
rect 400 98418 79570 98534
rect 400 98198 79959 98418
rect 430 98082 79959 98198
rect 400 97974 79959 98082
rect 400 97858 79570 97974
rect 400 97414 79959 97858
rect 400 97298 79570 97414
rect 400 96854 79959 97298
rect 430 96738 79570 96854
rect 400 96294 79959 96738
rect 400 96178 79570 96294
rect 400 95734 79959 96178
rect 400 95618 79570 95734
rect 400 95510 79959 95618
rect 430 95394 79959 95510
rect 400 95174 79959 95394
rect 400 95058 79570 95174
rect 400 94614 79959 95058
rect 400 94498 79570 94614
rect 400 94166 79959 94498
rect 430 94054 79959 94166
rect 430 94050 79570 94054
rect 400 93938 79570 94050
rect 400 93494 79959 93938
rect 400 93378 79570 93494
rect 400 92934 79959 93378
rect 400 92822 79570 92934
rect 430 92818 79570 92822
rect 430 92706 79959 92818
rect 400 92374 79959 92706
rect 400 92258 79570 92374
rect 400 91814 79959 92258
rect 400 91698 79570 91814
rect 400 91478 79959 91698
rect 430 91362 79959 91478
rect 400 91254 79959 91362
rect 400 91138 79570 91254
rect 400 90694 79959 91138
rect 400 90578 79570 90694
rect 400 90134 79959 90578
rect 430 90018 79570 90134
rect 400 89574 79959 90018
rect 400 89458 79570 89574
rect 400 89014 79959 89458
rect 400 88898 79570 89014
rect 400 88790 79959 88898
rect 430 88674 79959 88790
rect 400 88454 79959 88674
rect 400 88338 79570 88454
rect 400 87894 79959 88338
rect 400 87778 79570 87894
rect 400 87446 79959 87778
rect 430 87334 79959 87446
rect 430 87330 79570 87334
rect 400 87218 79570 87330
rect 400 86774 79959 87218
rect 400 86658 79570 86774
rect 400 86214 79959 86658
rect 400 86102 79570 86214
rect 430 86098 79570 86102
rect 430 85986 79959 86098
rect 400 85654 79959 85986
rect 400 85538 79570 85654
rect 400 85094 79959 85538
rect 400 84978 79570 85094
rect 400 84758 79959 84978
rect 430 84642 79959 84758
rect 400 84534 79959 84642
rect 400 84418 79570 84534
rect 400 83974 79959 84418
rect 400 83858 79570 83974
rect 400 83414 79959 83858
rect 430 83298 79570 83414
rect 400 82854 79959 83298
rect 400 82738 79570 82854
rect 400 82294 79959 82738
rect 400 82178 79570 82294
rect 400 82070 79959 82178
rect 430 81954 79959 82070
rect 400 81734 79959 81954
rect 400 81618 79570 81734
rect 400 81174 79959 81618
rect 400 81058 79570 81174
rect 400 80726 79959 81058
rect 430 80614 79959 80726
rect 430 80610 79570 80614
rect 400 80498 79570 80610
rect 400 80054 79959 80498
rect 400 79938 79570 80054
rect 400 79494 79959 79938
rect 400 79382 79570 79494
rect 430 79378 79570 79382
rect 430 79266 79959 79378
rect 400 78934 79959 79266
rect 400 78818 79570 78934
rect 400 78374 79959 78818
rect 400 78258 79570 78374
rect 400 78038 79959 78258
rect 430 77922 79959 78038
rect 400 77814 79959 77922
rect 400 77698 79570 77814
rect 400 77254 79959 77698
rect 400 77138 79570 77254
rect 400 76694 79959 77138
rect 430 76578 79570 76694
rect 400 76134 79959 76578
rect 400 76018 79570 76134
rect 400 75574 79959 76018
rect 400 75458 79570 75574
rect 400 75350 79959 75458
rect 430 75234 79959 75350
rect 400 75014 79959 75234
rect 400 74898 79570 75014
rect 400 74454 79959 74898
rect 400 74338 79570 74454
rect 400 74006 79959 74338
rect 430 73894 79959 74006
rect 430 73890 79570 73894
rect 400 73778 79570 73890
rect 400 73334 79959 73778
rect 400 73218 79570 73334
rect 400 72774 79959 73218
rect 400 72662 79570 72774
rect 430 72658 79570 72662
rect 430 72546 79959 72658
rect 400 72214 79959 72546
rect 400 72098 79570 72214
rect 400 71654 79959 72098
rect 400 71538 79570 71654
rect 400 71318 79959 71538
rect 430 71202 79959 71318
rect 400 71094 79959 71202
rect 400 70978 79570 71094
rect 400 70534 79959 70978
rect 400 70418 79570 70534
rect 400 69974 79959 70418
rect 430 69858 79570 69974
rect 400 69414 79959 69858
rect 400 69298 79570 69414
rect 400 68854 79959 69298
rect 400 68738 79570 68854
rect 400 68630 79959 68738
rect 430 68514 79959 68630
rect 400 68294 79959 68514
rect 400 68178 79570 68294
rect 400 67734 79959 68178
rect 400 67618 79570 67734
rect 400 67286 79959 67618
rect 430 67174 79959 67286
rect 430 67170 79570 67174
rect 400 67058 79570 67170
rect 400 66614 79959 67058
rect 400 66498 79570 66614
rect 400 66054 79959 66498
rect 400 65942 79570 66054
rect 430 65938 79570 65942
rect 430 65826 79959 65938
rect 400 65494 79959 65826
rect 400 65378 79570 65494
rect 400 64934 79959 65378
rect 400 64818 79570 64934
rect 400 64598 79959 64818
rect 430 64482 79959 64598
rect 400 64374 79959 64482
rect 400 64258 79570 64374
rect 400 63814 79959 64258
rect 400 63698 79570 63814
rect 400 63254 79959 63698
rect 430 63138 79570 63254
rect 400 62694 79959 63138
rect 400 62578 79570 62694
rect 400 62134 79959 62578
rect 400 62018 79570 62134
rect 400 61910 79959 62018
rect 430 61794 79959 61910
rect 400 61574 79959 61794
rect 400 61458 79570 61574
rect 400 61014 79959 61458
rect 400 60898 79570 61014
rect 400 60566 79959 60898
rect 430 60454 79959 60566
rect 430 60450 79570 60454
rect 400 60338 79570 60450
rect 400 59894 79959 60338
rect 400 59778 79570 59894
rect 400 59334 79959 59778
rect 400 59222 79570 59334
rect 430 59218 79570 59222
rect 430 59106 79959 59218
rect 400 58774 79959 59106
rect 400 58658 79570 58774
rect 400 58214 79959 58658
rect 400 58098 79570 58214
rect 400 57878 79959 58098
rect 430 57762 79959 57878
rect 400 57654 79959 57762
rect 400 57538 79570 57654
rect 400 57094 79959 57538
rect 400 56978 79570 57094
rect 400 56534 79959 56978
rect 430 56418 79570 56534
rect 400 55974 79959 56418
rect 400 55858 79570 55974
rect 400 55414 79959 55858
rect 400 55298 79570 55414
rect 400 55190 79959 55298
rect 430 55074 79959 55190
rect 400 54854 79959 55074
rect 400 54738 79570 54854
rect 400 54294 79959 54738
rect 400 54178 79570 54294
rect 400 53846 79959 54178
rect 430 53734 79959 53846
rect 430 53730 79570 53734
rect 400 53618 79570 53730
rect 400 53174 79959 53618
rect 400 53058 79570 53174
rect 400 52614 79959 53058
rect 400 52502 79570 52614
rect 430 52498 79570 52502
rect 430 52386 79959 52498
rect 400 52054 79959 52386
rect 400 51938 79570 52054
rect 400 51494 79959 51938
rect 400 51378 79570 51494
rect 400 51158 79959 51378
rect 430 51042 79959 51158
rect 400 50934 79959 51042
rect 400 50818 79570 50934
rect 400 50374 79959 50818
rect 400 50258 79570 50374
rect 400 49814 79959 50258
rect 430 49698 79570 49814
rect 400 49254 79959 49698
rect 400 49138 79570 49254
rect 400 48694 79959 49138
rect 400 48578 79570 48694
rect 400 48470 79959 48578
rect 430 48354 79959 48470
rect 400 48134 79959 48354
rect 400 48018 79570 48134
rect 400 47574 79959 48018
rect 400 47458 79570 47574
rect 400 47126 79959 47458
rect 430 47014 79959 47126
rect 430 47010 79570 47014
rect 400 46898 79570 47010
rect 400 46454 79959 46898
rect 400 46338 79570 46454
rect 400 45894 79959 46338
rect 400 45782 79570 45894
rect 430 45778 79570 45782
rect 430 45666 79959 45778
rect 400 45334 79959 45666
rect 400 45218 79570 45334
rect 400 44774 79959 45218
rect 400 44658 79570 44774
rect 400 44438 79959 44658
rect 430 44322 79959 44438
rect 400 44214 79959 44322
rect 400 44098 79570 44214
rect 400 43654 79959 44098
rect 400 43538 79570 43654
rect 400 43094 79959 43538
rect 430 42978 79570 43094
rect 400 42534 79959 42978
rect 400 42418 79570 42534
rect 400 41974 79959 42418
rect 400 41858 79570 41974
rect 400 41750 79959 41858
rect 430 41634 79959 41750
rect 400 41414 79959 41634
rect 400 41298 79570 41414
rect 400 40854 79959 41298
rect 400 40738 79570 40854
rect 400 40406 79959 40738
rect 430 40294 79959 40406
rect 430 40290 79570 40294
rect 400 40178 79570 40290
rect 400 39734 79959 40178
rect 400 39618 79570 39734
rect 400 39174 79959 39618
rect 400 39062 79570 39174
rect 430 39058 79570 39062
rect 430 38946 79959 39058
rect 400 38614 79959 38946
rect 400 38498 79570 38614
rect 400 38054 79959 38498
rect 400 37938 79570 38054
rect 400 37718 79959 37938
rect 430 37602 79959 37718
rect 400 37494 79959 37602
rect 400 37378 79570 37494
rect 400 36934 79959 37378
rect 400 36818 79570 36934
rect 400 36374 79959 36818
rect 430 36258 79570 36374
rect 400 35814 79959 36258
rect 400 35698 79570 35814
rect 400 35254 79959 35698
rect 400 35138 79570 35254
rect 400 35030 79959 35138
rect 430 34914 79959 35030
rect 400 34694 79959 34914
rect 400 34578 79570 34694
rect 400 34134 79959 34578
rect 400 34018 79570 34134
rect 400 33686 79959 34018
rect 430 33574 79959 33686
rect 430 33570 79570 33574
rect 400 33458 79570 33570
rect 400 33014 79959 33458
rect 400 32898 79570 33014
rect 400 32454 79959 32898
rect 400 32342 79570 32454
rect 430 32338 79570 32342
rect 430 32226 79959 32338
rect 400 31894 79959 32226
rect 400 31778 79570 31894
rect 400 31334 79959 31778
rect 400 31218 79570 31334
rect 400 30998 79959 31218
rect 430 30882 79959 30998
rect 400 30774 79959 30882
rect 400 30658 79570 30774
rect 400 30214 79959 30658
rect 400 30098 79570 30214
rect 400 29654 79959 30098
rect 430 29538 79570 29654
rect 400 29094 79959 29538
rect 400 28978 79570 29094
rect 400 28534 79959 28978
rect 400 28418 79570 28534
rect 400 28310 79959 28418
rect 430 28194 79959 28310
rect 400 27974 79959 28194
rect 400 27858 79570 27974
rect 400 27414 79959 27858
rect 400 27298 79570 27414
rect 400 26966 79959 27298
rect 430 26854 79959 26966
rect 430 26850 79570 26854
rect 400 26738 79570 26850
rect 400 26294 79959 26738
rect 400 26178 79570 26294
rect 400 25734 79959 26178
rect 400 25622 79570 25734
rect 430 25618 79570 25622
rect 430 25506 79959 25618
rect 400 25174 79959 25506
rect 400 25058 79570 25174
rect 400 24614 79959 25058
rect 400 24498 79570 24614
rect 400 24278 79959 24498
rect 430 24162 79959 24278
rect 400 24054 79959 24162
rect 400 23938 79570 24054
rect 400 23494 79959 23938
rect 400 23378 79570 23494
rect 400 22934 79959 23378
rect 430 22818 79570 22934
rect 400 22374 79959 22818
rect 400 22258 79570 22374
rect 400 21814 79959 22258
rect 400 21698 79570 21814
rect 400 21590 79959 21698
rect 430 21474 79959 21590
rect 400 21254 79959 21474
rect 400 21138 79570 21254
rect 400 20694 79959 21138
rect 400 20578 79570 20694
rect 400 20246 79959 20578
rect 430 20134 79959 20246
rect 430 20130 79570 20134
rect 400 20018 79570 20130
rect 400 19574 79959 20018
rect 400 19458 79570 19574
rect 400 19014 79959 19458
rect 400 18902 79570 19014
rect 430 18898 79570 18902
rect 430 18786 79959 18898
rect 400 18454 79959 18786
rect 400 18338 79570 18454
rect 400 17894 79959 18338
rect 400 17778 79570 17894
rect 400 17558 79959 17778
rect 430 17442 79959 17558
rect 400 17334 79959 17442
rect 400 17218 79570 17334
rect 400 16774 79959 17218
rect 400 16658 79570 16774
rect 400 16214 79959 16658
rect 430 16098 79570 16214
rect 400 15654 79959 16098
rect 400 15538 79570 15654
rect 400 15094 79959 15538
rect 400 14978 79570 15094
rect 400 14870 79959 14978
rect 430 14754 79959 14870
rect 400 14534 79959 14754
rect 400 14418 79570 14534
rect 400 13974 79959 14418
rect 400 13858 79570 13974
rect 400 13526 79959 13858
rect 430 13414 79959 13526
rect 430 13410 79570 13414
rect 400 13298 79570 13410
rect 400 12854 79959 13298
rect 400 12738 79570 12854
rect 400 12294 79959 12738
rect 400 12182 79570 12294
rect 430 12178 79570 12182
rect 430 12066 79959 12178
rect 400 11734 79959 12066
rect 400 11618 79570 11734
rect 400 11174 79959 11618
rect 400 11058 79570 11174
rect 400 10838 79959 11058
rect 430 10722 79959 10838
rect 400 10614 79959 10722
rect 400 10498 79570 10614
rect 400 10054 79959 10498
rect 400 9938 79570 10054
rect 400 9494 79959 9938
rect 430 9378 79570 9494
rect 400 8934 79959 9378
rect 400 8818 79570 8934
rect 400 8374 79959 8818
rect 400 8258 79570 8374
rect 400 8150 79959 8258
rect 430 8034 79959 8150
rect 400 7814 79959 8034
rect 400 7698 79570 7814
rect 400 7254 79959 7698
rect 400 7138 79570 7254
rect 400 6806 79959 7138
rect 430 6694 79959 6806
rect 430 6690 79570 6694
rect 400 6578 79570 6690
rect 400 6134 79959 6578
rect 400 6018 79570 6134
rect 400 5574 79959 6018
rect 400 5462 79570 5574
rect 430 5458 79570 5462
rect 430 5346 79959 5458
rect 400 5014 79959 5346
rect 400 4898 79570 5014
rect 400 4454 79959 4898
rect 400 4338 79570 4454
rect 400 4118 79959 4338
rect 430 4002 79959 4118
rect 400 3894 79959 4002
rect 400 3778 79570 3894
rect 400 3334 79959 3778
rect 400 3218 79570 3334
rect 400 2774 79959 3218
rect 430 2658 79959 2774
rect 400 1430 79959 2658
rect 430 1358 79959 1430
<< metal4 >>
rect 2224 1538 2384 138406
rect 9904 1538 10064 138406
rect 17584 1538 17744 138406
rect 25264 1538 25424 138406
rect 32944 1538 33104 138406
rect 40624 1538 40784 138406
rect 48304 1538 48464 138406
rect 55984 1538 56144 138406
rect 63664 1538 63824 138406
rect 71344 1538 71504 138406
rect 79024 1538 79184 138406
<< obsm4 >>
rect 3038 5217 9874 137919
rect 10094 5217 17554 137919
rect 17774 5217 25234 137919
rect 25454 5217 32914 137919
rect 33134 5217 40594 137919
rect 40814 5217 48274 137919
rect 48494 5217 55954 137919
rect 56174 5217 63634 137919
rect 63854 5217 71314 137919
rect 71534 5217 78994 137919
rect 79214 5217 79506 137919
<< labels >>
rlabel metal3 s 79600 3248 80000 3304 6 clk
port 1 nsew signal input
rlabel metal2 s 3584 139600 3640 140000 6 irq_in[0]
port 2 nsew signal input
rlabel metal2 s 10192 139600 10248 140000 6 irq_in[1]
port 3 nsew signal input
rlabel metal2 s 16800 139600 16856 140000 6 irq_in[2]
port 4 nsew signal input
rlabel metal2 s 23408 139600 23464 140000 6 irq_in[3]
port 5 nsew signal input
rlabel metal2 s 30016 139600 30072 140000 6 irq_oeb[0]
port 6 nsew signal output
rlabel metal2 s 36624 139600 36680 140000 6 irq_oeb[1]
port 7 nsew signal output
rlabel metal2 s 43232 139600 43288 140000 6 irq_oeb[2]
port 8 nsew signal output
rlabel metal2 s 49840 139600 49896 140000 6 irq_oeb[3]
port 9 nsew signal output
rlabel metal2 s 56448 139600 56504 140000 6 irq_out[0]
port 10 nsew signal output
rlabel metal2 s 63056 139600 63112 140000 6 irq_out[1]
port 11 nsew signal output
rlabel metal2 s 69664 139600 69720 140000 6 irq_out[2]
port 12 nsew signal output
rlabel metal2 s 76272 139600 76328 140000 6 irq_out[3]
port 13 nsew signal output
rlabel metal3 s 0 5376 400 5432 6 mem_addr[0]
port 14 nsew signal output
rlabel metal3 s 0 18816 400 18872 6 mem_addr[10]
port 15 nsew signal output
rlabel metal3 s 0 20160 400 20216 6 mem_addr[11]
port 16 nsew signal output
rlabel metal3 s 0 21504 400 21560 6 mem_addr[12]
port 17 nsew signal output
rlabel metal3 s 0 22848 400 22904 6 mem_addr[13]
port 18 nsew signal output
rlabel metal3 s 0 24192 400 24248 6 mem_addr[14]
port 19 nsew signal output
rlabel metal3 s 0 25536 400 25592 6 mem_addr[15]
port 20 nsew signal output
rlabel metal3 s 0 26880 400 26936 6 mem_addr[16]
port 21 nsew signal output
rlabel metal3 s 0 28224 400 28280 6 mem_addr[17]
port 22 nsew signal output
rlabel metal3 s 0 29568 400 29624 6 mem_addr[18]
port 23 nsew signal output
rlabel metal3 s 0 30912 400 30968 6 mem_addr[19]
port 24 nsew signal output
rlabel metal3 s 0 6720 400 6776 6 mem_addr[1]
port 25 nsew signal output
rlabel metal3 s 0 32256 400 32312 6 mem_addr[20]
port 26 nsew signal output
rlabel metal3 s 0 33600 400 33656 6 mem_addr[21]
port 27 nsew signal output
rlabel metal3 s 0 34944 400 35000 6 mem_addr[22]
port 28 nsew signal output
rlabel metal3 s 0 36288 400 36344 6 mem_addr[23]
port 29 nsew signal output
rlabel metal3 s 0 37632 400 37688 6 mem_addr[24]
port 30 nsew signal output
rlabel metal3 s 0 38976 400 39032 6 mem_addr[25]
port 31 nsew signal output
rlabel metal3 s 0 40320 400 40376 6 mem_addr[26]
port 32 nsew signal output
rlabel metal3 s 0 41664 400 41720 6 mem_addr[27]
port 33 nsew signal output
rlabel metal3 s 0 43008 400 43064 6 mem_addr[28]
port 34 nsew signal output
rlabel metal3 s 0 44352 400 44408 6 mem_addr[29]
port 35 nsew signal output
rlabel metal3 s 0 8064 400 8120 6 mem_addr[2]
port 36 nsew signal output
rlabel metal3 s 0 45696 400 45752 6 mem_addr[30]
port 37 nsew signal output
rlabel metal3 s 0 47040 400 47096 6 mem_addr[31]
port 38 nsew signal output
rlabel metal3 s 0 9408 400 9464 6 mem_addr[3]
port 39 nsew signal output
rlabel metal3 s 0 10752 400 10808 6 mem_addr[4]
port 40 nsew signal output
rlabel metal3 s 0 12096 400 12152 6 mem_addr[5]
port 41 nsew signal output
rlabel metal3 s 0 13440 400 13496 6 mem_addr[6]
port 42 nsew signal output
rlabel metal3 s 0 14784 400 14840 6 mem_addr[7]
port 43 nsew signal output
rlabel metal3 s 0 16128 400 16184 6 mem_addr[8]
port 44 nsew signal output
rlabel metal3 s 0 17472 400 17528 6 mem_addr[9]
port 45 nsew signal output
rlabel metal3 s 0 2688 400 2744 6 mem_instr
port 46 nsew signal output
rlabel metal3 s 0 96768 400 96824 6 mem_rdata[0]
port 47 nsew signal input
rlabel metal3 s 0 110208 400 110264 6 mem_rdata[10]
port 48 nsew signal input
rlabel metal3 s 0 111552 400 111608 6 mem_rdata[11]
port 49 nsew signal input
rlabel metal3 s 0 112896 400 112952 6 mem_rdata[12]
port 50 nsew signal input
rlabel metal3 s 0 114240 400 114296 6 mem_rdata[13]
port 51 nsew signal input
rlabel metal3 s 0 115584 400 115640 6 mem_rdata[14]
port 52 nsew signal input
rlabel metal3 s 0 116928 400 116984 6 mem_rdata[15]
port 53 nsew signal input
rlabel metal3 s 0 118272 400 118328 6 mem_rdata[16]
port 54 nsew signal input
rlabel metal3 s 0 119616 400 119672 6 mem_rdata[17]
port 55 nsew signal input
rlabel metal3 s 0 120960 400 121016 6 mem_rdata[18]
port 56 nsew signal input
rlabel metal3 s 0 122304 400 122360 6 mem_rdata[19]
port 57 nsew signal input
rlabel metal3 s 0 98112 400 98168 6 mem_rdata[1]
port 58 nsew signal input
rlabel metal3 s 0 123648 400 123704 6 mem_rdata[20]
port 59 nsew signal input
rlabel metal3 s 0 124992 400 125048 6 mem_rdata[21]
port 60 nsew signal input
rlabel metal3 s 0 126336 400 126392 6 mem_rdata[22]
port 61 nsew signal input
rlabel metal3 s 0 127680 400 127736 6 mem_rdata[23]
port 62 nsew signal input
rlabel metal3 s 0 129024 400 129080 6 mem_rdata[24]
port 63 nsew signal input
rlabel metal3 s 0 130368 400 130424 6 mem_rdata[25]
port 64 nsew signal input
rlabel metal3 s 0 131712 400 131768 6 mem_rdata[26]
port 65 nsew signal input
rlabel metal3 s 0 133056 400 133112 6 mem_rdata[27]
port 66 nsew signal input
rlabel metal3 s 0 134400 400 134456 6 mem_rdata[28]
port 67 nsew signal input
rlabel metal3 s 0 135744 400 135800 6 mem_rdata[29]
port 68 nsew signal input
rlabel metal3 s 0 99456 400 99512 6 mem_rdata[2]
port 69 nsew signal input
rlabel metal3 s 0 137088 400 137144 6 mem_rdata[30]
port 70 nsew signal input
rlabel metal3 s 0 138432 400 138488 6 mem_rdata[31]
port 71 nsew signal input
rlabel metal3 s 0 100800 400 100856 6 mem_rdata[3]
port 72 nsew signal input
rlabel metal3 s 0 102144 400 102200 6 mem_rdata[4]
port 73 nsew signal input
rlabel metal3 s 0 103488 400 103544 6 mem_rdata[5]
port 74 nsew signal input
rlabel metal3 s 0 104832 400 104888 6 mem_rdata[6]
port 75 nsew signal input
rlabel metal3 s 0 106176 400 106232 6 mem_rdata[7]
port 76 nsew signal input
rlabel metal3 s 0 107520 400 107576 6 mem_rdata[8]
port 77 nsew signal input
rlabel metal3 s 0 108864 400 108920 6 mem_rdata[9]
port 78 nsew signal input
rlabel metal3 s 0 4032 400 4088 6 mem_ready
port 79 nsew signal input
rlabel metal3 s 0 1344 400 1400 6 mem_valid
port 80 nsew signal output
rlabel metal3 s 0 48384 400 48440 6 mem_wdata[0]
port 81 nsew signal output
rlabel metal3 s 0 61824 400 61880 6 mem_wdata[10]
port 82 nsew signal output
rlabel metal3 s 0 63168 400 63224 6 mem_wdata[11]
port 83 nsew signal output
rlabel metal3 s 0 64512 400 64568 6 mem_wdata[12]
port 84 nsew signal output
rlabel metal3 s 0 65856 400 65912 6 mem_wdata[13]
port 85 nsew signal output
rlabel metal3 s 0 67200 400 67256 6 mem_wdata[14]
port 86 nsew signal output
rlabel metal3 s 0 68544 400 68600 6 mem_wdata[15]
port 87 nsew signal output
rlabel metal3 s 0 69888 400 69944 6 mem_wdata[16]
port 88 nsew signal output
rlabel metal3 s 0 71232 400 71288 6 mem_wdata[17]
port 89 nsew signal output
rlabel metal3 s 0 72576 400 72632 6 mem_wdata[18]
port 90 nsew signal output
rlabel metal3 s 0 73920 400 73976 6 mem_wdata[19]
port 91 nsew signal output
rlabel metal3 s 0 49728 400 49784 6 mem_wdata[1]
port 92 nsew signal output
rlabel metal3 s 0 75264 400 75320 6 mem_wdata[20]
port 93 nsew signal output
rlabel metal3 s 0 76608 400 76664 6 mem_wdata[21]
port 94 nsew signal output
rlabel metal3 s 0 77952 400 78008 6 mem_wdata[22]
port 95 nsew signal output
rlabel metal3 s 0 79296 400 79352 6 mem_wdata[23]
port 96 nsew signal output
rlabel metal3 s 0 80640 400 80696 6 mem_wdata[24]
port 97 nsew signal output
rlabel metal3 s 0 81984 400 82040 6 mem_wdata[25]
port 98 nsew signal output
rlabel metal3 s 0 83328 400 83384 6 mem_wdata[26]
port 99 nsew signal output
rlabel metal3 s 0 84672 400 84728 6 mem_wdata[27]
port 100 nsew signal output
rlabel metal3 s 0 86016 400 86072 6 mem_wdata[28]
port 101 nsew signal output
rlabel metal3 s 0 87360 400 87416 6 mem_wdata[29]
port 102 nsew signal output
rlabel metal3 s 0 51072 400 51128 6 mem_wdata[2]
port 103 nsew signal output
rlabel metal3 s 0 88704 400 88760 6 mem_wdata[30]
port 104 nsew signal output
rlabel metal3 s 0 90048 400 90104 6 mem_wdata[31]
port 105 nsew signal output
rlabel metal3 s 0 52416 400 52472 6 mem_wdata[3]
port 106 nsew signal output
rlabel metal3 s 0 53760 400 53816 6 mem_wdata[4]
port 107 nsew signal output
rlabel metal3 s 0 55104 400 55160 6 mem_wdata[5]
port 108 nsew signal output
rlabel metal3 s 0 56448 400 56504 6 mem_wdata[6]
port 109 nsew signal output
rlabel metal3 s 0 57792 400 57848 6 mem_wdata[7]
port 110 nsew signal output
rlabel metal3 s 0 59136 400 59192 6 mem_wdata[8]
port 111 nsew signal output
rlabel metal3 s 0 60480 400 60536 6 mem_wdata[9]
port 112 nsew signal output
rlabel metal3 s 0 91392 400 91448 6 mem_wstrb[0]
port 113 nsew signal output
rlabel metal3 s 0 92736 400 92792 6 mem_wstrb[1]
port 114 nsew signal output
rlabel metal3 s 0 94080 400 94136 6 mem_wstrb[2]
port 115 nsew signal output
rlabel metal3 s 0 95424 400 95480 6 mem_wstrb[3]
port 116 nsew signal output
rlabel metal3 s 79600 117488 80000 117544 6 pcpi_approx_mul_rd[0]
port 117 nsew signal input
rlabel metal3 s 79600 123088 80000 123144 6 pcpi_approx_mul_rd[10]
port 118 nsew signal input
rlabel metal3 s 79600 123648 80000 123704 6 pcpi_approx_mul_rd[11]
port 119 nsew signal input
rlabel metal3 s 79600 124208 80000 124264 6 pcpi_approx_mul_rd[12]
port 120 nsew signal input
rlabel metal3 s 79600 124768 80000 124824 6 pcpi_approx_mul_rd[13]
port 121 nsew signal input
rlabel metal3 s 79600 125328 80000 125384 6 pcpi_approx_mul_rd[14]
port 122 nsew signal input
rlabel metal3 s 79600 125888 80000 125944 6 pcpi_approx_mul_rd[15]
port 123 nsew signal input
rlabel metal3 s 79600 126448 80000 126504 6 pcpi_approx_mul_rd[16]
port 124 nsew signal input
rlabel metal3 s 79600 127008 80000 127064 6 pcpi_approx_mul_rd[17]
port 125 nsew signal input
rlabel metal3 s 79600 127568 80000 127624 6 pcpi_approx_mul_rd[18]
port 126 nsew signal input
rlabel metal3 s 79600 128128 80000 128184 6 pcpi_approx_mul_rd[19]
port 127 nsew signal input
rlabel metal3 s 79600 118048 80000 118104 6 pcpi_approx_mul_rd[1]
port 128 nsew signal input
rlabel metal3 s 79600 128688 80000 128744 6 pcpi_approx_mul_rd[20]
port 129 nsew signal input
rlabel metal3 s 79600 129248 80000 129304 6 pcpi_approx_mul_rd[21]
port 130 nsew signal input
rlabel metal3 s 79600 129808 80000 129864 6 pcpi_approx_mul_rd[22]
port 131 nsew signal input
rlabel metal3 s 79600 130368 80000 130424 6 pcpi_approx_mul_rd[23]
port 132 nsew signal input
rlabel metal3 s 79600 130928 80000 130984 6 pcpi_approx_mul_rd[24]
port 133 nsew signal input
rlabel metal3 s 79600 131488 80000 131544 6 pcpi_approx_mul_rd[25]
port 134 nsew signal input
rlabel metal3 s 79600 132048 80000 132104 6 pcpi_approx_mul_rd[26]
port 135 nsew signal input
rlabel metal3 s 79600 132608 80000 132664 6 pcpi_approx_mul_rd[27]
port 136 nsew signal input
rlabel metal3 s 79600 133168 80000 133224 6 pcpi_approx_mul_rd[28]
port 137 nsew signal input
rlabel metal3 s 79600 133728 80000 133784 6 pcpi_approx_mul_rd[29]
port 138 nsew signal input
rlabel metal3 s 79600 118608 80000 118664 6 pcpi_approx_mul_rd[2]
port 139 nsew signal input
rlabel metal3 s 79600 134288 80000 134344 6 pcpi_approx_mul_rd[30]
port 140 nsew signal input
rlabel metal3 s 79600 134848 80000 134904 6 pcpi_approx_mul_rd[31]
port 141 nsew signal input
rlabel metal3 s 79600 119168 80000 119224 6 pcpi_approx_mul_rd[3]
port 142 nsew signal input
rlabel metal3 s 79600 119728 80000 119784 6 pcpi_approx_mul_rd[4]
port 143 nsew signal input
rlabel metal3 s 79600 120288 80000 120344 6 pcpi_approx_mul_rd[5]
port 144 nsew signal input
rlabel metal3 s 79600 120848 80000 120904 6 pcpi_approx_mul_rd[6]
port 145 nsew signal input
rlabel metal3 s 79600 121408 80000 121464 6 pcpi_approx_mul_rd[7]
port 146 nsew signal input
rlabel metal3 s 79600 121968 80000 122024 6 pcpi_approx_mul_rd[8]
port 147 nsew signal input
rlabel metal3 s 79600 122528 80000 122584 6 pcpi_approx_mul_rd[9]
port 148 nsew signal input
rlabel metal3 s 79600 135408 80000 135464 6 pcpi_approx_mul_ready
port 149 nsew signal input
rlabel metal3 s 79600 135968 80000 136024 6 pcpi_approx_mul_wait
port 150 nsew signal input
rlabel metal3 s 79600 136528 80000 136584 6 pcpi_approx_mul_wr
port 151 nsew signal input
rlabel metal3 s 79600 78848 80000 78904 6 pcpi_div_rd[0]
port 152 nsew signal input
rlabel metal3 s 79600 84448 80000 84504 6 pcpi_div_rd[10]
port 153 nsew signal input
rlabel metal3 s 79600 85008 80000 85064 6 pcpi_div_rd[11]
port 154 nsew signal input
rlabel metal3 s 79600 85568 80000 85624 6 pcpi_div_rd[12]
port 155 nsew signal input
rlabel metal3 s 79600 86128 80000 86184 6 pcpi_div_rd[13]
port 156 nsew signal input
rlabel metal3 s 79600 86688 80000 86744 6 pcpi_div_rd[14]
port 157 nsew signal input
rlabel metal3 s 79600 87248 80000 87304 6 pcpi_div_rd[15]
port 158 nsew signal input
rlabel metal3 s 79600 87808 80000 87864 6 pcpi_div_rd[16]
port 159 nsew signal input
rlabel metal3 s 79600 88368 80000 88424 6 pcpi_div_rd[17]
port 160 nsew signal input
rlabel metal3 s 79600 88928 80000 88984 6 pcpi_div_rd[18]
port 161 nsew signal input
rlabel metal3 s 79600 89488 80000 89544 6 pcpi_div_rd[19]
port 162 nsew signal input
rlabel metal3 s 79600 79408 80000 79464 6 pcpi_div_rd[1]
port 163 nsew signal input
rlabel metal3 s 79600 90048 80000 90104 6 pcpi_div_rd[20]
port 164 nsew signal input
rlabel metal3 s 79600 90608 80000 90664 6 pcpi_div_rd[21]
port 165 nsew signal input
rlabel metal3 s 79600 91168 80000 91224 6 pcpi_div_rd[22]
port 166 nsew signal input
rlabel metal3 s 79600 91728 80000 91784 6 pcpi_div_rd[23]
port 167 nsew signal input
rlabel metal3 s 79600 92288 80000 92344 6 pcpi_div_rd[24]
port 168 nsew signal input
rlabel metal3 s 79600 92848 80000 92904 6 pcpi_div_rd[25]
port 169 nsew signal input
rlabel metal3 s 79600 93408 80000 93464 6 pcpi_div_rd[26]
port 170 nsew signal input
rlabel metal3 s 79600 93968 80000 94024 6 pcpi_div_rd[27]
port 171 nsew signal input
rlabel metal3 s 79600 94528 80000 94584 6 pcpi_div_rd[28]
port 172 nsew signal input
rlabel metal3 s 79600 95088 80000 95144 6 pcpi_div_rd[29]
port 173 nsew signal input
rlabel metal3 s 79600 79968 80000 80024 6 pcpi_div_rd[2]
port 174 nsew signal input
rlabel metal3 s 79600 95648 80000 95704 6 pcpi_div_rd[30]
port 175 nsew signal input
rlabel metal3 s 79600 96208 80000 96264 6 pcpi_div_rd[31]
port 176 nsew signal input
rlabel metal3 s 79600 80528 80000 80584 6 pcpi_div_rd[3]
port 177 nsew signal input
rlabel metal3 s 79600 81088 80000 81144 6 pcpi_div_rd[4]
port 178 nsew signal input
rlabel metal3 s 79600 81648 80000 81704 6 pcpi_div_rd[5]
port 179 nsew signal input
rlabel metal3 s 79600 82208 80000 82264 6 pcpi_div_rd[6]
port 180 nsew signal input
rlabel metal3 s 79600 82768 80000 82824 6 pcpi_div_rd[7]
port 181 nsew signal input
rlabel metal3 s 79600 83328 80000 83384 6 pcpi_div_rd[8]
port 182 nsew signal input
rlabel metal3 s 79600 83888 80000 83944 6 pcpi_div_rd[9]
port 183 nsew signal input
rlabel metal3 s 79600 97328 80000 97384 6 pcpi_div_ready
port 184 nsew signal input
rlabel metal3 s 79600 96768 80000 96824 6 pcpi_div_wait
port 185 nsew signal input
rlabel metal3 s 79600 78288 80000 78344 6 pcpi_div_wr
port 186 nsew signal input
rlabel metal3 s 79600 97888 80000 97944 6 pcpi_exact_mul_rd[0]
port 187 nsew signal input
rlabel metal3 s 79600 103488 80000 103544 6 pcpi_exact_mul_rd[10]
port 188 nsew signal input
rlabel metal3 s 79600 104048 80000 104104 6 pcpi_exact_mul_rd[11]
port 189 nsew signal input
rlabel metal3 s 79600 104608 80000 104664 6 pcpi_exact_mul_rd[12]
port 190 nsew signal input
rlabel metal3 s 79600 105168 80000 105224 6 pcpi_exact_mul_rd[13]
port 191 nsew signal input
rlabel metal3 s 79600 105728 80000 105784 6 pcpi_exact_mul_rd[14]
port 192 nsew signal input
rlabel metal3 s 79600 106288 80000 106344 6 pcpi_exact_mul_rd[15]
port 193 nsew signal input
rlabel metal3 s 79600 106848 80000 106904 6 pcpi_exact_mul_rd[16]
port 194 nsew signal input
rlabel metal3 s 79600 107408 80000 107464 6 pcpi_exact_mul_rd[17]
port 195 nsew signal input
rlabel metal3 s 79600 107968 80000 108024 6 pcpi_exact_mul_rd[18]
port 196 nsew signal input
rlabel metal3 s 79600 108528 80000 108584 6 pcpi_exact_mul_rd[19]
port 197 nsew signal input
rlabel metal3 s 79600 98448 80000 98504 6 pcpi_exact_mul_rd[1]
port 198 nsew signal input
rlabel metal3 s 79600 109088 80000 109144 6 pcpi_exact_mul_rd[20]
port 199 nsew signal input
rlabel metal3 s 79600 109648 80000 109704 6 pcpi_exact_mul_rd[21]
port 200 nsew signal input
rlabel metal3 s 79600 110208 80000 110264 6 pcpi_exact_mul_rd[22]
port 201 nsew signal input
rlabel metal3 s 79600 110768 80000 110824 6 pcpi_exact_mul_rd[23]
port 202 nsew signal input
rlabel metal3 s 79600 111328 80000 111384 6 pcpi_exact_mul_rd[24]
port 203 nsew signal input
rlabel metal3 s 79600 111888 80000 111944 6 pcpi_exact_mul_rd[25]
port 204 nsew signal input
rlabel metal3 s 79600 112448 80000 112504 6 pcpi_exact_mul_rd[26]
port 205 nsew signal input
rlabel metal3 s 79600 113008 80000 113064 6 pcpi_exact_mul_rd[27]
port 206 nsew signal input
rlabel metal3 s 79600 113568 80000 113624 6 pcpi_exact_mul_rd[28]
port 207 nsew signal input
rlabel metal3 s 79600 114128 80000 114184 6 pcpi_exact_mul_rd[29]
port 208 nsew signal input
rlabel metal3 s 79600 99008 80000 99064 6 pcpi_exact_mul_rd[2]
port 209 nsew signal input
rlabel metal3 s 79600 114688 80000 114744 6 pcpi_exact_mul_rd[30]
port 210 nsew signal input
rlabel metal3 s 79600 115248 80000 115304 6 pcpi_exact_mul_rd[31]
port 211 nsew signal input
rlabel metal3 s 79600 99568 80000 99624 6 pcpi_exact_mul_rd[3]
port 212 nsew signal input
rlabel metal3 s 79600 100128 80000 100184 6 pcpi_exact_mul_rd[4]
port 213 nsew signal input
rlabel metal3 s 79600 100688 80000 100744 6 pcpi_exact_mul_rd[5]
port 214 nsew signal input
rlabel metal3 s 79600 101248 80000 101304 6 pcpi_exact_mul_rd[6]
port 215 nsew signal input
rlabel metal3 s 79600 101808 80000 101864 6 pcpi_exact_mul_rd[7]
port 216 nsew signal input
rlabel metal3 s 79600 102368 80000 102424 6 pcpi_exact_mul_rd[8]
port 217 nsew signal input
rlabel metal3 s 79600 102928 80000 102984 6 pcpi_exact_mul_rd[9]
port 218 nsew signal input
rlabel metal3 s 79600 115808 80000 115864 6 pcpi_exact_mul_ready
port 219 nsew signal input
rlabel metal3 s 79600 116368 80000 116424 6 pcpi_exact_mul_wait
port 220 nsew signal input
rlabel metal3 s 79600 116928 80000 116984 6 pcpi_exact_mul_wr
port 221 nsew signal input
rlabel metal3 s 79600 4928 80000 4984 6 pcpi_insn[0]
port 222 nsew signal output
rlabel metal3 s 79600 10528 80000 10584 6 pcpi_insn[10]
port 223 nsew signal output
rlabel metal3 s 79600 11088 80000 11144 6 pcpi_insn[11]
port 224 nsew signal output
rlabel metal3 s 79600 11648 80000 11704 6 pcpi_insn[12]
port 225 nsew signal output
rlabel metal3 s 79600 12208 80000 12264 6 pcpi_insn[13]
port 226 nsew signal output
rlabel metal3 s 79600 12768 80000 12824 6 pcpi_insn[14]
port 227 nsew signal output
rlabel metal3 s 79600 13328 80000 13384 6 pcpi_insn[15]
port 228 nsew signal output
rlabel metal3 s 79600 13888 80000 13944 6 pcpi_insn[16]
port 229 nsew signal output
rlabel metal3 s 79600 14448 80000 14504 6 pcpi_insn[17]
port 230 nsew signal output
rlabel metal3 s 79600 15008 80000 15064 6 pcpi_insn[18]
port 231 nsew signal output
rlabel metal3 s 79600 15568 80000 15624 6 pcpi_insn[19]
port 232 nsew signal output
rlabel metal3 s 79600 5488 80000 5544 6 pcpi_insn[1]
port 233 nsew signal output
rlabel metal3 s 79600 16128 80000 16184 6 pcpi_insn[20]
port 234 nsew signal output
rlabel metal3 s 79600 16688 80000 16744 6 pcpi_insn[21]
port 235 nsew signal output
rlabel metal3 s 79600 17248 80000 17304 6 pcpi_insn[22]
port 236 nsew signal output
rlabel metal3 s 79600 17808 80000 17864 6 pcpi_insn[23]
port 237 nsew signal output
rlabel metal3 s 79600 18368 80000 18424 6 pcpi_insn[24]
port 238 nsew signal output
rlabel metal3 s 79600 18928 80000 18984 6 pcpi_insn[25]
port 239 nsew signal output
rlabel metal3 s 79600 19488 80000 19544 6 pcpi_insn[26]
port 240 nsew signal output
rlabel metal3 s 79600 20048 80000 20104 6 pcpi_insn[27]
port 241 nsew signal output
rlabel metal3 s 79600 20608 80000 20664 6 pcpi_insn[28]
port 242 nsew signal output
rlabel metal3 s 79600 21168 80000 21224 6 pcpi_insn[29]
port 243 nsew signal output
rlabel metal3 s 79600 6048 80000 6104 6 pcpi_insn[2]
port 244 nsew signal output
rlabel metal3 s 79600 21728 80000 21784 6 pcpi_insn[30]
port 245 nsew signal output
rlabel metal3 s 79600 22288 80000 22344 6 pcpi_insn[31]
port 246 nsew signal output
rlabel metal3 s 79600 6608 80000 6664 6 pcpi_insn[3]
port 247 nsew signal output
rlabel metal3 s 79600 7168 80000 7224 6 pcpi_insn[4]
port 248 nsew signal output
rlabel metal3 s 79600 7728 80000 7784 6 pcpi_insn[5]
port 249 nsew signal output
rlabel metal3 s 79600 8288 80000 8344 6 pcpi_insn[6]
port 250 nsew signal output
rlabel metal3 s 79600 8848 80000 8904 6 pcpi_insn[7]
port 251 nsew signal output
rlabel metal3 s 79600 9408 80000 9464 6 pcpi_insn[8]
port 252 nsew signal output
rlabel metal3 s 79600 9968 80000 10024 6 pcpi_insn[9]
port 253 nsew signal output
rlabel metal3 s 79600 59248 80000 59304 6 pcpi_mul_rd[0]
port 254 nsew signal input
rlabel metal3 s 79600 64848 80000 64904 6 pcpi_mul_rd[10]
port 255 nsew signal input
rlabel metal3 s 79600 65408 80000 65464 6 pcpi_mul_rd[11]
port 256 nsew signal input
rlabel metal3 s 79600 65968 80000 66024 6 pcpi_mul_rd[12]
port 257 nsew signal input
rlabel metal3 s 79600 66528 80000 66584 6 pcpi_mul_rd[13]
port 258 nsew signal input
rlabel metal3 s 79600 67088 80000 67144 6 pcpi_mul_rd[14]
port 259 nsew signal input
rlabel metal3 s 79600 67648 80000 67704 6 pcpi_mul_rd[15]
port 260 nsew signal input
rlabel metal3 s 79600 68208 80000 68264 6 pcpi_mul_rd[16]
port 261 nsew signal input
rlabel metal3 s 79600 68768 80000 68824 6 pcpi_mul_rd[17]
port 262 nsew signal input
rlabel metal3 s 79600 69328 80000 69384 6 pcpi_mul_rd[18]
port 263 nsew signal input
rlabel metal3 s 79600 69888 80000 69944 6 pcpi_mul_rd[19]
port 264 nsew signal input
rlabel metal3 s 79600 59808 80000 59864 6 pcpi_mul_rd[1]
port 265 nsew signal input
rlabel metal3 s 79600 70448 80000 70504 6 pcpi_mul_rd[20]
port 266 nsew signal input
rlabel metal3 s 79600 71008 80000 71064 6 pcpi_mul_rd[21]
port 267 nsew signal input
rlabel metal3 s 79600 71568 80000 71624 6 pcpi_mul_rd[22]
port 268 nsew signal input
rlabel metal3 s 79600 72128 80000 72184 6 pcpi_mul_rd[23]
port 269 nsew signal input
rlabel metal3 s 79600 72688 80000 72744 6 pcpi_mul_rd[24]
port 270 nsew signal input
rlabel metal3 s 79600 73248 80000 73304 6 pcpi_mul_rd[25]
port 271 nsew signal input
rlabel metal3 s 79600 73808 80000 73864 6 pcpi_mul_rd[26]
port 272 nsew signal input
rlabel metal3 s 79600 74368 80000 74424 6 pcpi_mul_rd[27]
port 273 nsew signal input
rlabel metal3 s 79600 74928 80000 74984 6 pcpi_mul_rd[28]
port 274 nsew signal input
rlabel metal3 s 79600 75488 80000 75544 6 pcpi_mul_rd[29]
port 275 nsew signal input
rlabel metal3 s 79600 60368 80000 60424 6 pcpi_mul_rd[2]
port 276 nsew signal input
rlabel metal3 s 79600 76048 80000 76104 6 pcpi_mul_rd[30]
port 277 nsew signal input
rlabel metal3 s 79600 76608 80000 76664 6 pcpi_mul_rd[31]
port 278 nsew signal input
rlabel metal3 s 79600 60928 80000 60984 6 pcpi_mul_rd[3]
port 279 nsew signal input
rlabel metal3 s 79600 61488 80000 61544 6 pcpi_mul_rd[4]
port 280 nsew signal input
rlabel metal3 s 79600 62048 80000 62104 6 pcpi_mul_rd[5]
port 281 nsew signal input
rlabel metal3 s 79600 62608 80000 62664 6 pcpi_mul_rd[6]
port 282 nsew signal input
rlabel metal3 s 79600 63168 80000 63224 6 pcpi_mul_rd[7]
port 283 nsew signal input
rlabel metal3 s 79600 63728 80000 63784 6 pcpi_mul_rd[8]
port 284 nsew signal input
rlabel metal3 s 79600 64288 80000 64344 6 pcpi_mul_rd[9]
port 285 nsew signal input
rlabel metal3 s 79600 77728 80000 77784 6 pcpi_mul_ready
port 286 nsew signal input
rlabel metal3 s 79600 77168 80000 77224 6 pcpi_mul_wait
port 287 nsew signal input
rlabel metal3 s 79600 58688 80000 58744 6 pcpi_mul_wr
port 288 nsew signal input
rlabel metal3 s 79600 22848 80000 22904 6 pcpi_rs1[0]
port 289 nsew signal output
rlabel metal3 s 79600 28448 80000 28504 6 pcpi_rs1[10]
port 290 nsew signal output
rlabel metal3 s 79600 29008 80000 29064 6 pcpi_rs1[11]
port 291 nsew signal output
rlabel metal3 s 79600 29568 80000 29624 6 pcpi_rs1[12]
port 292 nsew signal output
rlabel metal3 s 79600 30128 80000 30184 6 pcpi_rs1[13]
port 293 nsew signal output
rlabel metal3 s 79600 30688 80000 30744 6 pcpi_rs1[14]
port 294 nsew signal output
rlabel metal3 s 79600 31248 80000 31304 6 pcpi_rs1[15]
port 295 nsew signal output
rlabel metal3 s 79600 31808 80000 31864 6 pcpi_rs1[16]
port 296 nsew signal output
rlabel metal3 s 79600 32368 80000 32424 6 pcpi_rs1[17]
port 297 nsew signal output
rlabel metal3 s 79600 32928 80000 32984 6 pcpi_rs1[18]
port 298 nsew signal output
rlabel metal3 s 79600 33488 80000 33544 6 pcpi_rs1[19]
port 299 nsew signal output
rlabel metal3 s 79600 23408 80000 23464 6 pcpi_rs1[1]
port 300 nsew signal output
rlabel metal3 s 79600 34048 80000 34104 6 pcpi_rs1[20]
port 301 nsew signal output
rlabel metal3 s 79600 34608 80000 34664 6 pcpi_rs1[21]
port 302 nsew signal output
rlabel metal3 s 79600 35168 80000 35224 6 pcpi_rs1[22]
port 303 nsew signal output
rlabel metal3 s 79600 35728 80000 35784 6 pcpi_rs1[23]
port 304 nsew signal output
rlabel metal3 s 79600 36288 80000 36344 6 pcpi_rs1[24]
port 305 nsew signal output
rlabel metal3 s 79600 36848 80000 36904 6 pcpi_rs1[25]
port 306 nsew signal output
rlabel metal3 s 79600 37408 80000 37464 6 pcpi_rs1[26]
port 307 nsew signal output
rlabel metal3 s 79600 37968 80000 38024 6 pcpi_rs1[27]
port 308 nsew signal output
rlabel metal3 s 79600 38528 80000 38584 6 pcpi_rs1[28]
port 309 nsew signal output
rlabel metal3 s 79600 39088 80000 39144 6 pcpi_rs1[29]
port 310 nsew signal output
rlabel metal3 s 79600 23968 80000 24024 6 pcpi_rs1[2]
port 311 nsew signal output
rlabel metal3 s 79600 39648 80000 39704 6 pcpi_rs1[30]
port 312 nsew signal output
rlabel metal3 s 79600 40208 80000 40264 6 pcpi_rs1[31]
port 313 nsew signal output
rlabel metal3 s 79600 24528 80000 24584 6 pcpi_rs1[3]
port 314 nsew signal output
rlabel metal3 s 79600 25088 80000 25144 6 pcpi_rs1[4]
port 315 nsew signal output
rlabel metal3 s 79600 25648 80000 25704 6 pcpi_rs1[5]
port 316 nsew signal output
rlabel metal3 s 79600 26208 80000 26264 6 pcpi_rs1[6]
port 317 nsew signal output
rlabel metal3 s 79600 26768 80000 26824 6 pcpi_rs1[7]
port 318 nsew signal output
rlabel metal3 s 79600 27328 80000 27384 6 pcpi_rs1[8]
port 319 nsew signal output
rlabel metal3 s 79600 27888 80000 27944 6 pcpi_rs1[9]
port 320 nsew signal output
rlabel metal3 s 79600 40768 80000 40824 6 pcpi_rs2[0]
port 321 nsew signal output
rlabel metal3 s 79600 46368 80000 46424 6 pcpi_rs2[10]
port 322 nsew signal output
rlabel metal3 s 79600 46928 80000 46984 6 pcpi_rs2[11]
port 323 nsew signal output
rlabel metal3 s 79600 47488 80000 47544 6 pcpi_rs2[12]
port 324 nsew signal output
rlabel metal3 s 79600 48048 80000 48104 6 pcpi_rs2[13]
port 325 nsew signal output
rlabel metal3 s 79600 48608 80000 48664 6 pcpi_rs2[14]
port 326 nsew signal output
rlabel metal3 s 79600 49168 80000 49224 6 pcpi_rs2[15]
port 327 nsew signal output
rlabel metal3 s 79600 49728 80000 49784 6 pcpi_rs2[16]
port 328 nsew signal output
rlabel metal3 s 79600 50288 80000 50344 6 pcpi_rs2[17]
port 329 nsew signal output
rlabel metal3 s 79600 50848 80000 50904 6 pcpi_rs2[18]
port 330 nsew signal output
rlabel metal3 s 79600 51408 80000 51464 6 pcpi_rs2[19]
port 331 nsew signal output
rlabel metal3 s 79600 41328 80000 41384 6 pcpi_rs2[1]
port 332 nsew signal output
rlabel metal3 s 79600 51968 80000 52024 6 pcpi_rs2[20]
port 333 nsew signal output
rlabel metal3 s 79600 52528 80000 52584 6 pcpi_rs2[21]
port 334 nsew signal output
rlabel metal3 s 79600 53088 80000 53144 6 pcpi_rs2[22]
port 335 nsew signal output
rlabel metal3 s 79600 53648 80000 53704 6 pcpi_rs2[23]
port 336 nsew signal output
rlabel metal3 s 79600 54208 80000 54264 6 pcpi_rs2[24]
port 337 nsew signal output
rlabel metal3 s 79600 54768 80000 54824 6 pcpi_rs2[25]
port 338 nsew signal output
rlabel metal3 s 79600 55328 80000 55384 6 pcpi_rs2[26]
port 339 nsew signal output
rlabel metal3 s 79600 55888 80000 55944 6 pcpi_rs2[27]
port 340 nsew signal output
rlabel metal3 s 79600 56448 80000 56504 6 pcpi_rs2[28]
port 341 nsew signal output
rlabel metal3 s 79600 57008 80000 57064 6 pcpi_rs2[29]
port 342 nsew signal output
rlabel metal3 s 79600 41888 80000 41944 6 pcpi_rs2[2]
port 343 nsew signal output
rlabel metal3 s 79600 57568 80000 57624 6 pcpi_rs2[30]
port 344 nsew signal output
rlabel metal3 s 79600 58128 80000 58184 6 pcpi_rs2[31]
port 345 nsew signal output
rlabel metal3 s 79600 42448 80000 42504 6 pcpi_rs2[3]
port 346 nsew signal output
rlabel metal3 s 79600 43008 80000 43064 6 pcpi_rs2[4]
port 347 nsew signal output
rlabel metal3 s 79600 43568 80000 43624 6 pcpi_rs2[5]
port 348 nsew signal output
rlabel metal3 s 79600 44128 80000 44184 6 pcpi_rs2[6]
port 349 nsew signal output
rlabel metal3 s 79600 44688 80000 44744 6 pcpi_rs2[7]
port 350 nsew signal output
rlabel metal3 s 79600 45248 80000 45304 6 pcpi_rs2[8]
port 351 nsew signal output
rlabel metal3 s 79600 45808 80000 45864 6 pcpi_rs2[9]
port 352 nsew signal output
rlabel metal3 s 79600 4368 80000 4424 6 pcpi_valid
port 353 nsew signal output
rlabel metal3 s 79600 3808 80000 3864 6 resetn
port 354 nsew signal input
rlabel metal4 s 2224 1538 2384 138406 6 vdd
port 355 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 138406 6 vdd
port 355 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 138406 6 vdd
port 355 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 138406 6 vdd
port 355 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 138406 6 vdd
port 355 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 138406 6 vdd
port 355 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 138406 6 vss
port 356 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 138406 6 vss
port 356 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 138406 6 vss
port 356 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 138406 6 vss
port 356 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 138406 6 vss
port 356 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 80000 140000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 30558716
string GDS_FILE /home/luke/picosoc-w-approximation/openlane/cpu/runs/23_12_10_11_29/results/signoff/cpu.magic.gds
string GDS_START 546950
<< end >>


magic
tech gf180mcuD
magscale 1 10
timestamp 1702206088
<< metal1 >>
rect 24210 56702 24222 56754
rect 24274 56751 24286 56754
rect 24882 56751 24894 56754
rect 24274 56705 24894 56751
rect 24274 56702 24286 56705
rect 24882 56702 24894 56705
rect 24946 56702 24958 56754
rect 38322 56702 38334 56754
rect 38386 56751 38398 56754
rect 40226 56751 40238 56754
rect 38386 56705 40238 56751
rect 38386 56702 38398 56705
rect 40226 56702 40238 56705
rect 40290 56702 40302 56754
rect 50418 56702 50430 56754
rect 50482 56751 50494 56754
rect 51202 56751 51214 56754
rect 50482 56705 51214 56751
rect 50482 56702 50494 56705
rect 51202 56702 51214 56705
rect 51266 56702 51278 56754
rect 23986 56590 23998 56642
rect 24050 56639 24062 56642
rect 25106 56639 25118 56642
rect 24050 56593 25118 56639
rect 24050 56590 24062 56593
rect 25106 56590 25118 56593
rect 25170 56590 25182 56642
rect 1344 56474 58576 56508
rect 1344 56422 19838 56474
rect 19890 56422 19942 56474
rect 19994 56422 20046 56474
rect 20098 56422 50558 56474
rect 50610 56422 50662 56474
rect 50714 56422 50766 56474
rect 50818 56422 58576 56474
rect 1344 56388 58576 56422
rect 23438 56306 23490 56318
rect 23438 56242 23490 56254
rect 24894 56306 24946 56318
rect 24894 56242 24946 56254
rect 33182 56306 33234 56318
rect 33182 56242 33234 56254
rect 41022 56306 41074 56318
rect 41022 56242 41074 56254
rect 43038 56306 43090 56318
rect 43038 56242 43090 56254
rect 49758 56306 49810 56318
rect 49758 56242 49810 56254
rect 51214 56306 51266 56318
rect 51214 56242 51266 56254
rect 23662 56194 23714 56206
rect 23662 56130 23714 56142
rect 23998 56194 24050 56206
rect 31278 56194 31330 56206
rect 41358 56194 41410 56206
rect 24546 56142 24558 56194
rect 24610 56142 24622 56194
rect 35074 56142 35086 56194
rect 35138 56142 35150 56194
rect 38882 56142 38894 56194
rect 38946 56142 38958 56194
rect 40674 56142 40686 56194
rect 40738 56142 40750 56194
rect 23998 56130 24050 56142
rect 31278 56130 31330 56142
rect 41358 56130 41410 56142
rect 43710 56194 43762 56206
rect 43710 56130 43762 56142
rect 49982 56194 50034 56206
rect 49982 56130 50034 56142
rect 50318 56194 50370 56206
rect 51538 56142 51550 56194
rect 51602 56142 51614 56194
rect 50318 56130 50370 56142
rect 35422 56082 35474 56094
rect 39230 56082 39282 56094
rect 42590 56082 42642 56094
rect 27794 56030 27806 56082
rect 27858 56030 27870 56082
rect 30594 56030 30606 56082
rect 30658 56030 30670 56082
rect 31490 56030 31502 56082
rect 31554 56030 31566 56082
rect 32162 56030 32174 56082
rect 32226 56030 32238 56082
rect 38546 56030 38558 56082
rect 38610 56030 38622 56082
rect 40226 56030 40238 56082
rect 40290 56030 40302 56082
rect 41570 56030 41582 56082
rect 41634 56030 41646 56082
rect 35422 56018 35474 56030
rect 39230 56018 39282 56030
rect 42590 56018 42642 56030
rect 28590 55970 28642 55982
rect 25554 55918 25566 55970
rect 25618 55918 25630 55970
rect 28590 55906 28642 55918
rect 36206 55970 36258 55982
rect 36206 55906 36258 55918
rect 39790 55970 39842 55982
rect 39790 55906 39842 55918
rect 42142 55970 42194 55982
rect 42142 55906 42194 55918
rect 1344 55690 58576 55724
rect 1344 55638 4478 55690
rect 4530 55638 4582 55690
rect 4634 55638 4686 55690
rect 4738 55638 35198 55690
rect 35250 55638 35302 55690
rect 35354 55638 35406 55690
rect 35458 55638 58576 55690
rect 1344 55604 58576 55638
rect 24670 55522 24722 55534
rect 24670 55458 24722 55470
rect 24222 55410 24274 55422
rect 24222 55346 24274 55358
rect 28142 55410 28194 55422
rect 28142 55346 28194 55358
rect 28590 55410 28642 55422
rect 28590 55346 28642 55358
rect 30270 55410 30322 55422
rect 30270 55346 30322 55358
rect 31278 55410 31330 55422
rect 31278 55346 31330 55358
rect 33518 55410 33570 55422
rect 33518 55346 33570 55358
rect 37214 55410 37266 55422
rect 37214 55346 37266 55358
rect 42030 55410 42082 55422
rect 42030 55346 42082 55358
rect 50990 55410 51042 55422
rect 50990 55346 51042 55358
rect 29150 55298 29202 55310
rect 27010 55246 27022 55298
rect 27074 55246 27086 55298
rect 27458 55246 27470 55298
rect 27522 55246 27534 55298
rect 29150 55234 29202 55246
rect 29710 55298 29762 55310
rect 29710 55234 29762 55246
rect 30494 55298 30546 55310
rect 35646 55298 35698 55310
rect 39902 55298 39954 55310
rect 32498 55246 32510 55298
rect 32562 55246 32574 55298
rect 39442 55246 39454 55298
rect 39506 55246 39518 55298
rect 30494 55234 30546 55246
rect 35646 55234 35698 55246
rect 39902 55234 39954 55246
rect 40126 55298 40178 55310
rect 42478 55298 42530 55310
rect 41010 55246 41022 55298
rect 41074 55246 41086 55298
rect 40126 55234 40178 55246
rect 42478 55234 42530 55246
rect 35422 55186 35474 55198
rect 35422 55122 35474 55134
rect 36430 55186 36482 55198
rect 36430 55122 36482 55134
rect 41582 55186 41634 55198
rect 41582 55122 41634 55134
rect 27694 55074 27746 55086
rect 27694 55010 27746 55022
rect 30830 55074 30882 55086
rect 30830 55010 30882 55022
rect 31726 55074 31778 55086
rect 31726 55010 31778 55022
rect 32174 55074 32226 55086
rect 40798 55074 40850 55086
rect 35970 55022 35982 55074
rect 36034 55022 36046 55074
rect 40450 55022 40462 55074
rect 40514 55022 40526 55074
rect 32174 55010 32226 55022
rect 40798 55010 40850 55022
rect 1344 54906 58576 54940
rect 1344 54854 19838 54906
rect 19890 54854 19942 54906
rect 19994 54854 20046 54906
rect 20098 54854 50558 54906
rect 50610 54854 50662 54906
rect 50714 54854 50766 54906
rect 50818 54854 58576 54906
rect 1344 54820 58576 54854
rect 26238 54738 26290 54750
rect 26238 54674 26290 54686
rect 26462 54738 26514 54750
rect 26462 54674 26514 54686
rect 28926 54738 28978 54750
rect 28926 54674 28978 54686
rect 29822 54738 29874 54750
rect 29822 54674 29874 54686
rect 34190 54738 34242 54750
rect 34190 54674 34242 54686
rect 28478 54626 28530 54638
rect 28478 54562 28530 54574
rect 29150 54626 29202 54638
rect 29150 54562 29202 54574
rect 29486 54626 29538 54638
rect 32398 54626 32450 54638
rect 38782 54626 38834 54638
rect 30146 54574 30158 54626
rect 30210 54574 30222 54626
rect 36082 54574 36094 54626
rect 36146 54574 36158 54626
rect 37538 54574 37550 54626
rect 37602 54574 37614 54626
rect 29486 54562 29538 54574
rect 32398 54562 32450 54574
rect 38782 54562 38834 54574
rect 39902 54626 39954 54638
rect 39902 54562 39954 54574
rect 41022 54626 41074 54638
rect 41022 54562 41074 54574
rect 32286 54514 32338 54526
rect 32286 54450 32338 54462
rect 32622 54514 32674 54526
rect 33170 54462 33182 54514
rect 33234 54462 33246 54514
rect 36306 54462 36318 54514
rect 36370 54462 36382 54514
rect 40114 54462 40126 54514
rect 40178 54462 40190 54514
rect 32622 54450 32674 54462
rect 27470 54402 27522 54414
rect 26898 54350 26910 54402
rect 26962 54350 26974 54402
rect 27470 54338 27522 54350
rect 27918 54402 27970 54414
rect 27918 54338 27970 54350
rect 31838 54402 31890 54414
rect 37202 54350 37214 54402
rect 37266 54350 37278 54402
rect 31838 54338 31890 54350
rect 39230 54290 39282 54302
rect 39230 54226 39282 54238
rect 1344 54122 58576 54156
rect 1344 54070 4478 54122
rect 4530 54070 4582 54122
rect 4634 54070 4686 54122
rect 4738 54070 35198 54122
rect 35250 54070 35302 54122
rect 35354 54070 35406 54122
rect 35458 54070 58576 54122
rect 1344 54036 58576 54070
rect 22654 53842 22706 53854
rect 37214 53842 37266 53854
rect 25218 53790 25230 53842
rect 25282 53790 25294 53842
rect 33506 53790 33518 53842
rect 33570 53790 33582 53842
rect 35858 53790 35870 53842
rect 35922 53790 35934 53842
rect 22654 53778 22706 53790
rect 37214 53778 37266 53790
rect 13470 53730 13522 53742
rect 21982 53730 22034 53742
rect 30270 53730 30322 53742
rect 34638 53730 34690 53742
rect 39902 53730 39954 53742
rect 13682 53678 13694 53730
rect 13746 53678 13758 53730
rect 22306 53678 22318 53730
rect 22370 53678 22382 53730
rect 24994 53678 25006 53730
rect 25058 53678 25070 53730
rect 30706 53678 30718 53730
rect 30770 53678 30782 53730
rect 32834 53678 32846 53730
rect 32898 53678 32910 53730
rect 35746 53678 35758 53730
rect 35810 53678 35822 53730
rect 38770 53678 38782 53730
rect 38834 53678 38846 53730
rect 13470 53666 13522 53678
rect 21982 53666 22034 53678
rect 30270 53666 30322 53678
rect 34638 53666 34690 53678
rect 39902 53666 39954 53678
rect 40238 53730 40290 53742
rect 40238 53666 40290 53678
rect 14254 53618 14306 53630
rect 14254 53554 14306 53566
rect 21310 53618 21362 53630
rect 21310 53554 21362 53566
rect 21534 53618 21586 53630
rect 21534 53554 21586 53566
rect 23886 53618 23938 53630
rect 23886 53554 23938 53566
rect 24110 53618 24162 53630
rect 24110 53554 24162 53566
rect 24446 53618 24498 53630
rect 24446 53554 24498 53566
rect 25902 53618 25954 53630
rect 25902 53554 25954 53566
rect 31166 53618 31218 53630
rect 35086 53618 35138 53630
rect 39566 53618 39618 53630
rect 32386 53566 32398 53618
rect 32450 53566 32462 53618
rect 33282 53566 33294 53618
rect 33346 53566 33358 53618
rect 37650 53566 37662 53618
rect 37714 53566 37726 53618
rect 31166 53554 31218 53566
rect 35086 53554 35138 53566
rect 39566 53554 39618 53566
rect 42590 53618 42642 53630
rect 42590 53554 42642 53566
rect 43374 53618 43426 53630
rect 43374 53554 43426 53566
rect 44830 53618 44882 53630
rect 44830 53554 44882 53566
rect 47854 53618 47906 53630
rect 47854 53554 47906 53566
rect 21758 53506 21810 53518
rect 21758 53442 21810 53454
rect 22542 53506 22594 53518
rect 22542 53442 22594 53454
rect 23662 53506 23714 53518
rect 23662 53442 23714 53454
rect 24334 53506 24386 53518
rect 24334 53442 24386 53454
rect 29934 53506 29986 53518
rect 40014 53506 40066 53518
rect 39106 53454 39118 53506
rect 39170 53454 39182 53506
rect 29934 53442 29986 53454
rect 40014 53442 40066 53454
rect 42366 53506 42418 53518
rect 42366 53442 42418 53454
rect 42702 53506 42754 53518
rect 42702 53442 42754 53454
rect 42926 53506 42978 53518
rect 42926 53442 42978 53454
rect 43038 53506 43090 53518
rect 43038 53442 43090 53454
rect 43262 53506 43314 53518
rect 43262 53442 43314 53454
rect 44942 53506 44994 53518
rect 44942 53442 44994 53454
rect 45166 53506 45218 53518
rect 45166 53442 45218 53454
rect 1344 53338 58576 53372
rect 1344 53286 19838 53338
rect 19890 53286 19942 53338
rect 19994 53286 20046 53338
rect 20098 53286 50558 53338
rect 50610 53286 50662 53338
rect 50714 53286 50766 53338
rect 50818 53286 58576 53338
rect 1344 53252 58576 53286
rect 24782 53170 24834 53182
rect 13906 53118 13918 53170
rect 13970 53118 13982 53170
rect 24782 53106 24834 53118
rect 29150 53170 29202 53182
rect 29150 53106 29202 53118
rect 30046 53170 30098 53182
rect 41022 53170 41074 53182
rect 39330 53118 39342 53170
rect 39394 53118 39406 53170
rect 30046 53106 30098 53118
rect 41022 53106 41074 53118
rect 15598 53058 15650 53070
rect 12562 53006 12574 53058
rect 12626 53006 12638 53058
rect 15598 52994 15650 53006
rect 16158 53058 16210 53070
rect 21534 53058 21586 53070
rect 24558 53058 24610 53070
rect 31614 53058 31666 53070
rect 18050 53006 18062 53058
rect 18114 53006 18126 53058
rect 22418 53006 22430 53058
rect 22482 53006 22494 53058
rect 26450 53006 26462 53058
rect 26514 53006 26526 53058
rect 16158 52994 16210 53006
rect 21534 52994 21586 53006
rect 24558 52994 24610 53006
rect 31614 52994 31666 53006
rect 31838 53058 31890 53070
rect 36990 53058 37042 53070
rect 33394 53006 33406 53058
rect 33458 53006 33470 53058
rect 35410 53006 35422 53058
rect 35474 53006 35486 53058
rect 31838 52994 31890 53006
rect 36990 52994 37042 53006
rect 37102 53058 37154 53070
rect 37102 52994 37154 53006
rect 38782 53058 38834 53070
rect 38782 52994 38834 53006
rect 41134 53058 41186 53070
rect 41134 52994 41186 53006
rect 41358 53058 41410 53070
rect 49086 53058 49138 53070
rect 44258 53006 44270 53058
rect 44322 53006 44334 53058
rect 45714 53006 45726 53058
rect 45778 53006 45790 53058
rect 41358 52994 41410 53006
rect 49086 52994 49138 53006
rect 15486 52946 15538 52958
rect 24446 52946 24498 52958
rect 31390 52946 31442 52958
rect 37886 52946 37938 52958
rect 40910 52946 40962 52958
rect 42926 52946 42978 52958
rect 10434 52894 10446 52946
rect 10498 52894 10510 52946
rect 12786 52894 12798 52946
rect 12850 52894 12862 52946
rect 13458 52894 13470 52946
rect 13522 52894 13534 52946
rect 17378 52894 17390 52946
rect 17442 52894 17454 52946
rect 17938 52894 17950 52946
rect 18002 52894 18014 52946
rect 19618 52894 19630 52946
rect 19682 52894 19694 52946
rect 20626 52894 20638 52946
rect 20690 52894 20702 52946
rect 23650 52894 23662 52946
rect 23714 52894 23726 52946
rect 25666 52894 25678 52946
rect 25730 52894 25742 52946
rect 26226 52894 26238 52946
rect 26290 52894 26302 52946
rect 32050 52894 32062 52946
rect 32114 52894 32126 52946
rect 33842 52894 33854 52946
rect 33906 52894 33918 52946
rect 35298 52894 35310 52946
rect 35362 52894 35374 52946
rect 36754 52894 36766 52946
rect 36818 52894 36830 52946
rect 40114 52894 40126 52946
rect 40178 52894 40190 52946
rect 42690 52894 42702 52946
rect 42754 52894 42766 52946
rect 15486 52882 15538 52894
rect 24446 52882 24498 52894
rect 31390 52882 31442 52894
rect 37886 52882 37938 52894
rect 40910 52882 40962 52894
rect 42926 52882 42978 52894
rect 43374 52946 43426 52958
rect 48862 52946 48914 52958
rect 44482 52894 44494 52946
rect 44546 52894 44558 52946
rect 46946 52894 46958 52946
rect 47010 52894 47022 52946
rect 43374 52882 43426 52894
rect 48862 52882 48914 52894
rect 49198 52946 49250 52958
rect 49198 52882 49250 52894
rect 11118 52834 11170 52846
rect 10322 52782 10334 52834
rect 10386 52782 10398 52834
rect 11118 52770 11170 52782
rect 14926 52834 14978 52846
rect 20078 52834 20130 52846
rect 22094 52834 22146 52846
rect 18386 52782 18398 52834
rect 18450 52782 18462 52834
rect 19170 52782 19182 52834
rect 19234 52782 19246 52834
rect 20738 52782 20750 52834
rect 20802 52782 20814 52834
rect 14926 52770 14978 52782
rect 20078 52770 20130 52782
rect 22094 52770 22146 52782
rect 24110 52834 24162 52846
rect 24110 52770 24162 52782
rect 25342 52834 25394 52846
rect 29710 52834 29762 52846
rect 26338 52782 26350 52834
rect 26402 52782 26414 52834
rect 25342 52770 25394 52782
rect 29710 52770 29762 52782
rect 30606 52834 30658 52846
rect 30606 52770 30658 52782
rect 35982 52834 36034 52846
rect 35982 52770 36034 52782
rect 38446 52834 38498 52846
rect 38446 52770 38498 52782
rect 39678 52834 39730 52846
rect 39678 52770 39730 52782
rect 42030 52834 42082 52846
rect 42030 52770 42082 52782
rect 43598 52834 43650 52846
rect 49646 52834 49698 52846
rect 45154 52782 45166 52834
rect 45218 52782 45230 52834
rect 47618 52782 47630 52834
rect 47682 52782 47694 52834
rect 43598 52770 43650 52782
rect 49646 52770 49698 52782
rect 15598 52722 15650 52734
rect 39006 52722 39058 52734
rect 32386 52670 32398 52722
rect 32450 52670 32462 52722
rect 37538 52670 37550 52722
rect 37602 52670 37614 52722
rect 15598 52658 15650 52670
rect 39006 52658 39058 52670
rect 43934 52722 43986 52734
rect 43934 52658 43986 52670
rect 1344 52554 58576 52588
rect 1344 52502 4478 52554
rect 4530 52502 4582 52554
rect 4634 52502 4686 52554
rect 4738 52502 35198 52554
rect 35250 52502 35302 52554
rect 35354 52502 35406 52554
rect 35458 52502 58576 52554
rect 1344 52468 58576 52502
rect 37998 52386 38050 52398
rect 10994 52334 11006 52386
rect 11058 52334 11070 52386
rect 24658 52334 24670 52386
rect 24722 52334 24734 52386
rect 37998 52322 38050 52334
rect 17278 52274 17330 52286
rect 27134 52274 27186 52286
rect 10322 52222 10334 52274
rect 10386 52222 10398 52274
rect 14578 52222 14590 52274
rect 14642 52222 14654 52274
rect 16594 52222 16606 52274
rect 16658 52222 16670 52274
rect 26226 52222 26238 52274
rect 26290 52222 26302 52274
rect 17278 52210 17330 52222
rect 27134 52210 27186 52222
rect 31502 52274 31554 52286
rect 50878 52274 50930 52286
rect 38770 52222 38782 52274
rect 38834 52222 38846 52274
rect 43586 52222 43598 52274
rect 43650 52222 43662 52274
rect 45378 52222 45390 52274
rect 45442 52222 45454 52274
rect 31502 52210 31554 52222
rect 50878 52210 50930 52222
rect 7982 52162 8034 52174
rect 11790 52162 11842 52174
rect 7634 52110 7646 52162
rect 7698 52110 7710 52162
rect 10434 52110 10446 52162
rect 10498 52110 10510 52162
rect 7982 52098 8034 52110
rect 11790 52098 11842 52110
rect 12350 52162 12402 52174
rect 19742 52162 19794 52174
rect 22878 52162 22930 52174
rect 24222 52162 24274 52174
rect 29822 52162 29874 52174
rect 14130 52110 14142 52162
rect 14194 52110 14206 52162
rect 15138 52110 15150 52162
rect 15202 52110 15214 52162
rect 15698 52110 15710 52162
rect 15762 52110 15774 52162
rect 18610 52110 18622 52162
rect 18674 52110 18686 52162
rect 20178 52110 20190 52162
rect 20242 52110 20254 52162
rect 21298 52110 21310 52162
rect 21362 52110 21374 52162
rect 21858 52110 21870 52162
rect 21922 52110 21934 52162
rect 23090 52110 23102 52162
rect 23154 52110 23166 52162
rect 23314 52110 23326 52162
rect 23378 52110 23390 52162
rect 24434 52110 24446 52162
rect 24498 52110 24510 52162
rect 26002 52110 26014 52162
rect 26066 52110 26078 52162
rect 27346 52110 27358 52162
rect 27410 52110 27422 52162
rect 12350 52098 12402 52110
rect 19742 52098 19794 52110
rect 22878 52098 22930 52110
rect 24222 52098 24274 52110
rect 29822 52098 29874 52110
rect 29934 52162 29986 52174
rect 29934 52098 29986 52110
rect 30046 52162 30098 52174
rect 30942 52162 30994 52174
rect 36094 52162 36146 52174
rect 30258 52110 30270 52162
rect 30322 52110 30334 52162
rect 33506 52110 33518 52162
rect 33570 52110 33582 52162
rect 33954 52110 33966 52162
rect 34018 52110 34030 52162
rect 35522 52110 35534 52162
rect 35586 52110 35598 52162
rect 30046 52098 30098 52110
rect 30942 52098 30994 52110
rect 36094 52098 36146 52110
rect 36990 52162 37042 52174
rect 36990 52098 37042 52110
rect 37214 52162 37266 52174
rect 38334 52162 38386 52174
rect 37538 52110 37550 52162
rect 37602 52110 37614 52162
rect 37214 52098 37266 52110
rect 38334 52098 38386 52110
rect 38670 52162 38722 52174
rect 42478 52162 42530 52174
rect 40002 52110 40014 52162
rect 40066 52110 40078 52162
rect 41122 52110 41134 52162
rect 41186 52110 41198 52162
rect 38670 52098 38722 52110
rect 42478 52098 42530 52110
rect 42590 52162 42642 52174
rect 48078 52162 48130 52174
rect 42802 52110 42814 52162
rect 42866 52110 42878 52162
rect 43250 52110 43262 52162
rect 43314 52110 43326 52162
rect 45714 52110 45726 52162
rect 45778 52110 45790 52162
rect 46946 52110 46958 52162
rect 47010 52110 47022 52162
rect 42590 52098 42642 52110
rect 48078 52098 48130 52110
rect 48414 52162 48466 52174
rect 48850 52110 48862 52162
rect 48914 52110 48926 52162
rect 49298 52110 49310 52162
rect 49362 52110 49374 52162
rect 50194 52110 50206 52162
rect 50258 52110 50270 52162
rect 48414 52098 48466 52110
rect 8094 52050 8146 52062
rect 8094 51986 8146 51998
rect 12238 52050 12290 52062
rect 12238 51986 12290 51998
rect 12462 52050 12514 52062
rect 19294 52050 19346 52062
rect 14578 51998 14590 52050
rect 14642 51998 14654 52050
rect 17602 51998 17614 52050
rect 17666 51998 17678 52050
rect 12462 51986 12514 51998
rect 19294 51986 19346 51998
rect 19630 52050 19682 52062
rect 26686 52050 26738 52062
rect 21970 51998 21982 52050
rect 22034 51998 22046 52050
rect 19630 51986 19682 51998
rect 26686 51986 26738 51998
rect 27022 52050 27074 52062
rect 36318 52050 36370 52062
rect 32610 51998 32622 52050
rect 32674 51998 32686 52050
rect 27022 51986 27074 51998
rect 36318 51986 36370 51998
rect 36430 52050 36482 52062
rect 47630 52050 47682 52062
rect 37426 51998 37438 52050
rect 37490 51998 37502 52050
rect 39554 51998 39566 52050
rect 39618 51998 39630 52050
rect 41794 51998 41806 52050
rect 41858 51998 41870 52050
rect 36430 51986 36482 51998
rect 47630 51986 47682 51998
rect 48190 52050 48242 52062
rect 48190 51986 48242 51998
rect 48638 52050 48690 52062
rect 48638 51986 48690 51998
rect 30718 51938 30770 51950
rect 38446 51938 38498 51950
rect 21522 51886 21534 51938
rect 21586 51886 21598 51938
rect 32722 51886 32734 51938
rect 32786 51886 32798 51938
rect 30718 51874 30770 51886
rect 38446 51874 38498 51886
rect 38782 51938 38834 51950
rect 50418 51886 50430 51938
rect 50482 51886 50494 51938
rect 38782 51874 38834 51886
rect 1344 51770 58576 51804
rect 1344 51718 19838 51770
rect 19890 51718 19942 51770
rect 19994 51718 20046 51770
rect 20098 51718 50558 51770
rect 50610 51718 50662 51770
rect 50714 51718 50766 51770
rect 50818 51718 58576 51770
rect 1344 51684 58576 51718
rect 10446 51602 10498 51614
rect 10446 51538 10498 51550
rect 10894 51602 10946 51614
rect 10894 51538 10946 51550
rect 11118 51602 11170 51614
rect 20638 51602 20690 51614
rect 21646 51602 21698 51614
rect 16706 51550 16718 51602
rect 16770 51550 16782 51602
rect 21186 51550 21198 51602
rect 21250 51550 21262 51602
rect 11118 51538 11170 51550
rect 20638 51538 20690 51550
rect 21646 51538 21698 51550
rect 21870 51602 21922 51614
rect 21870 51538 21922 51550
rect 31054 51602 31106 51614
rect 31054 51538 31106 51550
rect 34638 51602 34690 51614
rect 34638 51538 34690 51550
rect 35646 51602 35698 51614
rect 36766 51602 36818 51614
rect 39454 51602 39506 51614
rect 36082 51550 36094 51602
rect 36146 51550 36158 51602
rect 39106 51550 39118 51602
rect 39170 51550 39182 51602
rect 35646 51538 35698 51550
rect 36766 51538 36818 51550
rect 39454 51538 39506 51550
rect 42926 51602 42978 51614
rect 42926 51538 42978 51550
rect 51550 51602 51602 51614
rect 51550 51538 51602 51550
rect 10222 51490 10274 51502
rect 20526 51490 20578 51502
rect 8306 51438 8318 51490
rect 8370 51438 8382 51490
rect 13234 51438 13246 51490
rect 13298 51438 13310 51490
rect 10222 51426 10274 51438
rect 20526 51426 20578 51438
rect 20862 51490 20914 51502
rect 20862 51426 20914 51438
rect 22542 51490 22594 51502
rect 22542 51426 22594 51438
rect 24446 51490 24498 51502
rect 24446 51426 24498 51438
rect 24558 51490 24610 51502
rect 24558 51426 24610 51438
rect 24782 51490 24834 51502
rect 24782 51426 24834 51438
rect 25566 51490 25618 51502
rect 25566 51426 25618 51438
rect 25678 51490 25730 51502
rect 30382 51490 30434 51502
rect 26338 51438 26350 51490
rect 26402 51438 26414 51490
rect 27570 51438 27582 51490
rect 27634 51438 27646 51490
rect 25678 51426 25730 51438
rect 30382 51426 30434 51438
rect 30494 51490 30546 51502
rect 30494 51426 30546 51438
rect 31614 51490 31666 51502
rect 31614 51426 31666 51438
rect 32510 51490 32562 51502
rect 32510 51426 32562 51438
rect 33070 51490 33122 51502
rect 33070 51426 33122 51438
rect 33406 51490 33458 51502
rect 33406 51426 33458 51438
rect 35534 51490 35586 51502
rect 42702 51490 42754 51502
rect 45502 51490 45554 51502
rect 37090 51438 37102 51490
rect 37154 51438 37166 51490
rect 37426 51438 37438 51490
rect 37490 51438 37502 51490
rect 43698 51438 43710 51490
rect 43762 51438 43774 51490
rect 35534 51426 35586 51438
rect 42702 51426 42754 51438
rect 45502 51426 45554 51438
rect 45614 51490 45666 51502
rect 45614 51426 45666 51438
rect 46958 51490 47010 51502
rect 51874 51438 51886 51490
rect 51938 51438 51950 51490
rect 46958 51426 47010 51438
rect 10110 51378 10162 51390
rect 6962 51326 6974 51378
rect 7026 51326 7038 51378
rect 7746 51326 7758 51378
rect 7810 51326 7822 51378
rect 10110 51314 10162 51326
rect 10782 51378 10834 51390
rect 10782 51314 10834 51326
rect 11790 51378 11842 51390
rect 16158 51378 16210 51390
rect 12002 51326 12014 51378
rect 12066 51326 12078 51378
rect 13570 51326 13582 51378
rect 13634 51326 13646 51378
rect 14466 51326 14478 51378
rect 14530 51326 14542 51378
rect 11790 51314 11842 51326
rect 16158 51314 16210 51326
rect 16382 51378 16434 51390
rect 19966 51378 20018 51390
rect 21534 51378 21586 51390
rect 29934 51378 29986 51390
rect 17938 51326 17950 51378
rect 18002 51326 18014 51378
rect 18946 51326 18958 51378
rect 19010 51326 19022 51378
rect 20290 51326 20302 51378
rect 20354 51326 20366 51378
rect 22194 51326 22206 51378
rect 22258 51326 22270 51378
rect 27346 51326 27358 51378
rect 27410 51326 27422 51378
rect 16382 51314 16434 51326
rect 19966 51314 20018 51326
rect 21534 51314 21586 51326
rect 29934 51314 29986 51326
rect 30718 51378 30770 51390
rect 34414 51378 34466 51390
rect 35086 51378 35138 51390
rect 32274 51326 32286 51378
rect 32338 51326 32350 51378
rect 34178 51326 34190 51378
rect 34242 51326 34254 51378
rect 34850 51326 34862 51378
rect 34914 51326 34926 51378
rect 30718 51314 30770 51326
rect 34414 51314 34466 51326
rect 35086 51314 35138 51326
rect 35758 51378 35810 51390
rect 37774 51378 37826 51390
rect 40910 51378 40962 51390
rect 36306 51326 36318 51378
rect 36370 51326 36382 51378
rect 38770 51326 38782 51378
rect 38834 51326 38846 51378
rect 35758 51314 35810 51326
rect 37774 51314 37826 51326
rect 40910 51314 40962 51326
rect 41358 51378 41410 51390
rect 41358 51314 41410 51326
rect 41806 51378 41858 51390
rect 43038 51378 43090 51390
rect 42466 51326 42478 51378
rect 42530 51326 42542 51378
rect 41806 51314 41858 51326
rect 43038 51314 43090 51326
rect 43486 51378 43538 51390
rect 45390 51378 45442 51390
rect 44146 51326 44158 51378
rect 44210 51326 44222 51378
rect 44706 51326 44718 51378
rect 44770 51326 44782 51378
rect 43486 51314 43538 51326
rect 45390 51314 45442 51326
rect 46286 51378 46338 51390
rect 46286 51314 46338 51326
rect 46510 51378 46562 51390
rect 46510 51314 46562 51326
rect 46622 51378 46674 51390
rect 46622 51314 46674 51326
rect 47854 51378 47906 51390
rect 47854 51314 47906 51326
rect 48750 51378 48802 51390
rect 50766 51378 50818 51390
rect 49074 51326 49086 51378
rect 49138 51326 49150 51378
rect 48750 51314 48802 51326
rect 50766 51314 50818 51326
rect 50990 51378 51042 51390
rect 50990 51314 51042 51326
rect 51326 51378 51378 51390
rect 51326 51314 51378 51326
rect 1822 51266 1874 51278
rect 26014 51266 26066 51278
rect 7970 51214 7982 51266
rect 8034 51214 8046 51266
rect 12338 51214 12350 51266
rect 12402 51214 12414 51266
rect 17490 51214 17502 51266
rect 17554 51214 17566 51266
rect 22306 51214 22318 51266
rect 22370 51214 22382 51266
rect 1822 51202 1874 51214
rect 26014 51202 26066 51214
rect 34526 51266 34578 51278
rect 34526 51202 34578 51214
rect 38558 51266 38610 51278
rect 38558 51202 38610 51214
rect 41134 51266 41186 51278
rect 41134 51202 41186 51214
rect 42814 51266 42866 51278
rect 42814 51202 42866 51214
rect 47294 51266 47346 51278
rect 49534 51266 49586 51278
rect 48962 51214 48974 51266
rect 49026 51214 49038 51266
rect 47294 51202 47346 51214
rect 49534 51202 49586 51214
rect 51102 51266 51154 51278
rect 51102 51202 51154 51214
rect 15822 51154 15874 51166
rect 25566 51154 25618 51166
rect 12450 51102 12462 51154
rect 12514 51102 12526 51154
rect 19170 51102 19182 51154
rect 19234 51102 19246 51154
rect 15822 51090 15874 51102
rect 25566 51090 25618 51102
rect 29710 51154 29762 51166
rect 29710 51090 29762 51102
rect 38222 51154 38274 51166
rect 38222 51090 38274 51102
rect 38334 51154 38386 51166
rect 38334 51090 38386 51102
rect 44158 51154 44210 51166
rect 49758 51154 49810 51166
rect 46050 51102 46062 51154
rect 46114 51102 46126 51154
rect 44158 51090 44210 51102
rect 49758 51090 49810 51102
rect 49982 51154 50034 51166
rect 49982 51090 50034 51102
rect 50430 51154 50482 51166
rect 50430 51090 50482 51102
rect 1344 50986 58576 51020
rect 1344 50934 4478 50986
rect 4530 50934 4582 50986
rect 4634 50934 4686 50986
rect 4738 50934 35198 50986
rect 35250 50934 35302 50986
rect 35354 50934 35406 50986
rect 35458 50934 58576 50986
rect 1344 50900 58576 50934
rect 8430 50818 8482 50830
rect 22542 50818 22594 50830
rect 12450 50766 12462 50818
rect 12514 50766 12526 50818
rect 17490 50766 17502 50818
rect 17554 50766 17566 50818
rect 38658 50766 38670 50818
rect 38722 50766 38734 50818
rect 8430 50754 8482 50766
rect 22542 50754 22594 50766
rect 7074 50654 7086 50706
rect 7138 50654 7150 50706
rect 8754 50654 8766 50706
rect 8818 50654 8830 50706
rect 14242 50654 14254 50706
rect 14306 50654 14318 50706
rect 17378 50654 17390 50706
rect 17442 50654 17454 50706
rect 24322 50654 24334 50706
rect 24386 50654 24398 50706
rect 27458 50654 27470 50706
rect 27522 50654 27534 50706
rect 32610 50654 32622 50706
rect 32674 50654 32686 50706
rect 37762 50654 37774 50706
rect 37826 50654 37838 50706
rect 39442 50654 39454 50706
rect 39506 50654 39518 50706
rect 41906 50654 41918 50706
rect 41970 50654 41982 50706
rect 47842 50654 47854 50706
rect 47906 50654 47918 50706
rect 48626 50654 48638 50706
rect 48690 50654 48702 50706
rect 50082 50654 50094 50706
rect 50146 50654 50158 50706
rect 8206 50594 8258 50606
rect 6850 50542 6862 50594
rect 6914 50542 6926 50594
rect 7186 50542 7198 50594
rect 7250 50542 7262 50594
rect 8206 50530 8258 50542
rect 9214 50594 9266 50606
rect 9214 50530 9266 50542
rect 11790 50594 11842 50606
rect 18174 50594 18226 50606
rect 12002 50542 12014 50594
rect 12066 50542 12078 50594
rect 13682 50542 13694 50594
rect 13746 50542 13758 50594
rect 15250 50542 15262 50594
rect 15314 50542 15326 50594
rect 16818 50542 16830 50594
rect 16882 50542 16894 50594
rect 11790 50530 11842 50542
rect 18174 50530 18226 50542
rect 20078 50594 20130 50606
rect 20078 50530 20130 50542
rect 20414 50594 20466 50606
rect 20414 50530 20466 50542
rect 22654 50594 22706 50606
rect 25678 50594 25730 50606
rect 30494 50594 30546 50606
rect 24210 50542 24222 50594
rect 24274 50542 24286 50594
rect 26674 50542 26686 50594
rect 26738 50542 26750 50594
rect 27010 50542 27022 50594
rect 27074 50542 27086 50594
rect 22654 50530 22706 50542
rect 25678 50530 25730 50542
rect 30494 50530 30546 50542
rect 31054 50594 31106 50606
rect 35086 50594 35138 50606
rect 33170 50542 33182 50594
rect 33234 50542 33246 50594
rect 34402 50542 34414 50594
rect 34466 50542 34478 50594
rect 31054 50530 31106 50542
rect 35086 50530 35138 50542
rect 36542 50594 36594 50606
rect 43150 50594 43202 50606
rect 37314 50542 37326 50594
rect 37378 50542 37390 50594
rect 38770 50542 38782 50594
rect 38834 50542 38846 50594
rect 40338 50542 40350 50594
rect 40402 50542 40414 50594
rect 41234 50542 41246 50594
rect 41298 50542 41310 50594
rect 36542 50530 36594 50542
rect 43150 50530 43202 50542
rect 43598 50594 43650 50606
rect 43598 50530 43650 50542
rect 43934 50594 43986 50606
rect 51662 50594 51714 50606
rect 44930 50542 44942 50594
rect 44994 50542 45006 50594
rect 47618 50542 47630 50594
rect 47682 50542 47694 50594
rect 48738 50542 48750 50594
rect 48802 50542 48814 50594
rect 49522 50542 49534 50594
rect 49586 50542 49598 50594
rect 43934 50530 43986 50542
rect 51662 50530 51714 50542
rect 51886 50594 51938 50606
rect 51886 50530 51938 50542
rect 1710 50482 1762 50494
rect 1710 50418 1762 50430
rect 2942 50482 2994 50494
rect 2942 50418 2994 50430
rect 3950 50482 4002 50494
rect 18398 50482 18450 50494
rect 5954 50430 5966 50482
rect 6018 50430 6030 50482
rect 7746 50430 7758 50482
rect 7810 50430 7822 50482
rect 3950 50418 4002 50430
rect 18398 50418 18450 50430
rect 18510 50482 18562 50494
rect 18510 50418 18562 50430
rect 21870 50482 21922 50494
rect 21870 50418 21922 50430
rect 21982 50482 22034 50494
rect 21982 50418 22034 50430
rect 22542 50482 22594 50494
rect 22542 50418 22594 50430
rect 24894 50482 24946 50494
rect 24894 50418 24946 50430
rect 25790 50482 25842 50494
rect 35422 50482 35474 50494
rect 27570 50430 27582 50482
rect 27634 50430 27646 50482
rect 32946 50430 32958 50482
rect 33010 50430 33022 50482
rect 33842 50430 33854 50482
rect 33906 50430 33918 50482
rect 25790 50418 25842 50430
rect 35422 50418 35474 50430
rect 36206 50482 36258 50494
rect 36206 50418 36258 50430
rect 36318 50482 36370 50494
rect 52670 50482 52722 50494
rect 37538 50430 37550 50482
rect 37602 50430 37614 50482
rect 43810 50430 43822 50482
rect 43874 50430 43886 50482
rect 45154 50430 45166 50482
rect 45218 50430 45230 50482
rect 45602 50430 45614 50482
rect 45666 50430 45678 50482
rect 36318 50418 36370 50430
rect 52670 50418 52722 50430
rect 52782 50482 52834 50494
rect 52782 50418 52834 50430
rect 53230 50482 53282 50494
rect 53230 50418 53282 50430
rect 2494 50370 2546 50382
rect 2034 50318 2046 50370
rect 2098 50318 2110 50370
rect 2494 50306 2546 50318
rect 3614 50370 3666 50382
rect 3614 50306 3666 50318
rect 5630 50370 5682 50382
rect 5630 50306 5682 50318
rect 20190 50370 20242 50382
rect 20190 50306 20242 50318
rect 21646 50370 21698 50382
rect 21646 50306 21698 50318
rect 26014 50370 26066 50382
rect 26014 50306 26066 50318
rect 42926 50370 42978 50382
rect 42926 50306 42978 50318
rect 51438 50370 51490 50382
rect 51438 50306 51490 50318
rect 51774 50370 51826 50382
rect 51774 50306 51826 50318
rect 53006 50370 53058 50382
rect 53006 50306 53058 50318
rect 53342 50370 53394 50382
rect 53342 50306 53394 50318
rect 1344 50202 58576 50236
rect 1344 50150 19838 50202
rect 19890 50150 19942 50202
rect 19994 50150 20046 50202
rect 20098 50150 50558 50202
rect 50610 50150 50662 50202
rect 50714 50150 50766 50202
rect 50818 50150 58576 50202
rect 1344 50116 58576 50150
rect 42254 50034 42306 50046
rect 47406 50034 47458 50046
rect 15698 49982 15710 50034
rect 15762 49982 15774 50034
rect 20850 49982 20862 50034
rect 20914 49982 20926 50034
rect 41794 49982 41806 50034
rect 41858 49982 41870 50034
rect 42578 49982 42590 50034
rect 42642 49982 42654 50034
rect 44930 49982 44942 50034
rect 44994 49982 45006 50034
rect 42254 49970 42306 49982
rect 47406 49970 47458 49982
rect 53902 50034 53954 50046
rect 53902 49970 53954 49982
rect 25790 49922 25842 49934
rect 53678 49922 53730 49934
rect 7410 49870 7422 49922
rect 7474 49870 7486 49922
rect 11330 49870 11342 49922
rect 11394 49870 11406 49922
rect 13570 49870 13582 49922
rect 13634 49870 13646 49922
rect 14130 49870 14142 49922
rect 14194 49870 14206 49922
rect 20178 49870 20190 49922
rect 20242 49870 20254 49922
rect 21634 49870 21646 49922
rect 21698 49870 21710 49922
rect 26898 49870 26910 49922
rect 26962 49870 26974 49922
rect 33394 49870 33406 49922
rect 33458 49870 33470 49922
rect 37650 49870 37662 49922
rect 37714 49870 37726 49922
rect 38882 49870 38894 49922
rect 38946 49870 38958 49922
rect 47730 49870 47742 49922
rect 47794 49870 47806 49922
rect 49522 49870 49534 49922
rect 49586 49870 49598 49922
rect 25790 49858 25842 49870
rect 53678 49858 53730 49870
rect 15374 49810 15426 49822
rect 20526 49810 20578 49822
rect 29822 49810 29874 49822
rect 8418 49758 8430 49810
rect 8482 49758 8494 49810
rect 11442 49758 11454 49810
rect 11506 49758 11518 49810
rect 12338 49758 12350 49810
rect 12402 49758 12414 49810
rect 13906 49758 13918 49810
rect 13970 49758 13982 49810
rect 19170 49758 19182 49810
rect 19234 49758 19246 49810
rect 19842 49758 19854 49810
rect 19906 49758 19918 49810
rect 22978 49758 22990 49810
rect 23042 49758 23054 49810
rect 27234 49758 27246 49810
rect 27298 49758 27310 49810
rect 27906 49758 27918 49810
rect 27970 49758 27982 49810
rect 15374 49746 15426 49758
rect 20526 49746 20578 49758
rect 29822 49746 29874 49758
rect 30158 49810 30210 49822
rect 30158 49746 30210 49758
rect 30382 49810 30434 49822
rect 30382 49746 30434 49758
rect 30606 49810 30658 49822
rect 32510 49810 32562 49822
rect 36318 49810 36370 49822
rect 41470 49810 41522 49822
rect 46622 49810 46674 49822
rect 32274 49758 32286 49810
rect 32338 49758 32350 49810
rect 34962 49758 34974 49810
rect 35026 49758 35038 49810
rect 36866 49758 36878 49810
rect 36930 49758 36942 49810
rect 37538 49758 37550 49810
rect 37602 49758 37614 49810
rect 38210 49758 38222 49810
rect 38274 49758 38286 49810
rect 39106 49758 39118 49810
rect 39170 49758 39182 49810
rect 43026 49758 43038 49810
rect 43090 49758 43102 49810
rect 43250 49758 43262 49810
rect 43314 49758 43326 49810
rect 44146 49758 44158 49810
rect 44210 49758 44222 49810
rect 44706 49758 44718 49810
rect 44770 49758 44782 49810
rect 30606 49746 30658 49758
rect 32510 49746 32562 49758
rect 36318 49746 36370 49758
rect 41470 49746 41522 49758
rect 46622 49746 46674 49758
rect 46734 49810 46786 49822
rect 46734 49746 46786 49758
rect 46958 49810 47010 49822
rect 51774 49810 51826 49822
rect 50418 49758 50430 49810
rect 50482 49758 50494 49810
rect 46958 49746 47010 49758
rect 51774 49746 51826 49758
rect 52110 49810 52162 49822
rect 52110 49746 52162 49758
rect 52334 49810 52386 49822
rect 52334 49746 52386 49758
rect 52782 49810 52834 49822
rect 52782 49746 52834 49758
rect 53006 49810 53058 49822
rect 53006 49746 53058 49758
rect 2046 49698 2098 49710
rect 2046 49634 2098 49646
rect 2494 49698 2546 49710
rect 2494 49634 2546 49646
rect 2830 49698 2882 49710
rect 2830 49634 2882 49646
rect 3390 49698 3442 49710
rect 3390 49634 3442 49646
rect 3726 49698 3778 49710
rect 3726 49634 3778 49646
rect 4174 49698 4226 49710
rect 4174 49634 4226 49646
rect 4622 49698 4674 49710
rect 8990 49698 9042 49710
rect 6850 49646 6862 49698
rect 6914 49646 6926 49698
rect 4622 49634 4674 49646
rect 8990 49634 9042 49646
rect 12910 49698 12962 49710
rect 12910 49634 12962 49646
rect 14590 49698 14642 49710
rect 23550 49698 23602 49710
rect 19618 49646 19630 49698
rect 19682 49646 19694 49698
rect 21410 49646 21422 49698
rect 21474 49646 21486 49698
rect 14590 49634 14642 49646
rect 23550 49634 23602 49646
rect 25902 49698 25954 49710
rect 25902 49634 25954 49646
rect 26014 49698 26066 49710
rect 26014 49634 26066 49646
rect 28590 49698 28642 49710
rect 51998 49698 52050 49710
rect 29362 49646 29374 49698
rect 29426 49646 29438 49698
rect 33170 49646 33182 49698
rect 33234 49646 33246 49698
rect 35746 49646 35758 49698
rect 35810 49646 35822 49698
rect 39218 49646 39230 49698
rect 39282 49646 39294 49698
rect 44034 49646 44046 49698
rect 44098 49646 44110 49698
rect 48962 49646 48974 49698
rect 49026 49646 49038 49698
rect 53890 49646 53902 49698
rect 53954 49646 53966 49698
rect 28590 49634 28642 49646
rect 51998 49634 52050 49646
rect 31054 49586 31106 49598
rect 47070 49586 47122 49598
rect 2034 49534 2046 49586
rect 2098 49583 2110 49586
rect 2370 49583 2382 49586
rect 2098 49537 2382 49583
rect 2098 49534 2110 49537
rect 2370 49534 2382 49537
rect 2434 49534 2446 49586
rect 31826 49534 31838 49586
rect 31890 49534 31902 49586
rect 36642 49534 36654 49586
rect 36706 49534 36718 49586
rect 31054 49522 31106 49534
rect 47070 49522 47122 49534
rect 51214 49586 51266 49598
rect 53330 49534 53342 49586
rect 53394 49534 53406 49586
rect 51214 49522 51266 49534
rect 1344 49418 58576 49452
rect 1344 49366 4478 49418
rect 4530 49366 4582 49418
rect 4634 49366 4686 49418
rect 4738 49366 35198 49418
rect 35250 49366 35302 49418
rect 35354 49366 35406 49418
rect 35458 49366 58576 49418
rect 1344 49332 58576 49366
rect 27582 49250 27634 49262
rect 7298 49198 7310 49250
rect 7362 49198 7374 49250
rect 19954 49198 19966 49250
rect 20018 49198 20030 49250
rect 27582 49186 27634 49198
rect 34750 49250 34802 49262
rect 34750 49186 34802 49198
rect 49534 49250 49586 49262
rect 49534 49186 49586 49198
rect 53118 49250 53170 49262
rect 53118 49186 53170 49198
rect 6974 49138 7026 49150
rect 21870 49138 21922 49150
rect 32734 49138 32786 49150
rect 7746 49086 7758 49138
rect 7810 49086 7822 49138
rect 15474 49086 15486 49138
rect 15538 49086 15550 49138
rect 16146 49086 16158 49138
rect 16210 49086 16222 49138
rect 24210 49086 24222 49138
rect 24274 49086 24286 49138
rect 6974 49074 7026 49086
rect 21870 49074 21922 49086
rect 32734 49074 32786 49086
rect 32846 49138 32898 49150
rect 32846 49074 32898 49086
rect 34302 49138 34354 49150
rect 34302 49074 34354 49086
rect 34526 49138 34578 49150
rect 34526 49074 34578 49086
rect 49086 49138 49138 49150
rect 53790 49138 53842 49150
rect 52770 49086 52782 49138
rect 52834 49086 52846 49138
rect 49086 49074 49138 49086
rect 53790 49074 53842 49086
rect 2382 49026 2434 49038
rect 2382 48962 2434 48974
rect 2942 49026 2994 49038
rect 2942 48962 2994 48974
rect 3278 49026 3330 49038
rect 3278 48962 3330 48974
rect 3950 49026 4002 49038
rect 3950 48962 4002 48974
rect 4846 49026 4898 49038
rect 4846 48962 4898 48974
rect 5182 49026 5234 49038
rect 5182 48962 5234 48974
rect 6190 49026 6242 49038
rect 6190 48962 6242 48974
rect 6526 49026 6578 49038
rect 6526 48962 6578 48974
rect 6750 49026 6802 49038
rect 13470 49026 13522 49038
rect 18510 49026 18562 49038
rect 9202 48974 9214 49026
rect 9266 48974 9278 49026
rect 11218 48974 11230 49026
rect 11282 48974 11294 49026
rect 13682 48974 13694 49026
rect 13746 48974 13758 49026
rect 14018 48974 14030 49026
rect 14082 48974 14094 49026
rect 15138 48974 15150 49026
rect 15202 48974 15214 49026
rect 16370 48974 16382 49026
rect 16434 48974 16446 49026
rect 6750 48962 6802 48974
rect 13470 48962 13522 48974
rect 18510 48962 18562 48974
rect 19294 49026 19346 49038
rect 19294 48962 19346 48974
rect 20190 49026 20242 49038
rect 22430 49026 22482 49038
rect 21970 48974 21982 49026
rect 22034 48974 22046 49026
rect 20190 48962 20242 48974
rect 22430 48962 22482 48974
rect 22654 49026 22706 49038
rect 23326 49026 23378 49038
rect 28254 49026 28306 49038
rect 22866 48974 22878 49026
rect 22930 48974 22942 49026
rect 23538 48974 23550 49026
rect 23602 48974 23614 49026
rect 24098 48974 24110 49026
rect 24162 48974 24174 49026
rect 26786 48974 26798 49026
rect 26850 48974 26862 49026
rect 27010 48974 27022 49026
rect 27074 48974 27086 49026
rect 28018 48974 28030 49026
rect 28082 48974 28094 49026
rect 22654 48962 22706 48974
rect 23326 48962 23378 48974
rect 28254 48962 28306 48974
rect 28590 49026 28642 49038
rect 28590 48962 28642 48974
rect 29822 49026 29874 49038
rect 33854 49026 33906 49038
rect 31042 48974 31054 49026
rect 31106 48974 31118 49026
rect 31490 48974 31502 49026
rect 31554 48974 31566 49026
rect 32498 48974 32510 49026
rect 32562 48974 32574 49026
rect 29822 48962 29874 48974
rect 33854 48962 33906 48974
rect 35198 49026 35250 49038
rect 35198 48962 35250 48974
rect 35534 49026 35586 49038
rect 37214 49026 37266 49038
rect 38334 49026 38386 49038
rect 46734 49026 46786 49038
rect 36082 48974 36094 49026
rect 36146 48974 36158 49026
rect 36978 48974 36990 49026
rect 37042 48974 37054 49026
rect 37650 48974 37662 49026
rect 37714 48974 37726 49026
rect 39554 48974 39566 49026
rect 39618 48974 39630 49026
rect 40674 48974 40686 49026
rect 40738 48974 40750 49026
rect 35534 48962 35586 48974
rect 37214 48962 37266 48974
rect 38334 48962 38386 48974
rect 46734 48962 46786 48974
rect 47294 49026 47346 49038
rect 47294 48962 47346 48974
rect 49422 49026 49474 49038
rect 50978 48974 50990 49026
rect 51042 48974 51054 49026
rect 51538 48974 51550 49026
rect 51602 48974 51614 49026
rect 49422 48962 49474 48974
rect 3838 48914 3890 48926
rect 3838 48850 3890 48862
rect 5854 48914 5906 48926
rect 5854 48850 5906 48862
rect 6302 48914 6354 48926
rect 11566 48914 11618 48926
rect 8194 48862 8206 48914
rect 8258 48862 8270 48914
rect 6302 48850 6354 48862
rect 11566 48850 11618 48862
rect 14702 48914 14754 48926
rect 14702 48850 14754 48862
rect 17054 48914 17106 48926
rect 17054 48850 17106 48862
rect 18846 48914 18898 48926
rect 18846 48850 18898 48862
rect 19406 48914 19458 48926
rect 19406 48850 19458 48862
rect 19518 48914 19570 48926
rect 19518 48850 19570 48862
rect 20750 48914 20802 48926
rect 20750 48850 20802 48862
rect 22542 48914 22594 48926
rect 28478 48914 28530 48926
rect 33182 48914 33234 48926
rect 24210 48862 24222 48914
rect 24274 48862 24286 48914
rect 30594 48862 30606 48914
rect 30658 48862 30670 48914
rect 31154 48862 31166 48914
rect 31218 48862 31230 48914
rect 31714 48862 31726 48914
rect 31778 48862 31790 48914
rect 22542 48850 22594 48862
rect 28478 48850 28530 48862
rect 33182 48850 33234 48862
rect 33406 48914 33458 48926
rect 46846 48914 46898 48926
rect 52894 48914 52946 48926
rect 35634 48862 35646 48914
rect 35698 48862 35710 48914
rect 35970 48862 35982 48914
rect 36034 48862 36046 48914
rect 37986 48862 37998 48914
rect 38050 48862 38062 48914
rect 39106 48862 39118 48914
rect 39170 48862 39182 48914
rect 41346 48862 41358 48914
rect 41410 48862 41422 48914
rect 50530 48862 50542 48914
rect 50594 48862 50606 48914
rect 33406 48850 33458 48862
rect 46846 48850 46898 48862
rect 52894 48850 52946 48862
rect 1710 48802 1762 48814
rect 2718 48802 2770 48814
rect 2034 48750 2046 48802
rect 2098 48750 2110 48802
rect 1710 48738 1762 48750
rect 2718 48738 2770 48750
rect 3166 48802 3218 48814
rect 3166 48738 3218 48750
rect 3614 48802 3666 48814
rect 3614 48738 3666 48750
rect 4510 48802 4562 48814
rect 4510 48738 4562 48750
rect 4958 48802 5010 48814
rect 4958 48738 5010 48750
rect 5518 48802 5570 48814
rect 5518 48738 5570 48750
rect 5742 48802 5794 48814
rect 5742 48738 5794 48750
rect 10558 48802 10610 48814
rect 10558 48738 10610 48750
rect 11454 48802 11506 48814
rect 11454 48738 11506 48750
rect 20526 48802 20578 48814
rect 20526 48738 20578 48750
rect 20862 48802 20914 48814
rect 20862 48738 20914 48750
rect 21534 48802 21586 48814
rect 21534 48738 21586 48750
rect 21758 48802 21810 48814
rect 33630 48802 33682 48814
rect 30146 48750 30158 48802
rect 30210 48750 30222 48802
rect 32050 48750 32062 48802
rect 32114 48750 32126 48802
rect 21758 48738 21810 48750
rect 33630 48738 33682 48750
rect 36542 48802 36594 48814
rect 36542 48738 36594 48750
rect 37326 48802 37378 48814
rect 37326 48738 37378 48750
rect 37438 48802 37490 48814
rect 37438 48738 37490 48750
rect 47070 48802 47122 48814
rect 47070 48738 47122 48750
rect 49534 48802 49586 48814
rect 53678 48802 53730 48814
rect 51426 48750 51438 48802
rect 51490 48750 51502 48802
rect 49534 48738 49586 48750
rect 53678 48738 53730 48750
rect 1344 48634 58576 48668
rect 1344 48582 19838 48634
rect 19890 48582 19942 48634
rect 19994 48582 20046 48634
rect 20098 48582 50558 48634
rect 50610 48582 50662 48634
rect 50714 48582 50766 48634
rect 50818 48582 58576 48634
rect 1344 48548 58576 48582
rect 18734 48466 18786 48478
rect 16706 48414 16718 48466
rect 16770 48414 16782 48466
rect 18734 48402 18786 48414
rect 19854 48466 19906 48478
rect 19854 48402 19906 48414
rect 20974 48466 21026 48478
rect 20974 48402 21026 48414
rect 21198 48466 21250 48478
rect 21198 48402 21250 48414
rect 22654 48466 22706 48478
rect 22654 48402 22706 48414
rect 30830 48466 30882 48478
rect 30830 48402 30882 48414
rect 32622 48466 32674 48478
rect 32622 48402 32674 48414
rect 35758 48466 35810 48478
rect 43710 48466 43762 48478
rect 50654 48466 50706 48478
rect 40226 48414 40238 48466
rect 40290 48414 40302 48466
rect 46050 48414 46062 48466
rect 46114 48414 46126 48466
rect 35758 48402 35810 48414
rect 43710 48402 43762 48414
rect 50654 48402 50706 48414
rect 53118 48466 53170 48478
rect 53118 48402 53170 48414
rect 53342 48466 53394 48478
rect 53342 48402 53394 48414
rect 2606 48354 2658 48366
rect 2146 48302 2158 48354
rect 2210 48302 2222 48354
rect 2606 48290 2658 48302
rect 2718 48354 2770 48366
rect 21982 48354 22034 48366
rect 9874 48302 9886 48354
rect 9938 48302 9950 48354
rect 10322 48302 10334 48354
rect 10386 48302 10398 48354
rect 11666 48302 11678 48354
rect 11730 48302 11742 48354
rect 15026 48302 15038 48354
rect 15090 48302 15102 48354
rect 2718 48290 2770 48302
rect 21982 48290 22034 48302
rect 22318 48354 22370 48366
rect 22318 48290 22370 48302
rect 25678 48354 25730 48366
rect 25678 48290 25730 48302
rect 25790 48354 25842 48366
rect 25790 48290 25842 48302
rect 26798 48354 26850 48366
rect 26798 48290 26850 48302
rect 29710 48354 29762 48366
rect 32286 48354 32338 48366
rect 31154 48302 31166 48354
rect 31218 48302 31230 48354
rect 29710 48290 29762 48302
rect 32286 48290 32338 48302
rect 32398 48354 32450 48366
rect 32398 48290 32450 48302
rect 34190 48354 34242 48366
rect 50878 48354 50930 48366
rect 36082 48302 36094 48354
rect 36146 48302 36158 48354
rect 37762 48302 37774 48354
rect 37826 48302 37838 48354
rect 38770 48302 38782 48354
rect 38834 48302 38846 48354
rect 40114 48302 40126 48354
rect 40178 48302 40190 48354
rect 41682 48302 41694 48354
rect 41746 48302 41758 48354
rect 44482 48302 44494 48354
rect 44546 48302 44558 48354
rect 46162 48302 46174 48354
rect 46226 48302 46238 48354
rect 34190 48290 34242 48302
rect 50878 48290 50930 48302
rect 50990 48354 51042 48366
rect 50990 48290 51042 48302
rect 3950 48242 4002 48254
rect 19294 48242 19346 48254
rect 21310 48242 21362 48254
rect 26238 48242 26290 48254
rect 1922 48190 1934 48242
rect 1986 48190 1998 48242
rect 3490 48190 3502 48242
rect 3554 48190 3566 48242
rect 4498 48190 4510 48242
rect 4562 48190 4574 48242
rect 5058 48190 5070 48242
rect 5122 48190 5134 48242
rect 6402 48190 6414 48242
rect 6466 48190 6478 48242
rect 7522 48190 7534 48242
rect 7586 48190 7598 48242
rect 7746 48190 7758 48242
rect 7810 48190 7822 48242
rect 9762 48190 9774 48242
rect 9826 48190 9838 48242
rect 12786 48190 12798 48242
rect 12850 48190 12862 48242
rect 16146 48190 16158 48242
rect 16210 48190 16222 48242
rect 18498 48190 18510 48242
rect 18562 48190 18574 48242
rect 19618 48190 19630 48242
rect 19682 48190 19694 48242
rect 21746 48190 21758 48242
rect 21810 48190 21822 48242
rect 3950 48178 4002 48190
rect 19294 48178 19346 48190
rect 21310 48178 21362 48190
rect 26238 48178 26290 48190
rect 26462 48242 26514 48254
rect 33518 48242 33570 48254
rect 30034 48190 30046 48242
rect 30098 48190 30110 48242
rect 26462 48178 26514 48190
rect 33518 48178 33570 48190
rect 33742 48242 33794 48254
rect 33742 48178 33794 48190
rect 34414 48242 34466 48254
rect 34414 48178 34466 48190
rect 34638 48242 34690 48254
rect 34638 48178 34690 48190
rect 34862 48242 34914 48254
rect 34862 48178 34914 48190
rect 35086 48242 35138 48254
rect 46846 48242 46898 48254
rect 36642 48190 36654 48242
rect 36706 48190 36718 48242
rect 37090 48190 37102 48242
rect 37154 48190 37166 48242
rect 38882 48190 38894 48242
rect 38946 48190 38958 48242
rect 42018 48190 42030 48242
rect 42082 48190 42094 48242
rect 43250 48190 43262 48242
rect 43314 48190 43326 48242
rect 47058 48190 47070 48242
rect 47122 48190 47134 48242
rect 53666 48190 53678 48242
rect 53730 48190 53742 48242
rect 35086 48178 35138 48190
rect 46846 48178 46898 48190
rect 4062 48130 4114 48142
rect 11006 48130 11058 48142
rect 26350 48130 26402 48142
rect 5954 48078 5966 48130
rect 6018 48078 6030 48130
rect 8306 48078 8318 48130
rect 8370 48078 8382 48130
rect 11442 48078 11454 48130
rect 11506 48078 11518 48130
rect 14690 48078 14702 48130
rect 14754 48078 14766 48130
rect 4062 48066 4114 48078
rect 11006 48066 11058 48078
rect 26350 48066 26402 48078
rect 29822 48130 29874 48142
rect 29822 48066 29874 48078
rect 33070 48130 33122 48142
rect 47742 48130 47794 48142
rect 37314 48078 37326 48130
rect 37378 48078 37390 48130
rect 44258 48078 44270 48130
rect 44322 48078 44334 48130
rect 33070 48066 33122 48078
rect 47742 48066 47794 48078
rect 53230 48130 53282 48142
rect 53230 48066 53282 48078
rect 2606 48018 2658 48030
rect 2606 47954 2658 47966
rect 14142 48018 14194 48030
rect 14142 47954 14194 47966
rect 19518 48018 19570 48030
rect 19518 47954 19570 47966
rect 25790 48018 25842 48030
rect 25790 47954 25842 47966
rect 33294 48018 33346 48030
rect 33294 47954 33346 47966
rect 1344 47850 58576 47884
rect 1344 47798 4478 47850
rect 4530 47798 4582 47850
rect 4634 47798 4686 47850
rect 4738 47798 35198 47850
rect 35250 47798 35302 47850
rect 35354 47798 35406 47850
rect 35458 47798 58576 47850
rect 1344 47764 58576 47798
rect 4286 47682 4338 47694
rect 3490 47630 3502 47682
rect 3554 47679 3566 47682
rect 3826 47679 3838 47682
rect 3554 47633 3838 47679
rect 3554 47630 3566 47633
rect 3826 47630 3838 47633
rect 3890 47630 3902 47682
rect 4286 47618 4338 47630
rect 4622 47682 4674 47694
rect 4622 47618 4674 47630
rect 5630 47682 5682 47694
rect 5630 47618 5682 47630
rect 5966 47682 6018 47694
rect 5966 47618 6018 47630
rect 32846 47682 32898 47694
rect 32846 47618 32898 47630
rect 3726 47570 3778 47582
rect 8318 47570 8370 47582
rect 21758 47570 21810 47582
rect 33406 47570 33458 47582
rect 7970 47518 7982 47570
rect 8034 47518 8046 47570
rect 11778 47518 11790 47570
rect 11842 47518 11854 47570
rect 14578 47518 14590 47570
rect 14642 47518 14654 47570
rect 17714 47518 17726 47570
rect 17778 47518 17790 47570
rect 23986 47518 23998 47570
rect 24050 47518 24062 47570
rect 31378 47518 31390 47570
rect 31442 47518 31454 47570
rect 41906 47518 41918 47570
rect 41970 47518 41982 47570
rect 47506 47518 47518 47570
rect 47570 47518 47582 47570
rect 51202 47518 51214 47570
rect 51266 47518 51278 47570
rect 3726 47506 3778 47518
rect 8318 47506 8370 47518
rect 21758 47506 21810 47518
rect 33406 47506 33458 47518
rect 1710 47458 1762 47470
rect 1710 47394 1762 47406
rect 2494 47458 2546 47470
rect 2494 47394 2546 47406
rect 2718 47458 2770 47470
rect 2718 47394 2770 47406
rect 4062 47458 4114 47470
rect 4062 47394 4114 47406
rect 5070 47458 5122 47470
rect 9774 47458 9826 47470
rect 17278 47458 17330 47470
rect 19630 47458 19682 47470
rect 7634 47406 7646 47458
rect 7698 47406 7710 47458
rect 10994 47406 11006 47458
rect 11058 47406 11070 47458
rect 12338 47406 12350 47458
rect 12402 47406 12414 47458
rect 13794 47406 13806 47458
rect 13858 47406 13870 47458
rect 14130 47406 14142 47458
rect 14194 47406 14206 47458
rect 15922 47406 15934 47458
rect 15986 47406 15998 47458
rect 16594 47406 16606 47458
rect 16658 47406 16670 47458
rect 17938 47406 17950 47458
rect 18002 47406 18014 47458
rect 5070 47394 5122 47406
rect 9774 47394 9826 47406
rect 17278 47394 17330 47406
rect 19630 47394 19682 47406
rect 19742 47458 19794 47470
rect 19742 47394 19794 47406
rect 21198 47458 21250 47470
rect 21198 47394 21250 47406
rect 21646 47458 21698 47470
rect 21646 47394 21698 47406
rect 22766 47458 22818 47470
rect 27022 47458 27074 47470
rect 30382 47458 30434 47470
rect 33518 47458 33570 47470
rect 38110 47458 38162 47470
rect 39230 47458 39282 47470
rect 43150 47458 43202 47470
rect 24210 47406 24222 47458
rect 24274 47406 24286 47458
rect 26002 47406 26014 47458
rect 26066 47406 26078 47458
rect 27346 47406 27358 47458
rect 27410 47406 27422 47458
rect 31042 47406 31054 47458
rect 31106 47406 31118 47458
rect 32050 47406 32062 47458
rect 32114 47406 32126 47458
rect 33170 47406 33182 47458
rect 33234 47406 33246 47458
rect 34962 47406 34974 47458
rect 35026 47406 35038 47458
rect 35410 47406 35422 47458
rect 35474 47406 35486 47458
rect 36306 47406 36318 47458
rect 36370 47406 36382 47458
rect 38322 47406 38334 47458
rect 38386 47406 38398 47458
rect 42130 47406 42142 47458
rect 42194 47406 42206 47458
rect 22766 47394 22818 47406
rect 27022 47394 27074 47406
rect 30382 47394 30434 47406
rect 33518 47394 33570 47406
rect 38110 47394 38162 47406
rect 39230 47394 39282 47406
rect 43150 47394 43202 47406
rect 44158 47458 44210 47470
rect 54126 47458 54178 47470
rect 49298 47406 49310 47458
rect 49362 47406 49374 47458
rect 51090 47406 51102 47458
rect 51154 47406 51166 47458
rect 53106 47406 53118 47458
rect 53170 47406 53182 47458
rect 54450 47406 54462 47458
rect 54514 47406 54526 47458
rect 44158 47394 44210 47406
rect 54126 47394 54178 47406
rect 5854 47346 5906 47358
rect 5854 47282 5906 47294
rect 6302 47346 6354 47358
rect 9550 47346 9602 47358
rect 6626 47294 6638 47346
rect 6690 47294 6702 47346
rect 6302 47282 6354 47294
rect 9550 47282 9602 47294
rect 9662 47346 9714 47358
rect 18622 47346 18674 47358
rect 10770 47294 10782 47346
rect 10834 47294 10846 47346
rect 14690 47294 14702 47346
rect 14754 47294 14766 47346
rect 15586 47294 15598 47346
rect 15650 47294 15662 47346
rect 9662 47282 9714 47294
rect 18622 47282 18674 47294
rect 19854 47346 19906 47358
rect 24782 47346 24834 47358
rect 20290 47294 20302 47346
rect 20354 47294 20366 47346
rect 19854 47282 19906 47294
rect 24782 47282 24834 47294
rect 25566 47346 25618 47358
rect 25566 47282 25618 47294
rect 30494 47346 30546 47358
rect 39006 47346 39058 47358
rect 31266 47294 31278 47346
rect 31330 47294 31342 47346
rect 35858 47294 35870 47346
rect 35922 47294 35934 47346
rect 30494 47282 30546 47294
rect 39006 47282 39058 47294
rect 39454 47346 39506 47358
rect 39454 47282 39506 47294
rect 39566 47346 39618 47358
rect 39566 47282 39618 47294
rect 42814 47346 42866 47358
rect 42814 47282 42866 47294
rect 43822 47346 43874 47358
rect 51662 47346 51714 47358
rect 48066 47294 48078 47346
rect 48130 47294 48142 47346
rect 49970 47294 49982 47346
rect 50034 47294 50046 47346
rect 52882 47294 52894 47346
rect 52946 47294 52958 47346
rect 43822 47282 43874 47294
rect 51662 47282 51714 47294
rect 3054 47234 3106 47246
rect 2034 47182 2046 47234
rect 2098 47182 2110 47234
rect 3054 47170 3106 47182
rect 3278 47234 3330 47246
rect 3278 47170 3330 47182
rect 3390 47234 3442 47246
rect 21870 47234 21922 47246
rect 10210 47182 10222 47234
rect 10274 47182 10286 47234
rect 3390 47170 3442 47182
rect 21870 47170 21922 47182
rect 22318 47234 22370 47246
rect 22318 47170 22370 47182
rect 23102 47234 23154 47246
rect 23102 47170 23154 47182
rect 23326 47234 23378 47246
rect 23326 47170 23378 47182
rect 23438 47234 23490 47246
rect 23438 47170 23490 47182
rect 30718 47234 30770 47246
rect 30718 47170 30770 47182
rect 33294 47234 33346 47246
rect 41470 47234 41522 47246
rect 43934 47234 43986 47246
rect 41122 47182 41134 47234
rect 41186 47182 41198 47234
rect 43474 47182 43486 47234
rect 43538 47182 43550 47234
rect 33294 47170 33346 47182
rect 41470 47170 41522 47182
rect 43934 47170 43986 47182
rect 1344 47066 58576 47100
rect 1344 47014 19838 47066
rect 19890 47014 19942 47066
rect 19994 47014 20046 47066
rect 20098 47014 50558 47066
rect 50610 47014 50662 47066
rect 50714 47014 50766 47066
rect 50818 47014 58576 47066
rect 1344 46980 58576 47014
rect 3838 46898 3890 46910
rect 12910 46898 12962 46910
rect 10882 46846 10894 46898
rect 10946 46846 10958 46898
rect 3838 46834 3890 46846
rect 12910 46834 12962 46846
rect 16046 46898 16098 46910
rect 22430 46898 22482 46910
rect 18050 46846 18062 46898
rect 18114 46846 18126 46898
rect 16046 46834 16098 46846
rect 22430 46834 22482 46846
rect 25790 46898 25842 46910
rect 25790 46834 25842 46846
rect 26014 46898 26066 46910
rect 43150 46898 43202 46910
rect 46062 46898 46114 46910
rect 26562 46846 26574 46898
rect 26626 46846 26638 46898
rect 45602 46846 45614 46898
rect 45666 46846 45678 46898
rect 26014 46834 26066 46846
rect 43150 46834 43202 46846
rect 46062 46834 46114 46846
rect 47966 46898 48018 46910
rect 51438 46898 51490 46910
rect 49074 46846 49086 46898
rect 49138 46846 49150 46898
rect 47966 46834 48018 46846
rect 51438 46834 51490 46846
rect 13806 46786 13858 46798
rect 4834 46734 4846 46786
rect 4898 46734 4910 46786
rect 5506 46734 5518 46786
rect 5570 46734 5582 46786
rect 6738 46734 6750 46786
rect 6802 46734 6814 46786
rect 10322 46734 10334 46786
rect 10386 46734 10398 46786
rect 10546 46734 10558 46786
rect 10610 46734 10622 46786
rect 13806 46722 13858 46734
rect 16270 46786 16322 46798
rect 16270 46722 16322 46734
rect 16382 46786 16434 46798
rect 16382 46722 16434 46734
rect 19406 46786 19458 46798
rect 19406 46722 19458 46734
rect 19630 46786 19682 46798
rect 19630 46722 19682 46734
rect 20302 46786 20354 46798
rect 20302 46722 20354 46734
rect 20750 46786 20802 46798
rect 22766 46786 22818 46798
rect 30942 46786 30994 46798
rect 21858 46734 21870 46786
rect 21922 46734 21934 46786
rect 24210 46734 24222 46786
rect 24274 46734 24286 46786
rect 27346 46734 27358 46786
rect 27410 46734 27422 46786
rect 29698 46734 29710 46786
rect 29762 46734 29774 46786
rect 20750 46722 20802 46734
rect 22766 46722 22818 46734
rect 30942 46722 30994 46734
rect 40014 46786 40066 46798
rect 40014 46722 40066 46734
rect 40126 46786 40178 46798
rect 40126 46722 40178 46734
rect 41246 46786 41298 46798
rect 41246 46722 41298 46734
rect 42030 46786 42082 46798
rect 47854 46786 47906 46798
rect 44146 46734 44158 46786
rect 44210 46734 44222 46786
rect 46386 46734 46398 46786
rect 46450 46734 46462 46786
rect 42030 46722 42082 46734
rect 47854 46722 47906 46734
rect 48190 46786 48242 46798
rect 51326 46786 51378 46798
rect 48962 46734 48974 46786
rect 49026 46734 49038 46786
rect 50418 46734 50430 46786
rect 50482 46734 50494 46786
rect 48190 46722 48242 46734
rect 51326 46722 51378 46734
rect 54126 46786 54178 46798
rect 54126 46722 54178 46734
rect 54238 46786 54290 46798
rect 54238 46722 54290 46734
rect 3054 46674 3106 46686
rect 3726 46674 3778 46686
rect 2370 46622 2382 46674
rect 2434 46622 2446 46674
rect 3378 46622 3390 46674
rect 3442 46622 3454 46674
rect 3054 46610 3106 46622
rect 3726 46610 3778 46622
rect 3950 46674 4002 46686
rect 12014 46674 12066 46686
rect 13358 46674 13410 46686
rect 4610 46622 4622 46674
rect 4674 46622 4686 46674
rect 6850 46622 6862 46674
rect 6914 46622 6926 46674
rect 7970 46622 7982 46674
rect 8034 46622 8046 46674
rect 10098 46622 10110 46674
rect 10162 46622 10174 46674
rect 12114 46622 12126 46674
rect 12178 46622 12190 46674
rect 3950 46610 4002 46622
rect 12014 46610 12066 46622
rect 13358 46610 13410 46622
rect 13470 46674 13522 46686
rect 13470 46610 13522 46622
rect 17726 46674 17778 46686
rect 17726 46610 17778 46622
rect 20078 46674 20130 46686
rect 20862 46674 20914 46686
rect 22206 46674 22258 46686
rect 20514 46622 20526 46674
rect 20578 46622 20590 46674
rect 21634 46622 21646 46674
rect 21698 46622 21710 46674
rect 20078 46610 20130 46622
rect 20862 46610 20914 46622
rect 22206 46610 22258 46622
rect 22542 46674 22594 46686
rect 26126 46674 26178 46686
rect 33070 46674 33122 46686
rect 41470 46674 41522 46686
rect 53006 46674 53058 46686
rect 23426 46622 23438 46674
rect 23490 46622 23502 46674
rect 23762 46622 23774 46674
rect 23826 46622 23838 46674
rect 25554 46622 25566 46674
rect 25618 46622 25630 46674
rect 26338 46622 26350 46674
rect 26402 46622 26414 46674
rect 26898 46622 26910 46674
rect 26962 46622 26974 46674
rect 29586 46622 29598 46674
rect 29650 46622 29662 46674
rect 33282 46622 33294 46674
rect 33346 46622 33358 46674
rect 34850 46622 34862 46674
rect 34914 46622 34926 46674
rect 36530 46622 36542 46674
rect 36594 46622 36606 46674
rect 36978 46622 36990 46674
rect 37042 46622 37054 46674
rect 40338 46622 40350 46674
rect 40402 46622 40414 46674
rect 41010 46622 41022 46674
rect 41074 46622 41086 46674
rect 41794 46622 41806 46674
rect 41858 46622 41870 46674
rect 42690 46622 42702 46674
rect 42754 46622 42766 46674
rect 42914 46622 42926 46674
rect 42978 46622 42990 46674
rect 45266 46622 45278 46674
rect 45330 46622 45342 46674
rect 52658 46622 52670 46674
rect 52722 46622 52734 46674
rect 53778 46622 53790 46674
rect 53842 46622 53854 46674
rect 22542 46610 22594 46622
rect 26126 46610 26178 46622
rect 33070 46610 33122 46622
rect 41470 46610 41522 46622
rect 53006 46610 53058 46622
rect 5854 46562 5906 46574
rect 13694 46562 13746 46574
rect 2594 46510 2606 46562
rect 2658 46510 2670 46562
rect 11890 46510 11902 46562
rect 11954 46510 11966 46562
rect 5854 46498 5906 46510
rect 13694 46498 13746 46510
rect 19854 46562 19906 46574
rect 31838 46562 31890 46574
rect 43710 46562 43762 46574
rect 53118 46562 53170 46574
rect 23650 46510 23662 46562
rect 23714 46510 23726 46562
rect 34962 46510 34974 46562
rect 35026 46510 35038 46562
rect 37538 46510 37550 46562
rect 37602 46510 37614 46562
rect 41906 46510 41918 46562
rect 41970 46510 41982 46562
rect 50866 46510 50878 46562
rect 50930 46510 50942 46562
rect 19854 46498 19906 46510
rect 31838 46498 31890 46510
rect 43710 46498 43762 46510
rect 53118 46498 53170 46510
rect 53454 46562 53506 46574
rect 53454 46498 53506 46510
rect 53566 46562 53618 46574
rect 53566 46498 53618 46510
rect 8990 46450 9042 46462
rect 43262 46450 43314 46462
rect 39554 46398 39566 46450
rect 39618 46398 39630 46450
rect 8990 46386 9042 46398
rect 43262 46386 43314 46398
rect 51438 46450 51490 46462
rect 51438 46386 51490 46398
rect 54238 46450 54290 46462
rect 54238 46386 54290 46398
rect 1344 46282 58576 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 58576 46282
rect 1344 46196 58576 46230
rect 31950 46114 32002 46126
rect 52782 46114 52834 46126
rect 22642 46062 22654 46114
rect 22706 46062 22718 46114
rect 32274 46062 32286 46114
rect 32338 46062 32350 46114
rect 33506 46062 33518 46114
rect 33570 46062 33582 46114
rect 31950 46050 32002 46062
rect 52782 46050 52834 46062
rect 22094 46002 22146 46014
rect 27134 46002 27186 46014
rect 31390 46002 31442 46014
rect 3042 45950 3054 46002
rect 3106 45950 3118 46002
rect 4162 45950 4174 46002
rect 4226 45950 4238 46002
rect 15698 45950 15710 46002
rect 15762 45950 15774 46002
rect 23090 45950 23102 46002
rect 23154 45950 23166 46002
rect 29250 45950 29262 46002
rect 29314 45950 29326 46002
rect 22094 45938 22146 45950
rect 27134 45938 27186 45950
rect 31390 45938 31442 45950
rect 31726 46002 31778 46014
rect 54798 46002 54850 46014
rect 32722 45950 32734 46002
rect 32786 45950 32798 46002
rect 48962 45950 48974 46002
rect 49026 45950 49038 46002
rect 54114 45950 54126 46002
rect 54178 45950 54190 46002
rect 31726 45938 31778 45950
rect 54798 45938 54850 45950
rect 1822 45890 1874 45902
rect 4510 45890 4562 45902
rect 6302 45890 6354 45902
rect 11118 45890 11170 45902
rect 13806 45890 13858 45902
rect 3154 45838 3166 45890
rect 3218 45838 3230 45890
rect 4946 45838 4958 45890
rect 5010 45838 5022 45890
rect 7634 45838 7646 45890
rect 7698 45838 7710 45890
rect 8418 45838 8430 45890
rect 8482 45838 8494 45890
rect 12898 45838 12910 45890
rect 12962 45838 12974 45890
rect 1822 45826 1874 45838
rect 4510 45826 4562 45838
rect 6302 45826 6354 45838
rect 11118 45826 11170 45838
rect 13806 45826 13858 45838
rect 13918 45890 13970 45902
rect 13918 45826 13970 45838
rect 14142 45890 14194 45902
rect 14142 45826 14194 45838
rect 22318 45890 22370 45902
rect 26014 45890 26066 45902
rect 24546 45838 24558 45890
rect 24610 45838 24622 45890
rect 22318 45826 22370 45838
rect 26014 45826 26066 45838
rect 27694 45890 27746 45902
rect 35870 45890 35922 45902
rect 30930 45838 30942 45890
rect 30994 45838 31006 45890
rect 33170 45838 33182 45890
rect 33234 45838 33246 45890
rect 33506 45838 33518 45890
rect 33570 45838 33582 45890
rect 34402 45838 34414 45890
rect 34466 45838 34478 45890
rect 35298 45838 35310 45890
rect 35362 45838 35374 45890
rect 27694 45826 27746 45838
rect 35870 45826 35922 45838
rect 36094 45890 36146 45902
rect 36094 45826 36146 45838
rect 38558 45890 38610 45902
rect 40910 45890 40962 45902
rect 38770 45838 38782 45890
rect 38834 45838 38846 45890
rect 38558 45826 38610 45838
rect 40910 45826 40962 45838
rect 41358 45890 41410 45902
rect 41358 45826 41410 45838
rect 41470 45890 41522 45902
rect 41470 45826 41522 45838
rect 41918 45890 41970 45902
rect 41918 45826 41970 45838
rect 42142 45890 42194 45902
rect 42142 45826 42194 45838
rect 43486 45890 43538 45902
rect 45054 45890 45106 45902
rect 43810 45838 43822 45890
rect 43874 45838 43886 45890
rect 43486 45826 43538 45838
rect 45054 45826 45106 45838
rect 45390 45890 45442 45902
rect 45390 45826 45442 45838
rect 47406 45890 47458 45902
rect 47406 45826 47458 45838
rect 47630 45890 47682 45902
rect 48738 45838 48750 45890
rect 48802 45838 48814 45890
rect 49634 45838 49646 45890
rect 49698 45838 49710 45890
rect 51762 45838 51774 45890
rect 51826 45838 51838 45890
rect 54338 45838 54350 45890
rect 54402 45838 54414 45890
rect 47630 45826 47682 45838
rect 2158 45778 2210 45790
rect 6414 45778 6466 45790
rect 5618 45726 5630 45778
rect 5682 45726 5694 45778
rect 2158 45714 2210 45726
rect 6414 45714 6466 45726
rect 6638 45778 6690 45790
rect 11902 45778 11954 45790
rect 7186 45726 7198 45778
rect 7250 45726 7262 45778
rect 6638 45714 6690 45726
rect 11902 45714 11954 45726
rect 14254 45778 14306 45790
rect 17838 45778 17890 45790
rect 16146 45726 16158 45778
rect 16210 45726 16222 45778
rect 17602 45726 17614 45778
rect 17666 45726 17678 45778
rect 14254 45714 14306 45726
rect 17838 45714 17890 45726
rect 18734 45778 18786 45790
rect 18734 45714 18786 45726
rect 21422 45778 21474 45790
rect 21422 45714 21474 45726
rect 21758 45778 21810 45790
rect 39790 45778 39842 45790
rect 23538 45726 23550 45778
rect 23602 45726 23614 45778
rect 29698 45726 29710 45778
rect 29762 45726 29774 45778
rect 35522 45726 35534 45778
rect 35586 45726 35598 45778
rect 36418 45726 36430 45778
rect 36482 45726 36494 45778
rect 21758 45714 21810 45726
rect 39790 45714 39842 45726
rect 40798 45778 40850 45790
rect 40798 45714 40850 45726
rect 43598 45778 43650 45790
rect 43598 45714 43650 45726
rect 44830 45778 44882 45790
rect 47518 45778 47570 45790
rect 52670 45778 52722 45790
rect 46162 45726 46174 45778
rect 46226 45726 46238 45778
rect 48850 45726 48862 45778
rect 48914 45726 48926 45778
rect 50978 45726 50990 45778
rect 51042 45726 51054 45778
rect 51538 45726 51550 45778
rect 51602 45726 51614 45778
rect 44830 45714 44882 45726
rect 47518 45714 47570 45726
rect 52670 45714 52722 45726
rect 52782 45778 52834 45790
rect 52782 45714 52834 45726
rect 5966 45666 6018 45678
rect 5966 45602 6018 45614
rect 9774 45666 9826 45678
rect 9774 45602 9826 45614
rect 12798 45666 12850 45678
rect 12798 45602 12850 45614
rect 19070 45666 19122 45678
rect 27022 45666 27074 45678
rect 25106 45614 25118 45666
rect 25170 45614 25182 45666
rect 26338 45614 26350 45666
rect 26402 45614 26414 45666
rect 19070 45602 19122 45614
rect 27022 45602 27074 45614
rect 27246 45666 27298 45678
rect 37102 45666 37154 45678
rect 40238 45666 40290 45678
rect 34626 45614 34638 45666
rect 34690 45614 34702 45666
rect 37426 45614 37438 45666
rect 37490 45614 37502 45666
rect 27246 45602 27298 45614
rect 37102 45602 37154 45614
rect 40238 45602 40290 45614
rect 40686 45666 40738 45678
rect 40686 45602 40738 45614
rect 41694 45666 41746 45678
rect 45054 45666 45106 45678
rect 43026 45614 43038 45666
rect 43090 45614 43102 45666
rect 41694 45602 41746 45614
rect 45054 45602 45106 45614
rect 45838 45666 45890 45678
rect 46946 45614 46958 45666
rect 47010 45614 47022 45666
rect 51314 45614 51326 45666
rect 51378 45614 51390 45666
rect 45838 45602 45890 45614
rect 1344 45498 58576 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 50558 45498
rect 50610 45446 50662 45498
rect 50714 45446 50766 45498
rect 50818 45446 58576 45498
rect 1344 45412 58576 45446
rect 2830 45330 2882 45342
rect 9774 45330 9826 45342
rect 4834 45278 4846 45330
rect 4898 45278 4910 45330
rect 2830 45266 2882 45278
rect 9774 45266 9826 45278
rect 16382 45330 16434 45342
rect 20078 45330 20130 45342
rect 26350 45330 26402 45342
rect 19506 45278 19518 45330
rect 19570 45278 19582 45330
rect 23650 45278 23662 45330
rect 23714 45278 23726 45330
rect 16382 45266 16434 45278
rect 20078 45266 20130 45278
rect 26350 45266 26402 45278
rect 26910 45330 26962 45342
rect 26910 45266 26962 45278
rect 27806 45330 27858 45342
rect 27806 45266 27858 45278
rect 32174 45330 32226 45342
rect 32174 45266 32226 45278
rect 38894 45330 38946 45342
rect 38894 45266 38946 45278
rect 45838 45330 45890 45342
rect 45838 45266 45890 45278
rect 47966 45330 48018 45342
rect 47966 45266 48018 45278
rect 48190 45330 48242 45342
rect 48190 45266 48242 45278
rect 48302 45330 48354 45342
rect 54798 45330 54850 45342
rect 52546 45278 52558 45330
rect 52610 45278 52622 45330
rect 48302 45266 48354 45278
rect 54798 45266 54850 45278
rect 16606 45218 16658 45230
rect 2034 45166 2046 45218
rect 2098 45166 2110 45218
rect 3938 45166 3950 45218
rect 4002 45166 4014 45218
rect 10770 45166 10782 45218
rect 10834 45166 10846 45218
rect 12562 45166 12574 45218
rect 12626 45166 12638 45218
rect 15586 45166 15598 45218
rect 15650 45166 15662 45218
rect 16606 45154 16658 45166
rect 16718 45218 16770 45230
rect 20414 45218 20466 45230
rect 17714 45166 17726 45218
rect 17778 45166 17790 45218
rect 16718 45154 16770 45166
rect 20414 45154 20466 45166
rect 26574 45218 26626 45230
rect 26574 45154 26626 45166
rect 27582 45218 27634 45230
rect 27582 45154 27634 45166
rect 32062 45218 32114 45230
rect 39118 45218 39170 45230
rect 34738 45166 34750 45218
rect 34802 45166 34814 45218
rect 36194 45166 36206 45218
rect 36258 45166 36270 45218
rect 38210 45166 38222 45218
rect 38274 45166 38286 45218
rect 32062 45154 32114 45166
rect 39118 45154 39170 45166
rect 45166 45218 45218 45230
rect 45166 45154 45218 45166
rect 47742 45218 47794 45230
rect 51650 45166 51662 45218
rect 51714 45166 51726 45218
rect 47742 45154 47794 45166
rect 2942 45106 2994 45118
rect 1810 45054 1822 45106
rect 1874 45054 1886 45106
rect 2942 45042 2994 45054
rect 3166 45106 3218 45118
rect 5294 45106 5346 45118
rect 19966 45106 20018 45118
rect 3378 45054 3390 45106
rect 3442 45054 3454 45106
rect 4050 45054 4062 45106
rect 4114 45054 4126 45106
rect 4722 45054 4734 45106
rect 4786 45054 4798 45106
rect 5506 45054 5518 45106
rect 5570 45054 5582 45106
rect 7186 45054 7198 45106
rect 7250 45054 7262 45106
rect 8530 45054 8542 45106
rect 8594 45054 8606 45106
rect 10994 45054 11006 45106
rect 11058 45054 11070 45106
rect 11330 45054 11342 45106
rect 11394 45054 11406 45106
rect 13570 45054 13582 45106
rect 13634 45054 13646 45106
rect 15922 45054 15934 45106
rect 15986 45054 15998 45106
rect 18946 45054 18958 45106
rect 19010 45054 19022 45106
rect 3166 45042 3218 45054
rect 5294 45042 5346 45054
rect 19966 45042 20018 45054
rect 20190 45106 20242 45118
rect 20190 45042 20242 45054
rect 23102 45106 23154 45118
rect 23102 45042 23154 45054
rect 23326 45106 23378 45118
rect 23326 45042 23378 45054
rect 26238 45106 26290 45118
rect 26238 45042 26290 45054
rect 26798 45106 26850 45118
rect 27470 45106 27522 45118
rect 27122 45054 27134 45106
rect 27186 45054 27198 45106
rect 26798 45042 26850 45054
rect 27470 45042 27522 45054
rect 33742 45106 33794 45118
rect 41694 45106 41746 45118
rect 44494 45106 44546 45118
rect 34850 45054 34862 45106
rect 34914 45054 34926 45106
rect 37426 45054 37438 45106
rect 37490 45054 37502 45106
rect 43698 45054 43710 45106
rect 43762 45054 43774 45106
rect 43922 45054 43934 45106
rect 43986 45054 43998 45106
rect 33742 45042 33794 45054
rect 41694 45042 41746 45054
rect 44494 45042 44546 45054
rect 44942 45106 44994 45118
rect 53006 45106 53058 45118
rect 49186 45054 49198 45106
rect 49250 45054 49262 45106
rect 49970 45054 49982 45106
rect 50034 45054 50046 45106
rect 51538 45054 51550 45106
rect 51602 45054 51614 45106
rect 52434 45054 52446 45106
rect 52498 45054 52510 45106
rect 44942 45042 44994 45054
rect 53006 45042 53058 45054
rect 53454 45106 53506 45118
rect 53454 45042 53506 45054
rect 53790 45106 53842 45118
rect 54574 45106 54626 45118
rect 54226 45054 54238 45106
rect 54290 45054 54302 45106
rect 53790 45042 53842 45054
rect 54574 45042 54626 45054
rect 3054 44994 3106 45006
rect 8990 44994 9042 45006
rect 33518 44994 33570 45006
rect 42254 44994 42306 45006
rect 45054 44994 45106 45006
rect 49086 44994 49138 45006
rect 7634 44942 7646 44994
rect 7698 44942 7710 44994
rect 9650 44942 9662 44994
rect 9714 44942 9726 44994
rect 10770 44942 10782 44994
rect 10834 44942 10846 44994
rect 12114 44942 12126 44994
rect 12178 44942 12190 44994
rect 17490 44942 17502 44994
rect 17554 44942 17566 44994
rect 33170 44942 33182 44994
rect 33234 44942 33246 44994
rect 34514 44942 34526 44994
rect 34578 44942 34590 44994
rect 35746 44942 35758 44994
rect 35810 44942 35822 44994
rect 43810 44942 43822 44994
rect 43874 44942 43886 44994
rect 46274 44942 46286 44994
rect 46338 44942 46350 44994
rect 3054 44930 3106 44942
rect 8990 44930 9042 44942
rect 33518 44930 33570 44942
rect 42254 44930 42306 44942
rect 45054 44930 45106 44942
rect 49086 44930 49138 44942
rect 54686 44994 54738 45006
rect 54686 44930 54738 44942
rect 9998 44882 10050 44894
rect 9998 44818 10050 44830
rect 14926 44882 14978 44894
rect 14926 44818 14978 44830
rect 15822 44882 15874 44894
rect 15822 44818 15874 44830
rect 32174 44882 32226 44894
rect 32174 44818 32226 44830
rect 38782 44882 38834 44894
rect 50094 44882 50146 44894
rect 44034 44830 44046 44882
rect 44098 44830 44110 44882
rect 38782 44818 38834 44830
rect 50094 44818 50146 44830
rect 1344 44714 58576 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 58576 44714
rect 1344 44628 58576 44662
rect 5630 44546 5682 44558
rect 21534 44546 21586 44558
rect 4834 44494 4846 44546
rect 4898 44494 4910 44546
rect 9986 44494 9998 44546
rect 10050 44494 10062 44546
rect 17378 44494 17390 44546
rect 17442 44494 17454 44546
rect 5630 44482 5682 44494
rect 21534 44482 21586 44494
rect 35758 44546 35810 44558
rect 35758 44482 35810 44494
rect 36206 44546 36258 44558
rect 36206 44482 36258 44494
rect 46734 44546 46786 44558
rect 46734 44482 46786 44494
rect 2382 44434 2434 44446
rect 7646 44434 7698 44446
rect 4274 44382 4286 44434
rect 4338 44382 4350 44434
rect 2382 44370 2434 44382
rect 7646 44370 7698 44382
rect 8878 44434 8930 44446
rect 12002 44382 12014 44434
rect 12066 44382 12078 44434
rect 14354 44382 14366 44434
rect 14418 44382 14430 44434
rect 17490 44382 17502 44434
rect 17554 44382 17566 44434
rect 23538 44382 23550 44434
rect 23602 44382 23614 44434
rect 34962 44382 34974 44434
rect 35026 44382 35038 44434
rect 35410 44382 35422 44434
rect 35474 44382 35486 44434
rect 40450 44382 40462 44434
rect 40514 44382 40526 44434
rect 44146 44382 44158 44434
rect 44210 44382 44222 44434
rect 45042 44382 45054 44434
rect 45106 44382 45118 44434
rect 47058 44382 47070 44434
rect 47122 44382 47134 44434
rect 47506 44382 47518 44434
rect 47570 44382 47582 44434
rect 8878 44370 8930 44382
rect 2606 44322 2658 44334
rect 6862 44322 6914 44334
rect 9550 44322 9602 44334
rect 19630 44322 19682 44334
rect 2930 44270 2942 44322
rect 2994 44270 3006 44322
rect 4610 44270 4622 44322
rect 4674 44270 4686 44322
rect 8418 44270 8430 44322
rect 8482 44270 8494 44322
rect 10882 44270 10894 44322
rect 10946 44270 10958 44322
rect 11778 44270 11790 44322
rect 11842 44270 11854 44322
rect 12338 44270 12350 44322
rect 12402 44270 12414 44322
rect 13794 44270 13806 44322
rect 13858 44270 13870 44322
rect 15810 44270 15822 44322
rect 15874 44270 15886 44322
rect 16818 44270 16830 44322
rect 16882 44270 16894 44322
rect 19394 44270 19406 44322
rect 19458 44270 19470 44322
rect 2606 44258 2658 44270
rect 6862 44258 6914 44270
rect 9550 44258 9602 44270
rect 19630 44258 19682 44270
rect 19854 44322 19906 44334
rect 19854 44258 19906 44270
rect 19966 44322 20018 44334
rect 21758 44322 21810 44334
rect 21298 44270 21310 44322
rect 21362 44270 21374 44322
rect 19966 44258 20018 44270
rect 21758 44258 21810 44270
rect 21870 44322 21922 44334
rect 36318 44322 36370 44334
rect 23090 44270 23102 44322
rect 23154 44270 23166 44322
rect 23874 44270 23886 44322
rect 23938 44270 23950 44322
rect 25778 44270 25790 44322
rect 25842 44270 25854 44322
rect 26786 44270 26798 44322
rect 26850 44270 26862 44322
rect 27682 44270 27694 44322
rect 27746 44270 27758 44322
rect 33394 44270 33406 44322
rect 33458 44270 33470 44322
rect 21870 44258 21922 44270
rect 36318 44258 36370 44270
rect 37326 44322 37378 44334
rect 50654 44322 50706 44334
rect 38658 44270 38670 44322
rect 38722 44270 38734 44322
rect 42130 44270 42142 44322
rect 42194 44270 42206 44322
rect 43698 44270 43710 44322
rect 43762 44270 43774 44322
rect 45154 44270 45166 44322
rect 45218 44270 45230 44322
rect 45490 44270 45502 44322
rect 45554 44270 45566 44322
rect 37326 44258 37378 44270
rect 50654 44258 50706 44270
rect 51662 44322 51714 44334
rect 51662 44258 51714 44270
rect 51774 44322 51826 44334
rect 54786 44270 54798 44322
rect 54850 44270 54862 44322
rect 55682 44270 55694 44322
rect 55746 44270 55758 44322
rect 51774 44258 51826 44270
rect 2718 44210 2770 44222
rect 2718 44146 2770 44158
rect 6302 44210 6354 44222
rect 6302 44146 6354 44158
rect 7198 44210 7250 44222
rect 7198 44146 7250 44158
rect 9326 44210 9378 44222
rect 9326 44146 9378 44158
rect 9438 44210 9490 44222
rect 26014 44210 26066 44222
rect 35534 44210 35586 44222
rect 23762 44158 23774 44210
rect 23826 44158 23838 44210
rect 28242 44158 28254 44210
rect 28306 44158 28318 44210
rect 32386 44158 32398 44210
rect 32450 44158 32462 44210
rect 34402 44158 34414 44210
rect 34466 44158 34478 44210
rect 9438 44146 9490 44158
rect 26014 44146 26066 44158
rect 35534 44146 35586 44158
rect 36206 44210 36258 44222
rect 36206 44146 36258 44158
rect 36990 44210 37042 44222
rect 46958 44210 47010 44222
rect 49646 44210 49698 44222
rect 38434 44158 38446 44210
rect 38498 44158 38510 44210
rect 39778 44158 39790 44210
rect 39842 44158 39854 44210
rect 40786 44158 40798 44210
rect 40850 44158 40862 44210
rect 42914 44158 42926 44210
rect 42978 44158 42990 44210
rect 44258 44158 44270 44210
rect 44322 44158 44334 44210
rect 47954 44158 47966 44210
rect 48018 44158 48030 44210
rect 49410 44158 49422 44210
rect 49474 44158 49486 44210
rect 36990 44146 37042 44158
rect 46958 44146 47010 44158
rect 49646 44146 49698 44158
rect 50766 44210 50818 44222
rect 50766 44146 50818 44158
rect 51886 44210 51938 44222
rect 53890 44158 53902 44210
rect 53954 44158 53966 44210
rect 55794 44158 55806 44210
rect 55858 44158 55870 44210
rect 51886 44146 51938 44158
rect 1710 44098 1762 44110
rect 3390 44098 3442 44110
rect 2034 44046 2046 44098
rect 2098 44046 2110 44098
rect 1710 44034 1762 44046
rect 3390 44034 3442 44046
rect 5742 44098 5794 44110
rect 5742 44034 5794 44046
rect 5854 44098 5906 44110
rect 7086 44098 7138 44110
rect 37102 44098 37154 44110
rect 50990 44098 51042 44110
rect 6626 44046 6638 44098
rect 6690 44046 6702 44098
rect 26562 44046 26574 44098
rect 26626 44046 26638 44098
rect 39666 44046 39678 44098
rect 39730 44046 39742 44098
rect 46050 44046 46062 44098
rect 46114 44046 46126 44098
rect 51202 44046 51214 44098
rect 51266 44046 51278 44098
rect 5854 44034 5906 44046
rect 7086 44034 7138 44046
rect 37102 44034 37154 44046
rect 50990 44034 51042 44046
rect 1344 43930 58576 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 50558 43930
rect 50610 43878 50662 43930
rect 50714 43878 50766 43930
rect 50818 43878 58576 43930
rect 1344 43844 58576 43878
rect 9550 43762 9602 43774
rect 3714 43710 3726 43762
rect 3778 43710 3790 43762
rect 9550 43698 9602 43710
rect 10782 43762 10834 43774
rect 20526 43762 20578 43774
rect 14018 43710 14030 43762
rect 14082 43710 14094 43762
rect 14802 43710 14814 43762
rect 14866 43710 14878 43762
rect 10782 43698 10834 43710
rect 20526 43698 20578 43710
rect 27918 43762 27970 43774
rect 27918 43698 27970 43710
rect 41694 43762 41746 43774
rect 41694 43698 41746 43710
rect 55246 43762 55298 43774
rect 55246 43698 55298 43710
rect 6078 43650 6130 43662
rect 4610 43598 4622 43650
rect 4674 43598 4686 43650
rect 6078 43586 6130 43598
rect 7534 43650 7586 43662
rect 16606 43650 16658 43662
rect 12562 43598 12574 43650
rect 12626 43598 12638 43650
rect 15586 43598 15598 43650
rect 15650 43598 15662 43650
rect 7534 43586 7586 43598
rect 16606 43586 16658 43598
rect 20078 43650 20130 43662
rect 25342 43650 25394 43662
rect 21634 43598 21646 43650
rect 21698 43598 21710 43650
rect 23874 43598 23886 43650
rect 23938 43598 23950 43650
rect 20078 43586 20130 43598
rect 25342 43586 25394 43598
rect 27246 43650 27298 43662
rect 27246 43586 27298 43598
rect 27470 43650 27522 43662
rect 27470 43586 27522 43598
rect 28814 43650 28866 43662
rect 28814 43586 28866 43598
rect 32174 43650 32226 43662
rect 32174 43586 32226 43598
rect 32286 43650 32338 43662
rect 32286 43586 32338 43598
rect 33070 43650 33122 43662
rect 34078 43650 34130 43662
rect 33394 43598 33406 43650
rect 33458 43598 33470 43650
rect 33070 43586 33122 43598
rect 34078 43586 34130 43598
rect 37326 43650 37378 43662
rect 37326 43586 37378 43598
rect 41134 43650 41186 43662
rect 41134 43586 41186 43598
rect 41470 43650 41522 43662
rect 46734 43650 46786 43662
rect 55022 43650 55074 43662
rect 42578 43598 42590 43650
rect 42642 43598 42654 43650
rect 51314 43598 51326 43650
rect 51378 43598 51390 43650
rect 41470 43586 41522 43598
rect 46734 43586 46786 43598
rect 55022 43586 55074 43598
rect 10110 43538 10162 43550
rect 20414 43538 20466 43550
rect 2706 43486 2718 43538
rect 2770 43486 2782 43538
rect 3490 43486 3502 43538
rect 3554 43486 3566 43538
rect 4050 43486 4062 43538
rect 4114 43486 4126 43538
rect 5058 43486 5070 43538
rect 5122 43486 5134 43538
rect 6850 43486 6862 43538
rect 6914 43486 6926 43538
rect 13458 43486 13470 43538
rect 13522 43486 13534 43538
rect 14578 43486 14590 43538
rect 14642 43486 14654 43538
rect 15698 43486 15710 43538
rect 15762 43486 15774 43538
rect 17938 43486 17950 43538
rect 18002 43486 18014 43538
rect 10110 43474 10162 43486
rect 20414 43474 20466 43486
rect 20750 43538 20802 43550
rect 25230 43538 25282 43550
rect 22530 43486 22542 43538
rect 22594 43486 22606 43538
rect 20750 43474 20802 43486
rect 25230 43474 25282 43486
rect 25566 43538 25618 43550
rect 25566 43474 25618 43486
rect 27134 43538 27186 43550
rect 27134 43474 27186 43486
rect 27582 43538 27634 43550
rect 27582 43474 27634 43486
rect 28030 43538 28082 43550
rect 28030 43474 28082 43486
rect 28254 43538 28306 43550
rect 31614 43538 31666 43550
rect 31378 43486 31390 43538
rect 31442 43486 31454 43538
rect 28254 43474 28306 43486
rect 31614 43474 31666 43486
rect 31950 43538 32002 43550
rect 54126 43538 54178 43550
rect 36194 43486 36206 43538
rect 36258 43486 36270 43538
rect 43922 43486 43934 43538
rect 43986 43486 43998 43538
rect 52434 43486 52446 43538
rect 52498 43486 52510 43538
rect 31950 43474 32002 43486
rect 54126 43474 54178 43486
rect 54350 43538 54402 43550
rect 54350 43474 54402 43486
rect 5518 43426 5570 43438
rect 2930 43374 2942 43426
rect 2994 43374 3006 43426
rect 5518 43362 5570 43374
rect 5854 43426 5906 43438
rect 5854 43362 5906 43374
rect 5966 43426 6018 43438
rect 8094 43426 8146 43438
rect 6738 43374 6750 43426
rect 6802 43374 6814 43426
rect 5966 43362 6018 43374
rect 8094 43362 8146 43374
rect 11342 43426 11394 43438
rect 11342 43362 11394 43374
rect 12126 43426 12178 43438
rect 12126 43362 12178 43374
rect 16270 43426 16322 43438
rect 18622 43426 18674 43438
rect 17714 43374 17726 43426
rect 17778 43374 17790 43426
rect 16270 43362 16322 43374
rect 18622 43362 18674 43374
rect 19182 43426 19234 43438
rect 19182 43362 19234 43374
rect 19406 43426 19458 43438
rect 19406 43362 19458 43374
rect 19742 43426 19794 43438
rect 26238 43426 26290 43438
rect 30718 43426 30770 43438
rect 36878 43426 36930 43438
rect 47294 43426 47346 43438
rect 21074 43374 21086 43426
rect 21138 43374 21150 43426
rect 28914 43374 28926 43426
rect 28978 43374 28990 43426
rect 36418 43374 36430 43426
rect 36482 43374 36494 43426
rect 41794 43374 41806 43426
rect 41858 43374 41870 43426
rect 42242 43374 42254 43426
rect 42306 43374 42318 43426
rect 50866 43374 50878 43426
rect 50930 43374 50942 43426
rect 53218 43374 53230 43426
rect 53282 43374 53294 43426
rect 19742 43362 19794 43374
rect 26238 43362 26290 43374
rect 30718 43362 30770 43374
rect 36878 43362 36930 43374
rect 47294 43362 47346 43374
rect 26350 43314 26402 43326
rect 3042 43262 3054 43314
rect 3106 43262 3118 43314
rect 26350 43250 26402 43262
rect 28590 43314 28642 43326
rect 28590 43250 28642 43262
rect 39678 43314 39730 43326
rect 39678 43250 39730 43262
rect 39790 43314 39842 43326
rect 39790 43250 39842 43262
rect 40014 43314 40066 43326
rect 40014 43250 40066 43262
rect 40126 43314 40178 43326
rect 45054 43314 45106 43326
rect 40898 43262 40910 43314
rect 40962 43311 40974 43314
rect 41122 43311 41134 43314
rect 40962 43265 41134 43311
rect 40962 43262 40974 43265
rect 41122 43262 41134 43265
rect 41186 43262 41198 43314
rect 40126 43250 40178 43262
rect 45054 43250 45106 43262
rect 48862 43314 48914 43326
rect 48862 43250 48914 43262
rect 48974 43314 49026 43326
rect 48974 43250 49026 43262
rect 49198 43314 49250 43326
rect 49198 43250 49250 43262
rect 49310 43314 49362 43326
rect 55358 43314 55410 43326
rect 54674 43262 54686 43314
rect 54738 43262 54750 43314
rect 49310 43250 49362 43262
rect 55358 43250 55410 43262
rect 1344 43146 58576 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 58576 43146
rect 1344 43060 58576 43094
rect 19406 42978 19458 42990
rect 43586 42926 43598 42978
rect 43650 42926 43662 42978
rect 46498 42926 46510 42978
rect 46562 42926 46574 42978
rect 54338 42926 54350 42978
rect 54402 42926 54414 42978
rect 19406 42914 19458 42926
rect 1934 42866 1986 42878
rect 19294 42866 19346 42878
rect 26798 42866 26850 42878
rect 5842 42814 5854 42866
rect 5906 42814 5918 42866
rect 12338 42814 12350 42866
rect 12402 42814 12414 42866
rect 15698 42814 15710 42866
rect 15762 42814 15774 42866
rect 23762 42814 23774 42866
rect 23826 42814 23838 42866
rect 1934 42802 1986 42814
rect 19294 42802 19346 42814
rect 26798 42802 26850 42814
rect 27246 42866 27298 42878
rect 48190 42866 48242 42878
rect 32162 42814 32174 42866
rect 32226 42814 32238 42866
rect 33730 42814 33742 42866
rect 33794 42814 33806 42866
rect 34514 42814 34526 42866
rect 34578 42814 34590 42866
rect 38994 42814 39006 42866
rect 39058 42814 39070 42866
rect 40562 42814 40574 42866
rect 40626 42814 40638 42866
rect 46162 42814 46174 42866
rect 46226 42814 46238 42866
rect 51202 42814 51214 42866
rect 51266 42814 51278 42866
rect 57138 42814 57150 42866
rect 57202 42814 57214 42866
rect 27246 42802 27298 42814
rect 48190 42802 48242 42814
rect 4622 42754 4674 42766
rect 11790 42754 11842 42766
rect 20862 42754 20914 42766
rect 4274 42702 4286 42754
rect 4338 42702 4350 42754
rect 7298 42702 7310 42754
rect 7362 42702 7374 42754
rect 9538 42702 9550 42754
rect 9602 42702 9614 42754
rect 11890 42702 11902 42754
rect 11954 42702 11966 42754
rect 13794 42702 13806 42754
rect 13858 42702 13870 42754
rect 14018 42702 14030 42754
rect 14082 42702 14094 42754
rect 14242 42702 14254 42754
rect 14306 42702 14318 42754
rect 4622 42690 4674 42702
rect 11790 42690 11842 42702
rect 20862 42690 20914 42702
rect 21870 42754 21922 42766
rect 26238 42754 26290 42766
rect 25330 42702 25342 42754
rect 25394 42702 25406 42754
rect 21870 42690 21922 42702
rect 26238 42690 26290 42702
rect 26910 42754 26962 42766
rect 26910 42690 26962 42702
rect 27470 42754 27522 42766
rect 36094 42754 36146 42766
rect 32386 42702 32398 42754
rect 32450 42702 32462 42754
rect 33506 42702 33518 42754
rect 33570 42702 33582 42754
rect 35074 42702 35086 42754
rect 35138 42702 35150 42754
rect 27470 42690 27522 42702
rect 36094 42690 36146 42702
rect 37102 42754 37154 42766
rect 37102 42690 37154 42702
rect 37886 42754 37938 42766
rect 44942 42754 44994 42766
rect 49870 42754 49922 42766
rect 51886 42754 51938 42766
rect 38882 42702 38894 42754
rect 38946 42702 38958 42754
rect 39778 42702 39790 42754
rect 39842 42702 39854 42754
rect 41346 42702 41358 42754
rect 41410 42702 41422 42754
rect 42354 42702 42366 42754
rect 42418 42702 42430 42754
rect 42690 42702 42702 42754
rect 42754 42702 42766 42754
rect 45378 42702 45390 42754
rect 45442 42702 45454 42754
rect 46386 42702 46398 42754
rect 46450 42702 46462 42754
rect 46834 42702 46846 42754
rect 46898 42702 46910 42754
rect 51426 42702 51438 42754
rect 51490 42702 51502 42754
rect 54114 42702 54126 42754
rect 54178 42702 54190 42754
rect 55234 42702 55246 42754
rect 55298 42702 55310 42754
rect 55682 42702 55694 42754
rect 55746 42702 55758 42754
rect 56690 42702 56702 42754
rect 56754 42702 56766 42754
rect 37886 42690 37938 42702
rect 44942 42690 44994 42702
rect 49870 42690 49922 42702
rect 51886 42690 51938 42702
rect 9326 42642 9378 42654
rect 17838 42642 17890 42654
rect 6290 42590 6302 42642
rect 6354 42590 6366 42642
rect 8530 42590 8542 42642
rect 8594 42590 8606 42642
rect 16258 42590 16270 42642
rect 16322 42590 16334 42642
rect 17602 42590 17614 42642
rect 17666 42590 17678 42642
rect 9326 42578 9378 42590
rect 17838 42578 17890 42590
rect 19182 42642 19234 42654
rect 19182 42578 19234 42590
rect 20526 42642 20578 42654
rect 20526 42578 20578 42590
rect 20638 42642 20690 42654
rect 20638 42578 20690 42590
rect 21310 42642 21362 42654
rect 21310 42578 21362 42590
rect 22094 42642 22146 42654
rect 22094 42578 22146 42590
rect 22206 42642 22258 42654
rect 30494 42642 30546 42654
rect 24210 42590 24222 42642
rect 24274 42590 24286 42642
rect 27794 42590 27806 42642
rect 27858 42590 27870 42642
rect 22206 42578 22258 42590
rect 30494 42578 30546 42590
rect 30606 42642 30658 42654
rect 30606 42578 30658 42590
rect 35758 42642 35810 42654
rect 35758 42578 35810 42590
rect 36990 42642 37042 42654
rect 36990 42578 37042 42590
rect 37774 42642 37826 42654
rect 48974 42642 49026 42654
rect 38322 42590 38334 42642
rect 38386 42590 38398 42642
rect 37774 42578 37826 42590
rect 48974 42578 49026 42590
rect 50318 42642 50370 42654
rect 50318 42578 50370 42590
rect 50654 42642 50706 42654
rect 50654 42578 50706 42590
rect 52670 42642 52722 42654
rect 52670 42578 52722 42590
rect 4958 42530 5010 42542
rect 4958 42466 5010 42478
rect 9774 42530 9826 42542
rect 9774 42466 9826 42478
rect 9886 42530 9938 42542
rect 9886 42466 9938 42478
rect 10110 42530 10162 42542
rect 12686 42530 12738 42542
rect 21646 42530 21698 42542
rect 10434 42478 10446 42530
rect 10498 42478 10510 42530
rect 14578 42478 14590 42530
rect 14642 42478 14654 42530
rect 10110 42466 10162 42478
rect 12686 42466 12738 42478
rect 21646 42466 21698 42478
rect 22654 42530 22706 42542
rect 26686 42530 26738 42542
rect 25778 42478 25790 42530
rect 25842 42478 25854 42530
rect 22654 42466 22706 42478
rect 26686 42466 26738 42478
rect 30830 42530 30882 42542
rect 30830 42466 30882 42478
rect 35982 42530 36034 42542
rect 35982 42466 36034 42478
rect 37550 42530 37602 42542
rect 37550 42466 37602 42478
rect 49870 42530 49922 42542
rect 49870 42466 49922 42478
rect 50430 42530 50482 42542
rect 52782 42530 52834 42542
rect 51650 42478 51662 42530
rect 51714 42478 51726 42530
rect 50430 42466 50482 42478
rect 52782 42466 52834 42478
rect 53006 42530 53058 42542
rect 53006 42466 53058 42478
rect 1344 42362 58576 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 50558 42362
rect 50610 42310 50662 42362
rect 50714 42310 50766 42362
rect 50818 42310 58576 42362
rect 1344 42276 58576 42310
rect 5294 42194 5346 42206
rect 5294 42130 5346 42142
rect 8654 42194 8706 42206
rect 16382 42194 16434 42206
rect 10546 42142 10558 42194
rect 10610 42142 10622 42194
rect 13346 42142 13358 42194
rect 13410 42142 13422 42194
rect 8654 42130 8706 42142
rect 16382 42130 16434 42142
rect 16606 42194 16658 42206
rect 16606 42130 16658 42142
rect 22878 42194 22930 42206
rect 22878 42130 22930 42142
rect 27134 42194 27186 42206
rect 27134 42130 27186 42142
rect 32174 42194 32226 42206
rect 32174 42130 32226 42142
rect 33854 42194 33906 42206
rect 36082 42142 36094 42194
rect 36146 42142 36158 42194
rect 36978 42142 36990 42194
rect 37042 42142 37054 42194
rect 40114 42142 40126 42194
rect 40178 42142 40190 42194
rect 43586 42142 43598 42194
rect 43650 42142 43662 42194
rect 33854 42130 33906 42142
rect 2494 42082 2546 42094
rect 2034 42030 2046 42082
rect 2098 42030 2110 42082
rect 2494 42018 2546 42030
rect 2606 42082 2658 42094
rect 8318 42082 8370 42094
rect 16718 42082 16770 42094
rect 31614 42082 31666 42094
rect 40910 42082 40962 42094
rect 6626 42030 6638 42082
rect 6690 42030 6702 42082
rect 9874 42030 9886 42082
rect 9938 42030 9950 42082
rect 11554 42030 11566 42082
rect 11618 42030 11630 42082
rect 18050 42030 18062 42082
rect 18114 42030 18126 42082
rect 34850 42030 34862 42082
rect 34914 42030 34926 42082
rect 36194 42030 36206 42082
rect 36258 42030 36270 42082
rect 37762 42030 37774 42082
rect 37826 42030 37838 42082
rect 39218 42030 39230 42082
rect 39282 42030 39294 42082
rect 2606 42018 2658 42030
rect 8318 42018 8370 42030
rect 16718 42018 16770 42030
rect 31614 42018 31666 42030
rect 40910 42018 40962 42030
rect 41022 42082 41074 42094
rect 42130 42030 42142 42082
rect 42194 42030 42206 42082
rect 43362 42030 43374 42082
rect 43426 42030 43438 42082
rect 47394 42030 47406 42082
rect 47458 42030 47470 42082
rect 49074 42030 49086 42082
rect 49138 42030 49150 42082
rect 54338 42030 54350 42082
rect 54402 42030 54414 42082
rect 41022 42018 41074 42030
rect 1710 41970 1762 41982
rect 4846 41970 4898 41982
rect 3602 41918 3614 41970
rect 3666 41918 3678 41970
rect 3938 41918 3950 41970
rect 4002 41918 4014 41970
rect 1710 41906 1762 41918
rect 4846 41906 4898 41918
rect 5406 41970 5458 41982
rect 5406 41906 5458 41918
rect 5518 41970 5570 41982
rect 13806 41970 13858 41982
rect 22094 41970 22146 41982
rect 6850 41918 6862 41970
rect 6914 41918 6926 41970
rect 7634 41918 7646 41970
rect 7698 41918 7710 41970
rect 8866 41918 8878 41970
rect 8930 41918 8942 41970
rect 9986 41918 9998 41970
rect 10050 41918 10062 41970
rect 10658 41918 10670 41970
rect 10722 41918 10734 41970
rect 12114 41918 12126 41970
rect 12178 41918 12190 41970
rect 12786 41918 12798 41970
rect 12850 41918 12862 41970
rect 14018 41918 14030 41970
rect 14082 41918 14094 41970
rect 14242 41918 14254 41970
rect 14306 41918 14318 41970
rect 15362 41918 15374 41970
rect 15426 41918 15438 41970
rect 18946 41918 18958 41970
rect 19010 41918 19022 41970
rect 5518 41906 5570 41918
rect 13806 41906 13858 41918
rect 22094 41906 22146 41918
rect 22206 41970 22258 41982
rect 22206 41906 22258 41918
rect 22542 41970 22594 41982
rect 24670 41970 24722 41982
rect 23090 41918 23102 41970
rect 23154 41918 23166 41970
rect 23314 41918 23326 41970
rect 23378 41918 23390 41970
rect 23986 41918 23998 41970
rect 24050 41918 24062 41970
rect 22542 41906 22594 41918
rect 24670 41906 24722 41918
rect 25790 41970 25842 41982
rect 31838 41970 31890 41982
rect 38558 41970 38610 41982
rect 26338 41918 26350 41970
rect 26402 41918 26414 41970
rect 28242 41918 28254 41970
rect 28306 41918 28318 41970
rect 29250 41918 29262 41970
rect 29314 41918 29326 41970
rect 36754 41918 36766 41970
rect 36818 41918 36830 41970
rect 37874 41918 37886 41970
rect 37938 41918 37950 41970
rect 38882 41918 38894 41970
rect 38946 41918 38958 41970
rect 39554 41918 39566 41970
rect 39618 41918 39630 41970
rect 40226 41918 40238 41970
rect 40290 41918 40302 41970
rect 44034 41918 44046 41970
rect 44098 41918 44110 41970
rect 44930 41918 44942 41970
rect 44994 41918 45006 41970
rect 45378 41918 45390 41970
rect 45442 41918 45454 41970
rect 47618 41918 47630 41970
rect 47682 41918 47694 41970
rect 48850 41918 48862 41970
rect 48914 41918 48926 41970
rect 49634 41918 49646 41970
rect 49698 41918 49710 41970
rect 51426 41918 51438 41970
rect 51490 41918 51502 41970
rect 52434 41918 52446 41970
rect 52498 41918 52510 41970
rect 54226 41918 54238 41970
rect 54290 41918 54302 41970
rect 25790 41906 25842 41918
rect 31838 41906 31890 41918
rect 38558 41906 38610 41918
rect 19630 41858 19682 41870
rect 4610 41806 4622 41858
rect 4674 41806 4686 41858
rect 15474 41806 15486 41858
rect 15538 41806 15550 41858
rect 17490 41806 17502 41858
rect 17554 41806 17566 41858
rect 19630 41794 19682 41806
rect 22430 41858 22482 41870
rect 25678 41858 25730 41870
rect 33294 41858 33346 41870
rect 41694 41858 41746 41870
rect 23874 41806 23886 41858
rect 23938 41806 23950 41858
rect 29138 41806 29150 41858
rect 29202 41806 29214 41858
rect 34290 41806 34302 41858
rect 34354 41806 34366 41858
rect 46162 41806 46174 41858
rect 46226 41806 46238 41858
rect 47394 41806 47406 41858
rect 47458 41806 47470 41858
rect 49522 41806 49534 41858
rect 49586 41806 49598 41858
rect 52882 41806 52894 41858
rect 52946 41806 52958 41858
rect 54898 41806 54910 41858
rect 54962 41806 54974 41858
rect 22430 41794 22482 41806
rect 25678 41794 25730 41806
rect 33294 41794 33346 41806
rect 41694 41794 41746 41806
rect 2494 41746 2546 41758
rect 23214 41746 23266 41758
rect 38894 41746 38946 41758
rect 15586 41694 15598 41746
rect 15650 41694 15662 41746
rect 27570 41694 27582 41746
rect 27634 41694 27646 41746
rect 2494 41682 2546 41694
rect 23214 41682 23266 41694
rect 38894 41682 38946 41694
rect 41022 41746 41074 41758
rect 50418 41694 50430 41746
rect 50482 41694 50494 41746
rect 41022 41682 41074 41694
rect 1344 41578 58576 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 58576 41578
rect 1344 41492 58576 41526
rect 14142 41410 14194 41422
rect 8306 41358 8318 41410
rect 8370 41407 8382 41410
rect 8866 41407 8878 41410
rect 8370 41361 8878 41407
rect 8370 41358 8382 41361
rect 8866 41358 8878 41361
rect 8930 41358 8942 41410
rect 14142 41346 14194 41358
rect 23662 41410 23714 41422
rect 23662 41346 23714 41358
rect 44046 41410 44098 41422
rect 44046 41346 44098 41358
rect 1934 41298 1986 41310
rect 8094 41298 8146 41310
rect 7186 41246 7198 41298
rect 7250 41246 7262 41298
rect 1934 41234 1986 41246
rect 8094 41234 8146 41246
rect 12350 41298 12402 41310
rect 20078 41298 20130 41310
rect 16706 41246 16718 41298
rect 16770 41246 16782 41298
rect 12350 41234 12402 41246
rect 20078 41234 20130 41246
rect 21534 41298 21586 41310
rect 21534 41234 21586 41246
rect 26014 41298 26066 41310
rect 26014 41234 26066 41246
rect 32174 41298 32226 41310
rect 34078 41298 34130 41310
rect 33394 41246 33406 41298
rect 33458 41246 33470 41298
rect 35858 41246 35870 41298
rect 35922 41246 35934 41298
rect 36306 41246 36318 41298
rect 36370 41246 36382 41298
rect 32174 41234 32226 41246
rect 34078 41234 34130 41246
rect 9550 41186 9602 41198
rect 4274 41134 4286 41186
rect 4338 41134 4350 41186
rect 4722 41134 4734 41186
rect 4786 41134 4798 41186
rect 5842 41134 5854 41186
rect 5906 41134 5918 41186
rect 6178 41134 6190 41186
rect 6242 41134 6254 41186
rect 7410 41134 7422 41186
rect 7474 41134 7486 41186
rect 9314 41134 9326 41186
rect 9378 41134 9390 41186
rect 9550 41122 9602 41134
rect 9662 41186 9714 41198
rect 17614 41186 17666 41198
rect 18734 41186 18786 41198
rect 21758 41186 21810 41198
rect 31950 41186 32002 41198
rect 34750 41186 34802 41198
rect 44942 41186 44994 41198
rect 10098 41134 10110 41186
rect 10162 41134 10174 41186
rect 10882 41134 10894 41186
rect 10946 41134 10958 41186
rect 11554 41134 11566 41186
rect 11618 41134 11630 41186
rect 11778 41134 11790 41186
rect 11842 41134 11854 41186
rect 14242 41134 14254 41186
rect 14306 41134 14318 41186
rect 14578 41134 14590 41186
rect 14642 41134 14654 41186
rect 15922 41134 15934 41186
rect 15986 41134 15998 41186
rect 17938 41134 17950 41186
rect 18002 41134 18014 41186
rect 18498 41134 18510 41186
rect 18562 41134 18574 41186
rect 19618 41134 19630 41186
rect 19682 41134 19694 41186
rect 22530 41134 22542 41186
rect 22594 41134 22606 41186
rect 22754 41134 22766 41186
rect 22818 41134 22830 41186
rect 23426 41134 23438 41186
rect 23490 41134 23502 41186
rect 32274 41134 32286 41186
rect 32338 41134 32350 41186
rect 33282 41134 33294 41186
rect 33346 41134 33358 41186
rect 35410 41134 35422 41186
rect 35474 41134 35486 41186
rect 36530 41134 36542 41186
rect 36594 41134 36606 41186
rect 38098 41134 38110 41186
rect 38162 41134 38174 41186
rect 39218 41134 39230 41186
rect 39282 41134 39294 41186
rect 41458 41134 41470 41186
rect 41522 41134 41534 41186
rect 42578 41134 42590 41186
rect 42642 41134 42654 41186
rect 45378 41134 45390 41186
rect 45442 41134 45454 41186
rect 47506 41134 47518 41186
rect 47570 41134 47582 41186
rect 48626 41134 48638 41186
rect 48690 41134 48702 41186
rect 50418 41134 50430 41186
rect 50482 41134 50494 41186
rect 51202 41134 51214 41186
rect 51266 41134 51278 41186
rect 51650 41134 51662 41186
rect 51714 41134 51726 41186
rect 54226 41134 54238 41186
rect 54290 41134 54302 41186
rect 55234 41134 55246 41186
rect 55298 41134 55310 41186
rect 9662 41122 9714 41134
rect 17614 41122 17666 41134
rect 18734 41122 18786 41134
rect 21758 41122 21810 41134
rect 31950 41122 32002 41134
rect 34750 41122 34802 41134
rect 44942 41122 44994 41134
rect 8542 41074 8594 41086
rect 12238 41074 12290 41086
rect 6738 41022 6750 41074
rect 6802 41022 6814 41074
rect 11666 41022 11678 41074
rect 11730 41022 11742 41074
rect 8542 41010 8594 41022
rect 12238 41010 12290 41022
rect 12462 41074 12514 41086
rect 18846 41074 18898 41086
rect 19966 41074 20018 41086
rect 13906 41022 13918 41074
rect 13970 41022 13982 41074
rect 16482 41022 16494 41074
rect 16546 41022 16558 41074
rect 19282 41022 19294 41074
rect 19346 41022 19358 41074
rect 12462 41010 12514 41022
rect 18846 41010 18898 41022
rect 19966 41010 20018 41022
rect 25118 41074 25170 41086
rect 25118 41010 25170 41022
rect 25566 41074 25618 41086
rect 25566 41010 25618 41022
rect 25678 41074 25730 41086
rect 25678 41010 25730 41022
rect 25902 41074 25954 41086
rect 25902 41010 25954 41022
rect 26238 41074 26290 41086
rect 26238 41010 26290 41022
rect 26462 41074 26514 41086
rect 26462 41010 26514 41022
rect 26798 41074 26850 41086
rect 26798 41010 26850 41022
rect 26910 41074 26962 41086
rect 26910 41010 26962 41022
rect 29486 41074 29538 41086
rect 29486 41010 29538 41022
rect 31166 41074 31218 41086
rect 31166 41010 31218 41022
rect 34638 41074 34690 41086
rect 44158 41074 44210 41086
rect 37314 41022 37326 41074
rect 37378 41022 37390 41074
rect 39330 41022 39342 41074
rect 39394 41022 39406 41074
rect 41010 41022 41022 41074
rect 41074 41022 41086 41074
rect 43474 41022 43486 41074
rect 43538 41022 43550 41074
rect 34638 41010 34690 41022
rect 44158 41010 44210 41022
rect 44830 41074 44882 41086
rect 47394 41022 47406 41074
rect 47458 41022 47470 41074
rect 53106 41022 53118 41074
rect 53170 41022 53182 41074
rect 55458 41022 55470 41074
rect 55522 41022 55534 41074
rect 44830 41010 44882 41022
rect 4958 40962 5010 40974
rect 8990 40962 9042 40974
rect 5730 40910 5742 40962
rect 5794 40910 5806 40962
rect 4958 40898 5010 40910
rect 8990 40898 9042 40910
rect 18174 40962 18226 40974
rect 18174 40898 18226 40910
rect 18286 40962 18338 40974
rect 18286 40898 18338 40910
rect 20190 40962 20242 40974
rect 25342 40962 25394 40974
rect 22082 40910 22094 40962
rect 22146 40910 22158 40962
rect 20190 40898 20242 40910
rect 25342 40898 25394 40910
rect 27134 40962 27186 40974
rect 27134 40898 27186 40910
rect 29150 40962 29202 40974
rect 29150 40898 29202 40910
rect 30830 40962 30882 40974
rect 30830 40898 30882 40910
rect 31838 40962 31890 40974
rect 31838 40898 31890 40910
rect 32510 40962 32562 40974
rect 32510 40898 32562 40910
rect 34414 40962 34466 40974
rect 34414 40898 34466 40910
rect 44046 40962 44098 40974
rect 51998 40962 52050 40974
rect 48738 40910 48750 40962
rect 48802 40910 48814 40962
rect 44046 40898 44098 40910
rect 51998 40898 52050 40910
rect 1344 40794 58576 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 50558 40794
rect 50610 40742 50662 40794
rect 50714 40742 50766 40794
rect 50818 40742 58576 40794
rect 1344 40708 58576 40742
rect 6078 40626 6130 40638
rect 5170 40574 5182 40626
rect 5234 40574 5246 40626
rect 6078 40562 6130 40574
rect 6862 40626 6914 40638
rect 6862 40562 6914 40574
rect 7198 40626 7250 40638
rect 7198 40562 7250 40574
rect 7422 40626 7474 40638
rect 11118 40626 11170 40638
rect 8530 40574 8542 40626
rect 8594 40574 8606 40626
rect 7422 40562 7474 40574
rect 11118 40562 11170 40574
rect 19518 40626 19570 40638
rect 19518 40562 19570 40574
rect 20526 40626 20578 40638
rect 25902 40626 25954 40638
rect 21858 40574 21870 40626
rect 21922 40574 21934 40626
rect 20526 40562 20578 40574
rect 25902 40562 25954 40574
rect 33406 40626 33458 40638
rect 33406 40562 33458 40574
rect 35310 40626 35362 40638
rect 35310 40562 35362 40574
rect 35422 40626 35474 40638
rect 35422 40562 35474 40574
rect 40910 40626 40962 40638
rect 40910 40562 40962 40574
rect 47630 40626 47682 40638
rect 50642 40574 50654 40626
rect 50706 40574 50718 40626
rect 47630 40562 47682 40574
rect 5854 40514 5906 40526
rect 5854 40450 5906 40462
rect 6302 40514 6354 40526
rect 6302 40450 6354 40462
rect 9102 40514 9154 40526
rect 18622 40514 18674 40526
rect 12002 40462 12014 40514
rect 12066 40462 12078 40514
rect 14578 40462 14590 40514
rect 14642 40462 14654 40514
rect 9102 40450 9154 40462
rect 18622 40450 18674 40462
rect 19070 40514 19122 40526
rect 19070 40450 19122 40462
rect 19294 40514 19346 40526
rect 19294 40450 19346 40462
rect 20414 40514 20466 40526
rect 25678 40514 25730 40526
rect 33854 40514 33906 40526
rect 22642 40462 22654 40514
rect 22706 40462 22718 40514
rect 27122 40462 27134 40514
rect 27186 40462 27198 40514
rect 30370 40462 30382 40514
rect 30434 40462 30446 40514
rect 35634 40462 35646 40514
rect 35698 40511 35710 40514
rect 35858 40511 35870 40514
rect 35698 40465 35870 40511
rect 35698 40462 35710 40465
rect 35858 40462 35870 40465
rect 35922 40462 35934 40514
rect 42466 40462 42478 40514
rect 42530 40462 42542 40514
rect 43026 40462 43038 40514
rect 43090 40462 43102 40514
rect 44034 40462 44046 40514
rect 44098 40462 44110 40514
rect 49186 40462 49198 40514
rect 49250 40462 49262 40514
rect 50754 40462 50766 40514
rect 50818 40462 50830 40514
rect 20414 40450 20466 40462
rect 25678 40450 25730 40462
rect 33854 40450 33906 40462
rect 5518 40402 5570 40414
rect 4274 40350 4286 40402
rect 4338 40350 4350 40402
rect 5518 40338 5570 40350
rect 6414 40402 6466 40414
rect 6414 40338 6466 40350
rect 6638 40402 6690 40414
rect 6638 40338 6690 40350
rect 6974 40402 7026 40414
rect 6974 40338 7026 40350
rect 7534 40402 7586 40414
rect 10558 40402 10610 40414
rect 16158 40402 16210 40414
rect 8306 40350 8318 40402
rect 8370 40350 8382 40402
rect 12338 40350 12350 40402
rect 12402 40350 12414 40402
rect 13234 40350 13246 40402
rect 13298 40350 13310 40402
rect 15586 40350 15598 40402
rect 15650 40350 15662 40402
rect 7534 40338 7586 40350
rect 10558 40338 10610 40350
rect 16158 40338 16210 40350
rect 18510 40402 18562 40414
rect 18510 40338 18562 40350
rect 18846 40402 18898 40414
rect 18846 40338 18898 40350
rect 19742 40402 19794 40414
rect 19742 40338 19794 40350
rect 19854 40402 19906 40414
rect 21310 40402 21362 40414
rect 24446 40402 24498 40414
rect 20178 40350 20190 40402
rect 20242 40350 20254 40402
rect 22866 40350 22878 40402
rect 22930 40350 22942 40402
rect 23762 40350 23774 40402
rect 23826 40350 23838 40402
rect 19854 40338 19906 40350
rect 21310 40338 21362 40350
rect 24446 40338 24498 40350
rect 25566 40402 25618 40414
rect 25566 40338 25618 40350
rect 26014 40402 26066 40414
rect 33294 40402 33346 40414
rect 26338 40350 26350 40402
rect 26402 40350 26414 40402
rect 29586 40350 29598 40402
rect 29650 40350 29662 40402
rect 26014 40338 26066 40350
rect 33294 40338 33346 40350
rect 34078 40402 34130 40414
rect 34078 40338 34130 40350
rect 35534 40402 35586 40414
rect 41470 40402 41522 40414
rect 37202 40350 37214 40402
rect 37266 40350 37278 40402
rect 38322 40350 38334 40402
rect 38386 40350 38398 40402
rect 38882 40350 38894 40402
rect 38946 40350 38958 40402
rect 35534 40338 35586 40350
rect 41470 40338 41522 40350
rect 43262 40402 43314 40414
rect 43262 40338 43314 40350
rect 43374 40402 43426 40414
rect 48190 40402 48242 40414
rect 54014 40402 54066 40414
rect 43586 40350 43598 40402
rect 43650 40350 43662 40402
rect 45378 40350 45390 40402
rect 45442 40350 45454 40402
rect 46946 40350 46958 40402
rect 47010 40350 47022 40402
rect 51538 40350 51550 40402
rect 51602 40350 51614 40402
rect 51762 40350 51774 40402
rect 51826 40350 51838 40402
rect 53218 40350 53230 40402
rect 53282 40350 53294 40402
rect 43374 40338 43426 40350
rect 48190 40338 48242 40350
rect 54014 40338 54066 40350
rect 54238 40402 54290 40414
rect 54674 40350 54686 40402
rect 54738 40350 54750 40402
rect 54238 40338 54290 40350
rect 4622 40290 4674 40302
rect 4622 40226 4674 40238
rect 4846 40290 4898 40302
rect 4846 40226 4898 40238
rect 16270 40290 16322 40302
rect 34414 40290 34466 40302
rect 46286 40290 46338 40302
rect 48974 40290 49026 40302
rect 29250 40238 29262 40290
rect 29314 40238 29326 40290
rect 32498 40238 32510 40290
rect 32562 40238 32574 40290
rect 36306 40238 36318 40290
rect 36370 40238 36382 40290
rect 38546 40238 38558 40290
rect 38610 40238 38622 40290
rect 39666 40238 39678 40290
rect 39730 40238 39742 40290
rect 45154 40238 45166 40290
rect 45218 40238 45230 40290
rect 47170 40238 47182 40290
rect 47234 40238 47246 40290
rect 16270 40226 16322 40238
rect 34414 40226 34466 40238
rect 46286 40226 46338 40238
rect 48974 40226 49026 40238
rect 51326 40290 51378 40302
rect 53678 40290 53730 40302
rect 53330 40238 53342 40290
rect 53394 40238 53406 40290
rect 51326 40226 51378 40238
rect 53678 40226 53730 40238
rect 1934 40178 1986 40190
rect 1934 40114 1986 40126
rect 21534 40178 21586 40190
rect 21534 40114 21586 40126
rect 33406 40178 33458 40190
rect 33406 40114 33458 40126
rect 1344 40010 58576 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 58576 40010
rect 1344 39924 58576 39958
rect 4286 39842 4338 39854
rect 2930 39790 2942 39842
rect 2994 39790 3006 39842
rect 4286 39778 4338 39790
rect 4622 39842 4674 39854
rect 24110 39842 24162 39854
rect 19506 39790 19518 39842
rect 19570 39790 19582 39842
rect 4622 39778 4674 39790
rect 24110 39778 24162 39790
rect 29822 39842 29874 39854
rect 29822 39778 29874 39790
rect 30158 39842 30210 39854
rect 30158 39778 30210 39790
rect 31614 39842 31666 39854
rect 31614 39778 31666 39790
rect 31950 39842 32002 39854
rect 31950 39778 32002 39790
rect 37662 39842 37714 39854
rect 37662 39778 37714 39790
rect 39790 39842 39842 39854
rect 39790 39778 39842 39790
rect 40126 39842 40178 39854
rect 40126 39778 40178 39790
rect 48302 39842 48354 39854
rect 48302 39778 48354 39790
rect 11118 39730 11170 39742
rect 2818 39678 2830 39730
rect 2882 39678 2894 39730
rect 11118 39666 11170 39678
rect 13694 39730 13746 39742
rect 13694 39666 13746 39678
rect 15486 39730 15538 39742
rect 15486 39666 15538 39678
rect 28702 39730 28754 39742
rect 38222 39730 38274 39742
rect 35858 39678 35870 39730
rect 35922 39678 35934 39730
rect 28702 39666 28754 39678
rect 38222 39666 38274 39678
rect 40574 39730 40626 39742
rect 49086 39730 49138 39742
rect 55134 39730 55186 39742
rect 44034 39678 44046 39730
rect 44098 39678 44110 39730
rect 51090 39678 51102 39730
rect 51154 39678 51166 39730
rect 40574 39666 40626 39678
rect 49086 39666 49138 39678
rect 55134 39666 55186 39678
rect 4062 39618 4114 39630
rect 9102 39618 9154 39630
rect 10894 39618 10946 39630
rect 1810 39566 1822 39618
rect 1874 39566 1886 39618
rect 3042 39566 3054 39618
rect 3106 39566 3118 39618
rect 3826 39566 3838 39618
rect 3890 39566 3902 39618
rect 6626 39566 6638 39618
rect 6690 39566 6702 39618
rect 7410 39566 7422 39618
rect 7474 39566 7486 39618
rect 8754 39566 8766 39618
rect 8818 39566 8830 39618
rect 10098 39566 10110 39618
rect 10162 39566 10174 39618
rect 4062 39554 4114 39566
rect 9102 39554 9154 39566
rect 10894 39554 10946 39566
rect 11342 39618 11394 39630
rect 11342 39554 11394 39566
rect 11454 39618 11506 39630
rect 17502 39618 17554 39630
rect 16818 39566 16830 39618
rect 16882 39566 16894 39618
rect 11454 39554 11506 39566
rect 17502 39554 17554 39566
rect 18958 39618 19010 39630
rect 18958 39554 19010 39566
rect 19182 39618 19234 39630
rect 19182 39554 19234 39566
rect 23998 39618 24050 39630
rect 33854 39618 33906 39630
rect 37774 39618 37826 39630
rect 24994 39566 25006 39618
rect 25058 39566 25070 39618
rect 27010 39566 27022 39618
rect 27074 39566 27086 39618
rect 30818 39566 30830 39618
rect 30882 39566 30894 39618
rect 32722 39566 32734 39618
rect 32786 39566 32798 39618
rect 34178 39566 34190 39618
rect 34242 39566 34254 39618
rect 35522 39566 35534 39618
rect 35586 39566 35598 39618
rect 23998 39554 24050 39566
rect 33854 39554 33906 39566
rect 37774 39554 37826 39566
rect 39454 39618 39506 39630
rect 47854 39618 47906 39630
rect 40898 39566 40910 39618
rect 40962 39566 40974 39618
rect 42130 39566 42142 39618
rect 42194 39566 42206 39618
rect 42802 39566 42814 39618
rect 42866 39566 42878 39618
rect 43586 39566 43598 39618
rect 43650 39566 43662 39618
rect 45938 39566 45950 39618
rect 46002 39566 46014 39618
rect 46610 39566 46622 39618
rect 46674 39566 46686 39618
rect 39454 39554 39506 39566
rect 47854 39554 47906 39566
rect 48078 39618 48130 39630
rect 48078 39554 48130 39566
rect 48862 39618 48914 39630
rect 48862 39554 48914 39566
rect 49310 39618 49362 39630
rect 49310 39554 49362 39566
rect 49422 39618 49474 39630
rect 49422 39554 49474 39566
rect 49982 39618 50034 39630
rect 49982 39554 50034 39566
rect 50206 39618 50258 39630
rect 50206 39554 50258 39566
rect 51550 39618 51602 39630
rect 51550 39554 51602 39566
rect 52222 39618 52274 39630
rect 52222 39554 52274 39566
rect 52670 39618 52722 39630
rect 55358 39618 55410 39630
rect 54114 39566 54126 39618
rect 54178 39566 54190 39618
rect 54562 39566 54574 39618
rect 54626 39566 54638 39618
rect 52670 39554 52722 39566
rect 55358 39554 55410 39566
rect 8094 39506 8146 39518
rect 6402 39454 6414 39506
rect 6466 39454 6478 39506
rect 8094 39442 8146 39454
rect 8542 39506 8594 39518
rect 17838 39506 17890 39518
rect 15810 39454 15822 39506
rect 15874 39454 15886 39506
rect 8542 39442 8594 39454
rect 17838 39442 17890 39454
rect 18174 39506 18226 39518
rect 18174 39442 18226 39454
rect 19854 39506 19906 39518
rect 19854 39442 19906 39454
rect 20190 39506 20242 39518
rect 20190 39442 20242 39454
rect 21646 39506 21698 39518
rect 21646 39442 21698 39454
rect 25566 39506 25618 39518
rect 36430 39506 36482 39518
rect 25778 39454 25790 39506
rect 25842 39454 25854 39506
rect 27122 39454 27134 39506
rect 27186 39454 27198 39506
rect 30930 39454 30942 39506
rect 30994 39454 31006 39506
rect 32498 39454 32510 39506
rect 32562 39454 32574 39506
rect 25566 39442 25618 39454
rect 36430 39442 36482 39454
rect 37102 39506 37154 39518
rect 37102 39442 37154 39454
rect 37214 39506 37266 39518
rect 37214 39442 37266 39454
rect 39902 39506 39954 39518
rect 51886 39506 51938 39518
rect 43698 39454 43710 39506
rect 43762 39454 43774 39506
rect 46834 39454 46846 39506
rect 46898 39454 46910 39506
rect 39902 39442 39954 39454
rect 51886 39442 51938 39454
rect 51998 39506 52050 39518
rect 54798 39506 54850 39518
rect 52994 39454 53006 39506
rect 53058 39454 53070 39506
rect 51998 39442 52050 39454
rect 54798 39442 54850 39454
rect 2046 39394 2098 39406
rect 2046 39330 2098 39342
rect 5182 39394 5234 39406
rect 5182 39330 5234 39342
rect 8990 39394 9042 39406
rect 8990 39330 9042 39342
rect 9438 39394 9490 39406
rect 9438 39330 9490 39342
rect 10446 39394 10498 39406
rect 10446 39330 10498 39342
rect 10558 39394 10610 39406
rect 10558 39330 10610 39342
rect 10670 39394 10722 39406
rect 10670 39330 10722 39342
rect 14926 39394 14978 39406
rect 14926 39330 14978 39342
rect 21310 39394 21362 39406
rect 21310 39330 21362 39342
rect 23774 39394 23826 39406
rect 23774 39330 23826 39342
rect 24110 39394 24162 39406
rect 24110 39330 24162 39342
rect 25230 39394 25282 39406
rect 25230 39330 25282 39342
rect 29486 39394 29538 39406
rect 29486 39330 29538 39342
rect 33294 39394 33346 39406
rect 33294 39330 33346 39342
rect 34414 39394 34466 39406
rect 34414 39330 34466 39342
rect 34526 39394 34578 39406
rect 34526 39330 34578 39342
rect 36878 39394 36930 39406
rect 36878 39330 36930 39342
rect 37662 39394 37714 39406
rect 48750 39394 48802 39406
rect 39106 39342 39118 39394
rect 39170 39342 39182 39394
rect 42690 39342 42702 39394
rect 42754 39342 42766 39394
rect 45378 39342 45390 39394
rect 45442 39342 45454 39394
rect 50530 39342 50542 39394
rect 50594 39342 50606 39394
rect 55682 39342 55694 39394
rect 55746 39342 55758 39394
rect 37662 39330 37714 39342
rect 48750 39330 48802 39342
rect 1344 39226 58576 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 50558 39226
rect 50610 39174 50662 39226
rect 50714 39174 50766 39226
rect 50818 39174 58576 39226
rect 1344 39140 58576 39174
rect 4174 39058 4226 39070
rect 4174 38994 4226 39006
rect 12126 39058 12178 39070
rect 12126 38994 12178 39006
rect 16046 39058 16098 39070
rect 16046 38994 16098 39006
rect 16270 39058 16322 39070
rect 16270 38994 16322 39006
rect 16942 39058 16994 39070
rect 16942 38994 16994 39006
rect 17390 39058 17442 39070
rect 17390 38994 17442 39006
rect 26014 39058 26066 39070
rect 26014 38994 26066 39006
rect 31166 39058 31218 39070
rect 31166 38994 31218 39006
rect 45614 39058 45666 39070
rect 45614 38994 45666 39006
rect 45838 39058 45890 39070
rect 45838 38994 45890 39006
rect 48862 39058 48914 39070
rect 48862 38994 48914 39006
rect 49086 39058 49138 39070
rect 49086 38994 49138 39006
rect 52446 39058 52498 39070
rect 52446 38994 52498 39006
rect 52782 39058 52834 39070
rect 52782 38994 52834 39006
rect 53566 39058 53618 39070
rect 53566 38994 53618 39006
rect 4734 38946 4786 38958
rect 11230 38946 11282 38958
rect 6290 38894 6302 38946
rect 6354 38894 6366 38946
rect 8306 38894 8318 38946
rect 8370 38894 8382 38946
rect 4734 38882 4786 38894
rect 11230 38882 11282 38894
rect 15934 38946 15986 38958
rect 15934 38882 15986 38894
rect 16382 38946 16434 38958
rect 18062 38946 18114 38958
rect 17714 38894 17726 38946
rect 17778 38894 17790 38946
rect 16382 38882 16434 38894
rect 18062 38882 18114 38894
rect 18174 38946 18226 38958
rect 18174 38882 18226 38894
rect 23998 38946 24050 38958
rect 23998 38882 24050 38894
rect 24222 38946 24274 38958
rect 24222 38882 24274 38894
rect 24334 38946 24386 38958
rect 24334 38882 24386 38894
rect 25342 38946 25394 38958
rect 25342 38882 25394 38894
rect 33294 38946 33346 38958
rect 33294 38882 33346 38894
rect 37102 38946 37154 38958
rect 37102 38882 37154 38894
rect 41918 38946 41970 38958
rect 45502 38946 45554 38958
rect 44482 38894 44494 38946
rect 44546 38894 44558 38946
rect 41918 38882 41970 38894
rect 45502 38882 45554 38894
rect 47742 38946 47794 38958
rect 49634 38894 49646 38946
rect 49698 38894 49710 38946
rect 50866 38894 50878 38946
rect 50930 38894 50942 38946
rect 51090 38894 51102 38946
rect 51154 38894 51166 38946
rect 53106 38894 53118 38946
rect 53170 38894 53182 38946
rect 54450 38894 54462 38946
rect 54514 38894 54526 38946
rect 47742 38882 47794 38894
rect 3838 38834 3890 38846
rect 2594 38782 2606 38834
rect 2658 38782 2670 38834
rect 3838 38770 3890 38782
rect 4622 38834 4674 38846
rect 10446 38834 10498 38846
rect 19966 38834 20018 38846
rect 7298 38782 7310 38834
rect 7362 38782 7374 38834
rect 10658 38782 10670 38834
rect 10722 38782 10734 38834
rect 13794 38782 13806 38834
rect 13858 38782 13870 38834
rect 15362 38782 15374 38834
rect 15426 38782 15438 38834
rect 19394 38782 19406 38834
rect 19458 38782 19470 38834
rect 4622 38770 4674 38782
rect 10446 38770 10498 38782
rect 19966 38770 20018 38782
rect 20414 38834 20466 38846
rect 20414 38770 20466 38782
rect 20638 38834 20690 38846
rect 20638 38770 20690 38782
rect 21534 38834 21586 38846
rect 21534 38770 21586 38782
rect 22430 38834 22482 38846
rect 22430 38770 22482 38782
rect 24558 38834 24610 38846
rect 36878 38834 36930 38846
rect 38558 38834 38610 38846
rect 41806 38834 41858 38846
rect 46286 38834 46338 38846
rect 33506 38782 33518 38834
rect 33570 38782 33582 38834
rect 37650 38782 37662 38834
rect 37714 38782 37726 38834
rect 41234 38782 41246 38834
rect 41298 38782 41310 38834
rect 43586 38782 43598 38834
rect 43650 38782 43662 38834
rect 44370 38782 44382 38834
rect 44434 38782 44446 38834
rect 24558 38770 24610 38782
rect 36878 38770 36930 38782
rect 38558 38770 38610 38782
rect 41806 38770 41858 38782
rect 46286 38770 46338 38782
rect 46398 38834 46450 38846
rect 48750 38834 48802 38846
rect 53454 38834 53506 38846
rect 46834 38782 46846 38834
rect 46898 38782 46910 38834
rect 49298 38782 49310 38834
rect 49362 38782 49374 38834
rect 51314 38782 51326 38834
rect 51378 38782 51390 38834
rect 46398 38770 46450 38782
rect 48750 38770 48802 38782
rect 53454 38770 53506 38782
rect 53790 38834 53842 38846
rect 54786 38782 54798 38834
rect 54850 38782 54862 38834
rect 55458 38782 55470 38834
rect 55522 38782 55534 38834
rect 53790 38770 53842 38782
rect 3054 38722 3106 38734
rect 2482 38670 2494 38722
rect 2546 38670 2558 38722
rect 3054 38658 3106 38670
rect 5406 38722 5458 38734
rect 14030 38722 14082 38734
rect 21310 38722 21362 38734
rect 5730 38670 5742 38722
rect 5794 38670 5806 38722
rect 19170 38670 19182 38722
rect 19234 38670 19246 38722
rect 20962 38670 20974 38722
rect 21026 38670 21038 38722
rect 5406 38658 5458 38670
rect 14030 38658 14082 38670
rect 21310 38658 21362 38670
rect 22206 38722 22258 38734
rect 22206 38658 22258 38670
rect 34078 38722 34130 38734
rect 34078 38658 34130 38670
rect 35982 38722 36034 38734
rect 35982 38658 36034 38670
rect 36542 38722 36594 38734
rect 47966 38722 48018 38734
rect 50206 38722 50258 38734
rect 37762 38670 37774 38722
rect 37826 38670 37838 38722
rect 42578 38670 42590 38722
rect 42642 38670 42654 38722
rect 49858 38670 49870 38722
rect 49922 38670 49934 38722
rect 36542 38658 36594 38670
rect 47966 38658 48018 38670
rect 50206 38658 50258 38670
rect 51886 38722 51938 38734
rect 54674 38670 54686 38722
rect 54738 38670 54750 38722
rect 51886 38658 51938 38670
rect 4510 38610 4562 38622
rect 4510 38546 4562 38558
rect 14254 38610 14306 38622
rect 14254 38546 14306 38558
rect 14366 38610 14418 38622
rect 14366 38546 14418 38558
rect 15038 38610 15090 38622
rect 15038 38546 15090 38558
rect 15374 38610 15426 38622
rect 15374 38546 15426 38558
rect 18174 38610 18226 38622
rect 18174 38546 18226 38558
rect 21870 38610 21922 38622
rect 47630 38610 47682 38622
rect 22754 38558 22766 38610
rect 22818 38558 22830 38610
rect 21870 38546 21922 38558
rect 47630 38546 47682 38558
rect 1344 38442 58576 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 58576 38442
rect 1344 38356 58576 38390
rect 6526 38274 6578 38286
rect 25902 38274 25954 38286
rect 43710 38274 43762 38286
rect 2706 38222 2718 38274
rect 2770 38222 2782 38274
rect 25106 38222 25118 38274
rect 25170 38222 25182 38274
rect 41682 38222 41694 38274
rect 41746 38222 41758 38274
rect 55570 38222 55582 38274
rect 55634 38222 55646 38274
rect 6526 38210 6578 38222
rect 25902 38210 25954 38222
rect 43710 38210 43762 38222
rect 8766 38162 8818 38174
rect 2930 38110 2942 38162
rect 2994 38110 3006 38162
rect 8766 38098 8818 38110
rect 13582 38162 13634 38174
rect 22206 38162 22258 38174
rect 14242 38110 14254 38162
rect 14306 38110 14318 38162
rect 15586 38110 15598 38162
rect 15650 38110 15662 38162
rect 17378 38110 17390 38162
rect 17442 38110 17454 38162
rect 13582 38098 13634 38110
rect 22206 38098 22258 38110
rect 26574 38162 26626 38174
rect 26574 38098 26626 38110
rect 28142 38162 28194 38174
rect 33058 38110 33070 38162
rect 33122 38110 33134 38162
rect 35298 38110 35310 38162
rect 35362 38110 35374 38162
rect 40338 38110 40350 38162
rect 40402 38110 40414 38162
rect 44034 38110 44046 38162
rect 44098 38110 44110 38162
rect 48178 38110 48190 38162
rect 48242 38110 48254 38162
rect 28142 38098 28194 38110
rect 4734 38050 4786 38062
rect 7870 38050 7922 38062
rect 9326 38050 9378 38062
rect 19742 38050 19794 38062
rect 24558 38050 24610 38062
rect 3042 37998 3054 38050
rect 3106 37998 3118 38050
rect 4386 37998 4398 38050
rect 4450 37998 4462 38050
rect 5730 37998 5742 38050
rect 5794 37998 5806 38050
rect 6290 37998 6302 38050
rect 6354 37998 6366 38050
rect 7074 37998 7086 38050
rect 7138 37998 7150 38050
rect 8306 37998 8318 38050
rect 8370 37998 8382 38050
rect 11330 37998 11342 38050
rect 11394 37998 11406 38050
rect 12226 37998 12238 38050
rect 12290 37998 12302 38050
rect 15250 37998 15262 38050
rect 15314 37998 15326 38050
rect 15922 37998 15934 38050
rect 15986 37998 15998 38050
rect 17042 37998 17054 38050
rect 17106 37998 17118 38050
rect 18722 37998 18734 38050
rect 18786 37998 18798 38050
rect 21410 37998 21422 38050
rect 21474 37998 21486 38050
rect 23538 37998 23550 38050
rect 23602 37998 23614 38050
rect 4734 37986 4786 37998
rect 7870 37986 7922 37998
rect 9326 37986 9378 37998
rect 19742 37986 19794 37998
rect 24558 37986 24610 37998
rect 24782 38050 24834 38062
rect 25678 38050 25730 38062
rect 36094 38050 36146 38062
rect 25442 37998 25454 38050
rect 25506 37998 25518 38050
rect 32386 37998 32398 38050
rect 32450 37998 32462 38050
rect 24782 37986 24834 37998
rect 25678 37986 25730 37998
rect 36094 37986 36146 37998
rect 36430 38050 36482 38062
rect 36430 37986 36482 37998
rect 36990 38050 37042 38062
rect 36990 37986 37042 37998
rect 37214 38050 37266 38062
rect 37214 37986 37266 37998
rect 37438 38050 37490 38062
rect 37438 37986 37490 37998
rect 37886 38050 37938 38062
rect 46398 38050 46450 38062
rect 40226 37998 40238 38050
rect 40290 37998 40302 38050
rect 41570 37998 41582 38050
rect 41634 37998 41646 38050
rect 45378 37998 45390 38050
rect 45442 37998 45454 38050
rect 37886 37986 37938 37998
rect 46398 37986 46450 37998
rect 46846 38050 46898 38062
rect 46846 37986 46898 37998
rect 47182 38050 47234 38062
rect 54462 38050 54514 38062
rect 47954 37998 47966 38050
rect 48018 37998 48030 38050
rect 48738 37998 48750 38050
rect 48802 37998 48814 38050
rect 50194 37998 50206 38050
rect 50258 37998 50270 38050
rect 51986 37998 51998 38050
rect 52050 37998 52062 38050
rect 53778 37998 53790 38050
rect 53842 37998 53854 38050
rect 55122 37998 55134 38050
rect 55186 37998 55198 38050
rect 47182 37986 47234 37998
rect 54462 37986 54514 37998
rect 4846 37938 4898 37950
rect 4846 37874 4898 37886
rect 9214 37938 9266 37950
rect 9214 37874 9266 37886
rect 9438 37938 9490 37950
rect 19070 37938 19122 37950
rect 21646 37938 21698 37950
rect 24222 37938 24274 37950
rect 11218 37886 11230 37938
rect 11282 37886 11294 37938
rect 20066 37886 20078 37938
rect 20130 37886 20142 37938
rect 22530 37886 22542 37938
rect 22594 37886 22606 37938
rect 9438 37874 9490 37886
rect 19070 37874 19122 37886
rect 21646 37874 21698 37886
rect 24222 37874 24274 37886
rect 26014 37938 26066 37950
rect 26014 37874 26066 37886
rect 29822 37938 29874 37950
rect 29822 37874 29874 37886
rect 43934 37938 43986 37950
rect 48290 37886 48302 37938
rect 48354 37886 48366 37938
rect 50082 37886 50094 37938
rect 50146 37886 50158 37938
rect 43934 37874 43986 37886
rect 1822 37826 1874 37838
rect 18958 37826 19010 37838
rect 9874 37774 9886 37826
rect 9938 37774 9950 37826
rect 12786 37774 12798 37826
rect 12850 37774 12862 37826
rect 1822 37762 1874 37774
rect 18958 37762 19010 37774
rect 29934 37826 29986 37838
rect 29934 37762 29986 37774
rect 30158 37826 30210 37838
rect 30158 37762 30210 37774
rect 30494 37826 30546 37838
rect 30494 37762 30546 37774
rect 35870 37826 35922 37838
rect 35870 37762 35922 37774
rect 36318 37826 36370 37838
rect 36318 37762 36370 37774
rect 37102 37826 37154 37838
rect 51886 37826 51938 37838
rect 38210 37774 38222 37826
rect 38274 37774 38286 37826
rect 45602 37774 45614 37826
rect 45666 37774 45678 37826
rect 37102 37762 37154 37774
rect 51886 37762 51938 37774
rect 1344 37658 58576 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 50558 37658
rect 50610 37606 50662 37658
rect 50714 37606 50766 37658
rect 50818 37606 58576 37658
rect 1344 37572 58576 37606
rect 5518 37490 5570 37502
rect 5518 37426 5570 37438
rect 9550 37490 9602 37502
rect 10782 37490 10834 37502
rect 27806 37490 27858 37502
rect 9874 37438 9886 37490
rect 9938 37438 9950 37490
rect 13458 37438 13470 37490
rect 13522 37438 13534 37490
rect 9550 37426 9602 37438
rect 10782 37426 10834 37438
rect 27806 37426 27858 37438
rect 31614 37490 31666 37502
rect 31614 37426 31666 37438
rect 33518 37490 33570 37502
rect 33518 37426 33570 37438
rect 33966 37490 34018 37502
rect 33966 37426 34018 37438
rect 35646 37490 35698 37502
rect 35646 37426 35698 37438
rect 37550 37490 37602 37502
rect 40338 37438 40350 37490
rect 40402 37438 40414 37490
rect 37550 37426 37602 37438
rect 4734 37378 4786 37390
rect 4734 37314 4786 37326
rect 4846 37378 4898 37390
rect 4846 37314 4898 37326
rect 5182 37378 5234 37390
rect 19966 37378 20018 37390
rect 6626 37326 6638 37378
rect 6690 37326 6702 37378
rect 12002 37326 12014 37378
rect 12066 37326 12078 37378
rect 14018 37326 14030 37378
rect 14082 37326 14094 37378
rect 14578 37326 14590 37378
rect 14642 37326 14654 37378
rect 15698 37326 15710 37378
rect 15762 37326 15774 37378
rect 18050 37326 18062 37378
rect 18114 37326 18126 37378
rect 5182 37314 5234 37326
rect 19966 37314 20018 37326
rect 20078 37378 20130 37390
rect 20078 37314 20130 37326
rect 21422 37378 21474 37390
rect 24446 37378 24498 37390
rect 22530 37326 22542 37378
rect 22594 37326 22606 37378
rect 21422 37314 21474 37326
rect 24446 37314 24498 37326
rect 26350 37378 26402 37390
rect 26350 37314 26402 37326
rect 26798 37378 26850 37390
rect 26798 37314 26850 37326
rect 27918 37378 27970 37390
rect 38558 37378 38610 37390
rect 34514 37326 34526 37378
rect 34578 37326 34590 37378
rect 34850 37326 34862 37378
rect 34914 37326 34926 37378
rect 27918 37314 27970 37326
rect 38558 37314 38610 37326
rect 46846 37378 46898 37390
rect 46846 37314 46898 37326
rect 47630 37378 47682 37390
rect 47630 37314 47682 37326
rect 55470 37378 55522 37390
rect 57810 37326 57822 37378
rect 57874 37326 57886 37378
rect 55470 37314 55522 37326
rect 5518 37266 5570 37278
rect 4162 37214 4174 37266
rect 4226 37214 4238 37266
rect 5518 37202 5570 37214
rect 5742 37266 5794 37278
rect 10894 37266 10946 37278
rect 21534 37266 21586 37278
rect 23886 37266 23938 37278
rect 6850 37214 6862 37266
rect 6914 37214 6926 37266
rect 7858 37214 7870 37266
rect 7922 37214 7934 37266
rect 12898 37214 12910 37266
rect 12962 37214 12974 37266
rect 13906 37214 13918 37266
rect 13970 37214 13982 37266
rect 15138 37214 15150 37266
rect 15202 37214 15214 37266
rect 15586 37214 15598 37266
rect 15650 37214 15662 37266
rect 19058 37214 19070 37266
rect 19122 37214 19134 37266
rect 21186 37214 21198 37266
rect 21250 37214 21262 37266
rect 22418 37214 22430 37266
rect 22482 37214 22494 37266
rect 23314 37214 23326 37266
rect 23378 37214 23390 37266
rect 5742 37202 5794 37214
rect 10894 37202 10946 37214
rect 21534 37202 21586 37214
rect 23886 37202 23938 37214
rect 24110 37266 24162 37278
rect 24110 37202 24162 37214
rect 25902 37266 25954 37278
rect 25902 37202 25954 37214
rect 26014 37266 26066 37278
rect 26014 37202 26066 37214
rect 26686 37266 26738 37278
rect 26686 37202 26738 37214
rect 26910 37266 26962 37278
rect 26910 37202 26962 37214
rect 27358 37266 27410 37278
rect 27358 37202 27410 37214
rect 27582 37266 27634 37278
rect 34302 37266 34354 37278
rect 28354 37214 28366 37266
rect 28418 37214 28430 37266
rect 27582 37202 27634 37214
rect 34302 37202 34354 37214
rect 37214 37266 37266 37278
rect 37214 37202 37266 37214
rect 37438 37266 37490 37278
rect 37438 37202 37490 37214
rect 37774 37266 37826 37278
rect 37774 37202 37826 37214
rect 38110 37266 38162 37278
rect 38110 37202 38162 37214
rect 38334 37266 38386 37278
rect 38334 37202 38386 37214
rect 39118 37266 39170 37278
rect 46734 37266 46786 37278
rect 42578 37214 42590 37266
rect 42642 37214 42654 37266
rect 43474 37214 43486 37266
rect 43538 37214 43550 37266
rect 44258 37214 44270 37266
rect 44322 37214 44334 37266
rect 44930 37214 44942 37266
rect 44994 37214 45006 37266
rect 39118 37202 39170 37214
rect 46734 37202 46786 37214
rect 47518 37266 47570 37278
rect 47518 37202 47570 37214
rect 48078 37266 48130 37278
rect 54798 37266 54850 37278
rect 50082 37214 50094 37266
rect 50146 37214 50158 37266
rect 50754 37214 50766 37266
rect 50818 37214 50830 37266
rect 52658 37214 52670 37266
rect 52722 37214 52734 37266
rect 54450 37214 54462 37266
rect 54514 37214 54526 37266
rect 48078 37202 48130 37214
rect 54798 37202 54850 37214
rect 55246 37266 55298 37278
rect 55246 37202 55298 37214
rect 58158 37266 58210 37278
rect 58158 37202 58210 37214
rect 19630 37154 19682 37166
rect 24334 37154 24386 37166
rect 11442 37102 11454 37154
rect 11506 37102 11518 37154
rect 15474 37102 15486 37154
rect 15538 37102 15550 37154
rect 17490 37102 17502 37154
rect 17554 37102 17566 37154
rect 22642 37102 22654 37154
rect 22706 37102 22718 37154
rect 19630 37090 19682 37102
rect 24334 37090 24386 37102
rect 25342 37154 25394 37166
rect 25342 37090 25394 37102
rect 26238 37154 26290 37166
rect 38446 37154 38498 37166
rect 29026 37102 29038 37154
rect 29090 37102 29102 37154
rect 31154 37102 31166 37154
rect 31218 37102 31230 37154
rect 26238 37090 26290 37102
rect 38446 37090 38498 37102
rect 38894 37154 38946 37166
rect 38894 37090 38946 37102
rect 39790 37154 39842 37166
rect 46174 37154 46226 37166
rect 42690 37102 42702 37154
rect 42754 37102 42766 37154
rect 43586 37102 43598 37154
rect 43650 37102 43662 37154
rect 39790 37090 39842 37102
rect 46174 37090 46226 37102
rect 47294 37154 47346 37166
rect 53902 37154 53954 37166
rect 48962 37102 48974 37154
rect 49026 37102 49038 37154
rect 52210 37102 52222 37154
rect 52274 37102 52286 37154
rect 47294 37090 47346 37102
rect 53902 37090 53954 37102
rect 55358 37154 55410 37166
rect 55358 37090 55410 37102
rect 56030 37154 56082 37166
rect 56030 37090 56082 37102
rect 57598 37154 57650 37166
rect 57598 37090 57650 37102
rect 1934 37042 1986 37054
rect 1934 36978 1986 36990
rect 4734 37042 4786 37054
rect 4734 36978 4786 36990
rect 8990 37042 9042 37054
rect 8990 36978 9042 36990
rect 11006 37042 11058 37054
rect 11006 36978 11058 36990
rect 20078 37042 20130 37054
rect 39454 37042 39506 37054
rect 21970 36990 21982 37042
rect 22034 36990 22046 37042
rect 20078 36978 20130 36990
rect 39454 36978 39506 36990
rect 40014 37042 40066 37054
rect 40014 36978 40066 36990
rect 46846 37042 46898 37054
rect 46846 36978 46898 36990
rect 48302 37042 48354 37054
rect 50306 36990 50318 37042
rect 50370 36990 50382 37042
rect 48302 36978 48354 36990
rect 1344 36874 58576 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 58576 36874
rect 1344 36788 58576 36822
rect 2606 36706 2658 36718
rect 2258 36654 2270 36706
rect 2322 36654 2334 36706
rect 2606 36642 2658 36654
rect 6750 36706 6802 36718
rect 6750 36642 6802 36654
rect 7086 36706 7138 36718
rect 7086 36642 7138 36654
rect 10334 36706 10386 36718
rect 11118 36706 11170 36718
rect 10770 36654 10782 36706
rect 10834 36654 10846 36706
rect 10334 36642 10386 36654
rect 11118 36642 11170 36654
rect 18510 36706 18562 36718
rect 18510 36642 18562 36654
rect 18622 36706 18674 36718
rect 18622 36642 18674 36654
rect 18958 36706 19010 36718
rect 18958 36642 19010 36654
rect 22766 36706 22818 36718
rect 22766 36642 22818 36654
rect 23102 36706 23154 36718
rect 23102 36642 23154 36654
rect 24782 36706 24834 36718
rect 24782 36642 24834 36654
rect 25118 36706 25170 36718
rect 25118 36642 25170 36654
rect 38110 36706 38162 36718
rect 38110 36642 38162 36654
rect 40574 36706 40626 36718
rect 40574 36642 40626 36654
rect 43486 36706 43538 36718
rect 53006 36706 53058 36718
rect 52658 36654 52670 36706
rect 52722 36654 52734 36706
rect 43486 36642 43538 36654
rect 53006 36642 53058 36654
rect 2830 36594 2882 36606
rect 6526 36594 6578 36606
rect 3266 36542 3278 36594
rect 3330 36542 3342 36594
rect 2830 36530 2882 36542
rect 6526 36530 6578 36542
rect 12910 36594 12962 36606
rect 12910 36530 12962 36542
rect 14366 36594 14418 36606
rect 14366 36530 14418 36542
rect 14702 36594 14754 36606
rect 14702 36530 14754 36542
rect 17166 36594 17218 36606
rect 17166 36530 17218 36542
rect 18734 36594 18786 36606
rect 29262 36594 29314 36606
rect 34414 36594 34466 36606
rect 19954 36542 19966 36594
rect 20018 36542 20030 36594
rect 26450 36542 26462 36594
rect 26514 36542 26526 36594
rect 28578 36542 28590 36594
rect 28642 36542 28654 36594
rect 33842 36542 33854 36594
rect 33906 36542 33918 36594
rect 18734 36530 18786 36542
rect 29262 36530 29314 36542
rect 34414 36530 34466 36542
rect 39902 36594 39954 36606
rect 39902 36530 39954 36542
rect 40462 36594 40514 36606
rect 44046 36594 44098 36606
rect 41682 36542 41694 36594
rect 41746 36542 41758 36594
rect 40462 36530 40514 36542
rect 44046 36530 44098 36542
rect 54126 36594 54178 36606
rect 54126 36530 54178 36542
rect 57934 36594 57986 36606
rect 57934 36530 57986 36542
rect 6190 36482 6242 36494
rect 3714 36430 3726 36482
rect 3778 36430 3790 36482
rect 4274 36430 4286 36482
rect 4338 36430 4350 36482
rect 6190 36418 6242 36430
rect 7422 36482 7474 36494
rect 7422 36418 7474 36430
rect 10222 36482 10274 36494
rect 10222 36418 10274 36430
rect 11342 36482 11394 36494
rect 11342 36418 11394 36430
rect 11678 36482 11730 36494
rect 11678 36418 11730 36430
rect 12350 36482 12402 36494
rect 12350 36418 12402 36430
rect 13806 36482 13858 36494
rect 18174 36482 18226 36494
rect 15138 36430 15150 36482
rect 15202 36430 15214 36482
rect 15586 36430 15598 36482
rect 15650 36430 15662 36482
rect 17938 36430 17950 36482
rect 18002 36430 18014 36482
rect 13806 36418 13858 36430
rect 18174 36418 18226 36430
rect 19182 36482 19234 36494
rect 20750 36482 20802 36494
rect 19842 36430 19854 36482
rect 19906 36430 19918 36482
rect 19182 36418 19234 36430
rect 20750 36418 20802 36430
rect 21310 36482 21362 36494
rect 21310 36418 21362 36430
rect 22990 36482 23042 36494
rect 29822 36482 29874 36494
rect 38222 36482 38274 36494
rect 45614 36482 45666 36494
rect 51214 36482 51266 36494
rect 53230 36482 53282 36494
rect 25666 36430 25678 36482
rect 25730 36430 25742 36482
rect 30930 36430 30942 36482
rect 30994 36430 31006 36482
rect 37314 36430 37326 36482
rect 37378 36430 37390 36482
rect 40226 36430 40238 36482
rect 40290 36430 40302 36482
rect 41346 36430 41358 36482
rect 41410 36430 41422 36482
rect 43026 36430 43038 36482
rect 43090 36430 43102 36482
rect 47282 36430 47294 36482
rect 47346 36430 47358 36482
rect 48402 36430 48414 36482
rect 48466 36430 48478 36482
rect 50530 36430 50542 36482
rect 50594 36430 50606 36482
rect 51538 36430 51550 36482
rect 51602 36430 51614 36482
rect 54226 36430 54238 36482
rect 54290 36430 54302 36482
rect 55234 36430 55246 36482
rect 55298 36430 55310 36482
rect 55570 36430 55582 36482
rect 55634 36430 55646 36482
rect 22990 36418 23042 36430
rect 29822 36418 29874 36430
rect 38222 36418 38274 36430
rect 45614 36418 45666 36430
rect 51214 36418 51266 36430
rect 53230 36418 53282 36430
rect 1710 36370 1762 36382
rect 1710 36306 1762 36318
rect 2046 36370 2098 36382
rect 4622 36370 4674 36382
rect 3602 36318 3614 36370
rect 3666 36318 3678 36370
rect 2046 36306 2098 36318
rect 4622 36306 4674 36318
rect 7646 36370 7698 36382
rect 7646 36306 7698 36318
rect 7758 36370 7810 36382
rect 25006 36370 25058 36382
rect 40910 36370 40962 36382
rect 49758 36370 49810 36382
rect 15810 36318 15822 36370
rect 15874 36318 15886 36370
rect 16146 36318 16158 36370
rect 16210 36318 16222 36370
rect 31602 36318 31614 36370
rect 31666 36318 31678 36370
rect 43362 36318 43374 36370
rect 43426 36318 43438 36370
rect 45938 36318 45950 36370
rect 46002 36318 46014 36370
rect 46834 36318 46846 36370
rect 46898 36318 46910 36370
rect 49074 36318 49086 36370
rect 49138 36318 49150 36370
rect 54114 36318 54126 36370
rect 54178 36318 54190 36370
rect 7758 36306 7810 36318
rect 25006 36306 25058 36318
rect 40910 36306 40962 36318
rect 49758 36306 49810 36318
rect 1822 36258 1874 36270
rect 1822 36194 1874 36206
rect 4734 36258 4786 36270
rect 4734 36194 4786 36206
rect 4846 36258 4898 36270
rect 4846 36194 4898 36206
rect 5630 36258 5682 36270
rect 5630 36194 5682 36206
rect 8206 36258 8258 36270
rect 8206 36194 8258 36206
rect 10334 36258 10386 36270
rect 10334 36194 10386 36206
rect 11790 36258 11842 36270
rect 11790 36194 11842 36206
rect 12014 36258 12066 36270
rect 23102 36258 23154 36270
rect 16370 36206 16382 36258
rect 16434 36206 16446 36258
rect 21634 36206 21646 36258
rect 21698 36206 21710 36258
rect 12014 36194 12066 36206
rect 23102 36194 23154 36206
rect 23774 36258 23826 36270
rect 23774 36194 23826 36206
rect 29150 36258 29202 36270
rect 29150 36194 29202 36206
rect 29374 36258 29426 36270
rect 29374 36194 29426 36206
rect 34862 36258 34914 36270
rect 34862 36194 34914 36206
rect 37550 36258 37602 36270
rect 37550 36194 37602 36206
rect 38110 36258 38162 36270
rect 38110 36194 38162 36206
rect 38670 36258 38722 36270
rect 38670 36194 38722 36206
rect 1344 36090 58576 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 50558 36090
rect 50610 36038 50662 36090
rect 50714 36038 50766 36090
rect 50818 36038 58576 36090
rect 1344 36004 58576 36038
rect 2606 35922 2658 35934
rect 2606 35858 2658 35870
rect 2718 35922 2770 35934
rect 5294 35922 5346 35934
rect 4946 35870 4958 35922
rect 5010 35870 5022 35922
rect 2718 35858 2770 35870
rect 5294 35858 5346 35870
rect 7310 35922 7362 35934
rect 12686 35922 12738 35934
rect 10882 35870 10894 35922
rect 10946 35870 10958 35922
rect 7310 35858 7362 35870
rect 12686 35858 12738 35870
rect 13022 35922 13074 35934
rect 13022 35858 13074 35870
rect 13582 35922 13634 35934
rect 13582 35858 13634 35870
rect 27358 35922 27410 35934
rect 27358 35858 27410 35870
rect 28142 35922 28194 35934
rect 28142 35858 28194 35870
rect 28926 35922 28978 35934
rect 28926 35858 28978 35870
rect 32174 35922 32226 35934
rect 32174 35858 32226 35870
rect 32398 35922 32450 35934
rect 32398 35858 32450 35870
rect 32958 35922 33010 35934
rect 32958 35858 33010 35870
rect 33182 35922 33234 35934
rect 33182 35858 33234 35870
rect 39678 35922 39730 35934
rect 39678 35858 39730 35870
rect 40014 35922 40066 35934
rect 40014 35858 40066 35870
rect 2382 35810 2434 35822
rect 2034 35758 2046 35810
rect 2098 35758 2110 35810
rect 2382 35746 2434 35758
rect 2942 35810 2994 35822
rect 2942 35746 2994 35758
rect 6862 35810 6914 35822
rect 17390 35810 17442 35822
rect 14466 35758 14478 35810
rect 14530 35758 14542 35810
rect 6862 35746 6914 35758
rect 17390 35746 17442 35758
rect 17614 35810 17666 35822
rect 17614 35746 17666 35758
rect 18958 35810 19010 35822
rect 18958 35746 19010 35758
rect 19182 35810 19234 35822
rect 19182 35746 19234 35758
rect 23662 35810 23714 35822
rect 23662 35746 23714 35758
rect 27694 35810 27746 35822
rect 27694 35746 27746 35758
rect 38222 35810 38274 35822
rect 50206 35810 50258 35822
rect 57822 35810 57874 35822
rect 44034 35758 44046 35810
rect 44098 35758 44110 35810
rect 45266 35758 45278 35810
rect 45330 35758 45342 35810
rect 49858 35758 49870 35810
rect 49922 35758 49934 35810
rect 50418 35758 50430 35810
rect 50482 35758 50494 35810
rect 51762 35758 51774 35810
rect 51826 35758 51838 35810
rect 55458 35758 55470 35810
rect 55522 35758 55534 35810
rect 38222 35746 38274 35758
rect 50206 35746 50258 35758
rect 57822 35746 57874 35758
rect 1710 35698 1762 35710
rect 1710 35634 1762 35646
rect 2830 35698 2882 35710
rect 4286 35698 4338 35710
rect 3714 35646 3726 35698
rect 3778 35646 3790 35698
rect 2830 35634 2882 35646
rect 4286 35634 4338 35646
rect 5630 35698 5682 35710
rect 6526 35698 6578 35710
rect 6066 35646 6078 35698
rect 6130 35646 6142 35698
rect 5630 35634 5682 35646
rect 6526 35634 6578 35646
rect 7198 35698 7250 35710
rect 12910 35698 12962 35710
rect 8642 35646 8654 35698
rect 8706 35646 8718 35698
rect 10658 35646 10670 35698
rect 10722 35646 10734 35698
rect 7198 35634 7250 35646
rect 12910 35634 12962 35646
rect 13470 35698 13522 35710
rect 13470 35634 13522 35646
rect 13806 35698 13858 35710
rect 17950 35698 18002 35710
rect 28030 35698 28082 35710
rect 14354 35646 14366 35698
rect 14418 35646 14430 35698
rect 15026 35646 15038 35698
rect 15090 35646 15102 35698
rect 15362 35646 15374 35698
rect 15426 35646 15438 35698
rect 16370 35646 16382 35698
rect 16434 35646 16446 35698
rect 25218 35646 25230 35698
rect 25282 35646 25294 35698
rect 13806 35634 13858 35646
rect 17950 35634 18002 35646
rect 7758 35586 7810 35598
rect 7758 35522 7810 35534
rect 9662 35586 9714 35598
rect 17838 35586 17890 35598
rect 21086 35586 21138 35598
rect 14242 35534 14254 35586
rect 14306 35534 14318 35586
rect 15698 35534 15710 35586
rect 15762 35534 15774 35586
rect 16034 35534 16046 35586
rect 16098 35534 16110 35586
rect 19282 35534 19294 35586
rect 19346 35534 19358 35586
rect 9662 35522 9714 35534
rect 17838 35522 17890 35534
rect 21086 35522 21138 35534
rect 23438 35586 23490 35598
rect 23438 35522 23490 35534
rect 24670 35586 24722 35598
rect 24670 35522 24722 35534
rect 7982 35474 8034 35486
rect 4386 35422 4398 35474
rect 4450 35422 4462 35474
rect 7982 35410 8034 35422
rect 8318 35474 8370 35486
rect 8318 35410 8370 35422
rect 8654 35474 8706 35486
rect 8654 35410 8706 35422
rect 8990 35474 9042 35486
rect 8990 35410 9042 35422
rect 13022 35474 13074 35486
rect 13022 35410 13074 35422
rect 23774 35474 23826 35486
rect 25233 35471 25279 35646
rect 28030 35634 28082 35646
rect 28254 35698 28306 35710
rect 28254 35634 28306 35646
rect 32510 35698 32562 35710
rect 32510 35634 32562 35646
rect 33294 35698 33346 35710
rect 38110 35698 38162 35710
rect 34850 35646 34862 35698
rect 34914 35646 34926 35698
rect 33294 35634 33346 35646
rect 38110 35634 38162 35646
rect 38446 35698 38498 35710
rect 38446 35634 38498 35646
rect 38558 35698 38610 35710
rect 41806 35698 41858 35710
rect 58158 35698 58210 35710
rect 41122 35646 41134 35698
rect 41186 35646 41198 35698
rect 42578 35646 42590 35698
rect 42642 35646 42654 35698
rect 49634 35646 49646 35698
rect 49698 35646 49710 35698
rect 51538 35646 51550 35698
rect 51602 35646 51614 35698
rect 54450 35646 54462 35698
rect 54514 35646 54526 35698
rect 55234 35646 55246 35698
rect 55298 35646 55310 35698
rect 38558 35634 38610 35646
rect 41806 35634 41858 35646
rect 58158 35634 58210 35646
rect 25342 35586 25394 35598
rect 25342 35522 25394 35534
rect 25790 35586 25842 35598
rect 25790 35522 25842 35534
rect 29374 35586 29426 35598
rect 29374 35522 29426 35534
rect 30494 35586 30546 35598
rect 30494 35522 30546 35534
rect 31950 35586 32002 35598
rect 31950 35522 32002 35534
rect 33854 35586 33906 35598
rect 33854 35522 33906 35534
rect 34190 35586 34242 35598
rect 39118 35586 39170 35598
rect 35522 35534 35534 35586
rect 35586 35534 35598 35586
rect 37650 35534 37662 35586
rect 37714 35534 37726 35586
rect 38210 35534 38222 35586
rect 38274 35534 38286 35586
rect 34190 35522 34242 35534
rect 39118 35522 39170 35534
rect 43710 35586 43762 35598
rect 43710 35522 43762 35534
rect 45726 35586 45778 35598
rect 45726 35522 45778 35534
rect 57598 35586 57650 35598
rect 57598 35522 57650 35534
rect 53118 35474 53170 35486
rect 25778 35471 25790 35474
rect 25233 35425 25790 35471
rect 25778 35422 25790 35425
rect 25842 35422 25854 35474
rect 28914 35422 28926 35474
rect 28978 35471 28990 35474
rect 29250 35471 29262 35474
rect 28978 35425 29262 35471
rect 28978 35422 28990 35425
rect 29250 35422 29262 35425
rect 29314 35422 29326 35474
rect 42802 35422 42814 35474
rect 42866 35422 42878 35474
rect 23774 35410 23826 35422
rect 53118 35410 53170 35422
rect 1344 35306 58576 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 58576 35306
rect 1344 35220 58576 35254
rect 4398 35138 4450 35150
rect 4398 35074 4450 35086
rect 9774 35138 9826 35150
rect 9774 35074 9826 35086
rect 10670 35138 10722 35150
rect 19070 35138 19122 35150
rect 17714 35086 17726 35138
rect 17778 35086 17790 35138
rect 10670 35074 10722 35086
rect 19070 35074 19122 35086
rect 33182 35138 33234 35150
rect 33182 35074 33234 35086
rect 34414 35138 34466 35150
rect 34414 35074 34466 35086
rect 34638 35138 34690 35150
rect 34638 35074 34690 35086
rect 35982 35138 36034 35150
rect 35982 35074 36034 35086
rect 37998 35138 38050 35150
rect 37998 35074 38050 35086
rect 39790 35138 39842 35150
rect 54350 35138 54402 35150
rect 43138 35086 43150 35138
rect 43202 35086 43214 35138
rect 39790 35074 39842 35086
rect 54350 35074 54402 35086
rect 54574 35138 54626 35150
rect 54574 35074 54626 35086
rect 4174 35026 4226 35038
rect 4174 34962 4226 34974
rect 4734 35026 4786 35038
rect 9550 35026 9602 35038
rect 16158 35026 16210 35038
rect 18846 35026 18898 35038
rect 6850 34974 6862 35026
rect 6914 34974 6926 35026
rect 8754 34974 8766 35026
rect 8818 34974 8830 35026
rect 13570 34974 13582 35026
rect 13634 34974 13646 35026
rect 17154 34974 17166 35026
rect 17218 34974 17230 35026
rect 4734 34962 4786 34974
rect 9550 34962 9602 34974
rect 16158 34962 16210 34974
rect 18846 34962 18898 34974
rect 20190 35026 20242 35038
rect 20190 34962 20242 34974
rect 21870 35026 21922 35038
rect 30494 35026 30546 35038
rect 27906 34974 27918 35026
rect 27970 34974 27982 35026
rect 21870 34962 21922 34974
rect 30494 34962 30546 34974
rect 30942 35026 30994 35038
rect 38782 35026 38834 35038
rect 32498 34974 32510 35026
rect 32562 34974 32574 35026
rect 30942 34962 30994 34974
rect 38782 34962 38834 34974
rect 39454 35026 39506 35038
rect 41806 35026 41858 35038
rect 52670 35026 52722 35038
rect 40338 34974 40350 35026
rect 40402 34974 40414 35026
rect 42578 34974 42590 35026
rect 42642 34974 42654 35026
rect 39454 34962 39506 34974
rect 41806 34962 41858 34974
rect 52670 34962 52722 34974
rect 5854 34914 5906 34926
rect 10558 34914 10610 34926
rect 15710 34914 15762 34926
rect 2594 34862 2606 34914
rect 2658 34862 2670 34914
rect 3154 34862 3166 34914
rect 3218 34862 3230 34914
rect 3602 34862 3614 34914
rect 3666 34862 3678 34914
rect 7298 34862 7310 34914
rect 7362 34862 7374 34914
rect 8306 34862 8318 34914
rect 8370 34862 8382 34914
rect 9202 34862 9214 34914
rect 9266 34862 9278 34914
rect 15138 34862 15150 34914
rect 15202 34862 15214 34914
rect 5854 34850 5906 34862
rect 10558 34850 10610 34862
rect 15710 34850 15762 34862
rect 16046 34914 16098 34926
rect 19742 34914 19794 34926
rect 16370 34862 16382 34914
rect 16434 34862 16446 34914
rect 17490 34862 17502 34914
rect 17554 34862 17566 34914
rect 19394 34862 19406 34914
rect 19458 34862 19470 34914
rect 16046 34850 16098 34862
rect 19742 34850 19794 34862
rect 19966 34914 20018 34926
rect 19966 34850 20018 34862
rect 20414 34914 20466 34926
rect 24222 34914 24274 34926
rect 23986 34862 23998 34914
rect 24050 34862 24062 34914
rect 20414 34850 20466 34862
rect 24222 34850 24274 34862
rect 24558 34914 24610 34926
rect 28478 34914 28530 34926
rect 24994 34862 25006 34914
rect 25058 34862 25070 34914
rect 24558 34850 24610 34862
rect 28478 34850 28530 34862
rect 29262 34914 29314 34926
rect 29262 34850 29314 34862
rect 29598 34914 29650 34926
rect 33966 34914 34018 34926
rect 33506 34862 33518 34914
rect 33570 34862 33582 34914
rect 29598 34850 29650 34862
rect 33966 34850 34018 34862
rect 35086 34914 35138 34926
rect 35086 34850 35138 34862
rect 38222 34914 38274 34926
rect 38222 34850 38274 34862
rect 40798 34914 40850 34926
rect 43822 34914 43874 34926
rect 41122 34862 41134 34914
rect 41186 34862 41198 34914
rect 42690 34862 42702 34914
rect 42754 34862 42766 34914
rect 40798 34850 40850 34862
rect 43822 34850 43874 34862
rect 44158 34914 44210 34926
rect 45726 34914 45778 34926
rect 49982 34914 50034 34926
rect 45266 34862 45278 34914
rect 45330 34862 45342 34914
rect 47058 34862 47070 34914
rect 47122 34862 47134 34914
rect 48514 34862 48526 34914
rect 48578 34862 48590 34914
rect 48850 34862 48862 34914
rect 48914 34862 48926 34914
rect 44158 34850 44210 34862
rect 45726 34850 45778 34862
rect 49982 34850 50034 34862
rect 51886 34914 51938 34926
rect 51886 34850 51938 34862
rect 52222 34914 52274 34926
rect 52222 34850 52274 34862
rect 53454 34914 53506 34926
rect 53454 34850 53506 34862
rect 53902 34914 53954 34926
rect 53902 34850 53954 34862
rect 54798 34914 54850 34926
rect 54798 34850 54850 34862
rect 7758 34802 7810 34814
rect 10670 34802 10722 34814
rect 28366 34802 28418 34814
rect 2034 34750 2046 34802
rect 2098 34750 2110 34802
rect 2482 34750 2494 34802
rect 2546 34750 2558 34802
rect 3826 34750 3838 34802
rect 3890 34750 3902 34802
rect 9090 34750 9102 34802
rect 9154 34750 9166 34802
rect 13906 34750 13918 34802
rect 13970 34750 13982 34802
rect 25778 34750 25790 34802
rect 25842 34750 25854 34802
rect 7758 34738 7810 34750
rect 10670 34738 10722 34750
rect 28366 34738 28418 34750
rect 29374 34802 29426 34814
rect 29374 34738 29426 34750
rect 29934 34802 29986 34814
rect 29934 34738 29986 34750
rect 30046 34802 30098 34814
rect 30046 34738 30098 34750
rect 30830 34802 30882 34814
rect 30830 34738 30882 34750
rect 31166 34802 31218 34814
rect 31166 34738 31218 34750
rect 31390 34802 31442 34814
rect 31390 34738 31442 34750
rect 32062 34802 32114 34814
rect 32062 34738 32114 34750
rect 33854 34802 33906 34814
rect 33854 34738 33906 34750
rect 35198 34802 35250 34814
rect 35198 34738 35250 34750
rect 35870 34802 35922 34814
rect 35870 34738 35922 34750
rect 37102 34802 37154 34814
rect 37102 34738 37154 34750
rect 37214 34802 37266 34814
rect 37214 34738 37266 34750
rect 39678 34802 39730 34814
rect 39678 34738 39730 34750
rect 39790 34802 39842 34814
rect 39790 34738 39842 34750
rect 44830 34802 44882 34814
rect 44830 34738 44882 34750
rect 46174 34802 46226 34814
rect 51998 34802 52050 34814
rect 53006 34802 53058 34814
rect 48962 34750 48974 34802
rect 49026 34750 49038 34802
rect 52770 34750 52782 34802
rect 52834 34750 52846 34802
rect 46174 34738 46226 34750
rect 51998 34738 52050 34750
rect 53006 34738 53058 34750
rect 1710 34690 1762 34702
rect 1710 34626 1762 34638
rect 6190 34690 6242 34702
rect 20526 34690 20578 34702
rect 10098 34638 10110 34690
rect 10162 34638 10174 34690
rect 6190 34626 6242 34638
rect 20526 34626 20578 34638
rect 20638 34690 20690 34702
rect 20638 34626 20690 34638
rect 21422 34690 21474 34702
rect 21422 34626 21474 34638
rect 24334 34690 24386 34702
rect 24334 34626 24386 34638
rect 24446 34690 24498 34702
rect 24446 34626 24498 34638
rect 28142 34690 28194 34702
rect 28142 34626 28194 34638
rect 29710 34690 29762 34702
rect 29710 34626 29762 34638
rect 32286 34690 32338 34702
rect 32286 34626 32338 34638
rect 32510 34690 32562 34702
rect 32510 34626 32562 34638
rect 33294 34690 33346 34702
rect 33294 34626 33346 34638
rect 34750 34690 34802 34702
rect 34750 34626 34802 34638
rect 35422 34690 35474 34702
rect 35422 34626 35474 34638
rect 35982 34690 36034 34702
rect 35982 34626 36034 34638
rect 36878 34690 36930 34702
rect 40238 34690 40290 34702
rect 37650 34638 37662 34690
rect 37714 34638 37726 34690
rect 36878 34626 36930 34638
rect 40238 34626 40290 34638
rect 40462 34690 40514 34702
rect 40462 34626 40514 34638
rect 41358 34690 41410 34702
rect 41358 34626 41410 34638
rect 43934 34690 43986 34702
rect 43934 34626 43986 34638
rect 46286 34690 46338 34702
rect 46286 34626 46338 34638
rect 46510 34690 46562 34702
rect 46510 34626 46562 34638
rect 49646 34690 49698 34702
rect 49646 34626 49698 34638
rect 49870 34690 49922 34702
rect 49870 34626 49922 34638
rect 53678 34690 53730 34702
rect 53678 34626 53730 34638
rect 1344 34522 58576 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 50558 34522
rect 50610 34470 50662 34522
rect 50714 34470 50766 34522
rect 50818 34470 58576 34522
rect 1344 34436 58576 34470
rect 4510 34354 4562 34366
rect 4510 34290 4562 34302
rect 5854 34354 5906 34366
rect 5854 34290 5906 34302
rect 7310 34354 7362 34366
rect 7310 34290 7362 34302
rect 7534 34354 7586 34366
rect 7534 34290 7586 34302
rect 8654 34354 8706 34366
rect 8654 34290 8706 34302
rect 9662 34354 9714 34366
rect 9662 34290 9714 34302
rect 10334 34354 10386 34366
rect 15598 34354 15650 34366
rect 15250 34302 15262 34354
rect 15314 34302 15326 34354
rect 10334 34290 10386 34302
rect 15598 34290 15650 34302
rect 26014 34354 26066 34366
rect 26014 34290 26066 34302
rect 26126 34354 26178 34366
rect 26126 34290 26178 34302
rect 26238 34354 26290 34366
rect 32958 34354 33010 34366
rect 27346 34302 27358 34354
rect 27410 34302 27422 34354
rect 26238 34290 26290 34302
rect 32958 34290 33010 34302
rect 35422 34354 35474 34366
rect 35422 34290 35474 34302
rect 37550 34354 37602 34366
rect 37550 34290 37602 34302
rect 41246 34354 41298 34366
rect 41246 34290 41298 34302
rect 42926 34354 42978 34366
rect 42926 34290 42978 34302
rect 43486 34354 43538 34366
rect 43486 34290 43538 34302
rect 44494 34354 44546 34366
rect 49310 34354 49362 34366
rect 53454 34354 53506 34366
rect 45602 34302 45614 34354
rect 45666 34302 45678 34354
rect 52770 34302 52782 34354
rect 52834 34302 52846 34354
rect 44494 34290 44546 34302
rect 49310 34290 49362 34302
rect 53454 34290 53506 34302
rect 7086 34242 7138 34254
rect 12350 34242 12402 34254
rect 5058 34190 5070 34242
rect 5122 34190 5134 34242
rect 9986 34190 9998 34242
rect 10050 34190 10062 34242
rect 10658 34190 10670 34242
rect 10722 34190 10734 34242
rect 7086 34178 7138 34190
rect 12350 34178 12402 34190
rect 14254 34242 14306 34254
rect 14254 34178 14306 34190
rect 15710 34242 15762 34254
rect 20862 34242 20914 34254
rect 19730 34190 19742 34242
rect 19794 34190 19806 34242
rect 15710 34178 15762 34190
rect 20862 34178 20914 34190
rect 25342 34242 25394 34254
rect 31278 34242 31330 34254
rect 30034 34190 30046 34242
rect 30098 34190 30110 34242
rect 25342 34178 25394 34190
rect 31278 34178 31330 34190
rect 31614 34242 31666 34254
rect 34974 34242 35026 34254
rect 33730 34190 33742 34242
rect 33794 34190 33806 34242
rect 31614 34178 31666 34190
rect 34974 34178 35026 34190
rect 40910 34242 40962 34254
rect 40910 34178 40962 34190
rect 41134 34242 41186 34254
rect 41134 34178 41186 34190
rect 42142 34242 42194 34254
rect 42142 34178 42194 34190
rect 43038 34242 43090 34254
rect 43038 34178 43090 34190
rect 43598 34242 43650 34254
rect 43598 34178 43650 34190
rect 44606 34242 44658 34254
rect 49198 34242 49250 34254
rect 53342 34242 53394 34254
rect 47506 34190 47518 34242
rect 47570 34190 47582 34242
rect 51986 34190 51998 34242
rect 52050 34190 52062 34242
rect 44606 34178 44658 34190
rect 49198 34178 49250 34190
rect 53342 34178 53394 34190
rect 4734 34130 4786 34142
rect 4274 34078 4286 34130
rect 4338 34078 4350 34130
rect 4734 34066 4786 34078
rect 5294 34130 5346 34142
rect 5294 34066 5346 34078
rect 5518 34130 5570 34142
rect 5518 34066 5570 34078
rect 6750 34130 6802 34142
rect 6750 34066 6802 34078
rect 7646 34130 7698 34142
rect 8430 34130 8482 34142
rect 8082 34078 8094 34130
rect 8146 34078 8158 34130
rect 7646 34066 7698 34078
rect 8430 34066 8482 34078
rect 8542 34130 8594 34142
rect 14142 34130 14194 34142
rect 11330 34078 11342 34130
rect 11394 34078 11406 34130
rect 13570 34078 13582 34130
rect 13634 34078 13646 34130
rect 8542 34066 8594 34078
rect 14142 34066 14194 34078
rect 14926 34130 14978 34142
rect 25118 34130 25170 34142
rect 20402 34078 20414 34130
rect 20466 34078 20478 34130
rect 21074 34078 21086 34130
rect 21138 34078 21150 34130
rect 24546 34078 24558 34130
rect 24610 34078 24622 34130
rect 14926 34066 14978 34078
rect 25118 34066 25170 34078
rect 25454 34130 25506 34142
rect 25454 34066 25506 34078
rect 26686 34130 26738 34142
rect 26686 34066 26738 34078
rect 27022 34130 27074 34142
rect 32062 34130 32114 34142
rect 30706 34078 30718 34130
rect 30770 34078 30782 34130
rect 27022 34066 27074 34078
rect 32062 34066 32114 34078
rect 32174 34130 32226 34142
rect 32174 34066 32226 34078
rect 32398 34130 32450 34142
rect 32398 34066 32450 34078
rect 32622 34130 32674 34142
rect 32622 34066 32674 34078
rect 33070 34130 33122 34142
rect 33070 34066 33122 34078
rect 33518 34130 33570 34142
rect 35198 34130 35250 34142
rect 41582 34130 41634 34142
rect 42590 34130 42642 34142
rect 33954 34078 33966 34130
rect 34018 34078 34030 34130
rect 35634 34078 35646 34130
rect 35698 34078 35710 34130
rect 39890 34078 39902 34130
rect 39954 34078 39966 34130
rect 41794 34078 41806 34130
rect 41858 34078 41870 34130
rect 33518 34066 33570 34078
rect 35198 34066 35250 34078
rect 41582 34066 41634 34078
rect 42590 34066 42642 34078
rect 43150 34130 43202 34142
rect 44158 34130 44210 34142
rect 43810 34078 43822 34130
rect 43874 34078 43886 34130
rect 43150 34066 43202 34078
rect 44158 34066 44210 34078
rect 44270 34130 44322 34142
rect 45950 34130 46002 34142
rect 49534 34130 49586 34142
rect 50654 34130 50706 34142
rect 53678 34130 53730 34142
rect 45378 34078 45390 34130
rect 45442 34078 45454 34130
rect 46610 34078 46622 34130
rect 46674 34078 46686 34130
rect 50306 34078 50318 34130
rect 50370 34078 50382 34130
rect 52434 34078 52446 34130
rect 52498 34078 52510 34130
rect 52994 34078 53006 34130
rect 53058 34078 53070 34130
rect 44270 34066 44322 34078
rect 45950 34066 46002 34078
rect 49534 34066 49586 34078
rect 50654 34066 50706 34078
rect 53678 34066 53730 34078
rect 12014 34018 12066 34030
rect 27918 34018 27970 34030
rect 6290 33966 6302 34018
rect 6354 33966 6366 34018
rect 11554 33966 11566 34018
rect 11618 33966 11630 34018
rect 17602 33966 17614 34018
rect 17666 33966 17678 34018
rect 21746 33966 21758 34018
rect 21810 33966 21822 34018
rect 23874 33966 23886 34018
rect 23938 33966 23950 34018
rect 12014 33954 12066 33966
rect 27918 33954 27970 33966
rect 33294 34018 33346 34030
rect 33294 33954 33346 33966
rect 35310 34018 35362 34030
rect 35310 33954 35362 33966
rect 36654 34018 36706 34030
rect 36654 33954 36706 33966
rect 39230 34018 39282 34030
rect 49758 34018 49810 34030
rect 40114 33966 40126 34018
rect 40178 33966 40190 34018
rect 41906 33966 41918 34018
rect 41970 33966 41982 34018
rect 48066 33966 48078 34018
rect 48130 33966 48142 34018
rect 39230 33954 39282 33966
rect 49758 33954 49810 33966
rect 1934 33906 1986 33918
rect 1934 33842 1986 33854
rect 12462 33906 12514 33918
rect 12462 33842 12514 33854
rect 1344 33738 58576 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 58576 33738
rect 1344 33652 58576 33686
rect 19518 33570 19570 33582
rect 19518 33506 19570 33518
rect 19854 33570 19906 33582
rect 19854 33506 19906 33518
rect 30606 33570 30658 33582
rect 30606 33506 30658 33518
rect 40350 33570 40402 33582
rect 40350 33506 40402 33518
rect 41022 33570 41074 33582
rect 41022 33506 41074 33518
rect 41806 33570 41858 33582
rect 41806 33506 41858 33518
rect 42142 33570 42194 33582
rect 42142 33506 42194 33518
rect 43822 33570 43874 33582
rect 43822 33506 43874 33518
rect 3614 33458 3666 33470
rect 3614 33394 3666 33406
rect 8430 33458 8482 33470
rect 8430 33394 8482 33406
rect 9326 33458 9378 33470
rect 19182 33458 19234 33470
rect 27806 33458 27858 33470
rect 9986 33406 9998 33458
rect 10050 33406 10062 33458
rect 12786 33406 12798 33458
rect 12850 33406 12862 33458
rect 14466 33406 14478 33458
rect 14530 33406 14542 33458
rect 23538 33406 23550 33458
rect 23602 33406 23614 33458
rect 9326 33394 9378 33406
rect 19182 33394 19234 33406
rect 27806 33394 27858 33406
rect 29262 33458 29314 33470
rect 40126 33458 40178 33470
rect 31938 33406 31950 33458
rect 32002 33406 32014 33458
rect 34402 33406 34414 33458
rect 34466 33406 34478 33458
rect 37090 33406 37102 33458
rect 37154 33406 37166 33458
rect 29262 33394 29314 33406
rect 40126 33394 40178 33406
rect 41134 33458 41186 33470
rect 46162 33406 46174 33458
rect 46226 33406 46238 33458
rect 48402 33406 48414 33458
rect 48466 33406 48478 33458
rect 51314 33406 51326 33458
rect 51378 33406 51390 33458
rect 54898 33406 54910 33458
rect 54962 33406 54974 33458
rect 57810 33406 57822 33458
rect 57874 33406 57886 33458
rect 41134 33394 41186 33406
rect 3502 33346 3554 33358
rect 3502 33282 3554 33294
rect 3838 33346 3890 33358
rect 15262 33346 15314 33358
rect 21758 33346 21810 33358
rect 31390 33346 31442 33358
rect 4050 33294 4062 33346
rect 4114 33294 4126 33346
rect 5954 33294 5966 33346
rect 6018 33294 6030 33346
rect 7074 33294 7086 33346
rect 7138 33294 7150 33346
rect 11554 33294 11566 33346
rect 11618 33294 11630 33346
rect 14354 33294 14366 33346
rect 14418 33294 14430 33346
rect 20626 33294 20638 33346
rect 20690 33294 20702 33346
rect 26786 33294 26798 33346
rect 26850 33294 26862 33346
rect 3838 33282 3890 33294
rect 15262 33282 15314 33294
rect 21758 33282 21810 33294
rect 31390 33282 31442 33294
rect 31614 33346 31666 33358
rect 35534 33346 35586 33358
rect 34514 33294 34526 33346
rect 34578 33294 34590 33346
rect 31614 33282 31666 33294
rect 35534 33282 35586 33294
rect 37886 33346 37938 33358
rect 37886 33282 37938 33294
rect 38558 33346 38610 33358
rect 38558 33282 38610 33294
rect 41918 33346 41970 33358
rect 45166 33346 45218 33358
rect 47518 33346 47570 33358
rect 42690 33294 42702 33346
rect 42754 33294 42766 33346
rect 42914 33294 42926 33346
rect 42978 33294 42990 33346
rect 43922 33294 43934 33346
rect 43986 33294 43998 33346
rect 46274 33294 46286 33346
rect 46338 33294 46350 33346
rect 47170 33294 47182 33346
rect 47234 33294 47246 33346
rect 48066 33294 48078 33346
rect 48130 33294 48142 33346
rect 49858 33294 49870 33346
rect 49922 33294 49934 33346
rect 53778 33294 53790 33346
rect 53842 33294 53854 33346
rect 54562 33294 54574 33346
rect 54626 33294 54638 33346
rect 55570 33294 55582 33346
rect 55634 33294 55646 33346
rect 41918 33282 41970 33294
rect 45166 33282 45218 33294
rect 47518 33282 47570 33294
rect 7758 33234 7810 33246
rect 30158 33234 30210 33246
rect 2034 33182 2046 33234
rect 2098 33182 2110 33234
rect 2706 33182 2718 33234
rect 2770 33182 2782 33234
rect 4946 33182 4958 33234
rect 5010 33182 5022 33234
rect 6178 33182 6190 33234
rect 6242 33182 6254 33234
rect 10434 33182 10446 33234
rect 10498 33182 10510 33234
rect 20514 33182 20526 33234
rect 20578 33182 20590 33234
rect 21410 33182 21422 33234
rect 21474 33182 21486 33234
rect 28130 33182 28142 33234
rect 28194 33182 28206 33234
rect 7758 33170 7810 33182
rect 30158 33170 30210 33182
rect 30494 33234 30546 33246
rect 30494 33170 30546 33182
rect 30606 33234 30658 33246
rect 30606 33170 30658 33182
rect 31054 33234 31106 33246
rect 31054 33170 31106 33182
rect 31166 33234 31218 33246
rect 31166 33170 31218 33182
rect 34862 33234 34914 33246
rect 34862 33170 34914 33182
rect 35870 33234 35922 33246
rect 35870 33170 35922 33182
rect 36094 33234 36146 33246
rect 36094 33170 36146 33182
rect 37326 33234 37378 33246
rect 37326 33170 37378 33182
rect 38334 33234 38386 33246
rect 38334 33170 38386 33182
rect 42254 33234 42306 33246
rect 54126 33234 54178 33246
rect 44818 33182 44830 33234
rect 44882 33182 44894 33234
rect 46050 33182 46062 33234
rect 46114 33182 46126 33234
rect 50754 33182 50766 33234
rect 50818 33182 50830 33234
rect 53106 33182 53118 33234
rect 53170 33182 53182 33234
rect 53554 33182 53566 33234
rect 53618 33182 53630 33234
rect 42254 33170 42306 33182
rect 54126 33170 54178 33182
rect 1710 33122 1762 33134
rect 1710 33058 1762 33070
rect 2382 33122 2434 33134
rect 7870 33122 7922 33134
rect 6514 33070 6526 33122
rect 6578 33070 6590 33122
rect 7298 33070 7310 33122
rect 7362 33070 7374 33122
rect 2382 33058 2434 33070
rect 7870 33058 7922 33070
rect 8094 33122 8146 33134
rect 8094 33058 8146 33070
rect 8878 33122 8930 33134
rect 8878 33058 8930 33070
rect 28478 33122 28530 33134
rect 28478 33058 28530 33070
rect 29710 33122 29762 33134
rect 29710 33058 29762 33070
rect 31950 33122 32002 33134
rect 31950 33058 32002 33070
rect 32174 33122 32226 33134
rect 32174 33058 32226 33070
rect 32734 33122 32786 33134
rect 32734 33058 32786 33070
rect 34974 33122 35026 33134
rect 34974 33058 35026 33070
rect 35198 33122 35250 33134
rect 35198 33058 35250 33070
rect 35758 33122 35810 33134
rect 35758 33058 35810 33070
rect 37102 33122 37154 33134
rect 37102 33058 37154 33070
rect 38222 33122 38274 33134
rect 40674 33070 40686 33122
rect 40738 33070 40750 33122
rect 49298 33070 49310 33122
rect 49362 33070 49374 33122
rect 53218 33070 53230 33122
rect 53282 33070 53294 33122
rect 38222 33058 38274 33070
rect 1344 32954 58576 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 50558 32954
rect 50610 32902 50662 32954
rect 50714 32902 50766 32954
rect 50818 32902 58576 32954
rect 1344 32868 58576 32902
rect 5518 32786 5570 32798
rect 9662 32786 9714 32798
rect 3266 32734 3278 32786
rect 3330 32734 3342 32786
rect 7074 32734 7086 32786
rect 7138 32734 7150 32786
rect 5518 32722 5570 32734
rect 9662 32722 9714 32734
rect 17838 32786 17890 32798
rect 17838 32722 17890 32734
rect 18734 32786 18786 32798
rect 18734 32722 18786 32734
rect 20526 32786 20578 32798
rect 20526 32722 20578 32734
rect 25454 32786 25506 32798
rect 42142 32786 42194 32798
rect 26562 32734 26574 32786
rect 26626 32734 26638 32786
rect 29810 32734 29822 32786
rect 29874 32734 29886 32786
rect 25454 32722 25506 32734
rect 42142 32722 42194 32734
rect 49646 32786 49698 32798
rect 49646 32722 49698 32734
rect 51662 32786 51714 32798
rect 51662 32722 51714 32734
rect 52222 32786 52274 32798
rect 56690 32734 56702 32786
rect 56754 32734 56766 32786
rect 52222 32722 52274 32734
rect 6190 32674 6242 32686
rect 2482 32622 2494 32674
rect 2546 32622 2558 32674
rect 5954 32622 5966 32674
rect 6018 32622 6030 32674
rect 6190 32610 6242 32622
rect 9550 32674 9602 32686
rect 9550 32610 9602 32622
rect 10110 32674 10162 32686
rect 10110 32610 10162 32622
rect 20862 32674 20914 32686
rect 42814 32674 42866 32686
rect 31042 32622 31054 32674
rect 31106 32622 31118 32674
rect 20862 32610 20914 32622
rect 42814 32610 42866 32622
rect 42926 32674 42978 32686
rect 49758 32674 49810 32686
rect 43698 32622 43710 32674
rect 43762 32622 43774 32674
rect 45154 32622 45166 32674
rect 45218 32622 45230 32674
rect 42926 32610 42978 32622
rect 49758 32610 49810 32622
rect 51550 32674 51602 32686
rect 51550 32610 51602 32622
rect 52670 32674 52722 32686
rect 52670 32610 52722 32622
rect 53006 32674 53058 32686
rect 53006 32610 53058 32622
rect 53230 32674 53282 32686
rect 57250 32622 57262 32674
rect 57314 32622 57326 32674
rect 53230 32610 53282 32622
rect 4958 32562 5010 32574
rect 2258 32510 2270 32562
rect 2322 32510 2334 32562
rect 3938 32510 3950 32562
rect 4002 32510 4014 32562
rect 4958 32498 5010 32510
rect 5854 32562 5906 32574
rect 5854 32498 5906 32510
rect 6638 32562 6690 32574
rect 6638 32498 6690 32510
rect 7422 32562 7474 32574
rect 7422 32498 7474 32510
rect 7646 32562 7698 32574
rect 10222 32562 10274 32574
rect 17390 32562 17442 32574
rect 18062 32562 18114 32574
rect 25118 32562 25170 32574
rect 8082 32510 8094 32562
rect 8146 32510 8158 32562
rect 8530 32510 8542 32562
rect 8594 32510 8606 32562
rect 11890 32510 11902 32562
rect 11954 32510 11966 32562
rect 13458 32510 13470 32562
rect 13522 32510 13534 32562
rect 14466 32510 14478 32562
rect 14530 32510 14542 32562
rect 15250 32510 15262 32562
rect 15314 32510 15326 32562
rect 17714 32510 17726 32562
rect 17778 32510 17790 32562
rect 21298 32510 21310 32562
rect 21362 32510 21374 32562
rect 24546 32510 24558 32562
rect 24610 32510 24622 32562
rect 7646 32498 7698 32510
rect 10222 32498 10274 32510
rect 17390 32498 17442 32510
rect 18062 32498 18114 32510
rect 25118 32498 25170 32510
rect 25454 32562 25506 32574
rect 25454 32498 25506 32510
rect 25790 32562 25842 32574
rect 28702 32562 28754 32574
rect 30718 32562 30770 32574
rect 42366 32562 42418 32574
rect 26338 32510 26350 32562
rect 26402 32510 26414 32562
rect 29026 32510 29038 32562
rect 29090 32510 29102 32562
rect 34738 32510 34750 32562
rect 34802 32510 34814 32562
rect 25790 32498 25842 32510
rect 28702 32498 28754 32510
rect 30718 32498 30770 32510
rect 42366 32498 42418 32510
rect 42590 32562 42642 32574
rect 51886 32562 51938 32574
rect 43810 32510 43822 32562
rect 43874 32510 43886 32562
rect 44706 32510 44718 32562
rect 44770 32510 44782 32562
rect 45266 32510 45278 32562
rect 45330 32510 45342 32562
rect 45826 32510 45838 32562
rect 45890 32510 45902 32562
rect 46610 32510 46622 32562
rect 46674 32510 46686 32562
rect 42590 32498 42642 32510
rect 51886 32498 51938 32510
rect 52110 32562 52162 32574
rect 52110 32498 52162 32510
rect 52446 32562 52498 32574
rect 54686 32562 54738 32574
rect 54450 32510 54462 32562
rect 54514 32510 54526 32562
rect 52446 32498 52498 32510
rect 54686 32498 54738 32510
rect 54910 32562 54962 32574
rect 56578 32510 56590 32562
rect 56642 32510 56654 32562
rect 57138 32510 57150 32562
rect 57202 32510 57214 32562
rect 54910 32498 54962 32510
rect 17950 32450 18002 32462
rect 27022 32450 27074 32462
rect 12338 32398 12350 32450
rect 12402 32398 12414 32450
rect 13570 32398 13582 32450
rect 13634 32398 13646 32450
rect 15138 32398 15150 32450
rect 15202 32398 15214 32450
rect 21746 32398 21758 32450
rect 21810 32398 21822 32450
rect 23874 32398 23886 32450
rect 23938 32398 23950 32450
rect 17950 32386 18002 32398
rect 27022 32386 27074 32398
rect 27470 32450 27522 32462
rect 27470 32386 27522 32398
rect 27918 32450 27970 32462
rect 27918 32386 27970 32398
rect 28254 32450 28306 32462
rect 28254 32386 28306 32398
rect 29486 32450 29538 32462
rect 29486 32386 29538 32398
rect 30382 32450 30434 32462
rect 30382 32386 30434 32398
rect 31502 32450 31554 32462
rect 31502 32386 31554 32398
rect 33182 32450 33234 32462
rect 52782 32450 52834 32462
rect 38322 32398 38334 32450
rect 38386 32398 38398 32450
rect 43922 32398 43934 32450
rect 43986 32398 43998 32450
rect 33182 32386 33234 32398
rect 52782 32386 52834 32398
rect 6862 32338 6914 32350
rect 9662 32338 9714 32350
rect 28366 32338 28418 32350
rect 8082 32286 8094 32338
rect 8146 32286 8158 32338
rect 27458 32286 27470 32338
rect 27522 32335 27534 32338
rect 27906 32335 27918 32338
rect 27522 32289 27918 32335
rect 27522 32286 27534 32289
rect 27906 32286 27918 32289
rect 27970 32286 27982 32338
rect 6862 32274 6914 32286
rect 9662 32274 9714 32286
rect 28366 32274 28418 32286
rect 30158 32338 30210 32350
rect 30158 32274 30210 32286
rect 42030 32338 42082 32350
rect 42030 32274 42082 32286
rect 49646 32338 49698 32350
rect 49646 32274 49698 32286
rect 1344 32170 58576 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 58576 32170
rect 1344 32084 58576 32118
rect 17502 32002 17554 32014
rect 17502 31938 17554 31950
rect 23886 32002 23938 32014
rect 27694 32002 27746 32014
rect 26562 31950 26574 32002
rect 26626 31950 26638 32002
rect 23886 31938 23938 31950
rect 27694 31938 27746 31950
rect 34974 32002 35026 32014
rect 34974 31938 35026 31950
rect 45278 32002 45330 32014
rect 45278 31938 45330 31950
rect 1934 31890 1986 31902
rect 1934 31826 1986 31838
rect 5630 31890 5682 31902
rect 5630 31826 5682 31838
rect 7982 31890 8034 31902
rect 7982 31826 8034 31838
rect 8654 31890 8706 31902
rect 13694 31890 13746 31902
rect 12002 31838 12014 31890
rect 12066 31838 12078 31890
rect 8654 31826 8706 31838
rect 13694 31826 13746 31838
rect 16382 31890 16434 31902
rect 19182 31890 19234 31902
rect 16818 31838 16830 31890
rect 16882 31838 16894 31890
rect 16382 31826 16434 31838
rect 19182 31826 19234 31838
rect 22206 31890 22258 31902
rect 22206 31826 22258 31838
rect 22766 31890 22818 31902
rect 22766 31826 22818 31838
rect 23662 31890 23714 31902
rect 23662 31826 23714 31838
rect 23998 31890 24050 31902
rect 23998 31826 24050 31838
rect 26126 31890 26178 31902
rect 26126 31826 26178 31838
rect 28030 31890 28082 31902
rect 32398 31890 32450 31902
rect 35086 31890 35138 31902
rect 45054 31890 45106 31902
rect 29586 31838 29598 31890
rect 29650 31838 29662 31890
rect 34626 31838 34638 31890
rect 34690 31838 34702 31890
rect 35970 31838 35982 31890
rect 36034 31838 36046 31890
rect 39890 31838 39902 31890
rect 39954 31838 39966 31890
rect 28030 31826 28082 31838
rect 32398 31826 32450 31838
rect 35086 31826 35138 31838
rect 45054 31826 45106 31838
rect 47966 31890 48018 31902
rect 51550 31890 51602 31902
rect 49186 31838 49198 31890
rect 49250 31838 49262 31890
rect 47966 31826 48018 31838
rect 51550 31826 51602 31838
rect 52110 31890 52162 31902
rect 52110 31826 52162 31838
rect 57934 31890 57986 31902
rect 57934 31826 57986 31838
rect 4622 31778 4674 31790
rect 4274 31726 4286 31778
rect 4338 31726 4350 31778
rect 4622 31714 4674 31726
rect 6190 31778 6242 31790
rect 6190 31714 6242 31726
rect 7422 31778 7474 31790
rect 7422 31714 7474 31726
rect 8542 31778 8594 31790
rect 8542 31714 8594 31726
rect 8878 31778 8930 31790
rect 8878 31714 8930 31726
rect 9662 31778 9714 31790
rect 9662 31714 9714 31726
rect 10110 31778 10162 31790
rect 10110 31714 10162 31726
rect 10334 31778 10386 31790
rect 13918 31778 13970 31790
rect 14926 31778 14978 31790
rect 11778 31726 11790 31778
rect 11842 31726 11854 31778
rect 14242 31726 14254 31778
rect 14306 31726 14318 31778
rect 14578 31726 14590 31778
rect 14642 31726 14654 31778
rect 10334 31714 10386 31726
rect 13918 31714 13970 31726
rect 14926 31714 14978 31726
rect 16158 31778 16210 31790
rect 16158 31714 16210 31726
rect 16606 31778 16658 31790
rect 16606 31714 16658 31726
rect 17726 31778 17778 31790
rect 17726 31714 17778 31726
rect 25118 31778 25170 31790
rect 25118 31714 25170 31726
rect 25454 31778 25506 31790
rect 25454 31714 25506 31726
rect 26014 31778 26066 31790
rect 26014 31714 26066 31726
rect 26350 31778 26402 31790
rect 28254 31778 28306 31790
rect 26562 31726 26574 31778
rect 26626 31726 26638 31778
rect 27682 31726 27694 31778
rect 27746 31726 27758 31778
rect 26350 31714 26402 31726
rect 28254 31714 28306 31726
rect 29374 31778 29426 31790
rect 33182 31778 33234 31790
rect 29810 31726 29822 31778
rect 29874 31726 29886 31778
rect 31042 31726 31054 31778
rect 31106 31726 31118 31778
rect 31938 31726 31950 31778
rect 32002 31726 32014 31778
rect 29374 31714 29426 31726
rect 33182 31714 33234 31726
rect 33854 31778 33906 31790
rect 33854 31714 33906 31726
rect 36430 31778 36482 31790
rect 40350 31778 40402 31790
rect 46622 31778 46674 31790
rect 37090 31726 37102 31778
rect 37154 31726 37166 31778
rect 45490 31726 45502 31778
rect 45554 31726 45566 31778
rect 36430 31714 36482 31726
rect 40350 31714 40402 31726
rect 46622 31714 46674 31726
rect 48190 31778 48242 31790
rect 51886 31778 51938 31790
rect 48738 31726 48750 31778
rect 48802 31726 48814 31778
rect 49074 31726 49086 31778
rect 49138 31726 49150 31778
rect 53442 31726 53454 31778
rect 53506 31726 53518 31778
rect 54114 31726 54126 31778
rect 54178 31726 54190 31778
rect 55570 31726 55582 31778
rect 55634 31726 55646 31778
rect 48190 31714 48242 31726
rect 51886 31714 51938 31726
rect 16830 31666 16882 31678
rect 4946 31614 4958 31666
rect 5010 31614 5022 31666
rect 11666 31614 11678 31666
rect 11730 31614 11742 31666
rect 16830 31602 16882 31614
rect 18174 31666 18226 31678
rect 18174 31602 18226 31614
rect 18734 31666 18786 31678
rect 18734 31602 18786 31614
rect 24446 31666 24498 31678
rect 24446 31602 24498 31614
rect 25230 31666 25282 31678
rect 25230 31602 25282 31614
rect 27358 31666 27410 31678
rect 33518 31666 33570 31678
rect 31154 31614 31166 31666
rect 31218 31614 31230 31666
rect 31490 31614 31502 31666
rect 31554 31614 31566 31666
rect 27358 31602 27410 31614
rect 33518 31602 33570 31614
rect 34190 31666 34242 31678
rect 35310 31666 35362 31678
rect 35870 31666 35922 31678
rect 44942 31666 44994 31678
rect 34290 31614 34302 31666
rect 34354 31614 34366 31666
rect 35634 31614 35646 31666
rect 35698 31614 35710 31666
rect 37762 31614 37774 31666
rect 37826 31614 37838 31666
rect 34190 31602 34242 31614
rect 35310 31602 35362 31614
rect 35870 31602 35922 31614
rect 44942 31602 44994 31614
rect 45950 31666 46002 31678
rect 45950 31602 46002 31614
rect 46062 31666 46114 31678
rect 46062 31602 46114 31614
rect 46510 31666 46562 31678
rect 46510 31602 46562 31614
rect 47070 31666 47122 31678
rect 47070 31602 47122 31614
rect 47182 31666 47234 31678
rect 49634 31614 49646 31666
rect 49698 31614 49710 31666
rect 54338 31614 54350 31666
rect 54402 31614 54414 31666
rect 47182 31602 47234 31614
rect 6862 31554 6914 31566
rect 6514 31502 6526 31554
rect 6578 31502 6590 31554
rect 6862 31490 6914 31502
rect 7086 31554 7138 31566
rect 7086 31490 7138 31502
rect 7310 31554 7362 31566
rect 7310 31490 7362 31502
rect 9326 31554 9378 31566
rect 9326 31490 9378 31502
rect 10222 31554 10274 31566
rect 10222 31490 10274 31502
rect 14814 31554 14866 31566
rect 14814 31490 14866 31502
rect 17054 31554 17106 31566
rect 17054 31490 17106 31502
rect 17950 31554 18002 31566
rect 17950 31490 18002 31502
rect 18062 31554 18114 31566
rect 18062 31490 18114 31502
rect 20302 31554 20354 31566
rect 20302 31490 20354 31502
rect 20750 31554 20802 31566
rect 20750 31490 20802 31502
rect 21310 31554 21362 31566
rect 23102 31554 23154 31566
rect 21634 31502 21646 31554
rect 21698 31502 21710 31554
rect 21310 31490 21362 31502
rect 23102 31490 23154 31502
rect 24782 31554 24834 31566
rect 32846 31554 32898 31566
rect 28578 31502 28590 31554
rect 28642 31502 28654 31554
rect 29586 31502 29598 31554
rect 29650 31502 29662 31554
rect 24782 31490 24834 31502
rect 32846 31490 32898 31502
rect 33406 31554 33458 31566
rect 33406 31490 33458 31502
rect 34078 31554 34130 31566
rect 34078 31490 34130 31502
rect 45726 31554 45778 31566
rect 45726 31490 45778 31502
rect 46286 31554 46338 31566
rect 46286 31490 46338 31502
rect 47406 31554 47458 31566
rect 47618 31502 47630 31554
rect 47682 31502 47694 31554
rect 52882 31502 52894 31554
rect 52946 31502 52958 31554
rect 47406 31490 47458 31502
rect 1344 31386 58576 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 50558 31386
rect 50610 31334 50662 31386
rect 50714 31334 50766 31386
rect 50818 31334 58576 31386
rect 1344 31300 58576 31334
rect 8094 31218 8146 31230
rect 8094 31154 8146 31166
rect 8878 31218 8930 31230
rect 21198 31218 21250 31230
rect 9762 31166 9774 31218
rect 9826 31166 9838 31218
rect 8878 31154 8930 31166
rect 21198 31154 21250 31166
rect 21310 31218 21362 31230
rect 21310 31154 21362 31166
rect 22094 31218 22146 31230
rect 22094 31154 22146 31166
rect 22318 31218 22370 31230
rect 22318 31154 22370 31166
rect 26574 31218 26626 31230
rect 32958 31218 33010 31230
rect 26898 31166 26910 31218
rect 26962 31166 26974 31218
rect 26574 31154 26626 31166
rect 32958 31154 33010 31166
rect 35982 31218 36034 31230
rect 35982 31154 36034 31166
rect 36430 31218 36482 31230
rect 36430 31154 36482 31166
rect 37550 31218 37602 31230
rect 37550 31154 37602 31166
rect 38558 31218 38610 31230
rect 38558 31154 38610 31166
rect 38670 31218 38722 31230
rect 38670 31154 38722 31166
rect 48974 31218 49026 31230
rect 48974 31154 49026 31166
rect 49310 31218 49362 31230
rect 49310 31154 49362 31166
rect 54798 31218 54850 31230
rect 54798 31154 54850 31166
rect 2606 31106 2658 31118
rect 2370 31054 2382 31106
rect 2434 31054 2446 31106
rect 2606 31042 2658 31054
rect 6750 31106 6802 31118
rect 12462 31106 12514 31118
rect 10210 31054 10222 31106
rect 10274 31054 10286 31106
rect 6750 31042 6802 31054
rect 12462 31042 12514 31054
rect 21086 31106 21138 31118
rect 23998 31106 24050 31118
rect 23650 31054 23662 31106
rect 23714 31054 23726 31106
rect 21086 31042 21138 31054
rect 23998 31042 24050 31054
rect 24558 31106 24610 31118
rect 24558 31042 24610 31054
rect 25230 31106 25282 31118
rect 25230 31042 25282 31054
rect 25342 31106 25394 31118
rect 39230 31106 39282 31118
rect 44494 31106 44546 31118
rect 25442 31054 25454 31106
rect 25506 31054 25518 31106
rect 34178 31054 34190 31106
rect 34242 31054 34254 31106
rect 35186 31054 35198 31106
rect 35250 31054 35262 31106
rect 35634 31054 35646 31106
rect 35698 31054 35710 31106
rect 42466 31054 42478 31106
rect 42530 31054 42542 31106
rect 43138 31054 43150 31106
rect 43202 31054 43214 31106
rect 25342 31042 25394 31054
rect 39230 31042 39282 31054
rect 44494 31042 44546 31054
rect 45838 31106 45890 31118
rect 45838 31042 45890 31054
rect 46846 31106 46898 31118
rect 46846 31042 46898 31054
rect 48750 31106 48802 31118
rect 48750 31042 48802 31054
rect 49198 31106 49250 31118
rect 49198 31042 49250 31054
rect 49534 31106 49586 31118
rect 51090 31054 51102 31106
rect 51154 31054 51166 31106
rect 49534 31042 49586 31054
rect 3054 30994 3106 31006
rect 5630 30994 5682 31006
rect 3490 30942 3502 30994
rect 3554 30942 3566 30994
rect 4498 30942 4510 30994
rect 4562 30942 4574 30994
rect 3054 30930 3106 30942
rect 5630 30930 5682 30942
rect 5854 30994 5906 31006
rect 5854 30930 5906 30942
rect 6078 30994 6130 31006
rect 6078 30930 6130 30942
rect 6526 30994 6578 31006
rect 8542 30994 8594 31006
rect 7074 30942 7086 30994
rect 7138 30942 7150 30994
rect 7634 30942 7646 30994
rect 7698 30942 7710 30994
rect 7858 30942 7870 30994
rect 7922 30942 7934 30994
rect 6526 30930 6578 30942
rect 8542 30930 8594 30942
rect 8766 30994 8818 31006
rect 16606 30994 16658 31006
rect 21422 30994 21474 31006
rect 8978 30942 8990 30994
rect 9042 30942 9054 30994
rect 9538 30942 9550 30994
rect 9602 30942 9614 30994
rect 10658 30942 10670 30994
rect 10722 30942 10734 30994
rect 11778 30942 11790 30994
rect 11842 30942 11854 30994
rect 16146 30942 16158 30994
rect 16210 30942 16222 30994
rect 20178 30942 20190 30994
rect 20242 30942 20254 30994
rect 20626 30942 20638 30994
rect 20690 30942 20702 30994
rect 8766 30930 8818 30942
rect 16606 30930 16658 30942
rect 21422 30930 21474 30942
rect 21646 30994 21698 31006
rect 21646 30930 21698 30942
rect 22990 30994 23042 31006
rect 22990 30930 23042 30942
rect 23326 30994 23378 31006
rect 23326 30930 23378 30942
rect 24334 30994 24386 31006
rect 38222 30994 38274 31006
rect 26002 30942 26014 30994
rect 26066 30942 26078 30994
rect 27234 30942 27246 30994
rect 27298 30942 27310 30994
rect 33058 30942 33070 30994
rect 33122 30942 33134 30994
rect 34066 30942 34078 30994
rect 34130 30942 34142 30994
rect 35074 30942 35086 30994
rect 35138 30942 35150 30994
rect 37314 30942 37326 30994
rect 37378 30942 37390 30994
rect 24334 30930 24386 30942
rect 38222 30930 38274 30942
rect 38446 30994 38498 31006
rect 38446 30930 38498 30942
rect 39118 30994 39170 31006
rect 42814 30994 42866 31006
rect 41346 30942 41358 30994
rect 41410 30942 41422 30994
rect 42242 30942 42254 30994
rect 42306 30942 42318 30994
rect 39118 30930 39170 30942
rect 42814 30930 42866 30942
rect 44382 30994 44434 31006
rect 44382 30930 44434 30942
rect 44606 30994 44658 31006
rect 44606 30930 44658 30942
rect 45054 30994 45106 31006
rect 45054 30930 45106 30942
rect 46286 30994 46338 31006
rect 46286 30930 46338 30942
rect 46622 30994 46674 31006
rect 48078 30994 48130 31006
rect 53006 30994 53058 31006
rect 54350 30994 54402 31006
rect 47618 30942 47630 30994
rect 47682 30942 47694 30994
rect 50194 30942 50206 30994
rect 50258 30942 50270 30994
rect 52658 30942 52670 30994
rect 52722 30942 52734 30994
rect 53778 30942 53790 30994
rect 53842 30942 53854 30994
rect 54114 30942 54126 30994
rect 54178 30942 54190 30994
rect 46622 30930 46674 30942
rect 48078 30930 48130 30942
rect 53006 30930 53058 30942
rect 54350 30930 54402 30942
rect 2270 30882 2322 30894
rect 2270 30818 2322 30830
rect 3278 30882 3330 30894
rect 5406 30882 5458 30894
rect 22206 30882 22258 30894
rect 3714 30830 3726 30882
rect 3778 30830 3790 30882
rect 4050 30830 4062 30882
rect 4114 30830 4126 30882
rect 12114 30830 12126 30882
rect 12178 30830 12190 30882
rect 13234 30830 13246 30882
rect 13298 30830 13310 30882
rect 15362 30830 15374 30882
rect 15426 30830 15438 30882
rect 17378 30830 17390 30882
rect 17442 30830 17454 30882
rect 19506 30830 19518 30882
rect 19570 30830 19582 30882
rect 3278 30818 3330 30830
rect 5406 30818 5458 30830
rect 22206 30818 22258 30830
rect 24110 30882 24162 30894
rect 39678 30882 39730 30894
rect 31826 30830 31838 30882
rect 31890 30830 31902 30882
rect 36306 30830 36318 30882
rect 36370 30830 36382 30882
rect 24110 30818 24162 30830
rect 39678 30818 39730 30830
rect 41022 30882 41074 30894
rect 46398 30882 46450 30894
rect 42354 30830 42366 30882
rect 42418 30830 42430 30882
rect 41022 30818 41074 30830
rect 46398 30818 46450 30830
rect 47182 30882 47234 30894
rect 51650 30830 51662 30882
rect 51714 30830 51726 30882
rect 54674 30830 54686 30882
rect 54738 30830 54750 30882
rect 47182 30818 47234 30830
rect 7086 30770 7138 30782
rect 7086 30706 7138 30718
rect 8206 30770 8258 30782
rect 36654 30770 36706 30782
rect 25778 30718 25790 30770
rect 25842 30718 25854 30770
rect 8206 30706 8258 30718
rect 36654 30706 36706 30718
rect 37662 30770 37714 30782
rect 37662 30706 37714 30718
rect 37998 30770 38050 30782
rect 37998 30706 38050 30718
rect 45278 30770 45330 30782
rect 45278 30706 45330 30718
rect 45614 30770 45666 30782
rect 55022 30770 55074 30782
rect 52546 30718 52558 30770
rect 52610 30718 52622 30770
rect 45614 30706 45666 30718
rect 55022 30706 55074 30718
rect 1344 30602 58576 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 58576 30602
rect 1344 30516 58576 30550
rect 16046 30434 16098 30446
rect 9986 30382 9998 30434
rect 10050 30382 10062 30434
rect 16046 30370 16098 30382
rect 19406 30434 19458 30446
rect 19406 30370 19458 30382
rect 28254 30434 28306 30446
rect 28254 30370 28306 30382
rect 31502 30434 31554 30446
rect 57934 30434 57986 30446
rect 45154 30382 45166 30434
rect 45218 30382 45230 30434
rect 31502 30370 31554 30382
rect 57934 30370 57986 30382
rect 26350 30322 26402 30334
rect 5954 30270 5966 30322
rect 6018 30270 6030 30322
rect 9650 30270 9662 30322
rect 9714 30270 9726 30322
rect 12450 30270 12462 30322
rect 12514 30270 12526 30322
rect 26350 30258 26402 30270
rect 28478 30322 28530 30334
rect 31838 30322 31890 30334
rect 37998 30322 38050 30334
rect 43374 30322 43426 30334
rect 29586 30270 29598 30322
rect 29650 30270 29662 30322
rect 37650 30270 37662 30322
rect 37714 30270 37726 30322
rect 42690 30270 42702 30322
rect 42754 30270 42766 30322
rect 28478 30258 28530 30270
rect 31838 30258 31890 30270
rect 37998 30258 38050 30270
rect 43374 30258 43426 30270
rect 43598 30322 43650 30334
rect 52670 30322 52722 30334
rect 43922 30270 43934 30322
rect 43986 30270 43998 30322
rect 45602 30270 45614 30322
rect 45666 30270 45678 30322
rect 51202 30270 51214 30322
rect 51266 30270 51278 30322
rect 54786 30270 54798 30322
rect 54850 30270 54862 30322
rect 43598 30258 43650 30270
rect 52670 30258 52722 30270
rect 4622 30210 4674 30222
rect 15710 30210 15762 30222
rect 26798 30210 26850 30222
rect 4274 30158 4286 30210
rect 4338 30158 4350 30210
rect 7410 30158 7422 30210
rect 7474 30158 7486 30210
rect 8978 30158 8990 30210
rect 9042 30158 9054 30210
rect 10098 30158 10110 30210
rect 10162 30158 10174 30210
rect 10882 30158 10894 30210
rect 10946 30158 10958 30210
rect 11442 30158 11454 30210
rect 11506 30158 11518 30210
rect 14466 30158 14478 30210
rect 14530 30158 14542 30210
rect 16818 30158 16830 30210
rect 16882 30158 16894 30210
rect 18274 30158 18286 30210
rect 18338 30158 18350 30210
rect 20178 30158 20190 30210
rect 20242 30158 20254 30210
rect 24546 30158 24558 30210
rect 24610 30158 24622 30210
rect 4622 30146 4674 30158
rect 15710 30146 15762 30158
rect 26798 30146 26850 30158
rect 27358 30210 27410 30222
rect 27358 30146 27410 30158
rect 28030 30210 28082 30222
rect 28030 30146 28082 30158
rect 29486 30210 29538 30222
rect 29486 30146 29538 30158
rect 30494 30210 30546 30222
rect 36318 30210 36370 30222
rect 39566 30210 39618 30222
rect 44270 30210 44322 30222
rect 46286 30210 46338 30222
rect 32274 30158 32286 30210
rect 32338 30158 32350 30210
rect 33282 30158 33294 30210
rect 33346 30158 33358 30210
rect 34514 30158 34526 30210
rect 34578 30158 34590 30210
rect 35298 30158 35310 30210
rect 35362 30158 35374 30210
rect 37202 30158 37214 30210
rect 37266 30158 37278 30210
rect 39778 30158 39790 30210
rect 39842 30158 39854 30210
rect 40562 30158 40574 30210
rect 40626 30158 40638 30210
rect 45714 30158 45726 30210
rect 45778 30158 45790 30210
rect 30494 30146 30546 30158
rect 36318 30146 36370 30158
rect 39566 30146 39618 30158
rect 44270 30146 44322 30158
rect 46286 30146 46338 30158
rect 47182 30210 47234 30222
rect 50318 30210 50370 30222
rect 47730 30158 47742 30210
rect 47794 30158 47806 30210
rect 48962 30158 48974 30210
rect 49026 30158 49038 30210
rect 49970 30158 49982 30210
rect 50034 30158 50046 30210
rect 50978 30158 50990 30210
rect 51042 30158 51054 30210
rect 53330 30158 53342 30210
rect 53394 30158 53406 30210
rect 55570 30158 55582 30210
rect 55634 30158 55646 30210
rect 47182 30146 47234 30158
rect 50318 30146 50370 30158
rect 8094 30098 8146 30110
rect 2482 30046 2494 30098
rect 2546 30046 2558 30098
rect 4946 30046 4958 30098
rect 5010 30046 5022 30098
rect 6514 30046 6526 30098
rect 6578 30046 6590 30098
rect 8094 30034 8146 30046
rect 14702 30098 14754 30110
rect 14702 30034 14754 30046
rect 15374 30098 15426 30110
rect 18510 30098 18562 30110
rect 16594 30046 16606 30098
rect 16658 30046 16670 30098
rect 15374 30034 15426 30046
rect 18510 30034 18562 30046
rect 19070 30098 19122 30110
rect 27582 30098 27634 30110
rect 20066 30046 20078 30098
rect 20130 30046 20142 30098
rect 23874 30046 23886 30098
rect 23938 30046 23950 30098
rect 19070 30034 19122 30046
rect 27582 30034 27634 30046
rect 30830 30098 30882 30110
rect 30830 30034 30882 30046
rect 31278 30098 31330 30110
rect 31278 30034 31330 30046
rect 32510 30098 32562 30110
rect 37774 30098 37826 30110
rect 47070 30098 47122 30110
rect 34402 30046 34414 30098
rect 34466 30046 34478 30098
rect 34962 30046 34974 30098
rect 35026 30046 35038 30098
rect 38546 30046 38558 30098
rect 38610 30046 38622 30098
rect 49858 30046 49870 30098
rect 49922 30046 49934 30098
rect 54226 30046 54238 30098
rect 54290 30046 54302 30098
rect 32510 30034 32562 30046
rect 37774 30034 37826 30046
rect 47070 30034 47122 30046
rect 20750 29986 20802 29998
rect 25230 29986 25282 29998
rect 29822 29986 29874 29998
rect 35758 29986 35810 29998
rect 38894 29986 38946 29998
rect 44046 29986 44098 29998
rect 21634 29934 21646 29986
rect 21698 29934 21710 29986
rect 25554 29934 25566 29986
rect 25618 29934 25630 29986
rect 27010 29934 27022 29986
rect 27074 29934 27086 29986
rect 34290 29934 34302 29986
rect 34354 29934 34366 29986
rect 36978 29934 36990 29986
rect 37042 29934 37054 29986
rect 43026 29934 43038 29986
rect 43090 29934 43102 29986
rect 20750 29922 20802 29934
rect 25230 29922 25282 29934
rect 29822 29922 29874 29934
rect 35758 29922 35810 29934
rect 38894 29922 38946 29934
rect 44046 29922 44098 29934
rect 46398 29986 46450 29998
rect 46398 29922 46450 29934
rect 46622 29986 46674 29998
rect 48962 29934 48974 29986
rect 49026 29934 49038 29986
rect 46622 29922 46674 29934
rect 1344 29818 58576 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 50558 29818
rect 50610 29766 50662 29818
rect 50714 29766 50766 29818
rect 50818 29766 58576 29818
rect 1344 29732 58576 29766
rect 7758 29650 7810 29662
rect 20078 29650 20130 29662
rect 8978 29598 8990 29650
rect 9042 29598 9054 29650
rect 7758 29586 7810 29598
rect 20078 29586 20130 29598
rect 23214 29650 23266 29662
rect 23214 29586 23266 29598
rect 23662 29650 23714 29662
rect 23662 29586 23714 29598
rect 24222 29650 24274 29662
rect 24222 29586 24274 29598
rect 24782 29650 24834 29662
rect 24782 29586 24834 29598
rect 25454 29650 25506 29662
rect 25454 29586 25506 29598
rect 28590 29650 28642 29662
rect 28590 29586 28642 29598
rect 28702 29650 28754 29662
rect 30046 29650 30098 29662
rect 29138 29598 29150 29650
rect 29202 29598 29214 29650
rect 28702 29586 28754 29598
rect 30046 29586 30098 29598
rect 31950 29650 32002 29662
rect 37998 29650 38050 29662
rect 32274 29598 32286 29650
rect 32338 29598 32350 29650
rect 34626 29598 34638 29650
rect 34690 29598 34702 29650
rect 31950 29586 32002 29598
rect 37998 29586 38050 29598
rect 40350 29650 40402 29662
rect 40350 29586 40402 29598
rect 40798 29650 40850 29662
rect 40798 29586 40850 29598
rect 45838 29650 45890 29662
rect 45838 29586 45890 29598
rect 46062 29650 46114 29662
rect 46062 29586 46114 29598
rect 7534 29538 7586 29550
rect 7534 29474 7586 29486
rect 8318 29538 8370 29550
rect 8318 29474 8370 29486
rect 14590 29538 14642 29550
rect 20302 29538 20354 29550
rect 16706 29486 16718 29538
rect 16770 29486 16782 29538
rect 14590 29474 14642 29486
rect 20302 29474 20354 29486
rect 20862 29538 20914 29550
rect 20862 29474 20914 29486
rect 22206 29538 22258 29550
rect 22206 29474 22258 29486
rect 23550 29538 23602 29550
rect 23550 29474 23602 29486
rect 26014 29538 26066 29550
rect 26014 29474 26066 29486
rect 26798 29538 26850 29550
rect 26798 29474 26850 29486
rect 30382 29538 30434 29550
rect 37550 29538 37602 29550
rect 44606 29538 44658 29550
rect 34738 29486 34750 29538
rect 34802 29486 34814 29538
rect 35522 29486 35534 29538
rect 35586 29486 35598 29538
rect 35970 29486 35982 29538
rect 36034 29486 36046 29538
rect 37314 29486 37326 29538
rect 37378 29486 37390 29538
rect 42018 29486 42030 29538
rect 42082 29486 42094 29538
rect 42690 29486 42702 29538
rect 42754 29486 42766 29538
rect 30382 29474 30434 29486
rect 37550 29474 37602 29486
rect 44606 29474 44658 29486
rect 46174 29538 46226 29550
rect 46174 29474 46226 29486
rect 5294 29426 5346 29438
rect 6414 29426 6466 29438
rect 7422 29426 7474 29438
rect 4274 29374 4286 29426
rect 4338 29374 4350 29426
rect 5506 29374 5518 29426
rect 5570 29374 5582 29426
rect 6626 29374 6638 29426
rect 6690 29374 6702 29426
rect 5294 29362 5346 29374
rect 6414 29362 6466 29374
rect 7422 29362 7474 29374
rect 7870 29426 7922 29438
rect 7870 29362 7922 29374
rect 8430 29426 8482 29438
rect 8430 29362 8482 29374
rect 8542 29426 8594 29438
rect 15598 29426 15650 29438
rect 21534 29426 21586 29438
rect 14354 29374 14366 29426
rect 14418 29374 14430 29426
rect 16594 29374 16606 29426
rect 16658 29374 16670 29426
rect 21298 29374 21310 29426
rect 21362 29374 21374 29426
rect 8542 29362 8594 29374
rect 15598 29362 15650 29374
rect 21534 29362 21586 29374
rect 22542 29426 22594 29438
rect 22542 29362 22594 29374
rect 22878 29426 22930 29438
rect 26350 29426 26402 29438
rect 25778 29374 25790 29426
rect 25842 29374 25854 29426
rect 22878 29362 22930 29374
rect 26350 29362 26402 29374
rect 26574 29426 26626 29438
rect 26574 29362 26626 29374
rect 27134 29426 27186 29438
rect 27134 29362 27186 29374
rect 27582 29426 27634 29438
rect 27582 29362 27634 29374
rect 27806 29426 27858 29438
rect 27806 29362 27858 29374
rect 28030 29426 28082 29438
rect 28030 29362 28082 29374
rect 28478 29426 28530 29438
rect 31614 29426 31666 29438
rect 37102 29426 37154 29438
rect 29362 29374 29374 29426
rect 29426 29374 29438 29426
rect 30594 29374 30606 29426
rect 30658 29374 30670 29426
rect 33394 29374 33406 29426
rect 33458 29374 33470 29426
rect 34626 29374 34638 29426
rect 34690 29374 34702 29426
rect 35298 29374 35310 29426
rect 35362 29374 35374 29426
rect 36194 29374 36206 29426
rect 36258 29374 36270 29426
rect 36754 29374 36766 29426
rect 36818 29374 36830 29426
rect 28478 29362 28530 29374
rect 31614 29362 31666 29374
rect 37102 29362 37154 29374
rect 37886 29426 37938 29438
rect 37886 29362 37938 29374
rect 38110 29426 38162 29438
rect 38110 29362 38162 29374
rect 38558 29426 38610 29438
rect 45502 29426 45554 29438
rect 40898 29374 40910 29426
rect 40962 29374 40974 29426
rect 41906 29374 41918 29426
rect 41970 29374 41982 29426
rect 42802 29374 42814 29426
rect 42866 29374 42878 29426
rect 45266 29374 45278 29426
rect 45330 29374 45342 29426
rect 38558 29362 38610 29374
rect 45502 29362 45554 29374
rect 15934 29314 15986 29326
rect 15934 29250 15986 29262
rect 18174 29314 18226 29326
rect 18174 29250 18226 29262
rect 19630 29314 19682 29326
rect 19630 29250 19682 29262
rect 26462 29314 26514 29326
rect 26462 29250 26514 29262
rect 27694 29314 27746 29326
rect 37438 29314 37490 29326
rect 31154 29262 31166 29314
rect 31218 29262 31230 29314
rect 27694 29250 27746 29262
rect 37438 29250 37490 29262
rect 39902 29314 39954 29326
rect 39902 29250 39954 29262
rect 1934 29202 1986 29214
rect 21758 29202 21810 29214
rect 6626 29150 6638 29202
rect 6690 29150 6702 29202
rect 1934 29138 1986 29150
rect 21758 29138 21810 29150
rect 21870 29202 21922 29214
rect 21870 29138 21922 29150
rect 1344 29034 58576 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 58576 29034
rect 1344 28948 58576 28982
rect 5630 28866 5682 28878
rect 5630 28802 5682 28814
rect 5966 28866 6018 28878
rect 5966 28802 6018 28814
rect 17390 28866 17442 28878
rect 17390 28802 17442 28814
rect 28478 28866 28530 28878
rect 41234 28814 41246 28866
rect 41298 28814 41310 28866
rect 28478 28802 28530 28814
rect 19070 28754 19122 28766
rect 20750 28754 20802 28766
rect 36430 28754 36482 28766
rect 2258 28702 2270 28754
rect 2322 28702 2334 28754
rect 13458 28702 13470 28754
rect 13522 28702 13534 28754
rect 15586 28702 15598 28754
rect 15650 28702 15662 28754
rect 19618 28702 19630 28754
rect 19682 28702 19694 28754
rect 29250 28702 29262 28754
rect 29314 28702 29326 28754
rect 31154 28702 31166 28754
rect 31218 28702 31230 28754
rect 19070 28690 19122 28702
rect 20750 28690 20802 28702
rect 36430 28690 36482 28702
rect 49758 28754 49810 28766
rect 49758 28690 49810 28702
rect 57934 28754 57986 28766
rect 57934 28690 57986 28702
rect 1934 28642 1986 28654
rect 1934 28578 1986 28590
rect 2718 28642 2770 28654
rect 2718 28578 2770 28590
rect 3054 28642 3106 28654
rect 17054 28642 17106 28654
rect 27694 28642 27746 28654
rect 30046 28642 30098 28654
rect 31614 28642 31666 28654
rect 16370 28590 16382 28642
rect 16434 28590 16446 28642
rect 17938 28590 17950 28642
rect 18002 28590 18014 28642
rect 26674 28590 26686 28642
rect 26738 28590 26750 28642
rect 28018 28590 28030 28642
rect 28082 28590 28094 28642
rect 29586 28590 29598 28642
rect 29650 28590 29662 28642
rect 30818 28590 30830 28642
rect 30882 28590 30894 28642
rect 3054 28578 3106 28590
rect 17054 28578 17106 28590
rect 27694 28578 27746 28590
rect 30046 28578 30098 28590
rect 31614 28578 31666 28590
rect 32174 28642 32226 28654
rect 32174 28578 32226 28590
rect 32510 28642 32562 28654
rect 32510 28578 32562 28590
rect 33294 28642 33346 28654
rect 33294 28578 33346 28590
rect 34526 28642 34578 28654
rect 34526 28578 34578 28590
rect 35086 28642 35138 28654
rect 35086 28578 35138 28590
rect 35310 28642 35362 28654
rect 35310 28578 35362 28590
rect 35982 28642 36034 28654
rect 35982 28578 36034 28590
rect 36990 28642 37042 28654
rect 36990 28578 37042 28590
rect 37662 28642 37714 28654
rect 37662 28578 37714 28590
rect 38670 28642 38722 28654
rect 38670 28578 38722 28590
rect 40350 28642 40402 28654
rect 42254 28642 42306 28654
rect 42926 28642 42978 28654
rect 41010 28590 41022 28642
rect 41074 28590 41086 28642
rect 41570 28590 41582 28642
rect 41634 28590 41646 28642
rect 42690 28590 42702 28642
rect 42754 28590 42766 28642
rect 40350 28578 40402 28590
rect 42254 28578 42306 28590
rect 42926 28578 42978 28590
rect 43710 28642 43762 28654
rect 50654 28642 50706 28654
rect 50306 28590 50318 28642
rect 50370 28590 50382 28642
rect 43710 28578 43762 28590
rect 50654 28578 50706 28590
rect 51102 28642 51154 28654
rect 51998 28642 52050 28654
rect 51762 28590 51774 28642
rect 51826 28590 51838 28642
rect 55570 28590 55582 28642
rect 55634 28590 55646 28642
rect 51102 28578 51154 28590
rect 51998 28578 52050 28590
rect 5854 28530 5906 28542
rect 19294 28530 19346 28542
rect 18050 28478 18062 28530
rect 18114 28478 18126 28530
rect 5854 28466 5906 28478
rect 19294 28466 19346 28478
rect 19518 28530 19570 28542
rect 27470 28530 27522 28542
rect 22082 28478 22094 28530
rect 22146 28478 22158 28530
rect 19518 28466 19570 28478
rect 27470 28466 27522 28478
rect 28366 28530 28418 28542
rect 34974 28530 35026 28542
rect 37998 28530 38050 28542
rect 33618 28478 33630 28530
rect 33682 28478 33694 28530
rect 37314 28478 37326 28530
rect 37378 28478 37390 28530
rect 28366 28466 28418 28478
rect 34974 28466 35026 28478
rect 37998 28466 38050 28478
rect 39342 28530 39394 28542
rect 39342 28466 39394 28478
rect 41806 28530 41858 28542
rect 41806 28466 41858 28478
rect 43150 28530 43202 28542
rect 43150 28466 43202 28478
rect 43262 28530 43314 28542
rect 43262 28466 43314 28478
rect 3390 28418 3442 28430
rect 3390 28354 3442 28366
rect 20190 28418 20242 28430
rect 20190 28354 20242 28366
rect 27582 28418 27634 28430
rect 27582 28354 27634 28366
rect 28478 28418 28530 28430
rect 28478 28354 28530 28366
rect 30382 28418 30434 28430
rect 30382 28354 30434 28366
rect 32846 28418 32898 28430
rect 32846 28354 32898 28366
rect 33966 28418 34018 28430
rect 33966 28354 34018 28366
rect 34750 28418 34802 28430
rect 34750 28354 34802 28366
rect 35758 28418 35810 28430
rect 35758 28354 35810 28366
rect 35870 28418 35922 28430
rect 35870 28354 35922 28366
rect 38558 28418 38610 28430
rect 38558 28354 38610 28366
rect 39118 28418 39170 28430
rect 39118 28354 39170 28366
rect 39230 28418 39282 28430
rect 39230 28354 39282 28366
rect 39902 28418 39954 28430
rect 39902 28354 39954 28366
rect 40798 28418 40850 28430
rect 40798 28354 40850 28366
rect 41694 28418 41746 28430
rect 41694 28354 41746 28366
rect 42142 28418 42194 28430
rect 42142 28354 42194 28366
rect 42366 28418 42418 28430
rect 42366 28354 42418 28366
rect 1344 28250 58576 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 50558 28250
rect 50610 28198 50662 28250
rect 50714 28198 50766 28250
rect 50818 28198 58576 28250
rect 1344 28164 58576 28198
rect 2046 28082 2098 28094
rect 2046 28018 2098 28030
rect 2718 28082 2770 28094
rect 2718 28018 2770 28030
rect 3614 28082 3666 28094
rect 3614 28018 3666 28030
rect 18062 28082 18114 28094
rect 18062 28018 18114 28030
rect 18510 28082 18562 28094
rect 18510 28018 18562 28030
rect 18734 28082 18786 28094
rect 22430 28082 22482 28094
rect 21634 28030 21646 28082
rect 21698 28030 21710 28082
rect 18734 28018 18786 28030
rect 22430 28018 22482 28030
rect 23326 28082 23378 28094
rect 23326 28018 23378 28030
rect 25566 28082 25618 28094
rect 25566 28018 25618 28030
rect 33294 28082 33346 28094
rect 36654 28082 36706 28094
rect 33618 28030 33630 28082
rect 33682 28030 33694 28082
rect 35410 28030 35422 28082
rect 35474 28030 35486 28082
rect 33294 28018 33346 28030
rect 36654 28018 36706 28030
rect 37102 28082 37154 28094
rect 37102 28018 37154 28030
rect 37326 28082 37378 28094
rect 37326 28018 37378 28030
rect 39230 28082 39282 28094
rect 39230 28018 39282 28030
rect 39342 28082 39394 28094
rect 39342 28018 39394 28030
rect 39790 28082 39842 28094
rect 39790 28018 39842 28030
rect 40014 28082 40066 28094
rect 52658 28030 52670 28082
rect 52722 28030 52734 28082
rect 40014 28018 40066 28030
rect 16270 27970 16322 27982
rect 16270 27906 16322 27918
rect 16606 27970 16658 27982
rect 16606 27906 16658 27918
rect 17614 27970 17666 27982
rect 22206 27970 22258 27982
rect 19058 27918 19070 27970
rect 19122 27918 19134 27970
rect 20290 27918 20302 27970
rect 20354 27918 20366 27970
rect 21746 27918 21758 27970
rect 21810 27918 21822 27970
rect 17614 27906 17666 27918
rect 22206 27906 22258 27918
rect 22654 27970 22706 27982
rect 24110 27970 24162 27982
rect 38446 27970 38498 27982
rect 44494 27970 44546 27982
rect 23650 27918 23662 27970
rect 23714 27918 23726 27970
rect 29362 27918 29374 27970
rect 29426 27918 29438 27970
rect 35186 27918 35198 27970
rect 35250 27918 35262 27970
rect 35858 27918 35870 27970
rect 35922 27918 35934 27970
rect 41682 27918 41694 27970
rect 41746 27918 41758 27970
rect 22654 27906 22706 27918
rect 24110 27906 24162 27918
rect 38446 27906 38498 27918
rect 44494 27906 44546 27918
rect 48750 27970 48802 27982
rect 53218 27918 53230 27970
rect 53282 27918 53294 27970
rect 48750 27906 48802 27918
rect 2382 27858 2434 27870
rect 1810 27806 1822 27858
rect 1874 27806 1886 27858
rect 2382 27794 2434 27806
rect 18398 27858 18450 27870
rect 18398 27794 18450 27806
rect 19294 27858 19346 27870
rect 23886 27858 23938 27870
rect 19618 27806 19630 27858
rect 19682 27806 19694 27858
rect 20178 27806 20190 27858
rect 20242 27806 20254 27858
rect 21186 27806 21198 27858
rect 21250 27806 21262 27858
rect 19294 27794 19346 27806
rect 23886 27794 23938 27806
rect 24222 27858 24274 27870
rect 24222 27794 24274 27806
rect 25678 27858 25730 27870
rect 30046 27858 30098 27870
rect 26114 27806 26126 27858
rect 26178 27806 26190 27858
rect 29586 27806 29598 27858
rect 29650 27806 29662 27858
rect 25678 27794 25730 27806
rect 30046 27794 30098 27806
rect 30942 27858 30994 27870
rect 37774 27858 37826 27870
rect 33954 27806 33966 27858
rect 34018 27806 34030 27858
rect 34962 27806 34974 27858
rect 35026 27806 35038 27858
rect 35970 27806 35982 27858
rect 36034 27806 36046 27858
rect 30942 27794 30994 27806
rect 37774 27794 37826 27806
rect 38222 27858 38274 27870
rect 38222 27794 38274 27806
rect 38558 27858 38610 27870
rect 38558 27794 38610 27806
rect 38782 27858 38834 27870
rect 38782 27794 38834 27806
rect 39454 27858 39506 27870
rect 39454 27794 39506 27806
rect 40462 27858 40514 27870
rect 40898 27806 40910 27858
rect 40962 27806 40974 27858
rect 45154 27806 45166 27858
rect 45218 27806 45230 27858
rect 46274 27806 46286 27858
rect 46338 27806 46350 27858
rect 47954 27806 47966 27858
rect 48018 27806 48030 27858
rect 49186 27806 49198 27858
rect 49250 27806 49262 27858
rect 50978 27806 50990 27858
rect 51042 27806 51054 27858
rect 51202 27806 51214 27858
rect 51266 27806 51278 27858
rect 51874 27806 51886 27858
rect 51938 27806 51950 27858
rect 52546 27806 52558 27858
rect 52610 27806 52622 27858
rect 53106 27806 53118 27858
rect 53170 27806 53182 27858
rect 40462 27794 40514 27806
rect 3166 27746 3218 27758
rect 3166 27682 3218 27694
rect 18958 27746 19010 27758
rect 24670 27746 24722 27758
rect 30606 27746 30658 27758
rect 32510 27746 32562 27758
rect 22530 27694 22542 27746
rect 22594 27694 22606 27746
rect 26786 27694 26798 27746
rect 26850 27694 26862 27746
rect 28914 27694 28926 27746
rect 28978 27694 28990 27746
rect 31378 27694 31390 27746
rect 31442 27694 31454 27746
rect 18958 27682 19010 27694
rect 24670 27682 24722 27694
rect 30606 27682 30658 27694
rect 32510 27682 32562 27694
rect 37214 27746 37266 27758
rect 37214 27682 37266 27694
rect 39902 27746 39954 27758
rect 57598 27746 57650 27758
rect 43810 27694 43822 27746
rect 43874 27694 43886 27746
rect 45378 27694 45390 27746
rect 45442 27694 45454 27746
rect 47618 27694 47630 27746
rect 47682 27694 47694 27746
rect 49074 27694 49086 27746
rect 49138 27694 49150 27746
rect 52098 27694 52110 27746
rect 52162 27694 52174 27746
rect 39902 27682 39954 27694
rect 57598 27682 57650 27694
rect 19966 27634 20018 27646
rect 19966 27570 20018 27582
rect 25566 27634 25618 27646
rect 45938 27582 45950 27634
rect 46002 27582 46014 27634
rect 25566 27570 25618 27582
rect 1344 27466 58576 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 58576 27466
rect 1344 27380 58576 27414
rect 18958 27298 19010 27310
rect 57934 27298 57986 27310
rect 22082 27246 22094 27298
rect 22146 27246 22158 27298
rect 18958 27234 19010 27246
rect 57934 27234 57986 27246
rect 20078 27186 20130 27198
rect 15138 27134 15150 27186
rect 15202 27134 15214 27186
rect 17266 27134 17278 27186
rect 17330 27134 17342 27186
rect 20078 27122 20130 27134
rect 20526 27186 20578 27198
rect 20526 27122 20578 27134
rect 22654 27186 22706 27198
rect 26574 27186 26626 27198
rect 22866 27134 22878 27186
rect 22930 27134 22942 27186
rect 24994 27134 25006 27186
rect 25058 27134 25070 27186
rect 22654 27122 22706 27134
rect 26574 27122 26626 27134
rect 27134 27186 27186 27198
rect 27134 27122 27186 27134
rect 27694 27186 27746 27198
rect 27694 27122 27746 27134
rect 28590 27186 28642 27198
rect 30382 27186 30434 27198
rect 29250 27134 29262 27186
rect 29314 27134 29326 27186
rect 28590 27122 28642 27134
rect 30382 27122 30434 27134
rect 32174 27186 32226 27198
rect 52670 27186 52722 27198
rect 32498 27134 32510 27186
rect 32562 27134 32574 27186
rect 37762 27134 37774 27186
rect 37826 27134 37838 27186
rect 39890 27134 39902 27186
rect 39954 27134 39966 27186
rect 41010 27134 41022 27186
rect 41074 27134 41086 27186
rect 43138 27134 43150 27186
rect 43202 27134 43214 27186
rect 47954 27134 47966 27186
rect 48018 27134 48030 27186
rect 51762 27134 51774 27186
rect 51826 27134 51838 27186
rect 32174 27122 32226 27134
rect 52670 27122 52722 27134
rect 1710 27074 1762 27086
rect 3166 27074 3218 27086
rect 2482 27022 2494 27074
rect 2546 27022 2558 27074
rect 1710 27010 1762 27022
rect 3166 27010 3218 27022
rect 3614 27074 3666 27086
rect 19070 27074 19122 27086
rect 6850 27022 6862 27074
rect 6914 27022 6926 27074
rect 7746 27022 7758 27074
rect 7810 27022 7822 27074
rect 17938 27022 17950 27074
rect 18002 27022 18014 27074
rect 3614 27010 3666 27022
rect 19070 27010 19122 27022
rect 19294 27074 19346 27086
rect 19294 27010 19346 27022
rect 19406 27074 19458 27086
rect 21534 27074 21586 27086
rect 21298 27022 21310 27074
rect 21362 27022 21374 27074
rect 19406 27010 19458 27022
rect 21534 27010 21586 27022
rect 21646 27074 21698 27086
rect 26014 27074 26066 27086
rect 25666 27022 25678 27074
rect 25730 27022 25742 27074
rect 21646 27010 21698 27022
rect 26014 27010 26066 27022
rect 27582 27074 27634 27086
rect 27582 27010 27634 27022
rect 28254 27074 28306 27086
rect 28254 27010 28306 27022
rect 29710 27074 29762 27086
rect 50990 27074 51042 27086
rect 53566 27074 53618 27086
rect 30818 27022 30830 27074
rect 30882 27022 30894 27074
rect 32610 27022 32622 27074
rect 32674 27022 32686 27074
rect 32834 27022 32846 27074
rect 32898 27022 32910 27074
rect 33954 27022 33966 27074
rect 34018 27022 34030 27074
rect 35298 27022 35310 27074
rect 35362 27022 35374 27074
rect 35970 27022 35982 27074
rect 36034 27022 36046 27074
rect 36978 27022 36990 27074
rect 37042 27022 37054 27074
rect 40338 27022 40350 27074
rect 40402 27022 40414 27074
rect 45490 27022 45502 27074
rect 45554 27022 45566 27074
rect 46610 27022 46622 27074
rect 46674 27022 46686 27074
rect 47394 27022 47406 27074
rect 47458 27022 47470 27074
rect 48066 27022 48078 27074
rect 48130 27022 48142 27074
rect 49074 27022 49086 27074
rect 49138 27022 49150 27074
rect 50194 27022 50206 27074
rect 50258 27022 50270 27074
rect 51874 27022 51886 27074
rect 51938 27022 51950 27074
rect 53106 27022 53118 27074
rect 53170 27022 53182 27074
rect 55570 27022 55582 27074
rect 55634 27022 55646 27074
rect 29710 27010 29762 27022
rect 50990 27010 51042 27022
rect 53566 27010 53618 27022
rect 2046 26962 2098 26974
rect 2046 26898 2098 26910
rect 2718 26962 2770 26974
rect 9102 26962 9154 26974
rect 6514 26910 6526 26962
rect 6578 26910 6590 26962
rect 2718 26898 2770 26910
rect 9102 26898 9154 26910
rect 18622 26962 18674 26974
rect 18622 26898 18674 26910
rect 26462 26962 26514 26974
rect 26462 26898 26514 26910
rect 33070 26962 33122 26974
rect 33070 26898 33122 26910
rect 33294 26962 33346 26974
rect 54350 26962 54402 26974
rect 35186 26910 35198 26962
rect 35250 26910 35262 26962
rect 36082 26910 36094 26962
rect 36146 26910 36158 26962
rect 45602 26910 45614 26962
rect 45666 26910 45678 26962
rect 48738 26910 48750 26962
rect 48802 26910 48814 26962
rect 49186 26910 49198 26962
rect 49250 26910 49262 26962
rect 33294 26898 33346 26910
rect 54350 26898 54402 26910
rect 54462 26962 54514 26974
rect 54462 26898 54514 26910
rect 54686 26962 54738 26974
rect 54686 26898 54738 26910
rect 54910 26962 54962 26974
rect 54910 26898 54962 26910
rect 26686 26850 26738 26862
rect 26686 26786 26738 26798
rect 27806 26850 27858 26862
rect 27806 26786 27858 26798
rect 31614 26850 31666 26862
rect 31614 26786 31666 26798
rect 33854 26850 33906 26862
rect 46498 26798 46510 26850
rect 46562 26798 46574 26850
rect 49970 26798 49982 26850
rect 50034 26798 50046 26850
rect 33854 26786 33906 26798
rect 1344 26682 58576 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 50558 26682
rect 50610 26630 50662 26682
rect 50714 26630 50766 26682
rect 50818 26630 58576 26682
rect 1344 26596 58576 26630
rect 2046 26514 2098 26526
rect 2046 26450 2098 26462
rect 2718 26514 2770 26526
rect 2718 26450 2770 26462
rect 3390 26514 3442 26526
rect 3390 26450 3442 26462
rect 12686 26514 12738 26526
rect 12686 26450 12738 26462
rect 14926 26514 14978 26526
rect 14926 26450 14978 26462
rect 15486 26514 15538 26526
rect 26462 26514 26514 26526
rect 25554 26462 25566 26514
rect 25618 26462 25630 26514
rect 15486 26450 15538 26462
rect 26462 26450 26514 26462
rect 26686 26514 26738 26526
rect 26686 26450 26738 26462
rect 28142 26514 28194 26526
rect 28142 26450 28194 26462
rect 28926 26514 28978 26526
rect 28926 26450 28978 26462
rect 29934 26514 29986 26526
rect 29934 26450 29986 26462
rect 31726 26514 31778 26526
rect 31726 26450 31778 26462
rect 41806 26514 41858 26526
rect 41806 26450 41858 26462
rect 42478 26514 42530 26526
rect 42478 26450 42530 26462
rect 47518 26514 47570 26526
rect 47518 26450 47570 26462
rect 51662 26514 51714 26526
rect 51662 26450 51714 26462
rect 52558 26514 52610 26526
rect 52558 26450 52610 26462
rect 55582 26514 55634 26526
rect 55582 26450 55634 26462
rect 4734 26402 4786 26414
rect 12462 26402 12514 26414
rect 5394 26350 5406 26402
rect 5458 26350 5470 26402
rect 6290 26350 6302 26402
rect 6354 26350 6366 26402
rect 4734 26338 4786 26350
rect 12462 26338 12514 26350
rect 13806 26402 13858 26414
rect 13806 26338 13858 26350
rect 14030 26402 14082 26414
rect 14030 26338 14082 26350
rect 18398 26402 18450 26414
rect 18398 26338 18450 26350
rect 26126 26402 26178 26414
rect 26126 26338 26178 26350
rect 27694 26402 27746 26414
rect 27694 26338 27746 26350
rect 29710 26402 29762 26414
rect 29710 26338 29762 26350
rect 30606 26402 30658 26414
rect 30606 26338 30658 26350
rect 30942 26402 30994 26414
rect 30942 26338 30994 26350
rect 31166 26402 31218 26414
rect 33518 26402 33570 26414
rect 32162 26350 32174 26402
rect 32226 26350 32238 26402
rect 31166 26338 31218 26350
rect 33518 26338 33570 26350
rect 41918 26402 41970 26414
rect 41918 26338 41970 26350
rect 42814 26402 42866 26414
rect 42814 26338 42866 26350
rect 45950 26402 46002 26414
rect 45950 26338 46002 26350
rect 50318 26402 50370 26414
rect 50318 26338 50370 26350
rect 51886 26402 51938 26414
rect 51886 26338 51938 26350
rect 51998 26402 52050 26414
rect 51998 26338 52050 26350
rect 52446 26402 52498 26414
rect 52446 26338 52498 26350
rect 52670 26402 52722 26414
rect 52670 26338 52722 26350
rect 53118 26402 53170 26414
rect 53118 26338 53170 26350
rect 54126 26402 54178 26414
rect 57810 26350 57822 26402
rect 57874 26350 57886 26402
rect 54126 26338 54178 26350
rect 2382 26290 2434 26302
rect 1810 26238 1822 26290
rect 1874 26238 1886 26290
rect 2382 26226 2434 26238
rect 3054 26290 3106 26302
rect 8206 26290 8258 26302
rect 5170 26238 5182 26290
rect 5234 26238 5246 26290
rect 6850 26238 6862 26290
rect 6914 26238 6926 26290
rect 7746 26238 7758 26290
rect 7810 26238 7822 26290
rect 3054 26226 3106 26238
rect 8206 26226 8258 26238
rect 9550 26290 9602 26302
rect 9550 26226 9602 26238
rect 9886 26290 9938 26302
rect 9886 26226 9938 26238
rect 10110 26290 10162 26302
rect 11454 26290 11506 26302
rect 11106 26238 11118 26290
rect 11170 26238 11182 26290
rect 10110 26226 10162 26238
rect 11454 26226 11506 26238
rect 11566 26290 11618 26302
rect 11566 26226 11618 26238
rect 12350 26290 12402 26302
rect 12350 26226 12402 26238
rect 13134 26290 13186 26302
rect 13134 26226 13186 26238
rect 14366 26290 14418 26302
rect 16494 26290 16546 26302
rect 14690 26238 14702 26290
rect 14754 26238 14766 26290
rect 14366 26226 14418 26238
rect 16494 26226 16546 26238
rect 18286 26290 18338 26302
rect 18286 26226 18338 26238
rect 18622 26290 18674 26302
rect 25118 26290 25170 26302
rect 25678 26290 25730 26302
rect 23650 26238 23662 26290
rect 23714 26238 23726 26290
rect 25442 26238 25454 26290
rect 25506 26238 25518 26290
rect 18622 26226 18674 26238
rect 25118 26226 25170 26238
rect 25678 26226 25730 26238
rect 27134 26290 27186 26302
rect 30158 26290 30210 26302
rect 27458 26238 27470 26290
rect 27522 26238 27534 26290
rect 27134 26226 27186 26238
rect 30158 26226 30210 26238
rect 30382 26290 30434 26302
rect 30382 26226 30434 26238
rect 30718 26290 30770 26302
rect 30718 26226 30770 26238
rect 31278 26290 31330 26302
rect 31278 26226 31330 26238
rect 31502 26290 31554 26302
rect 31502 26226 31554 26238
rect 31838 26290 31890 26302
rect 31838 26226 31890 26238
rect 32510 26290 32562 26302
rect 32510 26226 32562 26238
rect 33742 26290 33794 26302
rect 33742 26226 33794 26238
rect 34078 26290 34130 26302
rect 41582 26290 41634 26302
rect 46062 26290 46114 26302
rect 50094 26290 50146 26302
rect 34962 26238 34974 26290
rect 35026 26238 35038 26290
rect 43250 26238 43262 26290
rect 43314 26238 43326 26290
rect 44482 26238 44494 26290
rect 44546 26238 44558 26290
rect 45154 26238 45166 26290
rect 45218 26238 45230 26290
rect 47730 26238 47742 26290
rect 47794 26238 47806 26290
rect 49634 26238 49646 26290
rect 49698 26238 49710 26290
rect 34078 26226 34130 26238
rect 41582 26226 41634 26238
rect 46062 26226 46114 26238
rect 50094 26226 50146 26238
rect 50430 26290 50482 26302
rect 50430 26226 50482 26238
rect 52894 26290 52946 26302
rect 52894 26226 52946 26238
rect 53230 26290 53282 26302
rect 55358 26290 55410 26302
rect 54786 26238 54798 26290
rect 54850 26238 54862 26290
rect 53230 26226 53282 26238
rect 55358 26226 55410 26238
rect 55694 26290 55746 26302
rect 55694 26226 55746 26238
rect 55918 26290 55970 26302
rect 58158 26290 58210 26302
rect 56578 26238 56590 26290
rect 56642 26238 56654 26290
rect 55918 26226 55970 26238
rect 58158 26226 58210 26238
rect 3838 26178 3890 26190
rect 3838 26114 3890 26126
rect 4286 26178 4338 26190
rect 4286 26114 4338 26126
rect 9998 26178 10050 26190
rect 9998 26114 10050 26126
rect 12910 26178 12962 26190
rect 12910 26114 12962 26126
rect 18958 26178 19010 26190
rect 18958 26114 19010 26126
rect 19406 26178 19458 26190
rect 24222 26178 24274 26190
rect 20738 26126 20750 26178
rect 20802 26126 20814 26178
rect 22978 26126 22990 26178
rect 23042 26126 23054 26178
rect 19406 26114 19458 26126
rect 24222 26114 24274 26126
rect 25902 26178 25954 26190
rect 25902 26114 25954 26126
rect 26574 26178 26626 26190
rect 26574 26114 26626 26126
rect 29262 26178 29314 26190
rect 29262 26114 29314 26126
rect 30046 26178 30098 26190
rect 30046 26114 30098 26126
rect 33182 26178 33234 26190
rect 33182 26114 33234 26126
rect 33966 26178 34018 26190
rect 33966 26114 34018 26126
rect 34526 26178 34578 26190
rect 41022 26178 41074 26190
rect 44382 26178 44434 26190
rect 53790 26178 53842 26190
rect 57374 26178 57426 26190
rect 37090 26126 37102 26178
rect 37154 26126 37166 26178
rect 43698 26126 43710 26178
rect 43762 26126 43774 26178
rect 45266 26126 45278 26178
rect 45330 26126 45342 26178
rect 49410 26126 49422 26178
rect 49474 26126 49486 26178
rect 54562 26126 54574 26178
rect 54626 26126 54638 26178
rect 34526 26114 34578 26126
rect 41022 26114 41074 26126
rect 44382 26114 44434 26126
rect 53790 26114 53842 26126
rect 57374 26114 57426 26126
rect 13470 26066 13522 26078
rect 13470 26002 13522 26014
rect 14142 26066 14194 26078
rect 14142 26002 14194 26014
rect 15038 26066 15090 26078
rect 15038 26002 15090 26014
rect 16606 26066 16658 26078
rect 45950 26066 46002 26078
rect 18722 26014 18734 26066
rect 18786 26063 18798 26066
rect 19506 26063 19518 26066
rect 18786 26017 19518 26063
rect 18786 26014 18798 26017
rect 19506 26014 19518 26017
rect 19570 26014 19582 26066
rect 40786 26014 40798 26066
rect 40850 26063 40862 26066
rect 41458 26063 41470 26066
rect 40850 26017 41470 26063
rect 40850 26014 40862 26017
rect 41458 26014 41470 26017
rect 41522 26014 41534 26066
rect 16606 26002 16658 26014
rect 45950 26002 46002 26014
rect 47406 26066 47458 26078
rect 56590 26066 56642 26078
rect 49074 26014 49086 26066
rect 49138 26014 49150 26066
rect 47406 26002 47458 26014
rect 56590 26002 56642 26014
rect 56926 26066 56978 26078
rect 56926 26002 56978 26014
rect 1344 25898 58576 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 58576 25898
rect 1344 25812 58576 25846
rect 5966 25730 6018 25742
rect 5966 25666 6018 25678
rect 22990 25730 23042 25742
rect 22990 25666 23042 25678
rect 23214 25730 23266 25742
rect 23214 25666 23266 25678
rect 23774 25730 23826 25742
rect 52782 25730 52834 25742
rect 37762 25678 37774 25730
rect 37826 25727 37838 25730
rect 38210 25727 38222 25730
rect 37826 25681 38222 25727
rect 37826 25678 37838 25681
rect 38210 25678 38222 25681
rect 38274 25727 38286 25730
rect 38434 25727 38446 25730
rect 38274 25681 38446 25727
rect 38274 25678 38286 25681
rect 38434 25678 38446 25681
rect 38498 25678 38510 25730
rect 45490 25678 45502 25730
rect 45554 25678 45566 25730
rect 54674 25678 54686 25730
rect 54738 25678 54750 25730
rect 57474 25678 57486 25730
rect 57538 25678 57550 25730
rect 23774 25666 23826 25678
rect 52782 25666 52834 25678
rect 1934 25618 1986 25630
rect 20526 25618 20578 25630
rect 27470 25618 27522 25630
rect 38446 25618 38498 25630
rect 46958 25618 47010 25630
rect 6738 25566 6750 25618
rect 6802 25566 6814 25618
rect 13906 25566 13918 25618
rect 13970 25566 13982 25618
rect 24882 25566 24894 25618
rect 24946 25566 24958 25618
rect 27010 25566 27022 25618
rect 27074 25566 27086 25618
rect 29922 25566 29934 25618
rect 29986 25566 29998 25618
rect 33058 25566 33070 25618
rect 33122 25566 33134 25618
rect 35746 25566 35758 25618
rect 35810 25566 35822 25618
rect 46274 25566 46286 25618
rect 46338 25566 46350 25618
rect 1934 25554 1986 25566
rect 20526 25554 20578 25566
rect 27470 25554 27522 25566
rect 38446 25554 38498 25566
rect 46958 25554 47010 25566
rect 49982 25618 50034 25630
rect 55010 25566 55022 25618
rect 55074 25566 55086 25618
rect 49982 25554 50034 25566
rect 7534 25506 7586 25518
rect 4274 25454 4286 25506
rect 4338 25454 4350 25506
rect 4834 25454 4846 25506
rect 4898 25454 4910 25506
rect 5954 25454 5966 25506
rect 6018 25454 6030 25506
rect 6626 25454 6638 25506
rect 6690 25454 6702 25506
rect 7534 25442 7586 25454
rect 7870 25506 7922 25518
rect 9774 25506 9826 25518
rect 8866 25454 8878 25506
rect 8930 25454 8942 25506
rect 9426 25454 9438 25506
rect 9490 25454 9502 25506
rect 7870 25442 7922 25454
rect 9774 25442 9826 25454
rect 9998 25506 10050 25518
rect 9998 25442 10050 25454
rect 11454 25506 11506 25518
rect 11454 25442 11506 25454
rect 11678 25506 11730 25518
rect 14702 25506 14754 25518
rect 14018 25454 14030 25506
rect 14082 25454 14094 25506
rect 11678 25442 11730 25454
rect 14702 25442 14754 25454
rect 15038 25506 15090 25518
rect 18734 25506 18786 25518
rect 16594 25454 16606 25506
rect 16658 25454 16670 25506
rect 18162 25454 18174 25506
rect 18226 25454 18238 25506
rect 15038 25442 15090 25454
rect 18734 25442 18786 25454
rect 19518 25506 19570 25518
rect 19518 25442 19570 25454
rect 23662 25506 23714 25518
rect 27806 25506 27858 25518
rect 33406 25506 33458 25518
rect 37550 25506 37602 25518
rect 24210 25454 24222 25506
rect 24274 25454 24286 25506
rect 29250 25454 29262 25506
rect 29314 25454 29326 25506
rect 32610 25454 32622 25506
rect 32674 25454 32686 25506
rect 34178 25454 34190 25506
rect 34242 25454 34254 25506
rect 35074 25454 35086 25506
rect 35138 25454 35150 25506
rect 35970 25454 35982 25506
rect 36034 25454 36046 25506
rect 23662 25442 23714 25454
rect 27806 25442 27858 25454
rect 33406 25442 33458 25454
rect 37550 25442 37602 25454
rect 37998 25506 38050 25518
rect 37998 25442 38050 25454
rect 40238 25506 40290 25518
rect 41134 25506 41186 25518
rect 40674 25454 40686 25506
rect 40738 25454 40750 25506
rect 40238 25442 40290 25454
rect 41134 25442 41186 25454
rect 41582 25506 41634 25518
rect 41582 25442 41634 25454
rect 44830 25506 44882 25518
rect 44830 25442 44882 25454
rect 45166 25506 45218 25518
rect 46734 25506 46786 25518
rect 45938 25454 45950 25506
rect 46002 25454 46014 25506
rect 45166 25442 45218 25454
rect 46734 25442 46786 25454
rect 47182 25506 47234 25518
rect 47182 25442 47234 25454
rect 47630 25506 47682 25518
rect 47630 25442 47682 25454
rect 47966 25506 48018 25518
rect 49534 25506 49586 25518
rect 48626 25454 48638 25506
rect 48690 25454 48702 25506
rect 47966 25442 48018 25454
rect 49534 25442 49586 25454
rect 50206 25506 50258 25518
rect 50206 25442 50258 25454
rect 50318 25506 50370 25518
rect 50318 25442 50370 25454
rect 50654 25506 50706 25518
rect 50654 25442 50706 25454
rect 53566 25506 53618 25518
rect 53566 25442 53618 25454
rect 53902 25506 53954 25518
rect 54562 25454 54574 25506
rect 54626 25454 54638 25506
rect 55570 25454 55582 25506
rect 55634 25454 55646 25506
rect 53902 25442 53954 25454
rect 5630 25394 5682 25406
rect 5630 25330 5682 25342
rect 7198 25394 7250 25406
rect 7198 25330 7250 25342
rect 7646 25394 7698 25406
rect 10670 25394 10722 25406
rect 8418 25342 8430 25394
rect 8482 25342 8494 25394
rect 7646 25330 7698 25342
rect 10670 25330 10722 25342
rect 12350 25394 12402 25406
rect 18510 25394 18562 25406
rect 16258 25342 16270 25394
rect 16322 25342 16334 25394
rect 12350 25330 12402 25342
rect 18510 25330 18562 25342
rect 20078 25394 20130 25406
rect 33070 25394 33122 25406
rect 28130 25342 28142 25394
rect 28194 25342 28206 25394
rect 20078 25330 20130 25342
rect 33070 25330 33122 25342
rect 33182 25394 33234 25406
rect 37438 25394 37490 25406
rect 35186 25342 35198 25394
rect 35250 25342 35262 25394
rect 36194 25342 36206 25394
rect 36258 25342 36270 25394
rect 33182 25330 33234 25342
rect 37438 25330 37490 25342
rect 47406 25394 47458 25406
rect 47406 25330 47458 25342
rect 47854 25394 47906 25406
rect 47854 25330 47906 25342
rect 49758 25394 49810 25406
rect 49758 25330 49810 25342
rect 52782 25394 52834 25406
rect 52782 25330 52834 25342
rect 52894 25394 52946 25406
rect 52894 25330 52946 25342
rect 53678 25394 53730 25406
rect 53678 25330 53730 25342
rect 10782 25282 10834 25294
rect 5058 25230 5070 25282
rect 5122 25230 5134 25282
rect 9314 25230 9326 25282
rect 9378 25230 9390 25282
rect 10322 25230 10334 25282
rect 10386 25230 10398 25282
rect 10782 25218 10834 25230
rect 11006 25282 11058 25294
rect 12462 25282 12514 25294
rect 12002 25230 12014 25282
rect 12066 25230 12078 25282
rect 11006 25218 11058 25230
rect 12462 25218 12514 25230
rect 12574 25282 12626 25294
rect 12574 25218 12626 25230
rect 15150 25282 15202 25294
rect 15150 25218 15202 25230
rect 15374 25282 15426 25294
rect 19854 25282 19906 25294
rect 17602 25230 17614 25282
rect 17666 25230 17678 25282
rect 19058 25230 19070 25282
rect 19122 25230 19134 25282
rect 15374 25218 15426 25230
rect 19854 25218 19906 25230
rect 20190 25282 20242 25294
rect 20190 25218 20242 25230
rect 22878 25282 22930 25294
rect 37214 25282 37266 25294
rect 32162 25230 32174 25282
rect 32226 25230 32238 25282
rect 22878 25218 22930 25230
rect 37214 25218 37266 25230
rect 39006 25282 39058 25294
rect 39006 25218 39058 25230
rect 39454 25282 39506 25294
rect 39454 25218 39506 25230
rect 39902 25282 39954 25294
rect 39902 25218 39954 25230
rect 41694 25282 41746 25294
rect 41694 25218 41746 25230
rect 42142 25282 42194 25294
rect 42142 25218 42194 25230
rect 44942 25282 44994 25294
rect 50542 25282 50594 25294
rect 48850 25230 48862 25282
rect 48914 25230 48926 25282
rect 44942 25218 44994 25230
rect 50542 25218 50594 25230
rect 52110 25282 52162 25294
rect 52110 25218 52162 25230
rect 1344 25114 58576 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 50558 25114
rect 50610 25062 50662 25114
rect 50714 25062 50766 25114
rect 50818 25062 58576 25114
rect 1344 25028 58576 25062
rect 4286 24946 4338 24958
rect 4286 24882 4338 24894
rect 5406 24946 5458 24958
rect 5406 24882 5458 24894
rect 16718 24946 16770 24958
rect 16718 24882 16770 24894
rect 20862 24946 20914 24958
rect 20862 24882 20914 24894
rect 21646 24946 21698 24958
rect 21646 24882 21698 24894
rect 22206 24946 22258 24958
rect 22206 24882 22258 24894
rect 24110 24946 24162 24958
rect 24110 24882 24162 24894
rect 26462 24946 26514 24958
rect 27246 24946 27298 24958
rect 26462 24882 26514 24894
rect 26910 24890 26962 24902
rect 16270 24834 16322 24846
rect 3266 24782 3278 24834
rect 3330 24782 3342 24834
rect 16270 24770 16322 24782
rect 16606 24834 16658 24846
rect 27246 24882 27298 24894
rect 32174 24946 32226 24958
rect 32174 24882 32226 24894
rect 32510 24946 32562 24958
rect 32510 24882 32562 24894
rect 35422 24946 35474 24958
rect 46062 24946 46114 24958
rect 42578 24894 42590 24946
rect 42642 24894 42654 24946
rect 45602 24894 45614 24946
rect 45666 24894 45678 24946
rect 35422 24882 35474 24894
rect 46062 24882 46114 24894
rect 26910 24826 26962 24838
rect 27022 24834 27074 24846
rect 16606 24770 16658 24782
rect 27022 24770 27074 24782
rect 27694 24834 27746 24846
rect 27694 24770 27746 24782
rect 27806 24834 27858 24846
rect 27806 24770 27858 24782
rect 30270 24834 30322 24846
rect 30270 24770 30322 24782
rect 30382 24834 30434 24846
rect 30382 24770 30434 24782
rect 33518 24834 33570 24846
rect 34638 24834 34690 24846
rect 39902 24834 39954 24846
rect 34290 24782 34302 24834
rect 34354 24782 34366 24834
rect 35746 24782 35758 24834
rect 35810 24782 35822 24834
rect 33518 24770 33570 24782
rect 34638 24770 34690 24782
rect 39902 24770 39954 24782
rect 41022 24834 41074 24846
rect 43822 24834 43874 24846
rect 41682 24782 41694 24834
rect 41746 24782 41758 24834
rect 41022 24770 41074 24782
rect 43822 24770 43874 24782
rect 3054 24722 3106 24734
rect 3838 24722 3890 24734
rect 2034 24670 2046 24722
rect 2098 24670 2110 24722
rect 3378 24670 3390 24722
rect 3442 24670 3454 24722
rect 3054 24658 3106 24670
rect 3838 24658 3890 24670
rect 4734 24722 4786 24734
rect 4734 24658 4786 24670
rect 6302 24722 6354 24734
rect 9102 24722 9154 24734
rect 16942 24722 16994 24734
rect 20190 24722 20242 24734
rect 7858 24670 7870 24722
rect 7922 24670 7934 24722
rect 8082 24670 8094 24722
rect 8146 24670 8158 24722
rect 8306 24670 8318 24722
rect 8370 24670 8382 24722
rect 9762 24670 9774 24722
rect 9826 24670 9838 24722
rect 11778 24670 11790 24722
rect 11842 24670 11854 24722
rect 12674 24670 12686 24722
rect 12738 24670 12750 24722
rect 13570 24670 13582 24722
rect 13634 24670 13646 24722
rect 15586 24670 15598 24722
rect 15650 24670 15662 24722
rect 17266 24670 17278 24722
rect 17330 24670 17342 24722
rect 18050 24670 18062 24722
rect 18114 24670 18126 24722
rect 19282 24670 19294 24722
rect 19346 24670 19358 24722
rect 6302 24658 6354 24670
rect 9102 24658 9154 24670
rect 16942 24658 16994 24670
rect 20190 24658 20242 24670
rect 20526 24722 20578 24734
rect 20526 24658 20578 24670
rect 20862 24722 20914 24734
rect 20862 24658 20914 24670
rect 21198 24722 21250 24734
rect 21198 24658 21250 24670
rect 21422 24722 21474 24734
rect 21422 24658 21474 24670
rect 21758 24722 21810 24734
rect 21758 24658 21810 24670
rect 30046 24722 30098 24734
rect 32958 24722 33010 24734
rect 34862 24722 34914 24734
rect 30818 24670 30830 24722
rect 30882 24670 30894 24722
rect 33282 24670 33294 24722
rect 33346 24670 33358 24722
rect 34402 24670 34414 24722
rect 34466 24670 34478 24722
rect 30046 24658 30098 24670
rect 32958 24658 33010 24670
rect 34862 24658 34914 24670
rect 35198 24722 35250 24734
rect 40014 24722 40066 24734
rect 35634 24670 35646 24722
rect 35698 24670 35710 24722
rect 36306 24670 36318 24722
rect 36370 24670 36382 24722
rect 35198 24658 35250 24670
rect 40014 24658 40066 24670
rect 41134 24722 41186 24734
rect 49422 24722 49474 24734
rect 41570 24670 41582 24722
rect 41634 24670 41646 24722
rect 42466 24670 42478 24722
rect 42530 24670 42542 24722
rect 44258 24670 44270 24722
rect 44322 24670 44334 24722
rect 45378 24670 45390 24722
rect 45442 24670 45454 24722
rect 49074 24670 49086 24722
rect 49138 24670 49150 24722
rect 41134 24658 41186 24670
rect 49422 24658 49474 24670
rect 49982 24722 50034 24734
rect 49982 24658 50034 24670
rect 50318 24722 50370 24734
rect 50318 24658 50370 24670
rect 50654 24722 50706 24734
rect 50654 24658 50706 24670
rect 52110 24722 52162 24734
rect 52546 24670 52558 24722
rect 52610 24670 52622 24722
rect 53442 24670 53454 24722
rect 53506 24670 53518 24722
rect 57138 24670 57150 24722
rect 57202 24670 57214 24722
rect 52110 24658 52162 24670
rect 2494 24610 2546 24622
rect 2494 24546 2546 24558
rect 2830 24610 2882 24622
rect 2830 24546 2882 24558
rect 4510 24610 4562 24622
rect 4510 24546 4562 24558
rect 5742 24610 5794 24622
rect 5742 24546 5794 24558
rect 6078 24610 6130 24622
rect 18510 24610 18562 24622
rect 23662 24610 23714 24622
rect 10546 24558 10558 24610
rect 10610 24558 10622 24610
rect 11554 24558 11566 24610
rect 11618 24558 11630 24610
rect 13458 24558 13470 24610
rect 13522 24558 13534 24610
rect 15362 24558 15374 24610
rect 15426 24558 15438 24610
rect 19730 24558 19742 24610
rect 19794 24558 19806 24610
rect 6078 24546 6130 24558
rect 18510 24546 18562 24558
rect 23662 24546 23714 24558
rect 28366 24610 28418 24622
rect 33182 24610 33234 24622
rect 30370 24558 30382 24610
rect 30434 24558 30446 24610
rect 28366 24546 28418 24558
rect 33182 24546 33234 24558
rect 34750 24610 34802 24622
rect 49646 24610 49698 24622
rect 35970 24558 35982 24610
rect 36034 24558 36046 24610
rect 37090 24558 37102 24610
rect 37154 24558 37166 24610
rect 39218 24558 39230 24610
rect 39282 24558 39294 24610
rect 44146 24558 44158 24610
rect 44210 24558 44222 24610
rect 34750 24546 34802 24558
rect 49646 24546 49698 24558
rect 50430 24610 50482 24622
rect 56702 24610 56754 24622
rect 52994 24558 53006 24610
rect 53058 24558 53070 24610
rect 57362 24558 57374 24610
rect 57426 24558 57438 24610
rect 50430 24546 50482 24558
rect 56702 24546 56754 24558
rect 4958 24498 5010 24510
rect 4958 24434 5010 24446
rect 6526 24498 6578 24510
rect 6526 24434 6578 24446
rect 6750 24498 6802 24510
rect 6750 24434 6802 24446
rect 7198 24498 7250 24510
rect 27806 24498 27858 24510
rect 18274 24446 18286 24498
rect 18338 24446 18350 24498
rect 7198 24434 7250 24446
rect 27806 24434 27858 24446
rect 39902 24498 39954 24510
rect 39902 24434 39954 24446
rect 41246 24498 41298 24510
rect 55346 24446 55358 24498
rect 55410 24446 55422 24498
rect 41246 24434 41298 24446
rect 1344 24330 58576 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 58576 24330
rect 1344 24244 58576 24278
rect 3838 24162 3890 24174
rect 3838 24098 3890 24110
rect 17838 24162 17890 24174
rect 17838 24098 17890 24110
rect 18174 24162 18226 24174
rect 18174 24098 18226 24110
rect 18622 24162 18674 24174
rect 18622 24098 18674 24110
rect 20190 24162 20242 24174
rect 20190 24098 20242 24110
rect 24222 24162 24274 24174
rect 37102 24162 37154 24174
rect 34962 24110 34974 24162
rect 35026 24159 35038 24162
rect 35186 24159 35198 24162
rect 35026 24113 35198 24159
rect 35026 24110 35038 24113
rect 35186 24110 35198 24113
rect 35250 24110 35262 24162
rect 24222 24098 24274 24110
rect 37102 24098 37154 24110
rect 57934 24162 57986 24174
rect 57934 24098 57986 24110
rect 12910 24050 12962 24062
rect 2370 23998 2382 24050
rect 2434 23998 2446 24050
rect 9202 23998 9214 24050
rect 9266 23998 9278 24050
rect 10770 23998 10782 24050
rect 10834 23998 10846 24050
rect 12910 23986 12962 23998
rect 17166 24050 17218 24062
rect 17166 23986 17218 23998
rect 24446 24050 24498 24062
rect 24446 23986 24498 23998
rect 25118 24050 25170 24062
rect 33742 24050 33794 24062
rect 28354 23998 28366 24050
rect 28418 23998 28430 24050
rect 30034 23998 30046 24050
rect 30098 23998 30110 24050
rect 31714 23998 31726 24050
rect 31778 23998 31790 24050
rect 25118 23986 25170 23998
rect 33742 23986 33794 23998
rect 38222 24050 38274 24062
rect 44942 24050 44994 24062
rect 39778 23998 39790 24050
rect 39842 23998 39854 24050
rect 38222 23986 38274 23998
rect 44942 23986 44994 23998
rect 45838 24050 45890 24062
rect 45838 23986 45890 23998
rect 48414 24050 48466 24062
rect 48414 23986 48466 23998
rect 2830 23938 2882 23950
rect 4622 23938 4674 23950
rect 2034 23886 2046 23938
rect 2098 23886 2110 23938
rect 3378 23886 3390 23938
rect 3442 23886 3454 23938
rect 2830 23874 2882 23886
rect 4622 23874 4674 23886
rect 5854 23938 5906 23950
rect 5854 23874 5906 23886
rect 6526 23938 6578 23950
rect 7086 23938 7138 23950
rect 6850 23886 6862 23938
rect 6914 23886 6926 23938
rect 6526 23874 6578 23886
rect 7086 23874 7138 23886
rect 7534 23938 7586 23950
rect 7534 23874 7586 23886
rect 7870 23938 7922 23950
rect 7870 23874 7922 23886
rect 8206 23938 8258 23950
rect 14142 23938 14194 23950
rect 19742 23938 19794 23950
rect 8530 23886 8542 23938
rect 8594 23886 8606 23938
rect 12226 23886 12238 23938
rect 12290 23886 12302 23938
rect 13682 23886 13694 23938
rect 13746 23886 13758 23938
rect 15586 23886 15598 23938
rect 15650 23886 15662 23938
rect 16482 23886 16494 23938
rect 16546 23886 16558 23938
rect 8206 23874 8258 23886
rect 14142 23874 14194 23886
rect 19742 23874 19794 23886
rect 19966 23938 20018 23950
rect 29598 23938 29650 23950
rect 35870 23938 35922 23950
rect 23986 23886 23998 23938
rect 24050 23886 24062 23938
rect 25442 23886 25454 23938
rect 25506 23886 25518 23938
rect 30482 23886 30494 23938
rect 30546 23886 30558 23938
rect 31602 23886 31614 23938
rect 31666 23886 31678 23938
rect 34626 23886 34638 23938
rect 34690 23886 34702 23938
rect 19966 23874 20018 23886
rect 29598 23874 29650 23886
rect 35870 23874 35922 23886
rect 36990 23938 37042 23950
rect 36990 23874 37042 23886
rect 37774 23938 37826 23950
rect 41022 23938 41074 23950
rect 41918 23938 41970 23950
rect 39890 23886 39902 23938
rect 39954 23886 39966 23938
rect 41458 23886 41470 23938
rect 41522 23886 41534 23938
rect 37774 23874 37826 23886
rect 41022 23874 41074 23886
rect 41918 23874 41970 23886
rect 44270 23938 44322 23950
rect 46734 23938 46786 23950
rect 52110 23938 52162 23950
rect 46274 23886 46286 23938
rect 46338 23886 46350 23938
rect 47506 23886 47518 23938
rect 47570 23886 47582 23938
rect 49074 23886 49086 23938
rect 49138 23886 49150 23938
rect 49858 23886 49870 23938
rect 49922 23886 49934 23938
rect 53666 23886 53678 23938
rect 53730 23886 53742 23938
rect 55570 23886 55582 23938
rect 55634 23886 55646 23938
rect 44270 23874 44322 23886
rect 46734 23874 46786 23886
rect 52110 23874 52162 23886
rect 3166 23826 3218 23838
rect 14366 23826 14418 23838
rect 2930 23774 2942 23826
rect 2994 23774 3006 23826
rect 8866 23774 8878 23826
rect 8930 23774 8942 23826
rect 11218 23774 11230 23826
rect 11282 23774 11294 23826
rect 3166 23762 3218 23774
rect 14366 23762 14418 23774
rect 14478 23826 14530 23838
rect 18062 23826 18114 23838
rect 15474 23774 15486 23826
rect 15538 23774 15550 23826
rect 14478 23762 14530 23774
rect 18062 23762 18114 23774
rect 18510 23826 18562 23838
rect 18510 23762 18562 23774
rect 19406 23826 19458 23838
rect 19406 23762 19458 23774
rect 23326 23826 23378 23838
rect 23326 23762 23378 23774
rect 23438 23826 23490 23838
rect 23438 23762 23490 23774
rect 24558 23826 24610 23838
rect 29262 23826 29314 23838
rect 26226 23774 26238 23826
rect 26290 23774 26302 23826
rect 24558 23762 24610 23774
rect 29262 23762 29314 23774
rect 30158 23826 30210 23838
rect 30158 23762 30210 23774
rect 31278 23826 31330 23838
rect 37102 23826 37154 23838
rect 34402 23774 34414 23826
rect 34466 23774 34478 23826
rect 31278 23762 31330 23774
rect 37102 23762 37154 23774
rect 37662 23826 37714 23838
rect 37662 23762 37714 23774
rect 39342 23826 39394 23838
rect 39342 23762 39394 23774
rect 43934 23826 43986 23838
rect 43934 23762 43986 23774
rect 44046 23826 44098 23838
rect 50990 23826 51042 23838
rect 49970 23774 49982 23826
rect 50034 23774 50046 23826
rect 44046 23762 44098 23774
rect 50990 23762 51042 23774
rect 51214 23826 51266 23838
rect 51214 23762 51266 23774
rect 51438 23826 51490 23838
rect 55246 23826 55298 23838
rect 53442 23774 53454 23826
rect 53506 23774 53518 23826
rect 55010 23774 55022 23826
rect 55074 23774 55086 23826
rect 51438 23762 51490 23774
rect 55246 23762 55298 23774
rect 4062 23714 4114 23726
rect 4062 23650 4114 23662
rect 5182 23714 5234 23726
rect 5182 23650 5234 23662
rect 6190 23714 6242 23726
rect 6190 23650 6242 23662
rect 6974 23714 7026 23726
rect 6974 23650 7026 23662
rect 7198 23714 7250 23726
rect 7198 23650 7250 23662
rect 7870 23714 7922 23726
rect 7870 23650 7922 23662
rect 10446 23714 10498 23726
rect 18622 23714 18674 23726
rect 13906 23662 13918 23714
rect 13970 23662 13982 23714
rect 10446 23650 10498 23662
rect 18622 23650 18674 23662
rect 19518 23714 19570 23726
rect 19518 23650 19570 23662
rect 20526 23714 20578 23726
rect 20526 23650 20578 23662
rect 22542 23714 22594 23726
rect 23102 23714 23154 23726
rect 22866 23662 22878 23714
rect 22930 23662 22942 23714
rect 22542 23650 22594 23662
rect 23102 23650 23154 23662
rect 29374 23714 29426 23726
rect 29374 23650 29426 23662
rect 29822 23714 29874 23726
rect 29822 23650 29874 23662
rect 30046 23714 30098 23726
rect 30046 23650 30098 23662
rect 30942 23714 30994 23726
rect 30942 23650 30994 23662
rect 31166 23714 31218 23726
rect 31166 23650 31218 23662
rect 33294 23714 33346 23726
rect 33294 23650 33346 23662
rect 35198 23714 35250 23726
rect 35198 23650 35250 23662
rect 35982 23714 36034 23726
rect 35982 23650 36034 23662
rect 36206 23714 36258 23726
rect 36206 23650 36258 23662
rect 37438 23714 37490 23726
rect 50878 23714 50930 23726
rect 47730 23662 47742 23714
rect 47794 23662 47806 23714
rect 37438 23650 37490 23662
rect 50878 23650 50930 23662
rect 51774 23714 51826 23726
rect 51774 23650 51826 23662
rect 51998 23714 52050 23726
rect 51998 23650 52050 23662
rect 1344 23546 58576 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 50558 23546
rect 50610 23494 50662 23546
rect 50714 23494 50766 23546
rect 50818 23494 58576 23546
rect 1344 23460 58576 23494
rect 15486 23378 15538 23390
rect 27358 23378 27410 23390
rect 7298 23326 7310 23378
rect 7362 23326 7374 23378
rect 11666 23326 11678 23378
rect 11730 23326 11742 23378
rect 22306 23326 22318 23378
rect 22370 23326 22382 23378
rect 24098 23326 24110 23378
rect 24162 23326 24174 23378
rect 15486 23314 15538 23326
rect 27358 23314 27410 23326
rect 27470 23378 27522 23390
rect 27470 23314 27522 23326
rect 27806 23378 27858 23390
rect 27806 23314 27858 23326
rect 30046 23378 30098 23390
rect 30046 23314 30098 23326
rect 30830 23378 30882 23390
rect 30830 23314 30882 23326
rect 31054 23378 31106 23390
rect 31054 23314 31106 23326
rect 38558 23378 38610 23390
rect 38558 23314 38610 23326
rect 40238 23378 40290 23390
rect 40238 23314 40290 23326
rect 40462 23378 40514 23390
rect 40462 23314 40514 23326
rect 41022 23378 41074 23390
rect 41022 23314 41074 23326
rect 41470 23378 41522 23390
rect 41470 23314 41522 23326
rect 42142 23378 42194 23390
rect 42142 23314 42194 23326
rect 44046 23378 44098 23390
rect 44046 23314 44098 23326
rect 46734 23378 46786 23390
rect 56142 23378 56194 23390
rect 48066 23326 48078 23378
rect 48130 23326 48142 23378
rect 53890 23326 53902 23378
rect 53954 23326 53966 23378
rect 46734 23314 46786 23326
rect 56142 23314 56194 23326
rect 58158 23378 58210 23390
rect 58158 23314 58210 23326
rect 8766 23266 8818 23278
rect 13470 23266 13522 23278
rect 3714 23214 3726 23266
rect 3778 23214 3790 23266
rect 4722 23214 4734 23266
rect 4786 23214 4798 23266
rect 6850 23214 6862 23266
rect 6914 23214 6926 23266
rect 10658 23214 10670 23266
rect 10722 23214 10734 23266
rect 8766 23202 8818 23214
rect 13470 23202 13522 23214
rect 14926 23266 14978 23278
rect 14926 23202 14978 23214
rect 15710 23266 15762 23278
rect 15710 23202 15762 23214
rect 29822 23266 29874 23278
rect 40126 23266 40178 23278
rect 55806 23266 55858 23278
rect 35970 23214 35982 23266
rect 36034 23214 36046 23266
rect 47058 23214 47070 23266
rect 47122 23214 47134 23266
rect 52322 23214 52334 23266
rect 52386 23214 52398 23266
rect 55010 23214 55022 23266
rect 55074 23214 55086 23266
rect 29822 23202 29874 23214
rect 40126 23202 40178 23214
rect 55806 23202 55858 23214
rect 55918 23266 55970 23278
rect 55918 23202 55970 23214
rect 2270 23154 2322 23166
rect 7758 23154 7810 23166
rect 8654 23154 8706 23166
rect 11342 23154 11394 23166
rect 14814 23154 14866 23166
rect 4162 23102 4174 23154
rect 4226 23102 4238 23154
rect 4834 23102 4846 23154
rect 4898 23102 4910 23154
rect 7074 23102 7086 23154
rect 7138 23102 7150 23154
rect 8194 23102 8206 23154
rect 8258 23102 8270 23154
rect 9538 23102 9550 23154
rect 9602 23102 9614 23154
rect 10098 23102 10110 23154
rect 10162 23102 10174 23154
rect 12450 23102 12462 23154
rect 12514 23102 12526 23154
rect 12674 23102 12686 23154
rect 12738 23102 12750 23154
rect 13794 23102 13806 23154
rect 13858 23102 13870 23154
rect 2270 23090 2322 23102
rect 7758 23090 7810 23102
rect 8654 23090 8706 23102
rect 11342 23090 11394 23102
rect 14814 23090 14866 23102
rect 15822 23154 15874 23166
rect 15822 23090 15874 23102
rect 16158 23154 16210 23166
rect 16158 23090 16210 23102
rect 16718 23154 16770 23166
rect 21310 23154 21362 23166
rect 18162 23102 18174 23154
rect 18226 23102 18238 23154
rect 20850 23102 20862 23154
rect 20914 23102 20926 23154
rect 16718 23090 16770 23102
rect 21310 23090 21362 23102
rect 21982 23154 22034 23166
rect 21982 23090 22034 23102
rect 22542 23154 22594 23166
rect 22542 23090 22594 23102
rect 22878 23154 22930 23166
rect 22878 23090 22930 23102
rect 23102 23154 23154 23166
rect 23102 23090 23154 23102
rect 27582 23154 27634 23166
rect 27582 23090 27634 23102
rect 29710 23154 29762 23166
rect 29710 23090 29762 23102
rect 30718 23154 30770 23166
rect 30718 23090 30770 23102
rect 33966 23154 34018 23166
rect 33966 23090 34018 23102
rect 34414 23154 34466 23166
rect 34414 23090 34466 23102
rect 34638 23154 34690 23166
rect 40910 23154 40962 23166
rect 35298 23102 35310 23154
rect 35362 23102 35374 23154
rect 34638 23090 34690 23102
rect 40910 23090 40962 23102
rect 41246 23154 41298 23166
rect 41246 23090 41298 23102
rect 41582 23154 41634 23166
rect 41582 23090 41634 23102
rect 43038 23154 43090 23166
rect 43038 23090 43090 23102
rect 43710 23154 43762 23166
rect 43710 23090 43762 23102
rect 43934 23154 43986 23166
rect 43934 23090 43986 23102
rect 44270 23154 44322 23166
rect 44270 23090 44322 23102
rect 46398 23154 46450 23166
rect 54686 23154 54738 23166
rect 47394 23102 47406 23154
rect 47458 23102 47470 23154
rect 48178 23102 48190 23154
rect 48242 23102 48254 23154
rect 50418 23102 50430 23154
rect 50482 23102 50494 23154
rect 50866 23102 50878 23154
rect 50930 23102 50942 23154
rect 53554 23102 53566 23154
rect 53618 23102 53630 23154
rect 46398 23090 46450 23102
rect 54686 23090 54738 23102
rect 55246 23154 55298 23166
rect 55246 23090 55298 23102
rect 55470 23154 55522 23166
rect 57026 23102 57038 23154
rect 57090 23102 57102 23154
rect 55470 23090 55522 23102
rect 1822 23042 1874 23054
rect 1822 22978 1874 22990
rect 2830 23042 2882 23054
rect 18734 23042 18786 23054
rect 21758 23042 21810 23054
rect 4274 22990 4286 23042
rect 4338 22990 4350 23042
rect 10546 22990 10558 23042
rect 10610 22990 10622 23042
rect 12338 22990 12350 23042
rect 12402 22990 12414 23042
rect 14018 22990 14030 23042
rect 14082 22990 14094 23042
rect 20514 22990 20526 23042
rect 20578 22990 20590 23042
rect 2830 22978 2882 22990
rect 18734 22978 18786 22990
rect 21758 22978 21810 22990
rect 22766 23042 22818 23054
rect 22766 22978 22818 22990
rect 23550 23042 23602 23054
rect 23550 22978 23602 22990
rect 23774 23042 23826 23054
rect 23774 22978 23826 22990
rect 24670 23042 24722 23054
rect 24670 22978 24722 22990
rect 34526 23042 34578 23054
rect 42814 23042 42866 23054
rect 56702 23042 56754 23054
rect 38098 22990 38110 23042
rect 38162 22990 38174 23042
rect 50530 22990 50542 23042
rect 50594 22990 50606 23042
rect 52098 22990 52110 23042
rect 52162 22990 52174 23042
rect 57250 22990 57262 23042
rect 57314 22990 57326 23042
rect 34526 22978 34578 22990
rect 42814 22978 42866 22990
rect 56702 22978 56754 22990
rect 8766 22930 8818 22942
rect 8766 22866 8818 22878
rect 14926 22930 14978 22942
rect 14926 22866 14978 22878
rect 17838 22930 17890 22942
rect 17838 22866 17890 22878
rect 18174 22930 18226 22942
rect 51102 22930 51154 22942
rect 43362 22878 43374 22930
rect 43426 22878 43438 22930
rect 18174 22866 18226 22878
rect 51102 22866 51154 22878
rect 54462 22930 54514 22942
rect 54462 22866 54514 22878
rect 1344 22762 58576 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 58576 22762
rect 1344 22676 58576 22710
rect 8990 22594 9042 22606
rect 8990 22530 9042 22542
rect 12910 22594 12962 22606
rect 12910 22530 12962 22542
rect 13806 22594 13858 22606
rect 13806 22530 13858 22542
rect 22542 22594 22594 22606
rect 47854 22594 47906 22606
rect 28018 22542 28030 22594
rect 28082 22542 28094 22594
rect 49970 22542 49982 22594
rect 50034 22542 50046 22594
rect 56802 22542 56814 22594
rect 56866 22542 56878 22594
rect 22542 22530 22594 22542
rect 47854 22530 47906 22542
rect 5854 22482 5906 22494
rect 4498 22430 4510 22482
rect 4562 22430 4574 22482
rect 5854 22418 5906 22430
rect 14030 22482 14082 22494
rect 25118 22482 25170 22494
rect 23650 22430 23662 22482
rect 23714 22430 23726 22482
rect 14030 22418 14082 22430
rect 25118 22418 25170 22430
rect 26462 22482 26514 22494
rect 26462 22418 26514 22430
rect 29262 22482 29314 22494
rect 39566 22482 39618 22494
rect 37874 22430 37886 22482
rect 37938 22430 37950 22482
rect 29262 22418 29314 22430
rect 39566 22418 39618 22430
rect 41134 22482 41186 22494
rect 41134 22418 41186 22430
rect 42030 22482 42082 22494
rect 42030 22418 42082 22430
rect 45166 22482 45218 22494
rect 45166 22418 45218 22430
rect 47742 22482 47794 22494
rect 47742 22418 47794 22430
rect 50542 22482 50594 22494
rect 56578 22430 56590 22482
rect 56642 22430 56654 22482
rect 50542 22418 50594 22430
rect 21870 22370 21922 22382
rect 2482 22318 2494 22370
rect 2546 22318 2558 22370
rect 5058 22318 5070 22370
rect 5122 22318 5134 22370
rect 6738 22318 6750 22370
rect 6802 22318 6814 22370
rect 7634 22318 7646 22370
rect 7698 22318 7710 22370
rect 10658 22318 10670 22370
rect 10722 22318 10734 22370
rect 11666 22318 11678 22370
rect 11730 22318 11742 22370
rect 18162 22318 18174 22370
rect 18226 22318 18238 22370
rect 19058 22318 19070 22370
rect 19122 22318 19134 22370
rect 21870 22306 21922 22318
rect 22094 22370 22146 22382
rect 22094 22306 22146 22318
rect 22654 22370 22706 22382
rect 22654 22306 22706 22318
rect 23214 22370 23266 22382
rect 23214 22306 23266 22318
rect 25566 22370 25618 22382
rect 25566 22306 25618 22318
rect 26350 22370 26402 22382
rect 28254 22370 28306 22382
rect 27906 22318 27918 22370
rect 27970 22318 27982 22370
rect 26350 22306 26402 22318
rect 28254 22306 28306 22318
rect 30942 22370 30994 22382
rect 31726 22370 31778 22382
rect 31490 22318 31502 22370
rect 31554 22318 31566 22370
rect 30942 22306 30994 22318
rect 31726 22306 31778 22318
rect 32062 22370 32114 22382
rect 32062 22306 32114 22318
rect 34078 22370 34130 22382
rect 34078 22306 34130 22318
rect 34526 22370 34578 22382
rect 34526 22306 34578 22318
rect 35198 22370 35250 22382
rect 35198 22306 35250 22318
rect 35982 22370 36034 22382
rect 35982 22306 36034 22318
rect 36206 22370 36258 22382
rect 36206 22306 36258 22318
rect 36542 22370 36594 22382
rect 40462 22370 40514 22382
rect 45390 22370 45442 22382
rect 37426 22318 37438 22370
rect 37490 22318 37502 22370
rect 40002 22318 40014 22370
rect 40066 22318 40078 22370
rect 40898 22318 40910 22370
rect 40962 22318 40974 22370
rect 42578 22318 42590 22370
rect 42642 22318 42654 22370
rect 43586 22318 43598 22370
rect 43650 22318 43662 22370
rect 44818 22318 44830 22370
rect 44882 22318 44894 22370
rect 36542 22306 36594 22318
rect 40462 22306 40514 22318
rect 45390 22306 45442 22318
rect 46286 22370 46338 22382
rect 46286 22306 46338 22318
rect 47518 22370 47570 22382
rect 47518 22306 47570 22318
rect 50318 22370 50370 22382
rect 50318 22306 50370 22318
rect 51662 22370 51714 22382
rect 51662 22306 51714 22318
rect 51886 22370 51938 22382
rect 51886 22306 51938 22318
rect 52222 22370 52274 22382
rect 54910 22370 54962 22382
rect 53890 22318 53902 22370
rect 53954 22318 53966 22370
rect 54450 22318 54462 22370
rect 54514 22318 54526 22370
rect 52222 22306 52274 22318
rect 54910 22306 54962 22318
rect 55134 22370 55186 22382
rect 57150 22370 57202 22382
rect 56242 22318 56254 22370
rect 56306 22318 56318 22370
rect 56802 22318 56814 22370
rect 56866 22318 56878 22370
rect 57362 22318 57374 22370
rect 57426 22318 57438 22370
rect 55134 22306 55186 22318
rect 57150 22306 57202 22318
rect 22542 22258 22594 22270
rect 2706 22206 2718 22258
rect 2770 22206 2782 22258
rect 3602 22206 3614 22258
rect 3666 22206 3678 22258
rect 6626 22206 6638 22258
rect 6690 22206 6702 22258
rect 10546 22206 10558 22258
rect 10610 22206 10622 22258
rect 17938 22206 17950 22258
rect 18002 22206 18014 22258
rect 20402 22206 20414 22258
rect 20466 22206 20478 22258
rect 22542 22194 22594 22206
rect 23550 22258 23602 22270
rect 23550 22194 23602 22206
rect 24334 22258 24386 22270
rect 24334 22194 24386 22206
rect 24558 22258 24610 22270
rect 24558 22194 24610 22206
rect 26014 22258 26066 22270
rect 26014 22194 26066 22206
rect 26574 22258 26626 22270
rect 26574 22194 26626 22206
rect 28590 22258 28642 22270
rect 28590 22194 28642 22206
rect 33854 22258 33906 22270
rect 33854 22194 33906 22206
rect 34190 22258 34242 22270
rect 34190 22194 34242 22206
rect 34974 22258 35026 22270
rect 34974 22194 35026 22206
rect 36318 22258 36370 22270
rect 36318 22194 36370 22206
rect 36990 22258 37042 22270
rect 36990 22194 37042 22206
rect 41246 22258 41298 22270
rect 45950 22258 46002 22270
rect 43922 22206 43934 22258
rect 43986 22206 43998 22258
rect 41246 22194 41298 22206
rect 45950 22194 46002 22206
rect 46062 22258 46114 22270
rect 46062 22194 46114 22206
rect 51326 22258 51378 22270
rect 51326 22194 51378 22206
rect 51998 22258 52050 22270
rect 51998 22194 52050 22206
rect 52670 22258 52722 22270
rect 52670 22194 52722 22206
rect 53006 22258 53058 22270
rect 55470 22258 55522 22270
rect 53442 22206 53454 22258
rect 53506 22206 53518 22258
rect 53006 22194 53058 22206
rect 55470 22194 55522 22206
rect 23326 22146 23378 22158
rect 13458 22094 13470 22146
rect 13522 22094 13534 22146
rect 21522 22094 21534 22146
rect 21586 22094 21598 22146
rect 23326 22082 23378 22094
rect 23662 22146 23714 22158
rect 23662 22082 23714 22094
rect 24446 22146 24498 22158
rect 24446 22082 24498 22094
rect 27806 22146 27858 22158
rect 27806 22082 27858 22094
rect 31054 22146 31106 22158
rect 31054 22082 31106 22094
rect 31166 22146 31218 22158
rect 31166 22082 31218 22094
rect 31950 22146 32002 22158
rect 31950 22082 32002 22094
rect 34302 22146 34354 22158
rect 34302 22082 34354 22094
rect 35086 22146 35138 22158
rect 35086 22082 35138 22094
rect 47854 22146 47906 22158
rect 47854 22082 47906 22094
rect 51438 22146 51490 22158
rect 55134 22146 55186 22158
rect 54338 22094 54350 22146
rect 54402 22094 54414 22146
rect 51438 22082 51490 22094
rect 55134 22082 55186 22094
rect 1344 21978 58576 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 50558 21978
rect 50610 21926 50662 21978
rect 50714 21926 50766 21978
rect 50818 21926 58576 21978
rect 1344 21892 58576 21926
rect 1822 21810 1874 21822
rect 1822 21746 1874 21758
rect 9102 21810 9154 21822
rect 9102 21746 9154 21758
rect 11230 21810 11282 21822
rect 11790 21810 11842 21822
rect 11554 21758 11566 21810
rect 11618 21758 11630 21810
rect 11230 21746 11282 21758
rect 11790 21746 11842 21758
rect 12014 21810 12066 21822
rect 12014 21746 12066 21758
rect 33182 21810 33234 21822
rect 33182 21746 33234 21758
rect 33742 21810 33794 21822
rect 33742 21746 33794 21758
rect 34862 21810 34914 21822
rect 34862 21746 34914 21758
rect 38670 21810 38722 21822
rect 38670 21746 38722 21758
rect 39342 21810 39394 21822
rect 39342 21746 39394 21758
rect 39566 21810 39618 21822
rect 39566 21746 39618 21758
rect 39678 21810 39730 21822
rect 50990 21810 51042 21822
rect 41906 21758 41918 21810
rect 41970 21758 41982 21810
rect 47730 21758 47742 21810
rect 47794 21758 47806 21810
rect 49746 21758 49758 21810
rect 49810 21758 49822 21810
rect 39678 21746 39730 21758
rect 50990 21746 51042 21758
rect 51998 21810 52050 21822
rect 51998 21746 52050 21758
rect 53230 21810 53282 21822
rect 53230 21746 53282 21758
rect 54350 21810 54402 21822
rect 54674 21758 54686 21810
rect 54738 21758 54750 21810
rect 54350 21746 54402 21758
rect 16158 21698 16210 21710
rect 2034 21646 2046 21698
rect 2098 21646 2110 21698
rect 4274 21646 4286 21698
rect 4338 21646 4350 21698
rect 8194 21646 8206 21698
rect 8258 21646 8270 21698
rect 14466 21646 14478 21698
rect 14530 21646 14542 21698
rect 1698 21310 1710 21362
rect 1762 21359 1774 21362
rect 2049 21359 2095 21646
rect 16158 21634 16210 21646
rect 25678 21698 25730 21710
rect 25678 21634 25730 21646
rect 27022 21698 27074 21710
rect 27022 21634 27074 21646
rect 28590 21698 28642 21710
rect 35646 21698 35698 21710
rect 30258 21646 30270 21698
rect 30322 21646 30334 21698
rect 28590 21634 28642 21646
rect 35646 21634 35698 21646
rect 35870 21698 35922 21710
rect 35870 21634 35922 21646
rect 35982 21698 36034 21710
rect 35982 21634 36034 21646
rect 39902 21698 39954 21710
rect 45054 21698 45106 21710
rect 50766 21698 50818 21710
rect 41010 21646 41022 21698
rect 41074 21646 41086 21698
rect 46274 21646 46286 21698
rect 46338 21646 46350 21698
rect 39902 21634 39954 21646
rect 45054 21634 45106 21646
rect 50766 21634 50818 21646
rect 51886 21698 51938 21710
rect 51886 21634 51938 21646
rect 53006 21698 53058 21710
rect 53006 21634 53058 21646
rect 55918 21698 55970 21710
rect 56690 21646 56702 21698
rect 56754 21646 56766 21698
rect 55918 21634 55970 21646
rect 2270 21586 2322 21598
rect 2270 21522 2322 21534
rect 2494 21586 2546 21598
rect 2494 21522 2546 21534
rect 2718 21586 2770 21598
rect 2718 21522 2770 21534
rect 2830 21586 2882 21598
rect 8430 21586 8482 21598
rect 12126 21586 12178 21598
rect 27134 21586 27186 21598
rect 4498 21534 4510 21586
rect 4562 21534 4574 21586
rect 5618 21534 5630 21586
rect 5682 21534 5694 21586
rect 6850 21534 6862 21586
rect 6914 21534 6926 21586
rect 8642 21534 8654 21586
rect 8706 21534 8718 21586
rect 9426 21534 9438 21586
rect 9490 21534 9502 21586
rect 10322 21534 10334 21586
rect 10386 21534 10398 21586
rect 15474 21534 15486 21586
rect 15538 21534 15550 21586
rect 17602 21534 17614 21586
rect 17666 21534 17678 21586
rect 18722 21534 18734 21586
rect 18786 21534 18798 21586
rect 20290 21534 20302 21586
rect 20354 21534 20366 21586
rect 21298 21534 21310 21586
rect 21362 21534 21374 21586
rect 21746 21534 21758 21586
rect 21810 21534 21822 21586
rect 23538 21534 23550 21586
rect 23602 21534 23614 21586
rect 26338 21534 26350 21586
rect 26402 21534 26414 21586
rect 2830 21522 2882 21534
rect 8430 21522 8482 21534
rect 12126 21522 12178 21534
rect 27134 21522 27186 21534
rect 27470 21586 27522 21598
rect 33966 21586 34018 21598
rect 29474 21534 29486 21586
rect 29538 21534 29550 21586
rect 27470 21522 27522 21534
rect 33966 21522 34018 21534
rect 34414 21586 34466 21598
rect 34414 21522 34466 21534
rect 35086 21586 35138 21598
rect 35086 21522 35138 21534
rect 35534 21586 35586 21598
rect 35534 21522 35586 21534
rect 38558 21586 38610 21598
rect 38558 21522 38610 21534
rect 38894 21586 38946 21598
rect 38894 21522 38946 21534
rect 39006 21586 39058 21598
rect 39006 21522 39058 21534
rect 40238 21586 40290 21598
rect 52110 21586 52162 21598
rect 40898 21534 40910 21586
rect 40962 21534 40974 21586
rect 41794 21534 41806 21586
rect 41858 21534 41870 21586
rect 43698 21534 43710 21586
rect 43762 21534 43774 21586
rect 44370 21534 44382 21586
rect 44434 21534 44446 21586
rect 45266 21534 45278 21586
rect 45330 21534 45342 21586
rect 47282 21534 47294 21586
rect 47346 21534 47358 21586
rect 49522 21534 49534 21586
rect 49586 21534 49598 21586
rect 51202 21534 51214 21586
rect 51266 21534 51278 21586
rect 40238 21522 40290 21534
rect 52110 21522 52162 21534
rect 52558 21586 52610 21598
rect 52558 21522 52610 21534
rect 53566 21586 53618 21598
rect 54898 21534 54910 21586
rect 54962 21534 54974 21586
rect 55570 21534 55582 21586
rect 55634 21534 55646 21586
rect 56578 21534 56590 21586
rect 56642 21534 56654 21586
rect 57474 21534 57486 21586
rect 57538 21534 57550 21586
rect 53566 21522 53618 21534
rect 8094 21474 8146 21486
rect 12574 21474 12626 21486
rect 18174 21474 18226 21486
rect 24334 21474 24386 21486
rect 29150 21474 29202 21486
rect 33854 21474 33906 21486
rect 3266 21422 3278 21474
rect 3330 21422 3342 21474
rect 5170 21422 5182 21474
rect 5234 21422 5246 21474
rect 10098 21422 10110 21474
rect 10162 21422 10174 21474
rect 14018 21422 14030 21474
rect 14082 21422 14094 21474
rect 17714 21422 17726 21474
rect 17778 21422 17790 21474
rect 19170 21422 19182 21474
rect 19234 21422 19246 21474
rect 23650 21422 23662 21474
rect 23714 21422 23726 21474
rect 26002 21422 26014 21474
rect 26066 21422 26078 21474
rect 28690 21422 28702 21474
rect 28754 21422 28766 21474
rect 32386 21422 32398 21474
rect 32450 21422 32462 21474
rect 8094 21410 8146 21422
rect 12574 21410 12626 21422
rect 18174 21410 18226 21422
rect 24334 21410 24386 21422
rect 29150 21410 29202 21422
rect 33854 21410 33906 21422
rect 34974 21474 35026 21486
rect 34974 21410 35026 21422
rect 36430 21474 36482 21486
rect 36430 21410 36482 21422
rect 38334 21474 38386 21486
rect 38334 21410 38386 21422
rect 42478 21474 42530 21486
rect 45950 21474 46002 21486
rect 43922 21422 43934 21474
rect 43986 21422 43998 21474
rect 44594 21422 44606 21474
rect 44658 21422 44670 21474
rect 42478 21410 42530 21422
rect 45950 21410 46002 21422
rect 53342 21474 53394 21486
rect 55682 21422 55694 21474
rect 55746 21422 55758 21474
rect 56802 21422 56814 21474
rect 56866 21422 56878 21474
rect 53342 21410 53394 21422
rect 27694 21362 27746 21374
rect 28366 21362 28418 21374
rect 1762 21313 2095 21359
rect 1762 21310 1774 21313
rect 10434 21310 10446 21362
rect 10498 21310 10510 21362
rect 21746 21310 21758 21362
rect 21810 21310 21822 21362
rect 28018 21310 28030 21362
rect 28082 21310 28094 21362
rect 27694 21298 27746 21310
rect 28366 21298 28418 21310
rect 50654 21362 50706 21374
rect 50654 21298 50706 21310
rect 1344 21194 58576 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 58576 21194
rect 1344 21108 58576 21142
rect 7198 21026 7250 21038
rect 27470 21026 27522 21038
rect 15362 20974 15374 21026
rect 15426 21023 15438 21026
rect 15922 21023 15934 21026
rect 15426 20977 15934 21023
rect 15426 20974 15438 20977
rect 15922 20974 15934 20977
rect 15986 20974 15998 21026
rect 22866 20974 22878 21026
rect 22930 21023 22942 21026
rect 23426 21023 23438 21026
rect 22930 20977 23438 21023
rect 22930 20974 22942 20977
rect 23426 20974 23438 20977
rect 23490 20974 23502 21026
rect 7198 20962 7250 20974
rect 27470 20962 27522 20974
rect 36206 21026 36258 21038
rect 36206 20962 36258 20974
rect 44046 21026 44098 21038
rect 44046 20962 44098 20974
rect 46062 21026 46114 21038
rect 55806 21026 55858 21038
rect 51650 20974 51662 21026
rect 51714 20974 51726 21026
rect 46062 20962 46114 20974
rect 55806 20962 55858 20974
rect 2494 20914 2546 20926
rect 9102 20914 9154 20926
rect 13582 20914 13634 20926
rect 3266 20862 3278 20914
rect 3330 20862 3342 20914
rect 4834 20862 4846 20914
rect 4898 20862 4910 20914
rect 9874 20862 9886 20914
rect 9938 20862 9950 20914
rect 2494 20850 2546 20862
rect 9102 20850 9154 20862
rect 13582 20850 13634 20862
rect 15374 20914 15426 20926
rect 22878 20914 22930 20926
rect 27694 20914 27746 20926
rect 41358 20914 41410 20926
rect 57262 20914 57314 20926
rect 17266 20862 17278 20914
rect 17330 20862 17342 20914
rect 18610 20862 18622 20914
rect 18674 20862 18686 20914
rect 26002 20862 26014 20914
rect 26066 20862 26078 20914
rect 28018 20862 28030 20914
rect 28082 20862 28094 20914
rect 32498 20862 32510 20914
rect 32562 20862 32574 20914
rect 33618 20862 33630 20914
rect 33682 20862 33694 20914
rect 35746 20862 35758 20914
rect 35810 20862 35822 20914
rect 50418 20862 50430 20914
rect 50482 20862 50494 20914
rect 15374 20850 15426 20862
rect 22878 20850 22930 20862
rect 27694 20850 27746 20862
rect 41358 20850 41410 20862
rect 57262 20850 57314 20862
rect 1710 20802 1762 20814
rect 1710 20738 1762 20750
rect 3726 20802 3778 20814
rect 6190 20802 6242 20814
rect 4274 20750 4286 20802
rect 4338 20750 4350 20802
rect 3726 20738 3778 20750
rect 6190 20738 6242 20750
rect 6414 20802 6466 20814
rect 6414 20738 6466 20750
rect 6974 20802 7026 20814
rect 6974 20738 7026 20750
rect 7422 20802 7474 20814
rect 7422 20738 7474 20750
rect 7870 20802 7922 20814
rect 7870 20738 7922 20750
rect 8430 20802 8482 20814
rect 10894 20802 10946 20814
rect 22206 20802 22258 20814
rect 24558 20802 24610 20814
rect 36094 20802 36146 20814
rect 43374 20802 43426 20814
rect 46958 20802 47010 20814
rect 9314 20750 9326 20802
rect 9378 20750 9390 20802
rect 16818 20750 16830 20802
rect 16882 20750 16894 20802
rect 18050 20750 18062 20802
rect 18114 20750 18126 20802
rect 19058 20750 19070 20802
rect 19122 20750 19134 20802
rect 19394 20750 19406 20802
rect 19458 20750 19470 20802
rect 21746 20750 21758 20802
rect 21810 20750 21822 20802
rect 24210 20750 24222 20802
rect 24274 20750 24286 20802
rect 25218 20750 25230 20802
rect 25282 20750 25294 20802
rect 26898 20750 26910 20802
rect 26962 20750 26974 20802
rect 30706 20750 30718 20802
rect 30770 20750 30782 20802
rect 31266 20750 31278 20802
rect 31330 20750 31342 20802
rect 32386 20750 32398 20802
rect 32450 20750 32462 20802
rect 32834 20750 32846 20802
rect 32898 20750 32910 20802
rect 40002 20750 40014 20802
rect 40066 20750 40078 20802
rect 43698 20750 43710 20802
rect 43762 20750 43774 20802
rect 8430 20738 8482 20750
rect 10894 20738 10946 20750
rect 22206 20738 22258 20750
rect 24558 20738 24610 20750
rect 36094 20738 36146 20750
rect 43374 20738 43426 20750
rect 46958 20738 47010 20750
rect 49086 20802 49138 20814
rect 49086 20738 49138 20750
rect 51102 20802 51154 20814
rect 58158 20802 58210 20814
rect 56802 20750 56814 20802
rect 56866 20750 56878 20802
rect 57026 20750 57038 20802
rect 57090 20750 57102 20802
rect 51102 20738 51154 20750
rect 58158 20738 58210 20750
rect 2046 20690 2098 20702
rect 2046 20626 2098 20638
rect 3838 20690 3890 20702
rect 3838 20626 3890 20638
rect 8990 20690 9042 20702
rect 8990 20626 9042 20638
rect 9774 20690 9826 20702
rect 9774 20626 9826 20638
rect 10334 20690 10386 20702
rect 10334 20626 10386 20638
rect 10670 20690 10722 20702
rect 10670 20626 10722 20638
rect 11118 20690 11170 20702
rect 11118 20626 11170 20638
rect 11230 20690 11282 20702
rect 11230 20626 11282 20638
rect 11678 20690 11730 20702
rect 11678 20626 11730 20638
rect 12798 20690 12850 20702
rect 12798 20626 12850 20638
rect 12910 20690 12962 20702
rect 12910 20626 12962 20638
rect 21310 20690 21362 20702
rect 21310 20626 21362 20638
rect 27358 20690 27410 20702
rect 27358 20626 27410 20638
rect 27918 20690 27970 20702
rect 27918 20626 27970 20638
rect 29262 20690 29314 20702
rect 29262 20626 29314 20638
rect 29934 20690 29986 20702
rect 43934 20690 43986 20702
rect 31714 20638 31726 20690
rect 31778 20638 31790 20690
rect 32050 20638 32062 20690
rect 32114 20638 32126 20690
rect 39442 20638 39454 20690
rect 39506 20638 39518 20690
rect 41122 20638 41134 20690
rect 41186 20638 41198 20690
rect 29934 20626 29986 20638
rect 43934 20626 43986 20638
rect 45950 20690 46002 20702
rect 45950 20626 46002 20638
rect 46062 20690 46114 20702
rect 46062 20626 46114 20638
rect 46734 20690 46786 20702
rect 46734 20626 46786 20638
rect 47294 20690 47346 20702
rect 47294 20626 47346 20638
rect 49310 20690 49362 20702
rect 49310 20626 49362 20638
rect 49646 20690 49698 20702
rect 49646 20626 49698 20638
rect 50094 20690 50146 20702
rect 50094 20626 50146 20638
rect 50542 20690 50594 20702
rect 50542 20626 50594 20638
rect 50990 20690 51042 20702
rect 50990 20626 51042 20638
rect 51214 20690 51266 20702
rect 51214 20626 51266 20638
rect 55694 20690 55746 20702
rect 55694 20626 55746 20638
rect 55806 20690 55858 20702
rect 55806 20626 55858 20638
rect 57822 20690 57874 20702
rect 57822 20626 57874 20638
rect 2830 20578 2882 20590
rect 2830 20514 2882 20526
rect 4062 20578 4114 20590
rect 4062 20514 4114 20526
rect 4510 20578 4562 20590
rect 4510 20514 4562 20526
rect 4734 20578 4786 20590
rect 4734 20514 4786 20526
rect 4846 20578 4898 20590
rect 4846 20514 4898 20526
rect 5966 20578 6018 20590
rect 5966 20514 6018 20526
rect 6302 20578 6354 20590
rect 6302 20514 6354 20526
rect 8542 20578 8594 20590
rect 8542 20514 8594 20526
rect 8766 20578 8818 20590
rect 8766 20514 8818 20526
rect 9550 20578 9602 20590
rect 9550 20514 9602 20526
rect 9886 20578 9938 20590
rect 12686 20578 12738 20590
rect 12002 20526 12014 20578
rect 12066 20526 12078 20578
rect 9886 20514 9938 20526
rect 12686 20514 12738 20526
rect 15934 20578 15986 20590
rect 15934 20514 15986 20526
rect 23326 20578 23378 20590
rect 23326 20514 23378 20526
rect 27134 20578 27186 20590
rect 27134 20514 27186 20526
rect 29710 20578 29762 20590
rect 29710 20514 29762 20526
rect 29822 20578 29874 20590
rect 29822 20514 29874 20526
rect 36206 20578 36258 20590
rect 36206 20514 36258 20526
rect 37102 20578 37154 20590
rect 37102 20514 37154 20526
rect 46958 20578 47010 20590
rect 46958 20514 47010 20526
rect 48414 20578 48466 20590
rect 48414 20514 48466 20526
rect 48526 20578 48578 20590
rect 48526 20514 48578 20526
rect 48638 20578 48690 20590
rect 48638 20514 48690 20526
rect 50318 20578 50370 20590
rect 50318 20514 50370 20526
rect 1344 20410 58576 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 50558 20410
rect 50610 20358 50662 20410
rect 50714 20358 50766 20410
rect 50818 20358 58576 20410
rect 1344 20324 58576 20358
rect 6750 20242 6802 20254
rect 6750 20178 6802 20190
rect 24222 20242 24274 20254
rect 24222 20178 24274 20190
rect 31054 20242 31106 20254
rect 31054 20178 31106 20190
rect 33854 20242 33906 20254
rect 33854 20178 33906 20190
rect 40350 20242 40402 20254
rect 40350 20178 40402 20190
rect 56478 20242 56530 20254
rect 56478 20178 56530 20190
rect 58270 20242 58322 20254
rect 58270 20178 58322 20190
rect 5854 20130 5906 20142
rect 3266 20078 3278 20130
rect 3330 20078 3342 20130
rect 4946 20078 4958 20130
rect 5010 20078 5022 20130
rect 5854 20066 5906 20078
rect 7198 20130 7250 20142
rect 7198 20066 7250 20078
rect 7534 20130 7586 20142
rect 12462 20130 12514 20142
rect 10434 20078 10446 20130
rect 10498 20078 10510 20130
rect 7534 20066 7586 20078
rect 12462 20066 12514 20078
rect 12574 20130 12626 20142
rect 12574 20066 12626 20078
rect 13134 20130 13186 20142
rect 20078 20130 20130 20142
rect 23550 20130 23602 20142
rect 14466 20078 14478 20130
rect 14530 20078 14542 20130
rect 16482 20078 16494 20130
rect 16546 20078 16558 20130
rect 18162 20078 18174 20130
rect 18226 20078 18238 20130
rect 19282 20078 19294 20130
rect 19346 20078 19358 20130
rect 19618 20078 19630 20130
rect 19682 20078 19694 20130
rect 20402 20078 20414 20130
rect 20466 20078 20478 20130
rect 21186 20078 21198 20130
rect 21250 20078 21262 20130
rect 22866 20078 22878 20130
rect 22930 20078 22942 20130
rect 13134 20066 13186 20078
rect 20078 20066 20130 20078
rect 23550 20066 23602 20078
rect 24446 20130 24498 20142
rect 29374 20130 29426 20142
rect 25554 20078 25566 20130
rect 25618 20078 25630 20130
rect 28242 20078 28254 20130
rect 28306 20078 28318 20130
rect 24446 20066 24498 20078
rect 29374 20066 29426 20078
rect 29822 20130 29874 20142
rect 29822 20066 29874 20078
rect 30270 20130 30322 20142
rect 30270 20066 30322 20078
rect 31502 20130 31554 20142
rect 31502 20066 31554 20078
rect 31614 20130 31666 20142
rect 31614 20066 31666 20078
rect 32622 20130 32674 20142
rect 37774 20130 37826 20142
rect 40910 20130 40962 20142
rect 35186 20078 35198 20130
rect 35250 20078 35262 20130
rect 39778 20078 39790 20130
rect 39842 20127 39854 20130
rect 40114 20127 40126 20130
rect 39842 20081 40126 20127
rect 39842 20078 39854 20081
rect 40114 20078 40126 20081
rect 40178 20078 40190 20130
rect 32622 20066 32674 20078
rect 37774 20066 37826 20078
rect 40910 20066 40962 20078
rect 42478 20130 42530 20142
rect 42478 20066 42530 20078
rect 42926 20130 42978 20142
rect 42926 20066 42978 20078
rect 43822 20130 43874 20142
rect 43822 20066 43874 20078
rect 48750 20130 48802 20142
rect 48750 20066 48802 20078
rect 51326 20130 51378 20142
rect 56702 20130 56754 20142
rect 52882 20078 52894 20130
rect 52946 20078 52958 20130
rect 51326 20066 51378 20078
rect 56702 20066 56754 20078
rect 2606 20018 2658 20030
rect 6862 20018 6914 20030
rect 12238 20018 12290 20030
rect 2146 19966 2158 20018
rect 2210 19966 2222 20018
rect 3714 19966 3726 20018
rect 3778 19966 3790 20018
rect 5058 19966 5070 20018
rect 5122 19966 5134 20018
rect 6514 19966 6526 20018
rect 6578 19966 6590 20018
rect 9538 19966 9550 20018
rect 9602 19966 9614 20018
rect 10322 19966 10334 20018
rect 10386 19966 10398 20018
rect 11330 19966 11342 20018
rect 11394 19966 11406 20018
rect 2606 19954 2658 19966
rect 6862 19954 6914 19966
rect 12238 19954 12290 19966
rect 12910 20018 12962 20030
rect 24558 20018 24610 20030
rect 13458 19966 13470 20018
rect 13522 19966 13534 20018
rect 15362 19966 15374 20018
rect 15426 19966 15438 20018
rect 17378 19966 17390 20018
rect 17442 19966 17454 20018
rect 18386 19966 18398 20018
rect 18450 19966 18462 20018
rect 18946 19966 18958 20018
rect 19010 19966 19022 20018
rect 21634 19966 21646 20018
rect 21698 19966 21710 20018
rect 23090 19966 23102 20018
rect 23154 19966 23166 20018
rect 12910 19954 12962 19966
rect 24558 19954 24610 19966
rect 25230 20018 25282 20030
rect 29710 20018 29762 20030
rect 27458 19966 27470 20018
rect 27522 19966 27534 20018
rect 28130 19966 28142 20018
rect 28194 19966 28206 20018
rect 25230 19954 25282 19966
rect 29710 19954 29762 19966
rect 30046 20018 30098 20030
rect 30718 20018 30770 20030
rect 33070 20018 33122 20030
rect 40238 20018 40290 20030
rect 42366 20018 42418 20030
rect 30482 19966 30494 20018
rect 30546 19966 30558 20018
rect 30818 19966 30830 20018
rect 30882 19966 30894 20018
rect 33282 19966 33294 20018
rect 33346 19966 33358 20018
rect 33842 19966 33854 20018
rect 33906 19966 33918 20018
rect 34402 19966 34414 20018
rect 34466 19966 34478 20018
rect 41346 19966 41358 20018
rect 41410 19966 41422 20018
rect 30046 19954 30098 19966
rect 30718 19954 30770 19966
rect 33070 19954 33122 19966
rect 40238 19954 40290 19966
rect 42366 19954 42418 19966
rect 42702 20018 42754 20030
rect 43486 20018 43538 20030
rect 43138 19966 43150 20018
rect 43202 19966 43214 20018
rect 42702 19954 42754 19966
rect 43486 19954 43538 19966
rect 43598 20018 43650 20030
rect 43598 19954 43650 19966
rect 43934 20018 43986 20030
rect 43934 19954 43986 19966
rect 44158 20018 44210 20030
rect 44158 19954 44210 19966
rect 49086 20018 49138 20030
rect 50878 20018 50930 20030
rect 49298 19966 49310 20018
rect 49362 19966 49374 20018
rect 49086 19954 49138 19966
rect 50878 19954 50930 19966
rect 51102 20018 51154 20030
rect 51102 19954 51154 19966
rect 51550 20018 51602 20030
rect 56814 20018 56866 20030
rect 53106 19966 53118 20018
rect 53170 19966 53182 20018
rect 54226 19966 54238 20018
rect 54290 19966 54302 20018
rect 55010 19966 55022 20018
rect 55074 19966 55086 20018
rect 51550 19954 51602 19966
rect 56814 19954 56866 19966
rect 12014 19906 12066 19918
rect 9986 19854 9998 19906
rect 10050 19854 10062 19906
rect 11554 19854 11566 19906
rect 11618 19854 11630 19906
rect 12014 19842 12066 19854
rect 13022 19906 13074 19918
rect 43262 19906 43314 19918
rect 14018 19854 14030 19906
rect 14082 19854 14094 19906
rect 17826 19854 17838 19906
rect 17890 19854 17902 19906
rect 28018 19854 28030 19906
rect 28082 19854 28094 19906
rect 37314 19854 37326 19906
rect 37378 19854 37390 19906
rect 41682 19854 41694 19906
rect 41746 19854 41758 19906
rect 13022 19842 13074 19854
rect 43262 19842 43314 19854
rect 53790 19906 53842 19918
rect 54786 19854 54798 19906
rect 54850 19854 54862 19906
rect 53790 19842 53842 19854
rect 31726 19794 31778 19806
rect 48862 19794 48914 19806
rect 28914 19742 28926 19794
rect 28978 19791 28990 19794
rect 29474 19791 29486 19794
rect 28978 19745 29486 19791
rect 28978 19742 28990 19745
rect 29474 19742 29486 19745
rect 29538 19742 29550 19794
rect 33618 19742 33630 19794
rect 33682 19742 33694 19794
rect 31726 19730 31778 19742
rect 48862 19730 48914 19742
rect 1344 19626 58576 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 58576 19626
rect 1344 19540 58576 19574
rect 4622 19458 4674 19470
rect 4622 19394 4674 19406
rect 27806 19458 27858 19470
rect 27806 19394 27858 19406
rect 33070 19458 33122 19470
rect 33070 19394 33122 19406
rect 42366 19458 42418 19470
rect 42366 19394 42418 19406
rect 42814 19458 42866 19470
rect 42814 19394 42866 19406
rect 46286 19458 46338 19470
rect 46286 19394 46338 19406
rect 47518 19458 47570 19470
rect 47518 19394 47570 19406
rect 53006 19458 53058 19470
rect 53006 19394 53058 19406
rect 54126 19458 54178 19470
rect 55794 19406 55806 19458
rect 55858 19406 55870 19458
rect 54126 19394 54178 19406
rect 4958 19346 5010 19358
rect 14254 19346 14306 19358
rect 33630 19346 33682 19358
rect 10546 19294 10558 19346
rect 10610 19294 10622 19346
rect 11330 19294 11342 19346
rect 11394 19294 11406 19346
rect 17042 19294 17054 19346
rect 17106 19294 17118 19346
rect 17938 19294 17950 19346
rect 18002 19294 18014 19346
rect 19618 19294 19630 19346
rect 19682 19294 19694 19346
rect 21410 19294 21422 19346
rect 21474 19294 21486 19346
rect 23650 19294 23662 19346
rect 23714 19294 23726 19346
rect 29586 19294 29598 19346
rect 29650 19294 29662 19346
rect 4958 19282 5010 19294
rect 14254 19282 14306 19294
rect 33630 19282 33682 19294
rect 36990 19346 37042 19358
rect 38334 19346 38386 19358
rect 37426 19294 37438 19346
rect 37490 19294 37502 19346
rect 36990 19282 37042 19294
rect 38334 19282 38386 19294
rect 40574 19346 40626 19358
rect 40574 19282 40626 19294
rect 41022 19346 41074 19358
rect 41022 19282 41074 19294
rect 45278 19346 45330 19358
rect 45278 19282 45330 19294
rect 46622 19346 46674 19358
rect 46622 19282 46674 19294
rect 47182 19346 47234 19358
rect 51214 19346 51266 19358
rect 54910 19346 54962 19358
rect 50418 19294 50430 19346
rect 50482 19294 50494 19346
rect 54450 19294 54462 19346
rect 54514 19294 54526 19346
rect 47182 19282 47234 19294
rect 51214 19282 51266 19294
rect 54910 19282 54962 19294
rect 3950 19234 4002 19246
rect 1810 19182 1822 19234
rect 1874 19182 1886 19234
rect 3602 19182 3614 19234
rect 3666 19182 3678 19234
rect 3950 19170 4002 19182
rect 4398 19234 4450 19246
rect 6302 19234 6354 19246
rect 25006 19234 25058 19246
rect 6066 19182 6078 19234
rect 6130 19182 6142 19234
rect 6850 19182 6862 19234
rect 6914 19182 6926 19234
rect 8306 19182 8318 19234
rect 8370 19182 8382 19234
rect 8866 19182 8878 19234
rect 8930 19182 8942 19234
rect 10098 19182 10110 19234
rect 10162 19182 10174 19234
rect 11218 19182 11230 19234
rect 11282 19182 11294 19234
rect 14466 19182 14478 19234
rect 14530 19182 14542 19234
rect 16482 19182 16494 19234
rect 16546 19182 16558 19234
rect 18498 19182 18510 19234
rect 18562 19182 18574 19234
rect 19506 19182 19518 19234
rect 19570 19182 19582 19234
rect 20514 19182 20526 19234
rect 20578 19182 20590 19234
rect 21634 19182 21646 19234
rect 21698 19182 21710 19234
rect 22866 19182 22878 19234
rect 22930 19182 22942 19234
rect 24770 19182 24782 19234
rect 24834 19182 24846 19234
rect 4398 19170 4450 19182
rect 6302 19170 6354 19182
rect 25006 19170 25058 19182
rect 26014 19234 26066 19246
rect 26014 19170 26066 19182
rect 26126 19234 26178 19246
rect 28030 19234 28082 19246
rect 32734 19234 32786 19246
rect 39230 19234 39282 19246
rect 42590 19234 42642 19246
rect 43710 19234 43762 19246
rect 27570 19182 27582 19234
rect 27634 19182 27646 19234
rect 29138 19182 29150 19234
rect 29202 19182 29214 19234
rect 30034 19182 30046 19234
rect 30098 19182 30110 19234
rect 31602 19182 31614 19234
rect 31666 19182 31678 19234
rect 32162 19182 32174 19234
rect 32226 19182 32238 19234
rect 37650 19182 37662 19234
rect 37714 19182 37726 19234
rect 38770 19182 38782 19234
rect 38834 19182 38846 19234
rect 42018 19182 42030 19234
rect 42082 19182 42094 19234
rect 43474 19182 43486 19234
rect 43538 19182 43550 19234
rect 26126 19170 26178 19182
rect 28030 19170 28082 19182
rect 32734 19170 32786 19182
rect 39230 19170 39282 19182
rect 42590 19170 42642 19182
rect 43710 19170 43762 19182
rect 45166 19234 45218 19246
rect 45166 19170 45218 19182
rect 48414 19234 48466 19246
rect 53342 19234 53394 19246
rect 49634 19182 49646 19234
rect 49698 19182 49710 19234
rect 50754 19182 50766 19234
rect 50818 19182 50830 19234
rect 48414 19170 48466 19182
rect 53342 19170 53394 19182
rect 53902 19234 53954 19246
rect 57150 19234 57202 19246
rect 56130 19182 56142 19234
rect 56194 19182 56206 19234
rect 57474 19182 57486 19234
rect 57538 19182 57550 19234
rect 53902 19170 53954 19182
rect 57150 19170 57202 19182
rect 2046 19122 2098 19134
rect 2046 19058 2098 19070
rect 2382 19122 2434 19134
rect 2382 19058 2434 19070
rect 2718 19122 2770 19134
rect 2718 19058 2770 19070
rect 4062 19122 4114 19134
rect 4062 19058 4114 19070
rect 5742 19122 5794 19134
rect 5742 19058 5794 19070
rect 6414 19122 6466 19134
rect 6414 19058 6466 19070
rect 15038 19122 15090 19134
rect 25230 19122 25282 19134
rect 16594 19070 16606 19122
rect 16658 19070 16670 19122
rect 18722 19070 18734 19122
rect 18786 19070 18798 19122
rect 19730 19070 19742 19122
rect 19794 19070 19806 19122
rect 20402 19070 20414 19122
rect 20466 19070 20478 19122
rect 20738 19070 20750 19122
rect 20802 19070 20814 19122
rect 15038 19058 15090 19070
rect 25230 19058 25282 19070
rect 25566 19122 25618 19134
rect 25566 19058 25618 19070
rect 25790 19122 25842 19134
rect 25790 19058 25842 19070
rect 26686 19122 26738 19134
rect 32510 19122 32562 19134
rect 29250 19070 29262 19122
rect 29314 19070 29326 19122
rect 31490 19070 31502 19122
rect 31554 19070 31566 19122
rect 26686 19058 26738 19070
rect 32510 19058 32562 19070
rect 41806 19122 41858 19134
rect 41806 19058 41858 19070
rect 43822 19122 43874 19134
rect 46846 19122 46898 19134
rect 44258 19070 44270 19122
rect 44322 19070 44334 19122
rect 43822 19058 43874 19070
rect 46846 19058 46898 19070
rect 49422 19122 49474 19134
rect 49422 19058 49474 19070
rect 53566 19122 53618 19134
rect 53566 19058 53618 19070
rect 54798 19122 54850 19134
rect 54798 19058 54850 19070
rect 55022 19122 55074 19134
rect 55022 19058 55074 19070
rect 15934 19010 15986 19022
rect 15934 18946 15986 18958
rect 17502 19010 17554 19022
rect 17502 18946 17554 18958
rect 26798 19010 26850 19022
rect 26798 18946 26850 18958
rect 27022 19010 27074 19022
rect 27022 18946 27074 18958
rect 27694 19010 27746 19022
rect 40014 19010 40066 19022
rect 32050 18958 32062 19010
rect 32114 18958 32126 19010
rect 39666 18958 39678 19010
rect 39730 18958 39742 19010
rect 27694 18946 27746 18958
rect 40014 18946 40066 18958
rect 42254 19010 42306 19022
rect 44942 19010 44994 19022
rect 43138 18958 43150 19010
rect 43202 18958 43214 19010
rect 42254 18946 42306 18958
rect 44942 18946 44994 18958
rect 45390 19010 45442 19022
rect 45390 18946 45442 18958
rect 47406 19010 47458 19022
rect 47406 18946 47458 18958
rect 48526 19010 48578 19022
rect 48526 18946 48578 18958
rect 48750 19010 48802 19022
rect 48750 18946 48802 18958
rect 1344 18842 58576 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 50558 18842
rect 50610 18790 50662 18842
rect 50714 18790 50766 18842
rect 50818 18790 58576 18842
rect 1344 18756 58576 18790
rect 3390 18674 3442 18686
rect 3390 18610 3442 18622
rect 3726 18674 3778 18686
rect 15822 18674 15874 18686
rect 4050 18622 4062 18674
rect 4114 18622 4126 18674
rect 14242 18622 14254 18674
rect 14306 18622 14318 18674
rect 3726 18610 3778 18622
rect 15822 18610 15874 18622
rect 24558 18674 24610 18686
rect 24558 18610 24610 18622
rect 26574 18674 26626 18686
rect 26574 18610 26626 18622
rect 28590 18674 28642 18686
rect 28590 18610 28642 18622
rect 28814 18674 28866 18686
rect 28814 18610 28866 18622
rect 31390 18674 31442 18686
rect 31390 18610 31442 18622
rect 31502 18674 31554 18686
rect 33294 18674 33346 18686
rect 32386 18622 32398 18674
rect 32450 18622 32462 18674
rect 31502 18610 31554 18622
rect 33294 18610 33346 18622
rect 35422 18674 35474 18686
rect 35422 18610 35474 18622
rect 35870 18674 35922 18686
rect 35870 18610 35922 18622
rect 37214 18674 37266 18686
rect 42366 18674 42418 18686
rect 39106 18622 39118 18674
rect 39170 18622 39182 18674
rect 44930 18622 44942 18674
rect 44994 18622 45006 18674
rect 37214 18610 37266 18622
rect 42366 18610 42418 18622
rect 2046 18562 2098 18574
rect 3054 18562 3106 18574
rect 15150 18562 15202 18574
rect 2706 18510 2718 18562
rect 2770 18510 2782 18562
rect 6962 18510 6974 18562
rect 7026 18510 7038 18562
rect 10882 18510 10894 18562
rect 10946 18510 10958 18562
rect 13122 18510 13134 18562
rect 13186 18510 13198 18562
rect 2046 18498 2098 18510
rect 3054 18498 3106 18510
rect 15150 18498 15202 18510
rect 15710 18562 15762 18574
rect 15710 18498 15762 18510
rect 16830 18562 16882 18574
rect 24446 18562 24498 18574
rect 30494 18562 30546 18574
rect 18050 18510 18062 18562
rect 18114 18510 18126 18562
rect 21074 18510 21086 18562
rect 21138 18510 21150 18562
rect 23202 18510 23214 18562
rect 23266 18510 23278 18562
rect 23650 18510 23662 18562
rect 23714 18510 23726 18562
rect 26898 18510 26910 18562
rect 26962 18510 26974 18562
rect 27682 18510 27694 18562
rect 27746 18510 27758 18562
rect 16830 18498 16882 18510
rect 24446 18498 24498 18510
rect 30494 18498 30546 18510
rect 31278 18562 31330 18574
rect 36990 18562 37042 18574
rect 44158 18562 44210 18574
rect 35074 18510 35086 18562
rect 35138 18510 35150 18562
rect 37874 18510 37886 18562
rect 37938 18510 37950 18562
rect 39890 18510 39902 18562
rect 39954 18510 39966 18562
rect 31278 18498 31330 18510
rect 36990 18498 37042 18510
rect 44158 18498 44210 18510
rect 44270 18562 44322 18574
rect 47182 18562 47234 18574
rect 54126 18562 54178 18574
rect 46162 18510 46174 18562
rect 46226 18510 46238 18562
rect 51538 18510 51550 18562
rect 51602 18510 51614 18562
rect 44270 18498 44322 18510
rect 47182 18498 47234 18510
rect 54126 18498 54178 18510
rect 56590 18562 56642 18574
rect 56590 18498 56642 18510
rect 4510 18450 4562 18462
rect 1810 18398 1822 18450
rect 1874 18398 1886 18450
rect 2482 18398 2494 18450
rect 2546 18398 2558 18450
rect 4510 18386 4562 18398
rect 4734 18450 4786 18462
rect 4734 18386 4786 18398
rect 5070 18450 5122 18462
rect 5070 18386 5122 18398
rect 5294 18450 5346 18462
rect 5294 18386 5346 18398
rect 5518 18450 5570 18462
rect 9102 18450 9154 18462
rect 13694 18450 13746 18462
rect 5842 18398 5854 18450
rect 5906 18398 5918 18450
rect 7746 18398 7758 18450
rect 7810 18398 7822 18450
rect 11890 18398 11902 18450
rect 11954 18398 11966 18450
rect 13458 18398 13470 18450
rect 13522 18398 13534 18450
rect 5518 18386 5570 18398
rect 9102 18386 9154 18398
rect 13694 18386 13746 18398
rect 13806 18450 13858 18462
rect 13806 18386 13858 18398
rect 14590 18450 14642 18462
rect 14590 18386 14642 18398
rect 14814 18450 14866 18462
rect 14814 18386 14866 18398
rect 16046 18450 16098 18462
rect 16494 18450 16546 18462
rect 16258 18398 16270 18450
rect 16322 18398 16334 18450
rect 16046 18386 16098 18398
rect 16494 18386 16546 18398
rect 16718 18450 16770 18462
rect 24782 18450 24834 18462
rect 26238 18450 26290 18462
rect 28254 18450 28306 18462
rect 19282 18398 19294 18450
rect 19346 18398 19358 18450
rect 20962 18398 20974 18450
rect 21026 18398 21038 18450
rect 22754 18398 22766 18450
rect 22818 18398 22830 18450
rect 23874 18398 23886 18450
rect 23938 18398 23950 18450
rect 25666 18398 25678 18450
rect 25730 18398 25742 18450
rect 26002 18398 26014 18450
rect 26066 18398 26078 18450
rect 27458 18398 27470 18450
rect 27522 18398 27534 18450
rect 16718 18386 16770 18398
rect 24782 18386 24834 18398
rect 26238 18386 26290 18398
rect 28254 18386 28306 18398
rect 28926 18450 28978 18462
rect 28926 18386 28978 18398
rect 30606 18450 30658 18462
rect 30606 18386 30658 18398
rect 30830 18450 30882 18462
rect 30830 18386 30882 18398
rect 35982 18450 36034 18462
rect 37426 18398 37438 18450
rect 37490 18398 37502 18450
rect 38322 18398 38334 18450
rect 38386 18398 38398 18450
rect 38882 18398 38894 18450
rect 38946 18398 38958 18450
rect 40226 18398 40238 18450
rect 40290 18398 40302 18450
rect 41122 18398 41134 18450
rect 41186 18398 41198 18450
rect 42130 18398 42142 18450
rect 42194 18398 42206 18450
rect 43138 18398 43150 18450
rect 43202 18398 43214 18450
rect 45266 18398 45278 18450
rect 45330 18398 45342 18450
rect 47394 18398 47406 18450
rect 47458 18398 47470 18450
rect 47730 18398 47742 18450
rect 47794 18398 47806 18450
rect 48962 18398 48974 18450
rect 49026 18398 49038 18450
rect 50306 18398 50318 18450
rect 50370 18398 50382 18450
rect 52210 18398 52222 18450
rect 52274 18398 52286 18450
rect 53554 18398 53566 18450
rect 53618 18398 53630 18450
rect 54562 18398 54574 18450
rect 54626 18398 54638 18450
rect 57138 18398 57150 18450
rect 57202 18398 57214 18450
rect 35982 18386 36034 18398
rect 4846 18338 4898 18350
rect 15038 18338 15090 18350
rect 31838 18338 31890 18350
rect 6290 18286 6302 18338
rect 6354 18286 6366 18338
rect 10322 18286 10334 18338
rect 10386 18286 10398 18338
rect 17826 18286 17838 18338
rect 17890 18286 17902 18338
rect 20626 18286 20638 18338
rect 20690 18286 20702 18338
rect 4846 18274 4898 18286
rect 15038 18274 15090 18286
rect 31838 18274 31890 18286
rect 36430 18338 36482 18350
rect 36430 18274 36482 18286
rect 37326 18338 37378 18350
rect 41470 18338 41522 18350
rect 37874 18286 37886 18338
rect 37938 18286 37950 18338
rect 40338 18286 40350 18338
rect 40402 18286 40414 18338
rect 37326 18274 37378 18286
rect 41470 18274 41522 18286
rect 41694 18338 41746 18350
rect 41694 18274 41746 18286
rect 42702 18338 42754 18350
rect 46622 18338 46674 18350
rect 43026 18286 43038 18338
rect 43090 18286 43102 18338
rect 49074 18286 49086 18338
rect 49138 18286 49150 18338
rect 53442 18286 53454 18338
rect 53506 18286 53518 18338
rect 55010 18286 55022 18338
rect 55074 18286 55086 18338
rect 57474 18286 57486 18338
rect 57538 18286 57550 18338
rect 42702 18274 42754 18286
rect 46622 18274 46674 18286
rect 30494 18226 30546 18238
rect 30494 18162 30546 18174
rect 32062 18226 32114 18238
rect 32062 18162 32114 18174
rect 35870 18226 35922 18238
rect 35870 18162 35922 18174
rect 44158 18226 44210 18238
rect 50530 18174 50542 18226
rect 50594 18174 50606 18226
rect 44158 18162 44210 18174
rect 1344 18058 58576 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 58576 18058
rect 1344 17972 58576 18006
rect 9438 17890 9490 17902
rect 9438 17826 9490 17838
rect 9550 17890 9602 17902
rect 9550 17826 9602 17838
rect 14030 17890 14082 17902
rect 29262 17890 29314 17902
rect 37550 17890 37602 17902
rect 26114 17838 26126 17890
rect 26178 17838 26190 17890
rect 31490 17838 31502 17890
rect 31554 17838 31566 17890
rect 34850 17838 34862 17890
rect 34914 17838 34926 17890
rect 14030 17826 14082 17838
rect 29262 17826 29314 17838
rect 37550 17826 37602 17838
rect 5742 17778 5794 17790
rect 8654 17778 8706 17790
rect 6514 17726 6526 17778
rect 6578 17726 6590 17778
rect 5742 17714 5794 17726
rect 8654 17714 8706 17726
rect 10558 17778 10610 17790
rect 10558 17714 10610 17726
rect 12574 17778 12626 17790
rect 15934 17778 15986 17790
rect 15138 17726 15150 17778
rect 15202 17726 15214 17778
rect 12574 17714 12626 17726
rect 15934 17714 15986 17726
rect 20862 17778 20914 17790
rect 32734 17778 32786 17790
rect 42254 17778 42306 17790
rect 23314 17726 23326 17778
rect 23378 17726 23390 17778
rect 29698 17726 29710 17778
rect 29762 17726 29774 17778
rect 31154 17726 31166 17778
rect 31218 17726 31230 17778
rect 34290 17726 34302 17778
rect 34354 17726 34366 17778
rect 40786 17726 40798 17778
rect 40850 17726 40862 17778
rect 20862 17714 20914 17726
rect 32734 17714 32786 17726
rect 42254 17714 42306 17726
rect 45166 17778 45218 17790
rect 48526 17778 48578 17790
rect 47282 17726 47294 17778
rect 47346 17726 47358 17778
rect 45166 17714 45218 17726
rect 48526 17714 48578 17726
rect 55582 17778 55634 17790
rect 55582 17714 55634 17726
rect 1710 17666 1762 17678
rect 1710 17602 1762 17614
rect 3054 17666 3106 17678
rect 9214 17666 9266 17678
rect 19182 17666 19234 17678
rect 3938 17614 3950 17666
rect 4002 17614 4014 17666
rect 7970 17614 7982 17666
rect 8034 17614 8046 17666
rect 8978 17614 8990 17666
rect 9042 17614 9054 17666
rect 11890 17614 11902 17666
rect 11954 17614 11966 17666
rect 13458 17614 13470 17666
rect 13522 17614 13534 17666
rect 13682 17614 13694 17666
rect 13746 17614 13758 17666
rect 14466 17614 14478 17666
rect 14530 17614 14542 17666
rect 15474 17614 15486 17666
rect 15538 17614 15550 17666
rect 17154 17614 17166 17666
rect 17218 17614 17230 17666
rect 18610 17614 18622 17666
rect 18674 17614 18686 17666
rect 3054 17602 3106 17614
rect 9214 17602 9266 17614
rect 19182 17602 19234 17614
rect 19294 17666 19346 17678
rect 21646 17666 21698 17678
rect 22206 17666 22258 17678
rect 33070 17666 33122 17678
rect 19618 17614 19630 17666
rect 19682 17614 19694 17666
rect 21970 17614 21982 17666
rect 22034 17614 22046 17666
rect 22866 17614 22878 17666
rect 22930 17614 22942 17666
rect 24434 17614 24446 17666
rect 24498 17614 24510 17666
rect 25442 17614 25454 17666
rect 25506 17614 25518 17666
rect 25778 17614 25790 17666
rect 25842 17614 25854 17666
rect 29250 17614 29262 17666
rect 29314 17614 29326 17666
rect 29810 17614 29822 17666
rect 29874 17614 29886 17666
rect 31042 17614 31054 17666
rect 31106 17614 31118 17666
rect 19294 17602 19346 17614
rect 21646 17602 21698 17614
rect 22206 17602 22258 17614
rect 33070 17602 33122 17614
rect 33518 17666 33570 17678
rect 35646 17666 35698 17678
rect 38558 17666 38610 17678
rect 50878 17666 50930 17678
rect 34514 17614 34526 17666
rect 34578 17614 34590 17666
rect 35298 17614 35310 17666
rect 35362 17614 35374 17666
rect 35970 17614 35982 17666
rect 36034 17614 36046 17666
rect 38770 17614 38782 17666
rect 38834 17614 38846 17666
rect 40338 17614 40350 17666
rect 40402 17614 40414 17666
rect 41346 17614 41358 17666
rect 41410 17614 41422 17666
rect 42466 17614 42478 17666
rect 42530 17614 42542 17666
rect 45826 17614 45838 17666
rect 45890 17614 45902 17666
rect 56130 17614 56142 17666
rect 56194 17614 56206 17666
rect 57138 17614 57150 17666
rect 57202 17614 57214 17666
rect 33518 17602 33570 17614
rect 35646 17602 35698 17614
rect 38558 17602 38610 17614
rect 50878 17602 50930 17614
rect 2046 17554 2098 17566
rect 2046 17490 2098 17502
rect 2382 17554 2434 17566
rect 2382 17490 2434 17502
rect 2718 17554 2770 17566
rect 4510 17554 4562 17566
rect 14254 17554 14306 17566
rect 21310 17554 21362 17566
rect 3378 17502 3390 17554
rect 3442 17502 3454 17554
rect 4834 17502 4846 17554
rect 4898 17502 4910 17554
rect 6962 17502 6974 17554
rect 7026 17502 7038 17554
rect 10882 17502 10894 17554
rect 10946 17502 10958 17554
rect 17266 17502 17278 17554
rect 17330 17502 17342 17554
rect 19730 17502 19742 17554
rect 19794 17502 19806 17554
rect 20514 17502 20526 17554
rect 20578 17502 20590 17554
rect 2718 17490 2770 17502
rect 4510 17490 4562 17502
rect 14254 17490 14306 17502
rect 21310 17490 21362 17502
rect 22318 17554 22370 17566
rect 22318 17490 22370 17502
rect 37438 17554 37490 17566
rect 50990 17554 51042 17566
rect 46834 17502 46846 17554
rect 46898 17502 46910 17554
rect 48738 17502 48750 17554
rect 48802 17502 48814 17554
rect 50306 17502 50318 17554
rect 50370 17502 50382 17554
rect 57362 17502 57374 17554
rect 57426 17502 57438 17554
rect 37438 17490 37490 17502
rect 50990 17490 51042 17502
rect 13918 17442 13970 17454
rect 4162 17390 4174 17442
rect 4226 17390 4238 17442
rect 13918 17378 13970 17390
rect 16046 17442 16098 17454
rect 16046 17378 16098 17390
rect 16158 17442 16210 17454
rect 21422 17442 21474 17454
rect 17042 17390 17054 17442
rect 17106 17390 17118 17442
rect 16158 17378 16210 17390
rect 21422 17378 21474 17390
rect 35534 17442 35586 17454
rect 35534 17378 35586 17390
rect 35758 17442 35810 17454
rect 35758 17378 35810 17390
rect 36542 17442 36594 17454
rect 36542 17378 36594 17390
rect 37102 17442 37154 17454
rect 51214 17442 51266 17454
rect 50418 17390 50430 17442
rect 50482 17390 50494 17442
rect 37102 17378 37154 17390
rect 51214 17378 51266 17390
rect 1344 17274 58576 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 50558 17274
rect 50610 17222 50662 17274
rect 50714 17222 50766 17274
rect 50818 17222 58576 17274
rect 1344 17188 58576 17222
rect 2046 17106 2098 17118
rect 3054 17106 3106 17118
rect 2370 17054 2382 17106
rect 2434 17054 2446 17106
rect 2046 17042 2098 17054
rect 3054 17042 3106 17054
rect 3838 17106 3890 17118
rect 3838 17042 3890 17054
rect 4510 17106 4562 17118
rect 4510 17042 4562 17054
rect 4734 17106 4786 17118
rect 4734 17042 4786 17054
rect 6302 17106 6354 17118
rect 6302 17042 6354 17054
rect 6750 17106 6802 17118
rect 11790 17106 11842 17118
rect 7634 17054 7646 17106
rect 7698 17054 7710 17106
rect 6750 17042 6802 17054
rect 11790 17042 11842 17054
rect 12462 17106 12514 17118
rect 12462 17042 12514 17054
rect 14366 17106 14418 17118
rect 14366 17042 14418 17054
rect 14590 17106 14642 17118
rect 14590 17042 14642 17054
rect 20974 17106 21026 17118
rect 20974 17042 21026 17054
rect 28142 17106 28194 17118
rect 28142 17042 28194 17054
rect 28366 17106 28418 17118
rect 28366 17042 28418 17054
rect 28702 17106 28754 17118
rect 28702 17042 28754 17054
rect 28926 17106 28978 17118
rect 28926 17042 28978 17054
rect 34974 17106 35026 17118
rect 43598 17106 43650 17118
rect 35298 17054 35310 17106
rect 35362 17054 35374 17106
rect 38322 17054 38334 17106
rect 38386 17054 38398 17106
rect 47842 17054 47854 17106
rect 47906 17054 47918 17106
rect 53330 17054 53342 17106
rect 53394 17054 53406 17106
rect 56914 17054 56926 17106
rect 56978 17054 56990 17106
rect 34974 17042 35026 17054
rect 43598 17042 43650 17054
rect 5294 16994 5346 17006
rect 14142 16994 14194 17006
rect 27470 16994 27522 17006
rect 7746 16942 7758 16994
rect 7810 16942 7822 16994
rect 12114 16942 12126 16994
rect 12178 16942 12190 16994
rect 12786 16942 12798 16994
rect 12850 16942 12862 16994
rect 19506 16942 19518 16994
rect 19570 16942 19582 16994
rect 21746 16942 21758 16994
rect 21810 16942 21822 16994
rect 24322 16942 24334 16994
rect 24386 16942 24398 16994
rect 25554 16942 25566 16994
rect 25618 16942 25630 16994
rect 5294 16930 5346 16942
rect 14142 16930 14194 16942
rect 27470 16930 27522 16942
rect 37550 16994 37602 17006
rect 55022 16994 55074 17006
rect 39554 16942 39566 16994
rect 39618 16942 39630 16994
rect 41570 16942 41582 16994
rect 41634 16942 41646 16994
rect 43026 16942 43038 16994
rect 43090 16942 43102 16994
rect 46610 16942 46622 16994
rect 46674 16942 46686 16994
rect 47954 16942 47966 16994
rect 48018 16942 48030 16994
rect 52098 16942 52110 16994
rect 52162 16942 52174 16994
rect 57362 16942 57374 16994
rect 57426 16942 57438 16994
rect 37550 16930 37602 16942
rect 55022 16930 55074 16942
rect 3726 16882 3778 16894
rect 5854 16882 5906 16894
rect 13022 16882 13074 16894
rect 1810 16830 1822 16882
rect 1874 16830 1886 16882
rect 2594 16830 2606 16882
rect 2658 16830 2670 16882
rect 3266 16830 3278 16882
rect 3330 16830 3342 16882
rect 4274 16830 4286 16882
rect 4338 16830 4350 16882
rect 4946 16830 4958 16882
rect 5010 16830 5022 16882
rect 7522 16830 7534 16882
rect 7586 16830 7598 16882
rect 3726 16818 3778 16830
rect 5854 16818 5906 16830
rect 13022 16818 13074 16830
rect 13358 16882 13410 16894
rect 13358 16818 13410 16830
rect 13582 16882 13634 16894
rect 15374 16882 15426 16894
rect 16270 16882 16322 16894
rect 28030 16882 28082 16894
rect 15026 16830 15038 16882
rect 15090 16830 15102 16882
rect 15474 16830 15486 16882
rect 15538 16830 15550 16882
rect 18162 16830 18174 16882
rect 18226 16830 18238 16882
rect 18834 16830 18846 16882
rect 18898 16830 18910 16882
rect 19170 16830 19182 16882
rect 19234 16830 19246 16882
rect 22082 16830 22094 16882
rect 22146 16830 22158 16882
rect 22978 16830 22990 16882
rect 23042 16830 23054 16882
rect 26114 16830 26126 16882
rect 26178 16830 26190 16882
rect 26786 16830 26798 16882
rect 26850 16830 26862 16882
rect 13582 16818 13634 16830
rect 15374 16818 15426 16830
rect 16270 16818 16322 16830
rect 28030 16818 28082 16830
rect 28590 16882 28642 16894
rect 29486 16882 29538 16894
rect 34526 16882 34578 16894
rect 36206 16882 36258 16894
rect 29250 16830 29262 16882
rect 29314 16830 29326 16882
rect 31378 16830 31390 16882
rect 31442 16830 31454 16882
rect 35746 16830 35758 16882
rect 35810 16830 35822 16882
rect 28590 16818 28642 16830
rect 29486 16818 29538 16830
rect 34526 16818 34578 16830
rect 36206 16818 36258 16830
rect 36766 16882 36818 16894
rect 40462 16882 40514 16894
rect 54574 16882 54626 16894
rect 39778 16830 39790 16882
rect 39842 16830 39854 16882
rect 46834 16830 46846 16882
rect 46898 16830 46910 16882
rect 53218 16830 53230 16882
rect 53282 16830 53294 16882
rect 36766 16818 36818 16830
rect 40462 16818 40514 16830
rect 54574 16818 54626 16830
rect 54910 16882 54962 16894
rect 54910 16818 54962 16830
rect 55246 16882 55298 16894
rect 55246 16818 55298 16830
rect 55470 16882 55522 16894
rect 56018 16830 56030 16882
rect 56082 16830 56094 16882
rect 56690 16830 56702 16882
rect 56754 16830 56766 16882
rect 57810 16830 57822 16882
rect 57874 16830 57886 16882
rect 55470 16818 55522 16830
rect 4622 16770 4674 16782
rect 4622 16706 4674 16718
rect 13246 16770 13298 16782
rect 13246 16706 13298 16718
rect 14478 16770 14530 16782
rect 31838 16770 31890 16782
rect 31490 16718 31502 16770
rect 31554 16718 31566 16770
rect 14478 16706 14530 16718
rect 31838 16706 31890 16718
rect 38894 16770 38946 16782
rect 51662 16770 51714 16782
rect 39890 16718 39902 16770
rect 39954 16718 39966 16770
rect 41682 16718 41694 16770
rect 41746 16718 41758 16770
rect 38894 16706 38946 16718
rect 51662 16706 51714 16718
rect 3838 16658 3890 16670
rect 3838 16594 3890 16606
rect 29710 16658 29762 16670
rect 29710 16594 29762 16606
rect 29822 16658 29874 16670
rect 29822 16594 29874 16606
rect 34638 16658 34690 16670
rect 34638 16594 34690 16606
rect 37326 16658 37378 16670
rect 37326 16594 37378 16606
rect 37662 16658 37714 16670
rect 37662 16594 37714 16606
rect 38670 16658 38722 16670
rect 38670 16594 38722 16606
rect 55694 16658 55746 16670
rect 55694 16594 55746 16606
rect 1344 16490 58576 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 58576 16490
rect 1344 16404 58576 16438
rect 5854 16322 5906 16334
rect 5854 16258 5906 16270
rect 6190 16322 6242 16334
rect 6190 16258 6242 16270
rect 6974 16322 7026 16334
rect 18286 16322 18338 16334
rect 22990 16322 23042 16334
rect 14466 16270 14478 16322
rect 14530 16270 14542 16322
rect 19170 16270 19182 16322
rect 19234 16270 19246 16322
rect 6974 16258 7026 16270
rect 18286 16258 18338 16270
rect 22990 16258 23042 16270
rect 33294 16322 33346 16334
rect 33294 16258 33346 16270
rect 43486 16322 43538 16334
rect 43486 16258 43538 16270
rect 46510 16322 46562 16334
rect 46510 16258 46562 16270
rect 55582 16322 55634 16334
rect 55582 16258 55634 16270
rect 2494 16210 2546 16222
rect 2494 16146 2546 16158
rect 3502 16210 3554 16222
rect 22318 16210 22370 16222
rect 37998 16210 38050 16222
rect 53230 16210 53282 16222
rect 18946 16158 18958 16210
rect 19010 16158 19022 16210
rect 22642 16158 22654 16210
rect 22706 16158 22718 16210
rect 28018 16158 28030 16210
rect 28082 16158 28094 16210
rect 38770 16158 38782 16210
rect 38834 16158 38846 16210
rect 41122 16158 41134 16210
rect 41186 16158 41198 16210
rect 49186 16158 49198 16210
rect 49250 16158 49262 16210
rect 55346 16158 55358 16210
rect 55410 16158 55422 16210
rect 57922 16158 57934 16210
rect 57986 16158 57998 16210
rect 3502 16146 3554 16158
rect 22318 16146 22370 16158
rect 37998 16146 38050 16158
rect 53230 16146 53282 16158
rect 4286 16098 4338 16110
rect 4286 16034 4338 16046
rect 4510 16098 4562 16110
rect 4510 16034 4562 16046
rect 5630 16098 5682 16110
rect 7982 16098 8034 16110
rect 6626 16046 6638 16098
rect 6690 16046 6702 16098
rect 5630 16034 5682 16046
rect 7982 16034 8034 16046
rect 8654 16098 8706 16110
rect 8654 16034 8706 16046
rect 10782 16098 10834 16110
rect 13918 16098 13970 16110
rect 18846 16098 18898 16110
rect 20078 16098 20130 16110
rect 10994 16046 11006 16098
rect 11058 16046 11070 16098
rect 13682 16046 13694 16098
rect 13746 16046 13758 16098
rect 16034 16046 16046 16098
rect 16098 16046 16110 16098
rect 16930 16046 16942 16098
rect 16994 16046 17006 16098
rect 19170 16046 19182 16098
rect 19234 16046 19246 16098
rect 10782 16034 10834 16046
rect 13918 16034 13970 16046
rect 18846 16034 18898 16046
rect 20078 16034 20130 16046
rect 21422 16098 21474 16110
rect 24222 16098 24274 16110
rect 21634 16046 21646 16098
rect 21698 16046 21710 16098
rect 21422 16034 21474 16046
rect 24222 16034 24274 16046
rect 25118 16098 25170 16110
rect 25118 16034 25170 16046
rect 25790 16098 25842 16110
rect 26686 16098 26738 16110
rect 29822 16098 29874 16110
rect 26002 16046 26014 16098
rect 26066 16046 26078 16098
rect 27010 16046 27022 16098
rect 27074 16046 27086 16098
rect 27570 16046 27582 16098
rect 27634 16046 27646 16098
rect 25790 16034 25842 16046
rect 26686 16034 26738 16046
rect 29822 16034 29874 16046
rect 30046 16098 30098 16110
rect 30046 16034 30098 16046
rect 35534 16098 35586 16110
rect 35534 16034 35586 16046
rect 36206 16098 36258 16110
rect 36206 16034 36258 16046
rect 37102 16098 37154 16110
rect 41582 16098 41634 16110
rect 37314 16046 37326 16098
rect 37378 16046 37390 16098
rect 39778 16046 39790 16098
rect 39842 16046 39854 16098
rect 37102 16034 37154 16046
rect 41582 16034 41634 16046
rect 41918 16098 41970 16110
rect 51102 16098 51154 16110
rect 44034 16046 44046 16098
rect 44098 16046 44110 16098
rect 45266 16046 45278 16098
rect 45330 16046 45342 16098
rect 47842 16046 47854 16098
rect 47906 16046 47918 16098
rect 50754 16046 50766 16098
rect 50818 16046 50830 16098
rect 55122 16046 55134 16098
rect 55186 16046 55198 16098
rect 56130 16046 56142 16098
rect 56194 16046 56206 16098
rect 56466 16046 56478 16098
rect 56530 16046 56542 16098
rect 56802 16046 56814 16098
rect 56866 16046 56878 16098
rect 41918 16034 41970 16046
rect 51102 16034 51154 16046
rect 1710 15986 1762 15998
rect 1710 15922 1762 15934
rect 2046 15986 2098 15998
rect 4734 15986 4786 15998
rect 7534 15986 7586 15998
rect 3154 15934 3166 15986
rect 3218 15934 3230 15986
rect 3602 15934 3614 15986
rect 3666 15934 3678 15986
rect 3938 15934 3950 15986
rect 4002 15934 4014 15986
rect 5058 15934 5070 15986
rect 5122 15934 5134 15986
rect 2046 15922 2098 15934
rect 4734 15922 4786 15934
rect 7534 15922 7586 15934
rect 11678 15986 11730 15998
rect 11678 15922 11730 15934
rect 14030 15986 14082 15998
rect 20302 15986 20354 15998
rect 15922 15934 15934 15986
rect 15986 15934 15998 15986
rect 14030 15922 14082 15934
rect 20302 15922 20354 15934
rect 20414 15986 20466 15998
rect 20414 15922 20466 15934
rect 23326 15986 23378 15998
rect 24110 15986 24162 15998
rect 23650 15934 23662 15986
rect 23714 15934 23726 15986
rect 23326 15922 23378 15934
rect 24110 15922 24162 15934
rect 25230 15986 25282 15998
rect 33406 15986 33458 15998
rect 34974 15986 35026 15998
rect 35870 15986 35922 15998
rect 28130 15934 28142 15986
rect 28194 15934 28206 15986
rect 34402 15934 34414 15986
rect 34466 15934 34478 15986
rect 35298 15934 35310 15986
rect 35362 15934 35374 15986
rect 25230 15922 25282 15934
rect 33406 15922 33458 15934
rect 34974 15922 35026 15934
rect 35870 15922 35922 15934
rect 36094 15986 36146 15998
rect 41806 15986 41858 15998
rect 41010 15934 41022 15986
rect 41074 15934 41086 15986
rect 36094 15922 36146 15934
rect 41806 15922 41858 15934
rect 43374 15986 43426 15998
rect 50094 15986 50146 15998
rect 44258 15934 44270 15986
rect 44322 15934 44334 15986
rect 44930 15934 44942 15986
rect 44994 15934 45006 15986
rect 45490 15934 45502 15986
rect 45554 15934 45566 15986
rect 48962 15934 48974 15986
rect 49026 15934 49038 15986
rect 43374 15922 43426 15934
rect 50094 15922 50146 15934
rect 50990 15986 51042 15998
rect 50990 15922 51042 15934
rect 53566 15986 53618 15998
rect 53566 15922 53618 15934
rect 53678 15986 53730 15998
rect 53678 15922 53730 15934
rect 53902 15986 53954 15998
rect 53902 15922 53954 15934
rect 54238 15986 54290 15998
rect 54238 15922 54290 15934
rect 2830 15874 2882 15886
rect 2830 15810 2882 15822
rect 6862 15874 6914 15886
rect 6862 15810 6914 15822
rect 7198 15874 7250 15886
rect 7198 15810 7250 15822
rect 7422 15874 7474 15886
rect 7422 15810 7474 15822
rect 8318 15874 8370 15886
rect 22766 15874 22818 15886
rect 8978 15822 8990 15874
rect 9042 15822 9054 15874
rect 8318 15810 8370 15822
rect 22766 15810 22818 15822
rect 23886 15874 23938 15886
rect 23886 15810 23938 15822
rect 25454 15874 25506 15886
rect 33294 15874 33346 15886
rect 30370 15822 30382 15874
rect 30434 15822 30446 15874
rect 25454 15810 25506 15822
rect 33294 15810 33346 15822
rect 34078 15874 34130 15886
rect 34078 15810 34130 15822
rect 43486 15874 43538 15886
rect 54350 15874 54402 15886
rect 51538 15822 51550 15874
rect 51602 15822 51614 15874
rect 43486 15810 43538 15822
rect 54350 15810 54402 15822
rect 1344 15706 58576 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 50558 15706
rect 50610 15654 50662 15706
rect 50714 15654 50766 15706
rect 50818 15654 58576 15706
rect 1344 15620 58576 15654
rect 4958 15538 5010 15550
rect 4958 15474 5010 15486
rect 13246 15538 13298 15550
rect 13246 15474 13298 15486
rect 13582 15538 13634 15550
rect 31502 15538 31554 15550
rect 14914 15486 14926 15538
rect 14978 15486 14990 15538
rect 20626 15486 20638 15538
rect 20690 15486 20702 15538
rect 13582 15474 13634 15486
rect 31502 15474 31554 15486
rect 34638 15538 34690 15550
rect 39902 15538 39954 15550
rect 35634 15486 35646 15538
rect 35698 15486 35710 15538
rect 34638 15474 34690 15486
rect 39902 15474 39954 15486
rect 49982 15538 50034 15550
rect 49982 15474 50034 15486
rect 50542 15538 50594 15550
rect 50542 15474 50594 15486
rect 56478 15538 56530 15550
rect 56478 15474 56530 15486
rect 56590 15538 56642 15550
rect 56590 15474 56642 15486
rect 11678 15426 11730 15438
rect 6514 15374 6526 15426
rect 6578 15374 6590 15426
rect 10994 15374 11006 15426
rect 11058 15374 11070 15426
rect 11678 15362 11730 15374
rect 11790 15426 11842 15438
rect 11790 15362 11842 15374
rect 13358 15426 13410 15438
rect 27918 15426 27970 15438
rect 16482 15374 16494 15426
rect 16546 15374 16558 15426
rect 19394 15374 19406 15426
rect 19458 15374 19470 15426
rect 22418 15374 22430 15426
rect 22482 15374 22494 15426
rect 26002 15374 26014 15426
rect 26066 15374 26078 15426
rect 13358 15362 13410 15374
rect 27918 15362 27970 15374
rect 31054 15426 31106 15438
rect 31054 15362 31106 15374
rect 34862 15426 34914 15438
rect 49870 15426 49922 15438
rect 37762 15374 37774 15426
rect 37826 15374 37838 15426
rect 45938 15374 45950 15426
rect 46002 15374 46014 15426
rect 34862 15362 34914 15374
rect 49870 15362 49922 15374
rect 50430 15426 50482 15438
rect 55918 15426 55970 15438
rect 54002 15374 54014 15426
rect 54066 15374 54078 15426
rect 50430 15362 50482 15374
rect 55918 15362 55970 15374
rect 11454 15314 11506 15326
rect 4274 15262 4286 15314
rect 4338 15262 4350 15314
rect 7746 15262 7758 15314
rect 7810 15262 7822 15314
rect 10210 15262 10222 15314
rect 10274 15262 10286 15314
rect 10546 15262 10558 15314
rect 10610 15262 10622 15314
rect 11454 15250 11506 15262
rect 13918 15314 13970 15326
rect 29598 15314 29650 15326
rect 15138 15262 15150 15314
rect 15202 15262 15214 15314
rect 16034 15262 16046 15314
rect 16098 15262 16110 15314
rect 20290 15262 20302 15314
rect 20354 15262 20366 15314
rect 22530 15262 22542 15314
rect 22594 15262 22606 15314
rect 23426 15262 23438 15314
rect 23490 15262 23502 15314
rect 26338 15262 26350 15314
rect 26402 15262 26414 15314
rect 27234 15262 27246 15314
rect 27298 15262 27310 15314
rect 29250 15262 29262 15314
rect 29314 15262 29326 15314
rect 13918 15250 13970 15262
rect 29598 15250 29650 15262
rect 29710 15314 29762 15326
rect 30942 15314 30994 15326
rect 30370 15262 30382 15314
rect 30434 15262 30446 15314
rect 29710 15250 29762 15262
rect 30942 15250 30994 15262
rect 31278 15314 31330 15326
rect 31278 15250 31330 15262
rect 31614 15314 31666 15326
rect 31614 15250 31666 15262
rect 31838 15314 31890 15326
rect 34974 15314 35026 15326
rect 33730 15262 33742 15314
rect 33794 15262 33806 15314
rect 31838 15250 31890 15262
rect 34974 15250 35026 15262
rect 35982 15314 36034 15326
rect 37326 15314 37378 15326
rect 48750 15314 48802 15326
rect 50206 15314 50258 15326
rect 36866 15262 36878 15314
rect 36930 15262 36942 15314
rect 37650 15262 37662 15314
rect 37714 15262 37726 15314
rect 39442 15262 39454 15314
rect 39506 15262 39518 15314
rect 41458 15262 41470 15314
rect 41522 15262 41534 15314
rect 42914 15262 42926 15314
rect 42978 15262 42990 15314
rect 43922 15262 43934 15314
rect 43986 15262 43998 15314
rect 45714 15262 45726 15314
rect 45778 15262 45790 15314
rect 47506 15262 47518 15314
rect 47570 15262 47582 15314
rect 49074 15262 49086 15314
rect 49138 15262 49150 15314
rect 35982 15250 36034 15262
rect 37326 15250 37378 15262
rect 48750 15250 48802 15262
rect 50206 15250 50258 15262
rect 50766 15314 50818 15326
rect 50978 15262 50990 15314
rect 51042 15262 51054 15314
rect 52210 15262 52222 15314
rect 52274 15262 52286 15314
rect 52770 15262 52782 15314
rect 52834 15262 52846 15314
rect 55234 15262 55246 15314
rect 55298 15262 55310 15314
rect 56802 15262 56814 15314
rect 56866 15262 56878 15314
rect 57026 15262 57038 15314
rect 57090 15262 57102 15314
rect 50766 15250 50818 15262
rect 5518 15202 5570 15214
rect 34414 15202 34466 15214
rect 6066 15150 6078 15202
rect 6130 15150 6142 15202
rect 8754 15150 8766 15202
rect 8818 15150 8830 15202
rect 10994 15150 11006 15202
rect 11058 15150 11070 15202
rect 18834 15150 18846 15202
rect 18898 15150 18910 15202
rect 24658 15150 24670 15202
rect 24722 15150 24734 15202
rect 34066 15150 34078 15202
rect 34130 15150 34142 15202
rect 36530 15150 36542 15202
rect 36594 15150 36606 15202
rect 41122 15150 41134 15202
rect 41186 15150 41198 15202
rect 43586 15150 43598 15202
rect 43650 15150 43662 15202
rect 44370 15150 44382 15202
rect 44434 15150 44446 15202
rect 47282 15150 47294 15202
rect 47346 15150 47358 15202
rect 51650 15150 51662 15202
rect 51714 15150 51726 15202
rect 53778 15150 53790 15202
rect 53842 15150 53854 15202
rect 5518 15138 5570 15150
rect 34414 15138 34466 15150
rect 1934 15090 1986 15102
rect 49410 15038 49422 15090
rect 49474 15038 49486 15090
rect 1934 15026 1986 15038
rect 1344 14922 58576 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 58576 14922
rect 1344 14836 58576 14870
rect 6638 14754 6690 14766
rect 6638 14690 6690 14702
rect 6862 14754 6914 14766
rect 21310 14754 21362 14766
rect 17938 14702 17950 14754
rect 18002 14702 18014 14754
rect 6862 14690 6914 14702
rect 21310 14690 21362 14702
rect 29822 14754 29874 14766
rect 29822 14690 29874 14702
rect 33070 14754 33122 14766
rect 33070 14690 33122 14702
rect 39790 14754 39842 14766
rect 39790 14690 39842 14702
rect 43822 14754 43874 14766
rect 55134 14754 55186 14766
rect 48514 14702 48526 14754
rect 48578 14702 48590 14754
rect 52770 14702 52782 14754
rect 52834 14702 52846 14754
rect 43822 14690 43874 14702
rect 55134 14690 55186 14702
rect 2270 14642 2322 14654
rect 2270 14578 2322 14590
rect 3390 14642 3442 14654
rect 3390 14578 3442 14590
rect 3838 14642 3890 14654
rect 3838 14578 3890 14590
rect 4622 14642 4674 14654
rect 4622 14578 4674 14590
rect 4958 14642 5010 14654
rect 4958 14578 5010 14590
rect 6414 14642 6466 14654
rect 12910 14642 12962 14654
rect 20078 14642 20130 14654
rect 9538 14590 9550 14642
rect 9602 14590 9614 14642
rect 10770 14590 10782 14642
rect 10834 14590 10846 14642
rect 15586 14590 15598 14642
rect 15650 14590 15662 14642
rect 16258 14590 16270 14642
rect 16322 14590 16334 14642
rect 17826 14590 17838 14642
rect 17890 14590 17902 14642
rect 19282 14590 19294 14642
rect 19346 14590 19358 14642
rect 6414 14578 6466 14590
rect 12910 14578 12962 14590
rect 20078 14578 20130 14590
rect 22654 14642 22706 14654
rect 36990 14642 37042 14654
rect 55470 14642 55522 14654
rect 23538 14590 23550 14642
rect 23602 14590 23614 14642
rect 26898 14590 26910 14642
rect 26962 14590 26974 14642
rect 30818 14590 30830 14642
rect 30882 14590 30894 14642
rect 42466 14590 42478 14642
rect 42530 14590 42542 14642
rect 47394 14590 47406 14642
rect 47458 14590 47470 14642
rect 50754 14590 50766 14642
rect 50818 14590 50830 14642
rect 52882 14590 52894 14642
rect 52946 14590 52958 14642
rect 22654 14578 22706 14590
rect 36990 14578 37042 14590
rect 55470 14578 55522 14590
rect 2606 14530 2658 14542
rect 1810 14478 1822 14530
rect 1874 14478 1886 14530
rect 2606 14466 2658 14478
rect 8094 14530 8146 14542
rect 8094 14466 8146 14478
rect 8430 14530 8482 14542
rect 8430 14466 8482 14478
rect 8766 14530 8818 14542
rect 28366 14530 28418 14542
rect 8978 14478 8990 14530
rect 9042 14478 9054 14530
rect 9986 14478 9998 14530
rect 10050 14478 10062 14530
rect 15250 14478 15262 14530
rect 15314 14478 15326 14530
rect 16370 14478 16382 14530
rect 16434 14478 16446 14530
rect 16594 14478 16606 14530
rect 16658 14478 16670 14530
rect 17714 14478 17726 14530
rect 17778 14478 17790 14530
rect 19506 14478 19518 14530
rect 19570 14478 19582 14530
rect 21634 14478 21646 14530
rect 21698 14478 21710 14530
rect 23090 14478 23102 14530
rect 23154 14478 23166 14530
rect 23426 14478 23438 14530
rect 23490 14478 23502 14530
rect 24994 14478 25006 14530
rect 25058 14478 25070 14530
rect 25890 14478 25902 14530
rect 25954 14478 25966 14530
rect 26338 14478 26350 14530
rect 26402 14478 26414 14530
rect 8766 14466 8818 14478
rect 28366 14466 28418 14478
rect 28702 14530 28754 14542
rect 30046 14530 30098 14542
rect 32398 14530 32450 14542
rect 34526 14530 34578 14542
rect 29698 14478 29710 14530
rect 29762 14478 29774 14530
rect 30258 14478 30270 14530
rect 30322 14478 30334 14530
rect 31266 14478 31278 14530
rect 31330 14478 31342 14530
rect 33618 14478 33630 14530
rect 33682 14478 33694 14530
rect 28702 14466 28754 14478
rect 30046 14466 30098 14478
rect 32398 14466 32450 14478
rect 34526 14466 34578 14478
rect 34750 14530 34802 14542
rect 43710 14530 43762 14542
rect 38322 14478 38334 14530
rect 38386 14478 38398 14530
rect 41122 14478 41134 14530
rect 41186 14478 41198 14530
rect 43362 14478 43374 14530
rect 43426 14478 43438 14530
rect 34750 14466 34802 14478
rect 43710 14466 43762 14478
rect 44046 14530 44098 14542
rect 46174 14530 46226 14542
rect 54238 14530 54290 14542
rect 44258 14478 44270 14530
rect 44322 14478 44334 14530
rect 44930 14478 44942 14530
rect 44994 14478 45006 14530
rect 45378 14478 45390 14530
rect 45442 14478 45454 14530
rect 45714 14478 45726 14530
rect 45778 14478 45790 14530
rect 47506 14478 47518 14530
rect 47570 14478 47582 14530
rect 49298 14478 49310 14530
rect 49362 14478 49374 14530
rect 50418 14478 50430 14530
rect 50482 14478 50494 14530
rect 52994 14478 53006 14530
rect 53058 14478 53070 14530
rect 53218 14478 53230 14530
rect 53282 14478 53294 14530
rect 44046 14466 44098 14478
rect 46174 14466 46226 14478
rect 54238 14466 54290 14478
rect 54462 14530 54514 14542
rect 54462 14466 54514 14478
rect 54686 14530 54738 14542
rect 54686 14466 54738 14478
rect 55246 14530 55298 14542
rect 55246 14466 55298 14478
rect 55806 14530 55858 14542
rect 55806 14466 55858 14478
rect 56142 14530 56194 14542
rect 56142 14466 56194 14478
rect 2942 14418 2994 14430
rect 2942 14354 2994 14366
rect 8654 14418 8706 14430
rect 35422 14418 35474 14430
rect 10322 14366 10334 14418
rect 10386 14366 10398 14418
rect 11218 14366 11230 14418
rect 11282 14366 11294 14418
rect 12562 14366 12574 14418
rect 12626 14366 12638 14418
rect 30370 14366 30382 14418
rect 30434 14366 30446 14418
rect 33506 14366 33518 14418
rect 33570 14366 33582 14418
rect 8654 14354 8706 14366
rect 35422 14354 35474 14366
rect 36206 14418 36258 14430
rect 43038 14418 43090 14430
rect 37202 14366 37214 14418
rect 37266 14366 37278 14418
rect 38658 14366 38670 14418
rect 38722 14366 38734 14418
rect 42018 14366 42030 14418
rect 42082 14366 42094 14418
rect 36206 14354 36258 14366
rect 43038 14354 43090 14366
rect 55694 14418 55746 14430
rect 55694 14354 55746 14366
rect 56478 14418 56530 14430
rect 56478 14354 56530 14366
rect 7310 14306 7362 14318
rect 7310 14242 7362 14254
rect 8206 14306 8258 14318
rect 8206 14242 8258 14254
rect 21422 14306 21474 14318
rect 21422 14242 21474 14254
rect 28478 14306 28530 14318
rect 28478 14242 28530 14254
rect 29486 14306 29538 14318
rect 29486 14242 29538 14254
rect 32734 14306 32786 14318
rect 32734 14242 32786 14254
rect 32958 14306 33010 14318
rect 35534 14306 35586 14318
rect 33842 14254 33854 14306
rect 33906 14254 33918 14306
rect 35074 14254 35086 14306
rect 35138 14254 35150 14306
rect 32958 14242 33010 14254
rect 35534 14242 35586 14254
rect 35646 14306 35698 14318
rect 35646 14242 35698 14254
rect 36318 14306 36370 14318
rect 36318 14242 36370 14254
rect 36542 14306 36594 14318
rect 36542 14242 36594 14254
rect 43150 14306 43202 14318
rect 43150 14242 43202 14254
rect 56366 14306 56418 14318
rect 56366 14242 56418 14254
rect 1344 14138 58576 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 50558 14138
rect 50610 14086 50662 14138
rect 50714 14086 50766 14138
rect 50818 14086 58576 14138
rect 1344 14052 58576 14086
rect 2046 13970 2098 13982
rect 2046 13906 2098 13918
rect 2718 13970 2770 13982
rect 2718 13906 2770 13918
rect 3166 13970 3218 13982
rect 3166 13906 3218 13918
rect 3614 13970 3666 13982
rect 3614 13906 3666 13918
rect 5966 13970 6018 13982
rect 5966 13906 6018 13918
rect 6190 13970 6242 13982
rect 6190 13906 6242 13918
rect 8766 13970 8818 13982
rect 8766 13906 8818 13918
rect 10558 13970 10610 13982
rect 10558 13906 10610 13918
rect 17614 13970 17666 13982
rect 17614 13906 17666 13918
rect 24558 13970 24610 13982
rect 24558 13906 24610 13918
rect 26350 13970 26402 13982
rect 26350 13906 26402 13918
rect 28478 13970 28530 13982
rect 32510 13970 32562 13982
rect 31266 13918 31278 13970
rect 31330 13918 31342 13970
rect 28478 13906 28530 13918
rect 32510 13906 32562 13918
rect 48302 13970 48354 13982
rect 48302 13906 48354 13918
rect 53454 13970 53506 13982
rect 53454 13906 53506 13918
rect 54462 13970 54514 13982
rect 54462 13906 54514 13918
rect 55582 13970 55634 13982
rect 55582 13906 55634 13918
rect 1710 13858 1762 13870
rect 1710 13794 1762 13806
rect 8318 13858 8370 13870
rect 15262 13858 15314 13870
rect 11330 13806 11342 13858
rect 11394 13806 11406 13858
rect 13906 13806 13918 13858
rect 13970 13806 13982 13858
rect 8318 13794 8370 13806
rect 15262 13794 15314 13806
rect 15486 13858 15538 13870
rect 23886 13858 23938 13870
rect 23650 13806 23662 13858
rect 23714 13806 23726 13858
rect 15486 13794 15538 13806
rect 23886 13794 23938 13806
rect 26574 13858 26626 13870
rect 26574 13794 26626 13806
rect 28254 13858 28306 13870
rect 48750 13858 48802 13870
rect 55358 13858 55410 13870
rect 30258 13806 30270 13858
rect 30322 13806 30334 13858
rect 43586 13806 43598 13858
rect 43650 13806 43662 13858
rect 45826 13806 45838 13858
rect 45890 13806 45902 13858
rect 50754 13806 50766 13858
rect 50818 13806 50830 13858
rect 52658 13806 52670 13858
rect 52722 13806 52734 13858
rect 28254 13794 28306 13806
rect 48750 13794 48802 13806
rect 55358 13794 55410 13806
rect 2382 13746 2434 13758
rect 8542 13746 8594 13758
rect 6514 13694 6526 13746
rect 6578 13694 6590 13746
rect 2382 13682 2434 13694
rect 8542 13682 8594 13694
rect 8878 13746 8930 13758
rect 8878 13682 8930 13694
rect 9774 13746 9826 13758
rect 9774 13682 9826 13694
rect 9886 13746 9938 13758
rect 22430 13746 22482 13758
rect 10098 13694 10110 13746
rect 10162 13694 10174 13746
rect 11666 13694 11678 13746
rect 11730 13694 11742 13746
rect 12562 13694 12574 13746
rect 12626 13694 12638 13746
rect 9886 13682 9938 13694
rect 22430 13682 22482 13694
rect 22654 13746 22706 13758
rect 22654 13682 22706 13694
rect 23326 13746 23378 13758
rect 26238 13746 26290 13758
rect 27694 13746 27746 13758
rect 24098 13694 24110 13746
rect 24162 13694 24174 13746
rect 27234 13694 27246 13746
rect 27298 13694 27310 13746
rect 23326 13682 23378 13694
rect 26238 13682 26290 13694
rect 27694 13682 27746 13694
rect 27806 13746 27858 13758
rect 27806 13682 27858 13694
rect 28142 13746 28194 13758
rect 32398 13746 32450 13758
rect 30706 13694 30718 13746
rect 30770 13694 30782 13746
rect 31154 13694 31166 13746
rect 31218 13694 31230 13746
rect 28142 13682 28194 13694
rect 32398 13682 32450 13694
rect 33854 13746 33906 13758
rect 37550 13746 37602 13758
rect 39566 13746 39618 13758
rect 48974 13746 49026 13758
rect 34962 13694 34974 13746
rect 35026 13694 35038 13746
rect 35634 13694 35646 13746
rect 35698 13694 35710 13746
rect 36642 13694 36654 13746
rect 36706 13694 36718 13746
rect 37762 13694 37774 13746
rect 37826 13694 37838 13746
rect 41234 13694 41246 13746
rect 41298 13694 41310 13746
rect 41570 13694 41582 13746
rect 41634 13694 41646 13746
rect 44706 13694 44718 13746
rect 44770 13694 44782 13746
rect 47282 13694 47294 13746
rect 47346 13694 47358 13746
rect 47618 13694 47630 13746
rect 47682 13694 47694 13746
rect 33854 13682 33906 13694
rect 37550 13682 37602 13694
rect 39566 13682 39618 13694
rect 48974 13682 49026 13694
rect 49086 13746 49138 13758
rect 54350 13746 54402 13758
rect 51986 13694 51998 13746
rect 52050 13694 52062 13746
rect 53666 13694 53678 13746
rect 53730 13694 53742 13746
rect 49086 13682 49138 13694
rect 54350 13682 54402 13694
rect 54574 13746 54626 13758
rect 54574 13682 54626 13694
rect 55022 13746 55074 13758
rect 55022 13682 55074 13694
rect 55246 13746 55298 13758
rect 55246 13682 55298 13694
rect 4062 13634 4114 13646
rect 4062 13570 4114 13582
rect 6078 13634 6130 13646
rect 9550 13634 9602 13646
rect 22878 13634 22930 13646
rect 8754 13582 8766 13634
rect 8818 13582 8830 13634
rect 18050 13582 18062 13634
rect 18114 13582 18126 13634
rect 6078 13570 6130 13582
rect 9550 13570 9602 13582
rect 22878 13570 22930 13582
rect 23550 13634 23602 13646
rect 36866 13582 36878 13634
rect 36930 13582 36942 13634
rect 40114 13582 40126 13634
rect 40178 13582 40190 13634
rect 41458 13582 41470 13634
rect 41522 13582 41534 13634
rect 43138 13582 43150 13634
rect 43202 13582 43214 13634
rect 47954 13582 47966 13634
rect 48018 13582 48030 13634
rect 50194 13582 50206 13634
rect 50258 13582 50270 13634
rect 23550 13570 23602 13582
rect 15598 13522 15650 13534
rect 15598 13458 15650 13470
rect 39790 13522 39842 13534
rect 53342 13522 53394 13534
rect 41906 13470 41918 13522
rect 41970 13470 41982 13522
rect 39790 13458 39842 13470
rect 53342 13458 53394 13470
rect 1344 13354 58576 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 58576 13354
rect 1344 13268 58576 13302
rect 42366 13186 42418 13198
rect 53678 13186 53730 13198
rect 43474 13134 43486 13186
rect 43538 13134 43550 13186
rect 42366 13122 42418 13134
rect 53678 13122 53730 13134
rect 3166 13074 3218 13086
rect 3166 13010 3218 13022
rect 6302 13074 6354 13086
rect 28590 13074 28642 13086
rect 31390 13074 31442 13086
rect 39342 13074 39394 13086
rect 42478 13074 42530 13086
rect 55470 13074 55522 13086
rect 15026 13022 15038 13074
rect 15090 13022 15102 13074
rect 15922 13022 15934 13074
rect 15986 13022 15998 13074
rect 29250 13022 29262 13074
rect 29314 13022 29326 13074
rect 33170 13022 33182 13074
rect 33234 13022 33246 13074
rect 41122 13022 41134 13074
rect 41186 13022 41198 13074
rect 45714 13022 45726 13074
rect 45778 13022 45790 13074
rect 48962 13022 48974 13074
rect 49026 13022 49038 13074
rect 51650 13022 51662 13074
rect 51714 13022 51726 13074
rect 6302 13010 6354 13022
rect 28590 13010 28642 13022
rect 31390 13010 31442 13022
rect 39342 13010 39394 13022
rect 42478 13010 42530 13022
rect 55470 13010 55522 13022
rect 5742 12962 5794 12974
rect 2482 12910 2494 12962
rect 2546 12910 2558 12962
rect 5742 12898 5794 12910
rect 6750 12962 6802 12974
rect 6750 12898 6802 12910
rect 8990 12962 9042 12974
rect 8990 12898 9042 12910
rect 13694 12962 13746 12974
rect 18958 12962 19010 12974
rect 14578 12910 14590 12962
rect 14642 12910 14654 12962
rect 15250 12910 15262 12962
rect 15314 12910 15326 12962
rect 17378 12910 17390 12962
rect 17442 12910 17454 12962
rect 13694 12898 13746 12910
rect 18958 12898 19010 12910
rect 20414 12962 20466 12974
rect 38222 12962 38274 12974
rect 44158 12962 44210 12974
rect 47518 12962 47570 12974
rect 54574 12962 54626 12974
rect 21746 12910 21758 12962
rect 21810 12910 21822 12962
rect 23314 12910 23326 12962
rect 23378 12910 23390 12962
rect 23986 12910 23998 12962
rect 24050 12910 24062 12962
rect 27234 12910 27246 12962
rect 27298 12910 27310 12962
rect 27906 12910 27918 12962
rect 27970 12910 27982 12962
rect 34178 12910 34190 12962
rect 34242 12910 34254 12962
rect 35074 12910 35086 12962
rect 35138 12910 35150 12962
rect 40114 12910 40126 12962
rect 40178 12910 40190 12962
rect 41682 12910 41694 12962
rect 41746 12910 41758 12962
rect 45042 12910 45054 12962
rect 45106 12910 45118 12962
rect 46610 12910 46622 12962
rect 46674 12910 46686 12962
rect 48402 12910 48414 12962
rect 48466 12910 48478 12962
rect 48738 12910 48750 12962
rect 48802 12910 48814 12962
rect 50978 12910 50990 12962
rect 51042 12910 51054 12962
rect 52098 12910 52110 12962
rect 52162 12910 52174 12962
rect 54786 12910 54798 12962
rect 54850 12910 54862 12962
rect 20414 12898 20466 12910
rect 38222 12898 38274 12910
rect 44158 12898 44210 12910
rect 47518 12898 47570 12910
rect 54574 12898 54626 12910
rect 1710 12850 1762 12862
rect 1710 12786 1762 12798
rect 2046 12850 2098 12862
rect 2046 12786 2098 12798
rect 2718 12850 2770 12862
rect 2718 12786 2770 12798
rect 3614 12850 3666 12862
rect 3614 12786 3666 12798
rect 9326 12850 9378 12862
rect 12574 12850 12626 12862
rect 18062 12850 18114 12862
rect 9986 12798 9998 12850
rect 10050 12798 10062 12850
rect 14354 12798 14366 12850
rect 14418 12798 14430 12850
rect 16482 12798 16494 12850
rect 16546 12798 16558 12850
rect 9326 12786 9378 12798
rect 12574 12786 12626 12798
rect 18062 12786 18114 12798
rect 18734 12850 18786 12862
rect 18734 12786 18786 12798
rect 19294 12850 19346 12862
rect 19294 12786 19346 12798
rect 19966 12850 20018 12862
rect 19966 12786 20018 12798
rect 20078 12850 20130 12862
rect 24670 12850 24722 12862
rect 20738 12798 20750 12850
rect 20802 12798 20814 12850
rect 21634 12798 21646 12850
rect 21698 12798 21710 12850
rect 22082 12798 22094 12850
rect 22146 12798 22158 12850
rect 23090 12798 23102 12850
rect 23154 12798 23166 12850
rect 20078 12786 20130 12798
rect 24670 12786 24722 12798
rect 25790 12850 25842 12862
rect 25790 12786 25842 12798
rect 25902 12850 25954 12862
rect 25902 12786 25954 12798
rect 26126 12850 26178 12862
rect 38334 12850 38386 12862
rect 26674 12798 26686 12850
rect 26738 12798 26750 12850
rect 29474 12798 29486 12850
rect 29538 12798 29550 12850
rect 31154 12798 31166 12850
rect 31218 12798 31230 12850
rect 35298 12798 35310 12850
rect 35362 12798 35374 12850
rect 26126 12786 26178 12798
rect 38334 12786 38386 12798
rect 38558 12850 38610 12862
rect 43934 12850 43986 12862
rect 39666 12798 39678 12850
rect 39730 12798 39742 12850
rect 38558 12786 38610 12798
rect 43934 12786 43986 12798
rect 44046 12850 44098 12862
rect 53342 12850 53394 12862
rect 44818 12798 44830 12850
rect 44882 12798 44894 12850
rect 49410 12798 49422 12850
rect 49474 12798 49486 12850
rect 51090 12798 51102 12850
rect 51154 12798 51166 12850
rect 52994 12798 53006 12850
rect 53058 12798 53070 12850
rect 44046 12786 44098 12798
rect 53342 12786 53394 12798
rect 7086 12738 7138 12750
rect 7086 12674 7138 12686
rect 9662 12738 9714 12750
rect 19182 12738 19234 12750
rect 12898 12686 12910 12738
rect 12962 12686 12974 12738
rect 14018 12686 14030 12738
rect 14082 12686 14094 12738
rect 9662 12674 9714 12686
rect 19182 12674 19234 12686
rect 19742 12738 19794 12750
rect 19742 12674 19794 12686
rect 37102 12738 37154 12750
rect 37102 12674 37154 12686
rect 38782 12738 38834 12750
rect 38782 12674 38834 12686
rect 42590 12738 42642 12750
rect 42590 12674 42642 12686
rect 47630 12738 47682 12750
rect 47630 12674 47682 12686
rect 47854 12738 47906 12750
rect 47854 12674 47906 12686
rect 52670 12738 52722 12750
rect 52670 12674 52722 12686
rect 53566 12738 53618 12750
rect 53566 12674 53618 12686
rect 1344 12570 58576 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 50558 12570
rect 50610 12518 50662 12570
rect 50714 12518 50766 12570
rect 50818 12518 58576 12570
rect 1344 12484 58576 12518
rect 2046 12402 2098 12414
rect 2046 12338 2098 12350
rect 4958 12402 5010 12414
rect 37662 12402 37714 12414
rect 43374 12402 43426 12414
rect 51886 12402 51938 12414
rect 20626 12350 20638 12402
rect 20690 12350 20702 12402
rect 40114 12350 40126 12402
rect 40178 12350 40190 12402
rect 41794 12350 41806 12402
rect 41858 12350 41870 12402
rect 42690 12350 42702 12402
rect 42754 12350 42766 12402
rect 43698 12350 43710 12402
rect 43762 12350 43774 12402
rect 45042 12350 45054 12402
rect 45106 12350 45118 12402
rect 50754 12350 50766 12402
rect 50818 12350 50830 12402
rect 4958 12338 5010 12350
rect 37662 12338 37714 12350
rect 43374 12338 43426 12350
rect 51886 12338 51938 12350
rect 6414 12290 6466 12302
rect 18174 12290 18226 12302
rect 31054 12290 31106 12302
rect 38334 12290 38386 12302
rect 51662 12290 51714 12302
rect 8418 12238 8430 12290
rect 8482 12238 8494 12290
rect 16482 12238 16494 12290
rect 16546 12238 16558 12290
rect 18946 12238 18958 12290
rect 19010 12238 19022 12290
rect 23314 12238 23326 12290
rect 23378 12238 23390 12290
rect 36194 12238 36206 12290
rect 36258 12238 36270 12290
rect 36754 12238 36766 12290
rect 36818 12238 36830 12290
rect 38882 12238 38894 12290
rect 38946 12238 38958 12290
rect 39330 12238 39342 12290
rect 39394 12238 39406 12290
rect 39778 12238 39790 12290
rect 39842 12238 39854 12290
rect 44370 12238 44382 12290
rect 44434 12238 44446 12290
rect 44594 12238 44606 12290
rect 44658 12238 44670 12290
rect 48178 12238 48190 12290
rect 48242 12238 48254 12290
rect 6414 12226 6466 12238
rect 18174 12226 18226 12238
rect 31054 12226 31106 12238
rect 38334 12226 38386 12238
rect 51662 12226 51714 12238
rect 52110 12290 52162 12302
rect 52110 12226 52162 12238
rect 54798 12290 54850 12302
rect 54798 12226 54850 12238
rect 54910 12290 54962 12302
rect 54910 12226 54962 12238
rect 1710 12178 1762 12190
rect 1710 12114 1762 12126
rect 2494 12178 2546 12190
rect 2494 12114 2546 12126
rect 4846 12178 4898 12190
rect 4846 12114 4898 12126
rect 5182 12178 5234 12190
rect 6974 12178 7026 12190
rect 23774 12178 23826 12190
rect 37102 12178 37154 12190
rect 5954 12126 5966 12178
rect 6018 12126 6030 12178
rect 6178 12126 6190 12178
rect 6242 12126 6254 12178
rect 8754 12126 8766 12178
rect 8818 12126 8830 12178
rect 9762 12126 9774 12178
rect 9826 12126 9838 12178
rect 11330 12126 11342 12178
rect 11394 12126 11406 12178
rect 12338 12126 12350 12178
rect 12402 12126 12414 12178
rect 12786 12126 12798 12178
rect 12850 12126 12862 12178
rect 15250 12126 15262 12178
rect 15314 12126 15326 12178
rect 15922 12126 15934 12178
rect 15986 12126 15998 12178
rect 19170 12126 19182 12178
rect 19234 12126 19246 12178
rect 20178 12126 20190 12178
rect 20242 12126 20254 12178
rect 22082 12126 22094 12178
rect 22146 12126 22158 12178
rect 22530 12126 22542 12178
rect 22594 12126 22606 12178
rect 22978 12126 22990 12178
rect 23042 12126 23054 12178
rect 24322 12126 24334 12178
rect 24386 12126 24398 12178
rect 25442 12126 25454 12178
rect 25506 12126 25518 12178
rect 27010 12126 27022 12178
rect 27074 12126 27086 12178
rect 28018 12126 28030 12178
rect 28082 12126 28094 12178
rect 28578 12126 28590 12178
rect 28642 12126 28654 12178
rect 30370 12126 30382 12178
rect 30434 12126 30446 12178
rect 36418 12126 36430 12178
rect 36482 12126 36494 12178
rect 5182 12114 5234 12126
rect 6974 12114 7026 12126
rect 23774 12114 23826 12126
rect 37102 12114 37154 12126
rect 37550 12178 37602 12190
rect 37550 12114 37602 12126
rect 37886 12178 37938 12190
rect 38446 12178 38498 12190
rect 38098 12126 38110 12178
rect 38162 12126 38174 12178
rect 37886 12114 37938 12126
rect 38446 12114 38498 12126
rect 40238 12178 40290 12190
rect 40238 12114 40290 12126
rect 41358 12178 41410 12190
rect 47406 12178 47458 12190
rect 50206 12178 50258 12190
rect 41458 12126 41470 12178
rect 41522 12126 41534 12178
rect 42914 12126 42926 12178
rect 42978 12126 42990 12178
rect 44034 12126 44046 12178
rect 44098 12126 44110 12178
rect 47058 12126 47070 12178
rect 47122 12126 47134 12178
rect 47954 12126 47966 12178
rect 48018 12126 48030 12178
rect 49634 12126 49646 12178
rect 49698 12126 49710 12178
rect 41358 12114 41410 12126
rect 47406 12114 47458 12126
rect 50206 12114 50258 12126
rect 51550 12178 51602 12190
rect 52882 12126 52894 12178
rect 52946 12126 52958 12178
rect 53890 12126 53902 12178
rect 53954 12126 53966 12178
rect 51550 12114 51602 12126
rect 2942 12066 2994 12078
rect 2942 12002 2994 12014
rect 6750 12066 6802 12078
rect 14590 12066 14642 12078
rect 8978 12014 8990 12066
rect 9042 12014 9054 12066
rect 10210 12014 10222 12066
rect 10274 12014 10286 12066
rect 6750 12002 6802 12014
rect 14590 12002 14642 12014
rect 23998 12066 24050 12078
rect 47518 12066 47570 12078
rect 50430 12066 50482 12078
rect 25890 12014 25902 12066
rect 25954 12014 25966 12066
rect 27234 12014 27246 12066
rect 27298 12014 27310 12066
rect 30594 12014 30606 12066
rect 30658 12014 30670 12066
rect 36306 12014 36318 12066
rect 36370 12014 36382 12066
rect 41906 12014 41918 12066
rect 41970 12014 41982 12066
rect 49522 12014 49534 12066
rect 49586 12014 49598 12066
rect 53778 12014 53790 12066
rect 53842 12014 53854 12066
rect 23998 12002 24050 12014
rect 47518 12002 47570 12014
rect 50430 12002 50482 12014
rect 7310 11954 7362 11966
rect 17726 11954 17778 11966
rect 13010 11902 13022 11954
rect 13074 11902 13086 11954
rect 7310 11890 7362 11902
rect 17726 11890 17778 11902
rect 17838 11954 17890 11966
rect 17838 11890 17890 11902
rect 18062 11954 18114 11966
rect 54910 11954 54962 11966
rect 49074 11902 49086 11954
rect 49138 11902 49150 11954
rect 18062 11890 18114 11902
rect 54910 11890 54962 11902
rect 1344 11786 58576 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 58576 11786
rect 1344 11700 58576 11734
rect 6526 11618 6578 11630
rect 6526 11554 6578 11566
rect 11454 11618 11506 11630
rect 39902 11618 39954 11630
rect 48638 11618 48690 11630
rect 25554 11566 25566 11618
rect 25618 11566 25630 11618
rect 48066 11566 48078 11618
rect 48130 11566 48142 11618
rect 11454 11554 11506 11566
rect 39902 11554 39954 11566
rect 48638 11554 48690 11566
rect 15374 11506 15426 11518
rect 19294 11506 19346 11518
rect 34862 11506 34914 11518
rect 6850 11454 6862 11506
rect 6914 11454 6926 11506
rect 8642 11454 8654 11506
rect 8706 11454 8718 11506
rect 14242 11454 14254 11506
rect 14306 11454 14318 11506
rect 18274 11454 18286 11506
rect 18338 11454 18350 11506
rect 23874 11454 23886 11506
rect 23938 11454 23950 11506
rect 28018 11454 28030 11506
rect 28082 11454 28094 11506
rect 33170 11454 33182 11506
rect 33234 11454 33246 11506
rect 34066 11454 34078 11506
rect 34130 11454 34142 11506
rect 15374 11442 15426 11454
rect 19294 11442 19346 11454
rect 34862 11442 34914 11454
rect 40238 11506 40290 11518
rect 40238 11442 40290 11454
rect 44830 11506 44882 11518
rect 53678 11506 53730 11518
rect 47506 11454 47518 11506
rect 47570 11454 47582 11506
rect 52882 11454 52894 11506
rect 52946 11454 52958 11506
rect 44830 11442 44882 11454
rect 53678 11442 53730 11454
rect 5182 11394 5234 11406
rect 5182 11330 5234 11342
rect 5630 11394 5682 11406
rect 5630 11330 5682 11342
rect 5966 11394 6018 11406
rect 5966 11330 6018 11342
rect 6302 11394 6354 11406
rect 6302 11330 6354 11342
rect 7310 11394 7362 11406
rect 7310 11330 7362 11342
rect 7422 11394 7474 11406
rect 7422 11330 7474 11342
rect 7534 11394 7586 11406
rect 15710 11394 15762 11406
rect 19854 11394 19906 11406
rect 20750 11394 20802 11406
rect 32398 11394 32450 11406
rect 36206 11394 36258 11406
rect 40350 11394 40402 11406
rect 43822 11394 43874 11406
rect 10210 11342 10222 11394
rect 10274 11342 10286 11394
rect 12226 11342 12238 11394
rect 12290 11342 12302 11394
rect 12674 11342 12686 11394
rect 12738 11342 12750 11394
rect 13458 11342 13470 11394
rect 13522 11342 13534 11394
rect 17938 11342 17950 11394
rect 18002 11342 18014 11394
rect 20290 11342 20302 11394
rect 20354 11342 20366 11394
rect 21522 11342 21534 11394
rect 21586 11342 21598 11394
rect 24322 11342 24334 11394
rect 24386 11342 24398 11394
rect 25330 11342 25342 11394
rect 25394 11342 25406 11394
rect 27010 11342 27022 11394
rect 27074 11342 27086 11394
rect 27570 11342 27582 11394
rect 27634 11342 27646 11394
rect 32946 11342 32958 11394
rect 33010 11342 33022 11394
rect 34402 11342 34414 11394
rect 34466 11342 34478 11394
rect 37762 11342 37774 11394
rect 37826 11342 37838 11394
rect 38882 11342 38894 11394
rect 38946 11342 38958 11394
rect 40898 11342 40910 11394
rect 40962 11342 40974 11394
rect 7534 11330 7586 11342
rect 15710 11330 15762 11342
rect 19854 11330 19906 11342
rect 20750 11330 20802 11342
rect 32398 11330 32450 11342
rect 36206 11330 36258 11342
rect 40350 11330 40402 11342
rect 43822 11330 43874 11342
rect 44158 11394 44210 11406
rect 45490 11342 45502 11394
rect 45554 11342 45566 11394
rect 46386 11342 46398 11394
rect 46450 11342 46462 11394
rect 47618 11342 47630 11394
rect 47682 11342 47694 11394
rect 49970 11342 49982 11394
rect 50034 11342 50046 11394
rect 50754 11342 50766 11394
rect 50818 11342 50830 11394
rect 53218 11342 53230 11394
rect 53282 11342 53294 11394
rect 44158 11330 44210 11342
rect 1710 11282 1762 11294
rect 1710 11218 1762 11230
rect 2046 11282 2098 11294
rect 2046 11218 2098 11230
rect 5742 11282 5794 11294
rect 12910 11282 12962 11294
rect 7970 11230 7982 11282
rect 8034 11230 8046 11282
rect 8978 11230 8990 11282
rect 9042 11230 9054 11282
rect 5742 11218 5794 11230
rect 12910 11218 12962 11230
rect 13694 11282 13746 11294
rect 13694 11218 13746 11230
rect 13806 11282 13858 11294
rect 13806 11218 13858 11230
rect 16606 11282 16658 11294
rect 18734 11282 18786 11294
rect 36542 11282 36594 11294
rect 43934 11282 43986 11294
rect 54014 11282 54066 11294
rect 18050 11230 18062 11282
rect 18114 11230 18126 11282
rect 21858 11230 21870 11282
rect 21922 11230 21934 11282
rect 22418 11230 22430 11282
rect 22482 11230 22494 11282
rect 28018 11230 28030 11282
rect 28082 11230 28094 11282
rect 37314 11230 37326 11282
rect 37378 11230 37390 11282
rect 46722 11230 46734 11282
rect 46786 11230 46798 11282
rect 50866 11230 50878 11282
rect 50930 11230 50942 11282
rect 16606 11218 16658 11230
rect 18734 11218 18786 11230
rect 36542 11218 36594 11230
rect 43934 11218 43986 11230
rect 54014 11218 54066 11230
rect 2494 11170 2546 11182
rect 2494 11106 2546 11118
rect 17054 11170 17106 11182
rect 36318 11170 36370 11182
rect 22082 11118 22094 11170
rect 22146 11118 22158 11170
rect 17054 11106 17106 11118
rect 36318 11106 36370 11118
rect 54126 11170 54178 11182
rect 54126 11106 54178 11118
rect 1344 11002 58576 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 50558 11002
rect 50610 10950 50662 11002
rect 50714 10950 50766 11002
rect 50818 10950 58576 11002
rect 1344 10916 58576 10950
rect 2046 10834 2098 10846
rect 2046 10770 2098 10782
rect 5742 10834 5794 10846
rect 5742 10770 5794 10782
rect 6862 10834 6914 10846
rect 6862 10770 6914 10782
rect 7646 10834 7698 10846
rect 7646 10770 7698 10782
rect 10446 10834 10498 10846
rect 28142 10834 28194 10846
rect 47854 10834 47906 10846
rect 23202 10782 23214 10834
rect 23266 10782 23278 10834
rect 10446 10770 10498 10782
rect 28030 10778 28082 10790
rect 6078 10722 6130 10734
rect 6078 10658 6130 10670
rect 6190 10722 6242 10734
rect 6190 10658 6242 10670
rect 6974 10722 7026 10734
rect 6974 10658 7026 10670
rect 7198 10722 7250 10734
rect 11342 10722 11394 10734
rect 41234 10782 41246 10834
rect 41298 10782 41310 10834
rect 47282 10782 47294 10834
rect 47346 10782 47358 10834
rect 28142 10770 28194 10782
rect 47854 10770 47906 10782
rect 53230 10834 53282 10846
rect 53230 10770 53282 10782
rect 53342 10834 53394 10846
rect 53342 10770 53394 10782
rect 53902 10834 53954 10846
rect 53902 10770 53954 10782
rect 54238 10834 54290 10846
rect 55010 10782 55022 10834
rect 55074 10782 55086 10834
rect 54238 10770 54290 10782
rect 10770 10670 10782 10722
rect 10834 10670 10846 10722
rect 12450 10670 12462 10722
rect 12514 10670 12526 10722
rect 14914 10670 14926 10722
rect 14978 10670 14990 10722
rect 15362 10670 15374 10722
rect 15426 10670 15438 10722
rect 28030 10714 28082 10726
rect 30158 10722 30210 10734
rect 39566 10722 39618 10734
rect 46286 10722 46338 10734
rect 32498 10670 32510 10722
rect 32562 10670 32574 10722
rect 38210 10670 38222 10722
rect 38274 10670 38286 10722
rect 42466 10670 42478 10722
rect 42530 10670 42542 10722
rect 44706 10670 44718 10722
rect 44770 10670 44782 10722
rect 46050 10670 46062 10722
rect 46114 10670 46126 10722
rect 7198 10658 7250 10670
rect 11342 10658 11394 10670
rect 30158 10658 30210 10670
rect 39566 10658 39618 10670
rect 46286 10658 46338 10670
rect 49198 10722 49250 10734
rect 49198 10658 49250 10670
rect 53790 10722 53842 10734
rect 53790 10658 53842 10670
rect 1710 10610 1762 10622
rect 1710 10546 1762 10558
rect 6414 10610 6466 10622
rect 6414 10546 6466 10558
rect 6526 10610 6578 10622
rect 6526 10546 6578 10558
rect 9662 10610 9714 10622
rect 9662 10546 9714 10558
rect 10110 10610 10162 10622
rect 10110 10546 10162 10558
rect 11118 10610 11170 10622
rect 11118 10546 11170 10558
rect 11790 10610 11842 10622
rect 22654 10610 22706 10622
rect 13570 10558 13582 10610
rect 13634 10558 13646 10610
rect 15586 10558 15598 10610
rect 15650 10558 15662 10610
rect 16594 10558 16606 10610
rect 16658 10558 16670 10610
rect 17826 10558 17838 10610
rect 17890 10558 17902 10610
rect 18498 10558 18510 10610
rect 18562 10558 18574 10610
rect 19394 10558 19406 10610
rect 19458 10558 19470 10610
rect 20402 10558 20414 10610
rect 20466 10558 20478 10610
rect 20962 10558 20974 10610
rect 21026 10558 21038 10610
rect 11790 10546 11842 10558
rect 22654 10546 22706 10558
rect 22878 10610 22930 10622
rect 22878 10546 22930 10558
rect 28926 10610 28978 10622
rect 47518 10610 47570 10622
rect 29362 10558 29374 10610
rect 29426 10558 29438 10610
rect 29810 10558 29822 10610
rect 29874 10558 29886 10610
rect 30594 10558 30606 10610
rect 30658 10558 30670 10610
rect 33506 10558 33518 10610
rect 33570 10558 33582 10610
rect 34066 10558 34078 10610
rect 34130 10558 34142 10610
rect 35074 10558 35086 10610
rect 35138 10558 35150 10610
rect 36418 10558 36430 10610
rect 36482 10558 36494 10610
rect 38098 10558 38110 10610
rect 38162 10558 38174 10610
rect 38994 10558 39006 10610
rect 39058 10558 39070 10610
rect 39778 10558 39790 10610
rect 39842 10558 39854 10610
rect 40002 10558 40014 10610
rect 40066 10558 40078 10610
rect 41570 10558 41582 10610
rect 41634 10558 41646 10610
rect 44930 10558 44942 10610
rect 44994 10558 45006 10610
rect 47058 10558 47070 10610
rect 47122 10558 47134 10610
rect 28926 10546 28978 10558
rect 47518 10546 47570 10558
rect 47854 10610 47906 10622
rect 47854 10546 47906 10558
rect 48190 10610 48242 10622
rect 54014 10610 54066 10622
rect 49858 10558 49870 10610
rect 49922 10558 49934 10610
rect 48190 10546 48242 10558
rect 54014 10546 54066 10558
rect 54686 10610 54738 10622
rect 54686 10546 54738 10558
rect 2494 10498 2546 10510
rect 2494 10434 2546 10446
rect 11566 10498 11618 10510
rect 31950 10498 32002 10510
rect 12114 10446 12126 10498
rect 12178 10446 12190 10498
rect 15698 10446 15710 10498
rect 15762 10446 15774 10498
rect 30370 10446 30382 10498
rect 30434 10446 30446 10498
rect 36530 10446 36542 10498
rect 36594 10446 36606 10498
rect 38434 10446 38446 10498
rect 38498 10446 38510 10498
rect 43026 10446 43038 10498
rect 43090 10446 43102 10498
rect 50082 10446 50094 10498
rect 50146 10446 50158 10498
rect 11566 10434 11618 10446
rect 31950 10434 32002 10446
rect 9774 10386 9826 10398
rect 9774 10322 9826 10334
rect 9998 10386 10050 10398
rect 28142 10386 28194 10398
rect 20514 10334 20526 10386
rect 20578 10334 20590 10386
rect 9998 10322 10050 10334
rect 28142 10322 28194 10334
rect 32174 10386 32226 10398
rect 39454 10386 39506 10398
rect 37426 10334 37438 10386
rect 37490 10334 37502 10386
rect 32174 10322 32226 10334
rect 39454 10322 39506 10334
rect 53454 10386 53506 10398
rect 53454 10322 53506 10334
rect 1344 10218 58576 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 58576 10218
rect 1344 10132 58576 10166
rect 14366 10050 14418 10062
rect 14366 9986 14418 9998
rect 23998 10050 24050 10062
rect 23998 9986 24050 9998
rect 26910 10050 26962 10062
rect 54450 9998 54462 10050
rect 54514 9998 54526 10050
rect 26910 9986 26962 9998
rect 7086 9938 7138 9950
rect 6626 9886 6638 9938
rect 6690 9886 6702 9938
rect 7086 9874 7138 9886
rect 8430 9938 8482 9950
rect 8430 9874 8482 9886
rect 10446 9938 10498 9950
rect 28478 9938 28530 9950
rect 31390 9938 31442 9950
rect 32958 9938 33010 9950
rect 38894 9938 38946 9950
rect 43934 9938 43986 9950
rect 20178 9886 20190 9938
rect 20242 9886 20254 9938
rect 29250 9886 29262 9938
rect 29314 9886 29326 9938
rect 32274 9886 32286 9938
rect 32338 9886 32350 9938
rect 34850 9886 34862 9938
rect 34914 9886 34926 9938
rect 37090 9886 37102 9938
rect 37154 9886 37166 9938
rect 43138 9886 43150 9938
rect 43202 9886 43214 9938
rect 10446 9874 10498 9886
rect 28478 9874 28530 9886
rect 31390 9874 31442 9886
rect 32958 9874 33010 9886
rect 38894 9874 38946 9886
rect 43934 9874 43986 9886
rect 44830 9938 44882 9950
rect 44830 9874 44882 9886
rect 53454 9938 53506 9950
rect 53454 9874 53506 9886
rect 12798 9826 12850 9838
rect 6402 9774 6414 9826
rect 6466 9774 6478 9826
rect 9986 9774 9998 9826
rect 10050 9774 10062 9826
rect 12798 9762 12850 9774
rect 14142 9826 14194 9838
rect 17054 9826 17106 9838
rect 25902 9826 25954 9838
rect 32622 9826 32674 9838
rect 15362 9774 15374 9826
rect 15426 9774 15438 9826
rect 16258 9774 16270 9826
rect 16322 9774 16334 9826
rect 18722 9774 18734 9826
rect 18786 9774 18798 9826
rect 19282 9774 19294 9826
rect 19346 9774 19358 9826
rect 20514 9774 20526 9826
rect 20578 9774 20590 9826
rect 23426 9774 23438 9826
rect 23490 9774 23502 9826
rect 26450 9774 26462 9826
rect 26514 9774 26526 9826
rect 30706 9774 30718 9826
rect 30770 9774 30782 9826
rect 14142 9762 14194 9774
rect 17054 9762 17106 9774
rect 25902 9762 25954 9774
rect 32622 9762 32674 9774
rect 32734 9826 32786 9838
rect 32734 9762 32786 9774
rect 33070 9826 33122 9838
rect 33070 9762 33122 9774
rect 33406 9826 33458 9838
rect 35086 9826 35138 9838
rect 34738 9774 34750 9826
rect 34802 9774 34814 9826
rect 33406 9762 33458 9774
rect 35086 9762 35138 9774
rect 35422 9826 35474 9838
rect 35422 9762 35474 9774
rect 37550 9826 37602 9838
rect 37550 9762 37602 9774
rect 38222 9826 38274 9838
rect 38222 9762 38274 9774
rect 38446 9826 38498 9838
rect 38446 9762 38498 9774
rect 39454 9826 39506 9838
rect 53118 9826 53170 9838
rect 40786 9774 40798 9826
rect 40850 9774 40862 9826
rect 41570 9774 41582 9826
rect 41634 9774 41646 9826
rect 43474 9774 43486 9826
rect 43538 9774 43550 9826
rect 45266 9774 45278 9826
rect 45330 9774 45342 9826
rect 39454 9762 39506 9774
rect 53118 9762 53170 9774
rect 53678 9826 53730 9838
rect 53678 9762 53730 9774
rect 53902 9826 53954 9838
rect 53902 9762 53954 9774
rect 54126 9826 54178 9838
rect 54126 9762 54178 9774
rect 7646 9714 7698 9726
rect 7646 9650 7698 9662
rect 7758 9714 7810 9726
rect 12686 9714 12738 9726
rect 8866 9662 8878 9714
rect 8930 9662 8942 9714
rect 7758 9650 7810 9662
rect 12686 9650 12738 9662
rect 14478 9714 14530 9726
rect 14478 9650 14530 9662
rect 14702 9714 14754 9726
rect 16942 9714 16994 9726
rect 15810 9662 15822 9714
rect 15874 9662 15886 9714
rect 14702 9650 14754 9662
rect 16942 9650 16994 9662
rect 17838 9714 17890 9726
rect 17838 9650 17890 9662
rect 17950 9714 18002 9726
rect 17950 9650 18002 9662
rect 21422 9714 21474 9726
rect 21422 9650 21474 9662
rect 21534 9714 21586 9726
rect 24782 9714 24834 9726
rect 23650 9662 23662 9714
rect 23714 9662 23726 9714
rect 21534 9650 21586 9662
rect 24782 9650 24834 9662
rect 24894 9714 24946 9726
rect 26238 9714 26290 9726
rect 26002 9662 26014 9714
rect 26066 9662 26078 9714
rect 24894 9650 24946 9662
rect 26238 9650 26290 9662
rect 28366 9714 28418 9726
rect 28366 9650 28418 9662
rect 28590 9714 28642 9726
rect 35758 9714 35810 9726
rect 51998 9714 52050 9726
rect 29474 9662 29486 9714
rect 29538 9662 29550 9714
rect 34514 9662 34526 9714
rect 34578 9662 34590 9714
rect 37874 9662 37886 9714
rect 37938 9662 37950 9714
rect 40562 9662 40574 9714
rect 40626 9662 40638 9714
rect 28590 9650 28642 9662
rect 35758 9650 35810 9662
rect 51998 9650 52050 9662
rect 53230 9714 53282 9726
rect 53230 9650 53282 9662
rect 7982 9602 8034 9614
rect 7982 9538 8034 9550
rect 12462 9602 12514 9614
rect 16718 9602 16770 9614
rect 16370 9550 16382 9602
rect 16434 9550 16446 9602
rect 12462 9538 12514 9550
rect 16718 9538 16770 9550
rect 18174 9602 18226 9614
rect 18174 9538 18226 9550
rect 21198 9602 21250 9614
rect 21198 9538 21250 9550
rect 24110 9602 24162 9614
rect 24110 9538 24162 9550
rect 24222 9602 24274 9614
rect 24222 9538 24274 9550
rect 24558 9602 24610 9614
rect 24558 9538 24610 9550
rect 32062 9602 32114 9614
rect 32062 9538 32114 9550
rect 32286 9602 32338 9614
rect 32286 9538 32338 9550
rect 35422 9602 35474 9614
rect 35422 9538 35474 9550
rect 38782 9602 38834 9614
rect 38782 9538 38834 9550
rect 39006 9602 39058 9614
rect 51662 9602 51714 9614
rect 42018 9550 42030 9602
rect 42082 9550 42094 9602
rect 39006 9538 39058 9550
rect 51662 9538 51714 9550
rect 51886 9602 51938 9614
rect 51886 9538 51938 9550
rect 1344 9434 58576 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 50558 9434
rect 50610 9382 50662 9434
rect 50714 9382 50766 9434
rect 50818 9382 58576 9434
rect 1344 9348 58576 9382
rect 5630 9266 5682 9278
rect 5630 9202 5682 9214
rect 7422 9266 7474 9278
rect 18734 9266 18786 9278
rect 14242 9214 14254 9266
rect 14306 9214 14318 9266
rect 15810 9214 15822 9266
rect 15874 9214 15886 9266
rect 7422 9202 7474 9214
rect 18734 9202 18786 9214
rect 19182 9266 19234 9278
rect 26126 9266 26178 9278
rect 19506 9214 19518 9266
rect 19570 9214 19582 9266
rect 19182 9202 19234 9214
rect 26126 9202 26178 9214
rect 27694 9266 27746 9278
rect 27694 9202 27746 9214
rect 30606 9266 30658 9278
rect 30606 9202 30658 9214
rect 30830 9266 30882 9278
rect 36094 9266 36146 9278
rect 38782 9266 38834 9278
rect 34290 9214 34302 9266
rect 34354 9214 34366 9266
rect 35186 9214 35198 9266
rect 35250 9214 35262 9266
rect 38322 9214 38334 9266
rect 38386 9214 38398 9266
rect 30830 9202 30882 9214
rect 36094 9202 36146 9214
rect 38782 9202 38834 9214
rect 43374 9266 43426 9278
rect 47070 9266 47122 9278
rect 44818 9214 44830 9266
rect 44882 9214 44894 9266
rect 43374 9202 43426 9214
rect 47070 9202 47122 9214
rect 48862 9266 48914 9278
rect 52882 9214 52894 9266
rect 52946 9214 52958 9266
rect 48862 9202 48914 9214
rect 2046 9154 2098 9166
rect 6526 9154 6578 9166
rect 6178 9102 6190 9154
rect 6242 9102 6254 9154
rect 2046 9090 2098 9102
rect 6526 9090 6578 9102
rect 6750 9154 6802 9166
rect 6750 9090 6802 9102
rect 7086 9154 7138 9166
rect 7086 9090 7138 9102
rect 8654 9154 8706 9166
rect 27470 9154 27522 9166
rect 30158 9154 30210 9166
rect 8978 9102 8990 9154
rect 9042 9102 9054 9154
rect 12562 9102 12574 9154
rect 12626 9102 12638 9154
rect 15138 9102 15150 9154
rect 15202 9102 15214 9154
rect 15474 9102 15486 9154
rect 15538 9102 15550 9154
rect 20626 9102 20638 9154
rect 20690 9102 20702 9154
rect 22866 9102 22878 9154
rect 22930 9102 22942 9154
rect 28242 9102 28254 9154
rect 28306 9102 28318 9154
rect 8654 9090 8706 9102
rect 27470 9090 27522 9102
rect 30158 9090 30210 9102
rect 31166 9154 31218 9166
rect 33182 9154 33234 9166
rect 36542 9154 36594 9166
rect 31826 9102 31838 9154
rect 31890 9102 31902 9154
rect 35298 9102 35310 9154
rect 35362 9102 35374 9154
rect 31166 9090 31218 9102
rect 33182 9090 33234 9102
rect 36542 9090 36594 9102
rect 37214 9154 37266 9166
rect 37214 9090 37266 9102
rect 37662 9154 37714 9166
rect 37662 9090 37714 9102
rect 37774 9154 37826 9166
rect 37774 9090 37826 9102
rect 38670 9154 38722 9166
rect 38670 9090 38722 9102
rect 39006 9154 39058 9166
rect 39006 9090 39058 9102
rect 39230 9154 39282 9166
rect 39230 9090 39282 9102
rect 40350 9154 40402 9166
rect 40350 9090 40402 9102
rect 42254 9154 42306 9166
rect 47182 9154 47234 9166
rect 43922 9102 43934 9154
rect 43986 9102 43998 9154
rect 46050 9102 46062 9154
rect 46114 9102 46126 9154
rect 42254 9090 42306 9102
rect 47182 9090 47234 9102
rect 49758 9154 49810 9166
rect 49758 9090 49810 9102
rect 50654 9154 50706 9166
rect 52098 9102 52110 9154
rect 52162 9102 52174 9154
rect 50654 9090 50706 9102
rect 1710 9042 1762 9054
rect 7982 9042 8034 9054
rect 5954 8990 5966 9042
rect 6018 8990 6030 9042
rect 1710 8978 1762 8990
rect 7982 8978 8034 8990
rect 9550 9042 9602 9054
rect 9550 8978 9602 8990
rect 9886 9042 9938 9054
rect 9886 8978 9938 8990
rect 10110 9042 10162 9054
rect 25230 9042 25282 9054
rect 13010 8990 13022 9042
rect 13074 8990 13086 9042
rect 13794 8990 13806 9042
rect 13858 8990 13870 9042
rect 14802 8990 14814 9042
rect 14866 8990 14878 9042
rect 17714 8990 17726 9042
rect 17778 8990 17790 9042
rect 17938 8990 17950 9042
rect 18002 8990 18014 9042
rect 21634 8990 21646 9042
rect 21698 8990 21710 9042
rect 23650 8990 23662 9042
rect 23714 8990 23726 9042
rect 24434 8990 24446 9042
rect 24498 8990 24510 9042
rect 10110 8978 10162 8990
rect 25230 8978 25282 8990
rect 25454 9042 25506 9054
rect 25454 8978 25506 8990
rect 27358 9042 27410 9054
rect 30494 9042 30546 9054
rect 28578 8990 28590 9042
rect 28642 8990 28654 9042
rect 29474 8990 29486 9042
rect 29538 8990 29550 9042
rect 27358 8978 27410 8990
rect 30494 8978 30546 8990
rect 32174 9042 32226 9054
rect 32174 8978 32226 8990
rect 33742 9042 33794 9054
rect 33742 8978 33794 8990
rect 33966 9042 34018 9054
rect 35870 9042 35922 9054
rect 35634 8990 35646 9042
rect 35698 8990 35710 9042
rect 33966 8978 34018 8990
rect 35870 8978 35922 8990
rect 36206 9042 36258 9054
rect 37886 9042 37938 9054
rect 36978 8990 36990 9042
rect 37042 8990 37054 9042
rect 36206 8978 36258 8990
rect 37886 8978 37938 8990
rect 40910 9042 40962 9054
rect 40910 8978 40962 8990
rect 41022 9042 41074 9054
rect 41022 8978 41074 8990
rect 41134 9042 41186 9054
rect 41134 8978 41186 8990
rect 41358 9042 41410 9054
rect 42366 9042 42418 9054
rect 41794 8990 41806 9042
rect 41858 8990 41870 9042
rect 42018 8990 42030 9042
rect 42082 8990 42094 9042
rect 41358 8978 41410 8990
rect 42366 8978 42418 8990
rect 42814 9042 42866 9054
rect 42814 8978 42866 8990
rect 43262 9042 43314 9054
rect 43262 8978 43314 8990
rect 43486 9042 43538 9054
rect 45726 9042 45778 9054
rect 44146 8990 44158 9042
rect 44210 8990 44222 9042
rect 44706 8990 44718 9042
rect 44770 8990 44782 9042
rect 43486 8978 43538 8990
rect 45726 8978 45778 8990
rect 46846 9042 46898 9054
rect 51214 9042 51266 9054
rect 48738 8990 48750 9042
rect 48802 8990 48814 9042
rect 49970 8990 49982 9042
rect 50034 8990 50046 9042
rect 46846 8978 46898 8990
rect 51214 8978 51266 8990
rect 51438 9042 51490 9054
rect 51438 8978 51490 8990
rect 51550 9042 51602 9054
rect 51550 8978 51602 8990
rect 51774 9042 51826 9054
rect 52546 8990 52558 9042
rect 52610 8990 52622 9042
rect 52882 8990 52894 9042
rect 52946 8990 52958 9042
rect 51774 8978 51826 8990
rect 2494 8930 2546 8942
rect 2494 8866 2546 8878
rect 6974 8930 7026 8942
rect 6974 8866 7026 8878
rect 9998 8930 10050 8942
rect 17490 8878 17502 8930
rect 17554 8878 17566 8930
rect 20066 8878 20078 8930
rect 20130 8878 20142 8930
rect 23986 8878 23998 8930
rect 24050 8878 24062 8930
rect 24322 8878 24334 8930
rect 24386 8878 24398 8930
rect 31154 8878 31166 8930
rect 31218 8878 31230 8930
rect 9998 8866 10050 8878
rect 25678 8818 25730 8830
rect 25678 8754 25730 8766
rect 31390 8818 31442 8830
rect 31390 8754 31442 8766
rect 33070 8818 33122 8830
rect 33070 8754 33122 8766
rect 33406 8818 33458 8830
rect 33406 8754 33458 8766
rect 39902 8818 39954 8830
rect 39902 8754 39954 8766
rect 40014 8818 40066 8830
rect 40014 8754 40066 8766
rect 40238 8818 40290 8830
rect 40238 8754 40290 8766
rect 48974 8818 49026 8830
rect 48974 8754 49026 8766
rect 49198 8818 49250 8830
rect 49198 8754 49250 8766
rect 50430 8818 50482 8830
rect 50430 8754 50482 8766
rect 50766 8818 50818 8830
rect 50766 8754 50818 8766
rect 1344 8650 58576 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 58576 8650
rect 1344 8564 58576 8598
rect 7422 8482 7474 8494
rect 7422 8418 7474 8430
rect 19182 8482 19234 8494
rect 19182 8418 19234 8430
rect 26910 8482 26962 8494
rect 39454 8482 39506 8494
rect 34402 8430 34414 8482
rect 34466 8430 34478 8482
rect 42578 8430 42590 8482
rect 42642 8430 42654 8482
rect 44258 8430 44270 8482
rect 44322 8430 44334 8482
rect 26910 8418 26962 8430
rect 39454 8418 39506 8430
rect 6526 8370 6578 8382
rect 14478 8370 14530 8382
rect 22094 8370 22146 8382
rect 29374 8370 29426 8382
rect 7746 8318 7758 8370
rect 7810 8318 7822 8370
rect 8194 8318 8206 8370
rect 8258 8318 8270 8370
rect 11666 8318 11678 8370
rect 11730 8318 11742 8370
rect 15922 8318 15934 8370
rect 15986 8318 15998 8370
rect 22866 8318 22878 8370
rect 22930 8318 22942 8370
rect 24098 8318 24110 8370
rect 24162 8318 24174 8370
rect 6526 8306 6578 8318
rect 14478 8306 14530 8318
rect 22094 8306 22146 8318
rect 29374 8306 29426 8318
rect 29710 8370 29762 8382
rect 42926 8370 42978 8382
rect 31042 8318 31054 8370
rect 31106 8318 31118 8370
rect 33506 8318 33518 8370
rect 33570 8318 33582 8370
rect 36418 8318 36430 8370
rect 36482 8318 36494 8370
rect 37090 8318 37102 8370
rect 37154 8318 37166 8370
rect 29710 8306 29762 8318
rect 42926 8306 42978 8318
rect 43150 8370 43202 8382
rect 43150 8306 43202 8318
rect 44942 8370 44994 8382
rect 52558 8370 52610 8382
rect 46162 8318 46174 8370
rect 46226 8318 46238 8370
rect 48850 8318 48862 8370
rect 48914 8318 48926 8370
rect 49410 8318 49422 8370
rect 49474 8318 49486 8370
rect 44942 8306 44994 8318
rect 52558 8306 52610 8318
rect 6750 8258 6802 8270
rect 6750 8194 6802 8206
rect 7086 8258 7138 8270
rect 11006 8258 11058 8270
rect 13582 8258 13634 8270
rect 15262 8258 15314 8270
rect 9650 8206 9662 8258
rect 9714 8206 9726 8258
rect 11218 8206 11230 8258
rect 11282 8206 11294 8258
rect 11778 8206 11790 8258
rect 11842 8206 11854 8258
rect 13794 8206 13806 8258
rect 13858 8206 13870 8258
rect 7086 8194 7138 8206
rect 11006 8194 11058 8206
rect 13582 8194 13634 8206
rect 15262 8194 15314 8206
rect 15374 8258 15426 8270
rect 20526 8258 20578 8270
rect 16930 8206 16942 8258
rect 16994 8206 17006 8258
rect 17826 8206 17838 8258
rect 17890 8206 17902 8258
rect 20066 8206 20078 8258
rect 20130 8206 20142 8258
rect 15374 8194 15426 8206
rect 20526 8194 20578 8206
rect 20750 8258 20802 8270
rect 20750 8194 20802 8206
rect 21310 8258 21362 8270
rect 22430 8258 22482 8270
rect 34078 8258 34130 8270
rect 35758 8258 35810 8270
rect 41134 8258 41186 8270
rect 44718 8258 44770 8270
rect 21522 8206 21534 8258
rect 21586 8206 21598 8258
rect 25554 8206 25566 8258
rect 25618 8206 25630 8258
rect 27458 8206 27470 8258
rect 27522 8206 27534 8258
rect 28354 8206 28366 8258
rect 28418 8206 28430 8258
rect 34290 8206 34302 8258
rect 34354 8206 34366 8258
rect 35522 8206 35534 8258
rect 35586 8206 35598 8258
rect 38546 8206 38558 8258
rect 38610 8206 38622 8258
rect 40786 8206 40798 8258
rect 40850 8206 40862 8258
rect 43474 8206 43486 8258
rect 43538 8206 43550 8258
rect 21310 8194 21362 8206
rect 22430 8194 22482 8206
rect 34078 8194 34130 8206
rect 35758 8194 35810 8206
rect 41134 8194 41186 8206
rect 44718 8194 44770 8206
rect 45054 8258 45106 8270
rect 45054 8194 45106 8206
rect 45278 8258 45330 8270
rect 53006 8258 53058 8270
rect 47282 8206 47294 8258
rect 47346 8206 47358 8258
rect 49746 8206 49758 8258
rect 49810 8206 49822 8258
rect 50866 8206 50878 8258
rect 50930 8206 50942 8258
rect 45278 8194 45330 8206
rect 53006 8194 53058 8206
rect 53230 8258 53282 8270
rect 53230 8194 53282 8206
rect 53454 8258 53506 8270
rect 53454 8194 53506 8206
rect 53902 8258 53954 8270
rect 53902 8194 53954 8206
rect 54014 8258 54066 8270
rect 54014 8194 54066 8206
rect 7646 8146 7698 8158
rect 12686 8146 12738 8158
rect 8642 8094 8654 8146
rect 8706 8094 8718 8146
rect 12338 8094 12350 8146
rect 12402 8094 12414 8146
rect 7646 8082 7698 8094
rect 12686 8082 12738 8094
rect 12798 8146 12850 8158
rect 12798 8082 12850 8094
rect 15486 8146 15538 8158
rect 23438 8146 23490 8158
rect 16706 8094 16718 8146
rect 16770 8094 16782 8146
rect 15486 8082 15538 8094
rect 23438 8082 23490 8094
rect 23550 8146 23602 8158
rect 29150 8146 29202 8158
rect 32846 8146 32898 8158
rect 24546 8094 24558 8146
rect 24610 8094 24622 8146
rect 27570 8094 27582 8146
rect 27634 8094 27646 8146
rect 31154 8094 31166 8146
rect 31218 8094 31230 8146
rect 23550 8082 23602 8094
rect 29150 8082 29202 8094
rect 32846 8082 32898 8094
rect 36094 8146 36146 8158
rect 43710 8146 43762 8158
rect 37650 8094 37662 8146
rect 37714 8094 37726 8146
rect 40450 8094 40462 8146
rect 40514 8094 40526 8146
rect 36094 8082 36146 8094
rect 43710 8082 43762 8094
rect 43822 8146 43874 8158
rect 54238 8146 54290 8158
rect 48290 8094 48302 8146
rect 48354 8094 48366 8146
rect 51426 8094 51438 8146
rect 51490 8094 51502 8146
rect 43822 8082 43874 8094
rect 54238 8082 54290 8094
rect 6974 8034 7026 8046
rect 6974 7970 7026 7982
rect 13022 8034 13074 8046
rect 13022 7970 13074 7982
rect 23214 8034 23266 8046
rect 36318 8034 36370 8046
rect 41694 8034 41746 8046
rect 28466 7982 28478 8034
rect 28530 7982 28542 8034
rect 40226 7982 40238 8034
rect 40290 7982 40302 8034
rect 23214 7970 23266 7982
rect 36318 7970 36370 7982
rect 41694 7970 41746 7982
rect 53790 8034 53842 8046
rect 53790 7970 53842 7982
rect 1344 7866 58576 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 50558 7866
rect 50610 7814 50662 7866
rect 50714 7814 50766 7866
rect 50818 7814 58576 7866
rect 1344 7780 58576 7814
rect 8766 7698 8818 7710
rect 8766 7634 8818 7646
rect 8878 7698 8930 7710
rect 8878 7634 8930 7646
rect 8990 7698 9042 7710
rect 8990 7634 9042 7646
rect 10446 7698 10498 7710
rect 10446 7634 10498 7646
rect 12798 7698 12850 7710
rect 12798 7634 12850 7646
rect 14142 7698 14194 7710
rect 14142 7634 14194 7646
rect 14926 7698 14978 7710
rect 14926 7634 14978 7646
rect 15374 7698 15426 7710
rect 15374 7634 15426 7646
rect 25342 7698 25394 7710
rect 25342 7634 25394 7646
rect 25678 7698 25730 7710
rect 25678 7634 25730 7646
rect 26798 7698 26850 7710
rect 32622 7698 32674 7710
rect 27570 7646 27582 7698
rect 27634 7646 27646 7698
rect 26798 7634 26850 7646
rect 32622 7634 32674 7646
rect 34190 7698 34242 7710
rect 45726 7698 45778 7710
rect 48302 7698 48354 7710
rect 34850 7646 34862 7698
rect 34914 7646 34926 7698
rect 47618 7646 47630 7698
rect 47682 7646 47694 7698
rect 34190 7634 34242 7646
rect 45726 7634 45778 7646
rect 48302 7634 48354 7646
rect 49534 7698 49586 7710
rect 49534 7634 49586 7646
rect 53342 7698 53394 7710
rect 53342 7634 53394 7646
rect 11790 7586 11842 7598
rect 11790 7522 11842 7534
rect 11902 7586 11954 7598
rect 11902 7522 11954 7534
rect 12350 7586 12402 7598
rect 12350 7522 12402 7534
rect 19406 7586 19458 7598
rect 26574 7586 26626 7598
rect 30158 7586 30210 7598
rect 20514 7534 20526 7586
rect 20578 7534 20590 7586
rect 24434 7534 24446 7586
rect 24498 7534 24510 7586
rect 26002 7534 26014 7586
rect 26066 7534 26078 7586
rect 27794 7534 27806 7586
rect 27858 7534 27870 7586
rect 28018 7534 28030 7586
rect 28082 7534 28094 7586
rect 19406 7522 19458 7534
rect 26574 7522 26626 7534
rect 30158 7522 30210 7534
rect 33070 7586 33122 7598
rect 39342 7586 39394 7598
rect 37090 7534 37102 7586
rect 37154 7534 37166 7586
rect 33070 7522 33122 7534
rect 39342 7522 39394 7534
rect 47070 7586 47122 7598
rect 47070 7522 47122 7534
rect 47182 7586 47234 7598
rect 47182 7522 47234 7534
rect 48078 7586 48130 7598
rect 48078 7522 48130 7534
rect 50206 7586 50258 7598
rect 50206 7522 50258 7534
rect 50430 7586 50482 7598
rect 50430 7522 50482 7534
rect 50542 7586 50594 7598
rect 51202 7534 51214 7586
rect 51266 7534 51278 7586
rect 50542 7522 50594 7534
rect 9550 7474 9602 7486
rect 8418 7422 8430 7474
rect 8482 7422 8494 7474
rect 9550 7410 9602 7422
rect 9998 7474 10050 7486
rect 9998 7410 10050 7422
rect 10782 7474 10834 7486
rect 10782 7410 10834 7422
rect 11006 7474 11058 7486
rect 11006 7410 11058 7422
rect 11566 7474 11618 7486
rect 11566 7410 11618 7422
rect 15262 7474 15314 7486
rect 15262 7410 15314 7422
rect 15598 7474 15650 7486
rect 16382 7474 16434 7486
rect 16034 7422 16046 7474
rect 16098 7422 16110 7474
rect 15598 7410 15650 7422
rect 16382 7410 16434 7422
rect 16606 7474 16658 7486
rect 19966 7474 20018 7486
rect 26350 7474 26402 7486
rect 18162 7422 18174 7474
rect 18226 7422 18238 7474
rect 18610 7422 18622 7474
rect 18674 7422 18686 7474
rect 20290 7422 20302 7474
rect 20354 7422 20366 7474
rect 22754 7422 22766 7474
rect 22818 7422 22830 7474
rect 24098 7422 24110 7474
rect 24162 7422 24174 7474
rect 16606 7410 16658 7422
rect 19966 7410 20018 7422
rect 26350 7410 26402 7422
rect 27022 7474 27074 7486
rect 27022 7410 27074 7422
rect 27246 7474 27298 7486
rect 30270 7474 30322 7486
rect 31726 7474 31778 7486
rect 29138 7422 29150 7474
rect 29202 7422 29214 7474
rect 30594 7422 30606 7474
rect 30658 7422 30670 7474
rect 27246 7410 27298 7422
rect 30270 7410 30322 7422
rect 31726 7410 31778 7422
rect 31950 7474 32002 7486
rect 31950 7410 32002 7422
rect 33294 7474 33346 7486
rect 33294 7410 33346 7422
rect 33742 7474 33794 7486
rect 35870 7474 35922 7486
rect 34626 7422 34638 7474
rect 34690 7422 34702 7474
rect 35634 7422 35646 7474
rect 35698 7422 35710 7474
rect 33742 7410 33794 7422
rect 35870 7410 35922 7422
rect 36206 7474 36258 7486
rect 36206 7410 36258 7422
rect 36318 7474 36370 7486
rect 39230 7474 39282 7486
rect 37202 7422 37214 7474
rect 37266 7422 37278 7474
rect 37538 7422 37550 7474
rect 37602 7422 37614 7474
rect 38546 7422 38558 7474
rect 38610 7422 38622 7474
rect 36318 7410 36370 7422
rect 39230 7410 39282 7422
rect 39454 7474 39506 7486
rect 46062 7474 46114 7486
rect 47966 7474 48018 7486
rect 39890 7422 39902 7474
rect 39954 7422 39966 7474
rect 41122 7422 41134 7474
rect 41186 7422 41198 7474
rect 42914 7422 42926 7474
rect 42978 7422 42990 7474
rect 43922 7422 43934 7474
rect 43986 7422 43998 7474
rect 46834 7422 46846 7474
rect 46898 7422 46910 7474
rect 39454 7410 39506 7422
rect 46062 7410 46114 7422
rect 47966 7410 48018 7422
rect 48750 7474 48802 7486
rect 48750 7410 48802 7422
rect 48974 7474 49026 7486
rect 49422 7474 49474 7486
rect 49298 7422 49310 7474
rect 49362 7422 49374 7474
rect 48974 7410 49026 7422
rect 49422 7410 49474 7422
rect 49646 7474 49698 7486
rect 52434 7422 52446 7474
rect 52498 7422 52510 7474
rect 49646 7410 49698 7422
rect 18734 7362 18786 7374
rect 14242 7310 14254 7362
rect 14306 7310 14318 7362
rect 20850 7310 20862 7362
rect 20914 7310 20926 7362
rect 22418 7310 22430 7362
rect 22482 7310 22494 7362
rect 28914 7310 28926 7362
rect 28978 7310 28990 7362
rect 41234 7310 41246 7362
rect 41298 7310 41310 7362
rect 43586 7310 43598 7362
rect 43650 7310 43662 7362
rect 44370 7310 44382 7362
rect 44434 7310 44446 7362
rect 50978 7310 50990 7362
rect 51042 7310 51054 7362
rect 18734 7298 18786 7310
rect 9774 7250 9826 7262
rect 12238 7250 12290 7262
rect 11330 7198 11342 7250
rect 11394 7198 11406 7250
rect 9774 7186 9826 7198
rect 12238 7186 12290 7198
rect 13918 7250 13970 7262
rect 32174 7250 32226 7262
rect 29250 7198 29262 7250
rect 29314 7198 29326 7250
rect 13918 7186 13970 7198
rect 32174 7186 32226 7198
rect 33518 7250 33570 7262
rect 35298 7198 35310 7250
rect 35362 7198 35374 7250
rect 33518 7186 33570 7198
rect 1344 7082 58576 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 58576 7082
rect 1344 6996 58576 7030
rect 10670 6914 10722 6926
rect 37438 6914 37490 6926
rect 15474 6862 15486 6914
rect 15538 6862 15550 6914
rect 10670 6850 10722 6862
rect 37438 6850 37490 6862
rect 37886 6914 37938 6926
rect 37886 6850 37938 6862
rect 44830 6914 44882 6926
rect 44830 6850 44882 6862
rect 52782 6914 52834 6926
rect 52782 6850 52834 6862
rect 52894 6914 52946 6926
rect 52894 6850 52946 6862
rect 53230 6914 53282 6926
rect 53230 6850 53282 6862
rect 11342 6802 11394 6814
rect 18062 6802 18114 6814
rect 36990 6802 37042 6814
rect 10994 6750 11006 6802
rect 11058 6750 11070 6802
rect 11666 6750 11678 6802
rect 11730 6750 11742 6802
rect 13570 6750 13582 6802
rect 13634 6750 13646 6802
rect 16482 6750 16494 6802
rect 16546 6750 16558 6802
rect 22194 6750 22206 6802
rect 22258 6750 22270 6802
rect 23986 6750 23998 6802
rect 24050 6750 24062 6802
rect 11342 6738 11394 6750
rect 18062 6738 18114 6750
rect 36990 6738 37042 6750
rect 37214 6802 37266 6814
rect 37214 6738 37266 6750
rect 40350 6802 40402 6814
rect 44942 6802 44994 6814
rect 41570 6750 41582 6802
rect 41634 6750 41646 6802
rect 44146 6750 44158 6802
rect 44210 6750 44222 6802
rect 50754 6750 50766 6802
rect 50818 6750 50830 6802
rect 40350 6738 40402 6750
rect 44942 6738 44994 6750
rect 9326 6690 9378 6702
rect 9326 6626 9378 6638
rect 9662 6690 9714 6702
rect 9662 6626 9714 6638
rect 12462 6690 12514 6702
rect 17278 6690 17330 6702
rect 14018 6638 14030 6690
rect 14082 6638 14094 6690
rect 15138 6638 15150 6690
rect 15202 6638 15214 6690
rect 16370 6638 16382 6690
rect 16434 6638 16446 6690
rect 12462 6626 12514 6638
rect 17278 6626 17330 6638
rect 17950 6690 18002 6702
rect 17950 6626 18002 6638
rect 18510 6690 18562 6702
rect 18510 6626 18562 6638
rect 18734 6690 18786 6702
rect 22542 6690 22594 6702
rect 24558 6690 24610 6702
rect 25454 6690 25506 6702
rect 22082 6638 22094 6690
rect 22146 6638 22158 6690
rect 22978 6638 22990 6690
rect 23042 6638 23054 6690
rect 24098 6638 24110 6690
rect 24162 6638 24174 6690
rect 24770 6638 24782 6690
rect 24834 6638 24846 6690
rect 18734 6626 18786 6638
rect 22542 6626 22594 6638
rect 24558 6626 24610 6638
rect 25454 6626 25506 6638
rect 28142 6690 28194 6702
rect 28142 6626 28194 6638
rect 31390 6690 31442 6702
rect 32398 6690 32450 6702
rect 53118 6690 53170 6702
rect 31826 6638 31838 6690
rect 31890 6638 31902 6690
rect 32722 6638 32734 6690
rect 32786 6638 32798 6690
rect 34290 6638 34302 6690
rect 34354 6638 34366 6690
rect 38994 6638 39006 6690
rect 39058 6638 39070 6690
rect 42690 6638 42702 6690
rect 42754 6638 42766 6690
rect 46386 6638 46398 6690
rect 46450 6638 46462 6690
rect 47282 6638 47294 6690
rect 47346 6638 47358 6690
rect 50642 6638 50654 6690
rect 50706 6638 50718 6690
rect 51426 6638 51438 6690
rect 51490 6638 51502 6690
rect 31390 6626 31442 6638
rect 32398 6626 32450 6638
rect 53118 6626 53170 6638
rect 9438 6578 9490 6590
rect 9438 6514 9490 6526
rect 10894 6578 10946 6590
rect 10894 6514 10946 6526
rect 11566 6578 11618 6590
rect 11566 6514 11618 6526
rect 12350 6578 12402 6590
rect 12350 6514 12402 6526
rect 19854 6578 19906 6590
rect 19854 6514 19906 6526
rect 20190 6578 20242 6590
rect 20190 6514 20242 6526
rect 20302 6578 20354 6590
rect 27806 6578 27858 6590
rect 23650 6526 23662 6578
rect 23714 6526 23726 6578
rect 20302 6514 20354 6526
rect 27806 6514 27858 6526
rect 27918 6578 27970 6590
rect 27918 6514 27970 6526
rect 30494 6578 30546 6590
rect 36094 6578 36146 6590
rect 40686 6578 40738 6590
rect 33618 6526 33630 6578
rect 33682 6526 33694 6578
rect 34514 6526 34526 6578
rect 34578 6526 34590 6578
rect 38546 6526 38558 6578
rect 38610 6526 38622 6578
rect 40114 6526 40126 6578
rect 40178 6526 40190 6578
rect 30494 6514 30546 6526
rect 36094 6514 36146 6526
rect 40686 6514 40738 6526
rect 41022 6578 41074 6590
rect 49534 6578 49586 6590
rect 43474 6526 43486 6578
rect 43538 6526 43550 6578
rect 46834 6526 46846 6578
rect 46898 6526 46910 6578
rect 50306 6526 50318 6578
rect 50370 6526 50382 6578
rect 41022 6514 41074 6526
rect 49534 6514 49586 6526
rect 12126 6466 12178 6478
rect 12126 6402 12178 6414
rect 12574 6466 12626 6478
rect 12574 6402 12626 6414
rect 17726 6466 17778 6478
rect 17726 6402 17778 6414
rect 18174 6466 18226 6478
rect 20526 6466 20578 6478
rect 19058 6414 19070 6466
rect 19122 6414 19134 6466
rect 18174 6402 18226 6414
rect 20526 6402 20578 6414
rect 31054 6466 31106 6478
rect 31054 6402 31106 6414
rect 36430 6466 36482 6478
rect 36430 6402 36482 6414
rect 45054 6466 45106 6478
rect 45054 6402 45106 6414
rect 45614 6466 45666 6478
rect 49982 6466 50034 6478
rect 47394 6414 47406 6466
rect 47458 6414 47470 6466
rect 45614 6402 45666 6414
rect 49982 6402 50034 6414
rect 1344 6298 58576 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 50558 6298
rect 50610 6246 50662 6298
rect 50714 6246 50766 6298
rect 50818 6246 58576 6298
rect 1344 6212 58576 6246
rect 12238 6130 12290 6142
rect 12238 6066 12290 6078
rect 16270 6130 16322 6142
rect 16270 6066 16322 6078
rect 16494 6130 16546 6142
rect 42702 6130 42754 6142
rect 35858 6078 35870 6130
rect 35922 6078 35934 6130
rect 40002 6078 40014 6130
rect 40066 6078 40078 6130
rect 41906 6078 41918 6130
rect 41970 6078 41982 6130
rect 16494 6066 16546 6078
rect 42702 6066 42754 6078
rect 46062 6130 46114 6142
rect 46062 6066 46114 6078
rect 48862 6130 48914 6142
rect 51886 6130 51938 6142
rect 51650 6078 51662 6130
rect 51714 6078 51726 6130
rect 48862 6066 48914 6078
rect 51886 6066 51938 6078
rect 52670 6130 52722 6142
rect 52670 6066 52722 6078
rect 12350 6018 12402 6030
rect 12350 5954 12402 5966
rect 13806 6018 13858 6030
rect 13806 5954 13858 5966
rect 16158 6018 16210 6030
rect 16158 5954 16210 5966
rect 34190 6018 34242 6030
rect 38670 6018 38722 6030
rect 52110 6018 52162 6030
rect 34962 5966 34974 6018
rect 35026 5966 35038 6018
rect 41010 5966 41022 6018
rect 41074 5966 41086 6018
rect 49298 5966 49310 6018
rect 49362 5966 49374 6018
rect 34190 5954 34242 5966
rect 38670 5954 38722 5966
rect 52110 5954 52162 5966
rect 52222 6018 52274 6030
rect 52222 5954 52274 5966
rect 12910 5906 12962 5918
rect 29486 5906 29538 5918
rect 13122 5854 13134 5906
rect 13186 5854 13198 5906
rect 19058 5854 19070 5906
rect 19122 5854 19134 5906
rect 20850 5854 20862 5906
rect 20914 5854 20926 5906
rect 21634 5854 21646 5906
rect 21698 5854 21710 5906
rect 12910 5842 12962 5854
rect 29486 5842 29538 5854
rect 30046 5906 30098 5918
rect 30942 5906 30994 5918
rect 33070 5906 33122 5918
rect 30482 5854 30494 5906
rect 30546 5854 30558 5906
rect 31378 5854 31390 5906
rect 31442 5854 31454 5906
rect 30046 5842 30098 5854
rect 30942 5842 30994 5854
rect 33070 5842 33122 5854
rect 34078 5906 34130 5918
rect 34078 5842 34130 5854
rect 34414 5906 34466 5918
rect 43150 5906 43202 5918
rect 36082 5854 36094 5906
rect 36146 5854 36158 5906
rect 36530 5854 36542 5906
rect 36594 5854 36606 5906
rect 37762 5854 37774 5906
rect 37826 5854 37838 5906
rect 39330 5854 39342 5906
rect 39394 5854 39406 5906
rect 40226 5854 40238 5906
rect 40290 5854 40302 5906
rect 41346 5854 41358 5906
rect 41410 5854 41422 5906
rect 41794 5854 41806 5906
rect 41858 5854 41870 5906
rect 34414 5842 34466 5854
rect 43150 5842 43202 5854
rect 43374 5906 43426 5918
rect 43374 5842 43426 5854
rect 43598 5906 43650 5918
rect 45950 5906 46002 5918
rect 44034 5854 44046 5906
rect 44098 5854 44110 5906
rect 44594 5854 44606 5906
rect 44658 5854 44670 5906
rect 45378 5854 45390 5906
rect 45442 5854 45454 5906
rect 43598 5842 43650 5854
rect 45950 5842 46002 5854
rect 48974 5906 49026 5918
rect 51326 5906 51378 5918
rect 49970 5854 49982 5906
rect 50034 5854 50046 5906
rect 50418 5854 50430 5906
rect 50482 5854 50494 5906
rect 48974 5842 49026 5854
rect 51326 5842 51378 5854
rect 29262 5794 29314 5806
rect 19170 5742 19182 5794
rect 19234 5742 19246 5794
rect 21858 5742 21870 5794
rect 21922 5742 21934 5794
rect 29262 5730 29314 5742
rect 31838 5794 31890 5806
rect 31838 5730 31890 5742
rect 32622 5794 32674 5806
rect 42478 5794 42530 5806
rect 46622 5794 46674 5806
rect 33506 5742 33518 5794
rect 33570 5742 33582 5794
rect 39554 5742 39566 5794
rect 39618 5742 39630 5794
rect 45154 5742 45166 5794
rect 45218 5742 45230 5794
rect 32622 5730 32674 5742
rect 42478 5730 42530 5742
rect 46622 5730 46674 5742
rect 47070 5794 47122 5806
rect 47070 5730 47122 5742
rect 46062 5682 46114 5694
rect 22306 5630 22318 5682
rect 22370 5630 22382 5682
rect 46062 5618 46114 5630
rect 48862 5682 48914 5694
rect 48862 5618 48914 5630
rect 1344 5514 58576 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 58576 5514
rect 1344 5428 58576 5462
rect 20750 5346 20802 5358
rect 20750 5282 20802 5294
rect 22094 5346 22146 5358
rect 31166 5346 31218 5358
rect 22418 5294 22430 5346
rect 22482 5294 22494 5346
rect 22094 5282 22146 5294
rect 31166 5282 31218 5294
rect 47518 5346 47570 5358
rect 47518 5282 47570 5294
rect 21870 5234 21922 5246
rect 17938 5182 17950 5234
rect 18002 5182 18014 5234
rect 21870 5170 21922 5182
rect 30942 5234 30994 5246
rect 30942 5170 30994 5182
rect 33518 5234 33570 5246
rect 37438 5234 37490 5246
rect 45614 5234 45666 5246
rect 46958 5234 47010 5246
rect 35858 5182 35870 5234
rect 35922 5182 35934 5234
rect 40114 5182 40126 5234
rect 40178 5182 40190 5234
rect 41794 5182 41806 5234
rect 41858 5182 41870 5234
rect 45938 5182 45950 5234
rect 46002 5182 46014 5234
rect 49522 5182 49534 5234
rect 49586 5182 49598 5234
rect 33518 5170 33570 5182
rect 37438 5170 37490 5182
rect 45614 5170 45666 5182
rect 46958 5170 47010 5182
rect 29710 5122 29762 5134
rect 31950 5122 32002 5134
rect 19394 5070 19406 5122
rect 19458 5070 19470 5122
rect 28354 5070 28366 5122
rect 28418 5070 28430 5122
rect 31602 5070 31614 5122
rect 31666 5070 31678 5122
rect 29710 5058 29762 5070
rect 31950 5058 32002 5070
rect 32174 5122 32226 5134
rect 43486 5122 43538 5134
rect 32498 5070 32510 5122
rect 32562 5070 32574 5122
rect 35746 5070 35758 5122
rect 35810 5070 35822 5122
rect 36418 5070 36430 5122
rect 36482 5070 36494 5122
rect 39442 5070 39454 5122
rect 39506 5070 39518 5122
rect 40562 5070 40574 5122
rect 40626 5070 40638 5122
rect 42242 5070 42254 5122
rect 42306 5070 42318 5122
rect 43026 5070 43038 5122
rect 43090 5070 43102 5122
rect 32174 5058 32226 5070
rect 43486 5058 43538 5070
rect 43598 5122 43650 5134
rect 43598 5058 43650 5070
rect 43934 5122 43986 5134
rect 43934 5058 43986 5070
rect 44830 5122 44882 5134
rect 47182 5122 47234 5134
rect 46050 5070 46062 5122
rect 46114 5070 46126 5122
rect 44830 5058 44882 5070
rect 47182 5058 47234 5070
rect 47742 5122 47794 5134
rect 47742 5058 47794 5070
rect 49086 5122 49138 5134
rect 49086 5058 49138 5070
rect 49982 5122 50034 5134
rect 49982 5058 50034 5070
rect 28590 5010 28642 5022
rect 18386 4958 18398 5010
rect 18450 4958 18462 5010
rect 28590 4946 28642 4958
rect 30046 5010 30098 5022
rect 44158 5010 44210 5022
rect 31714 4958 31726 5010
rect 31778 4958 31790 5010
rect 30046 4946 30098 4958
rect 44158 4946 44210 4958
rect 44270 5010 44322 5022
rect 47966 5010 48018 5022
rect 45154 4958 45166 5010
rect 45218 4958 45230 5010
rect 44270 4946 44322 4958
rect 47966 4946 48018 4958
rect 48078 5010 48130 5022
rect 50306 4958 50318 5010
rect 50370 4958 50382 5010
rect 48078 4946 48130 4958
rect 29374 4898 29426 4910
rect 29374 4834 29426 4846
rect 30382 4898 30434 4910
rect 30382 4834 30434 4846
rect 35982 4898 36034 4910
rect 35982 4834 36034 4846
rect 36206 4898 36258 4910
rect 36206 4834 36258 4846
rect 43262 4898 43314 4910
rect 43262 4834 43314 4846
rect 43374 4898 43426 4910
rect 43374 4834 43426 4846
rect 1344 4730 58576 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 50558 4730
rect 50610 4678 50662 4730
rect 50714 4678 50766 4730
rect 50818 4678 58576 4730
rect 1344 4644 58576 4678
rect 27694 4562 27746 4574
rect 27694 4498 27746 4510
rect 32622 4562 32674 4574
rect 40350 4562 40402 4574
rect 43822 4562 43874 4574
rect 45390 4562 45442 4574
rect 37762 4510 37774 4562
rect 37826 4510 37838 4562
rect 41682 4510 41694 4562
rect 41746 4510 41758 4562
rect 44706 4510 44718 4562
rect 44770 4510 44782 4562
rect 46050 4510 46062 4562
rect 46114 4510 46126 4562
rect 32622 4498 32674 4510
rect 40350 4498 40402 4510
rect 43822 4498 43874 4510
rect 45390 4498 45442 4510
rect 31950 4450 32002 4462
rect 46398 4450 46450 4462
rect 31714 4398 31726 4450
rect 31778 4398 31790 4450
rect 33954 4398 33966 4450
rect 34018 4398 34030 4450
rect 34850 4398 34862 4450
rect 34914 4398 34926 4450
rect 36642 4398 36654 4450
rect 36706 4398 36718 4450
rect 38994 4398 39006 4450
rect 39058 4398 39070 4450
rect 40898 4398 40910 4450
rect 40962 4398 40974 4450
rect 31950 4386 32002 4398
rect 46398 4386 46450 4398
rect 31614 4338 31666 4350
rect 42254 4338 42306 4350
rect 28802 4286 28814 4338
rect 28866 4286 28878 4338
rect 32162 4286 32174 4338
rect 32226 4286 32238 4338
rect 34402 4286 34414 4338
rect 34466 4286 34478 4338
rect 36306 4286 36318 4338
rect 36370 4286 36382 4338
rect 36978 4286 36990 4338
rect 37042 4286 37054 4338
rect 39218 4286 39230 4338
rect 39282 4286 39294 4338
rect 41122 4286 41134 4338
rect 41186 4286 41198 4338
rect 31614 4274 31666 4286
rect 42254 4274 42306 4286
rect 42478 4338 42530 4350
rect 42478 4274 42530 4286
rect 42702 4338 42754 4350
rect 42702 4274 42754 4286
rect 43150 4338 43202 4350
rect 43150 4274 43202 4286
rect 43262 4338 43314 4350
rect 43262 4274 43314 4286
rect 43486 4338 43538 4350
rect 43486 4274 43538 4286
rect 44382 4338 44434 4350
rect 44930 4286 44942 4338
rect 44994 4286 45006 4338
rect 45602 4286 45614 4338
rect 45666 4286 45678 4338
rect 44382 4274 44434 4286
rect 25342 4226 25394 4238
rect 25342 4162 25394 4174
rect 28254 4226 28306 4238
rect 42030 4226 42082 4238
rect 34962 4174 34974 4226
rect 35026 4174 35038 4226
rect 28254 4162 28306 4174
rect 42030 4162 42082 4174
rect 46846 4226 46898 4238
rect 46846 4162 46898 4174
rect 47294 4226 47346 4238
rect 47294 4162 47346 4174
rect 47742 4226 47794 4238
rect 47742 4162 47794 4174
rect 48190 4226 48242 4238
rect 48190 4162 48242 4174
rect 48862 4226 48914 4238
rect 48862 4162 48914 4174
rect 49758 4226 49810 4238
rect 49758 4162 49810 4174
rect 29486 4114 29538 4126
rect 29486 4050 29538 4062
rect 1344 3946 58576 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 58576 3946
rect 1344 3860 58576 3894
rect 40014 3778 40066 3790
rect 40014 3714 40066 3726
rect 41134 3778 41186 3790
rect 41458 3726 41470 3778
rect 41522 3726 41534 3778
rect 41134 3714 41186 3726
rect 26798 3666 26850 3678
rect 26798 3602 26850 3614
rect 29262 3666 29314 3678
rect 29262 3602 29314 3614
rect 32398 3666 32450 3678
rect 32398 3602 32450 3614
rect 36990 3666 37042 3678
rect 36990 3602 37042 3614
rect 40350 3666 40402 3678
rect 40350 3602 40402 3614
rect 40910 3666 40962 3678
rect 40910 3602 40962 3614
rect 41806 3666 41858 3678
rect 41806 3602 41858 3614
rect 49310 3666 49362 3678
rect 49310 3602 49362 3614
rect 24894 3554 24946 3566
rect 39790 3554 39842 3566
rect 43934 3554 43986 3566
rect 45950 3554 46002 3566
rect 27682 3502 27694 3554
rect 27746 3502 27758 3554
rect 31154 3502 31166 3554
rect 31218 3502 31230 3554
rect 34626 3502 34638 3554
rect 34690 3502 34702 3554
rect 35298 3502 35310 3554
rect 35362 3502 35374 3554
rect 36418 3502 36430 3554
rect 36482 3502 36494 3554
rect 39106 3502 39118 3554
rect 39170 3502 39182 3554
rect 42242 3502 42254 3554
rect 42306 3502 42318 3554
rect 44482 3502 44494 3554
rect 44546 3502 44558 3554
rect 45154 3502 45166 3554
rect 45218 3502 45230 3554
rect 24894 3490 24946 3502
rect 39790 3490 39842 3502
rect 43934 3490 43986 3502
rect 45950 3490 46002 3502
rect 46622 3554 46674 3566
rect 49982 3554 50034 3566
rect 47618 3502 47630 3554
rect 47682 3502 47694 3554
rect 48178 3502 48190 3554
rect 48242 3502 48254 3554
rect 46622 3490 46674 3502
rect 49982 3490 50034 3502
rect 22206 3442 22258 3454
rect 22206 3378 22258 3390
rect 22430 3442 22482 3454
rect 24558 3442 24610 3454
rect 22754 3390 22766 3442
rect 22818 3390 22830 3442
rect 22430 3378 22482 3390
rect 24558 3378 24610 3390
rect 28366 3442 28418 3454
rect 28366 3378 28418 3390
rect 28702 3442 28754 3454
rect 28702 3378 28754 3390
rect 35086 3442 35138 3454
rect 42702 3442 42754 3454
rect 38882 3390 38894 3442
rect 38946 3390 38958 3442
rect 35086 3378 35138 3390
rect 42702 3378 42754 3390
rect 43038 3442 43090 3454
rect 43038 3378 43090 3390
rect 43598 3442 43650 3454
rect 44942 3442 44994 3454
rect 46286 3442 46338 3454
rect 44258 3390 44270 3442
rect 44322 3390 44334 3442
rect 45602 3390 45614 3442
rect 45666 3390 45678 3442
rect 43598 3378 43650 3390
rect 44942 3378 44994 3390
rect 46286 3378 46338 3390
rect 47406 3442 47458 3454
rect 47406 3378 47458 3390
rect 48414 3442 48466 3454
rect 48414 3378 48466 3390
rect 50318 3442 50370 3454
rect 50318 3378 50370 3390
rect 19742 3330 19794 3342
rect 19742 3266 19794 3278
rect 48862 3330 48914 3342
rect 48862 3266 48914 3278
rect 1344 3162 58576 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 50558 3162
rect 50610 3110 50662 3162
rect 50714 3110 50766 3162
rect 50818 3110 58576 3162
rect 1344 3076 58576 3110
<< via1 >>
rect 24222 56702 24274 56754
rect 24894 56702 24946 56754
rect 38334 56702 38386 56754
rect 40238 56702 40290 56754
rect 50430 56702 50482 56754
rect 51214 56702 51266 56754
rect 23998 56590 24050 56642
rect 25118 56590 25170 56642
rect 19838 56422 19890 56474
rect 19942 56422 19994 56474
rect 20046 56422 20098 56474
rect 50558 56422 50610 56474
rect 50662 56422 50714 56474
rect 50766 56422 50818 56474
rect 23438 56254 23490 56306
rect 24894 56254 24946 56306
rect 33182 56254 33234 56306
rect 41022 56254 41074 56306
rect 43038 56254 43090 56306
rect 49758 56254 49810 56306
rect 51214 56254 51266 56306
rect 23662 56142 23714 56194
rect 23998 56142 24050 56194
rect 24558 56142 24610 56194
rect 31278 56142 31330 56194
rect 35086 56142 35138 56194
rect 38894 56142 38946 56194
rect 40686 56142 40738 56194
rect 41358 56142 41410 56194
rect 43710 56142 43762 56194
rect 49982 56142 50034 56194
rect 50318 56142 50370 56194
rect 51550 56142 51602 56194
rect 27806 56030 27858 56082
rect 30606 56030 30658 56082
rect 31502 56030 31554 56082
rect 32174 56030 32226 56082
rect 35422 56030 35474 56082
rect 38558 56030 38610 56082
rect 39230 56030 39282 56082
rect 40238 56030 40290 56082
rect 41582 56030 41634 56082
rect 42590 56030 42642 56082
rect 25566 55918 25618 55970
rect 28590 55918 28642 55970
rect 36206 55918 36258 55970
rect 39790 55918 39842 55970
rect 42142 55918 42194 55970
rect 4478 55638 4530 55690
rect 4582 55638 4634 55690
rect 4686 55638 4738 55690
rect 35198 55638 35250 55690
rect 35302 55638 35354 55690
rect 35406 55638 35458 55690
rect 24670 55470 24722 55522
rect 24222 55358 24274 55410
rect 28142 55358 28194 55410
rect 28590 55358 28642 55410
rect 30270 55358 30322 55410
rect 31278 55358 31330 55410
rect 33518 55358 33570 55410
rect 37214 55358 37266 55410
rect 42030 55358 42082 55410
rect 50990 55358 51042 55410
rect 27022 55246 27074 55298
rect 27470 55246 27522 55298
rect 29150 55246 29202 55298
rect 29710 55246 29762 55298
rect 30494 55246 30546 55298
rect 32510 55246 32562 55298
rect 35646 55246 35698 55298
rect 39454 55246 39506 55298
rect 39902 55246 39954 55298
rect 40126 55246 40178 55298
rect 41022 55246 41074 55298
rect 42478 55246 42530 55298
rect 35422 55134 35474 55186
rect 36430 55134 36482 55186
rect 41582 55134 41634 55186
rect 27694 55022 27746 55074
rect 30830 55022 30882 55074
rect 31726 55022 31778 55074
rect 32174 55022 32226 55074
rect 35982 55022 36034 55074
rect 40462 55022 40514 55074
rect 40798 55022 40850 55074
rect 19838 54854 19890 54906
rect 19942 54854 19994 54906
rect 20046 54854 20098 54906
rect 50558 54854 50610 54906
rect 50662 54854 50714 54906
rect 50766 54854 50818 54906
rect 26238 54686 26290 54738
rect 26462 54686 26514 54738
rect 28926 54686 28978 54738
rect 29822 54686 29874 54738
rect 34190 54686 34242 54738
rect 28478 54574 28530 54626
rect 29150 54574 29202 54626
rect 29486 54574 29538 54626
rect 30158 54574 30210 54626
rect 32398 54574 32450 54626
rect 36094 54574 36146 54626
rect 37550 54574 37602 54626
rect 38782 54574 38834 54626
rect 39902 54574 39954 54626
rect 41022 54574 41074 54626
rect 32286 54462 32338 54514
rect 32622 54462 32674 54514
rect 33182 54462 33234 54514
rect 36318 54462 36370 54514
rect 40126 54462 40178 54514
rect 26910 54350 26962 54402
rect 27470 54350 27522 54402
rect 27918 54350 27970 54402
rect 31838 54350 31890 54402
rect 37214 54350 37266 54402
rect 39230 54238 39282 54290
rect 4478 54070 4530 54122
rect 4582 54070 4634 54122
rect 4686 54070 4738 54122
rect 35198 54070 35250 54122
rect 35302 54070 35354 54122
rect 35406 54070 35458 54122
rect 22654 53790 22706 53842
rect 25230 53790 25282 53842
rect 33518 53790 33570 53842
rect 35870 53790 35922 53842
rect 37214 53790 37266 53842
rect 13470 53678 13522 53730
rect 13694 53678 13746 53730
rect 21982 53678 22034 53730
rect 22318 53678 22370 53730
rect 25006 53678 25058 53730
rect 30270 53678 30322 53730
rect 30718 53678 30770 53730
rect 32846 53678 32898 53730
rect 34638 53678 34690 53730
rect 35758 53678 35810 53730
rect 38782 53678 38834 53730
rect 39902 53678 39954 53730
rect 40238 53678 40290 53730
rect 14254 53566 14306 53618
rect 21310 53566 21362 53618
rect 21534 53566 21586 53618
rect 23886 53566 23938 53618
rect 24110 53566 24162 53618
rect 24446 53566 24498 53618
rect 25902 53566 25954 53618
rect 31166 53566 31218 53618
rect 32398 53566 32450 53618
rect 33294 53566 33346 53618
rect 35086 53566 35138 53618
rect 37662 53566 37714 53618
rect 39566 53566 39618 53618
rect 42590 53566 42642 53618
rect 43374 53566 43426 53618
rect 44830 53566 44882 53618
rect 47854 53566 47906 53618
rect 21758 53454 21810 53506
rect 22542 53454 22594 53506
rect 23662 53454 23714 53506
rect 24334 53454 24386 53506
rect 29934 53454 29986 53506
rect 39118 53454 39170 53506
rect 40014 53454 40066 53506
rect 42366 53454 42418 53506
rect 42702 53454 42754 53506
rect 42926 53454 42978 53506
rect 43038 53454 43090 53506
rect 43262 53454 43314 53506
rect 44942 53454 44994 53506
rect 45166 53454 45218 53506
rect 19838 53286 19890 53338
rect 19942 53286 19994 53338
rect 20046 53286 20098 53338
rect 50558 53286 50610 53338
rect 50662 53286 50714 53338
rect 50766 53286 50818 53338
rect 13918 53118 13970 53170
rect 24782 53118 24834 53170
rect 29150 53118 29202 53170
rect 30046 53118 30098 53170
rect 39342 53118 39394 53170
rect 41022 53118 41074 53170
rect 12574 53006 12626 53058
rect 15598 53006 15650 53058
rect 16158 53006 16210 53058
rect 18062 53006 18114 53058
rect 21534 53006 21586 53058
rect 22430 53006 22482 53058
rect 24558 53006 24610 53058
rect 26462 53006 26514 53058
rect 31614 53006 31666 53058
rect 31838 53006 31890 53058
rect 33406 53006 33458 53058
rect 35422 53006 35474 53058
rect 36990 53006 37042 53058
rect 37102 53006 37154 53058
rect 38782 53006 38834 53058
rect 41134 53006 41186 53058
rect 41358 53006 41410 53058
rect 44270 53006 44322 53058
rect 45726 53006 45778 53058
rect 49086 53006 49138 53058
rect 10446 52894 10498 52946
rect 12798 52894 12850 52946
rect 13470 52894 13522 52946
rect 15486 52894 15538 52946
rect 17390 52894 17442 52946
rect 17950 52894 18002 52946
rect 19630 52894 19682 52946
rect 20638 52894 20690 52946
rect 23662 52894 23714 52946
rect 24446 52894 24498 52946
rect 25678 52894 25730 52946
rect 26238 52894 26290 52946
rect 31390 52894 31442 52946
rect 32062 52894 32114 52946
rect 33854 52894 33906 52946
rect 35310 52894 35362 52946
rect 36766 52894 36818 52946
rect 37886 52894 37938 52946
rect 40126 52894 40178 52946
rect 40910 52894 40962 52946
rect 42702 52894 42754 52946
rect 42926 52894 42978 52946
rect 43374 52894 43426 52946
rect 44494 52894 44546 52946
rect 46958 52894 47010 52946
rect 48862 52894 48914 52946
rect 49198 52894 49250 52946
rect 10334 52782 10386 52834
rect 11118 52782 11170 52834
rect 14926 52782 14978 52834
rect 18398 52782 18450 52834
rect 19182 52782 19234 52834
rect 20078 52782 20130 52834
rect 20750 52782 20802 52834
rect 22094 52782 22146 52834
rect 24110 52782 24162 52834
rect 25342 52782 25394 52834
rect 26350 52782 26402 52834
rect 29710 52782 29762 52834
rect 30606 52782 30658 52834
rect 35982 52782 36034 52834
rect 38446 52782 38498 52834
rect 39678 52782 39730 52834
rect 42030 52782 42082 52834
rect 43598 52782 43650 52834
rect 45166 52782 45218 52834
rect 47630 52782 47682 52834
rect 49646 52782 49698 52834
rect 15598 52670 15650 52722
rect 32398 52670 32450 52722
rect 37550 52670 37602 52722
rect 39006 52670 39058 52722
rect 43934 52670 43986 52722
rect 4478 52502 4530 52554
rect 4582 52502 4634 52554
rect 4686 52502 4738 52554
rect 35198 52502 35250 52554
rect 35302 52502 35354 52554
rect 35406 52502 35458 52554
rect 11006 52334 11058 52386
rect 24670 52334 24722 52386
rect 37998 52334 38050 52386
rect 10334 52222 10386 52274
rect 14590 52222 14642 52274
rect 16606 52222 16658 52274
rect 17278 52222 17330 52274
rect 26238 52222 26290 52274
rect 27134 52222 27186 52274
rect 31502 52222 31554 52274
rect 38782 52222 38834 52274
rect 43598 52222 43650 52274
rect 45390 52222 45442 52274
rect 50878 52222 50930 52274
rect 7646 52110 7698 52162
rect 7982 52110 8034 52162
rect 10446 52110 10498 52162
rect 11790 52110 11842 52162
rect 12350 52110 12402 52162
rect 14142 52110 14194 52162
rect 15150 52110 15202 52162
rect 15710 52110 15762 52162
rect 18622 52110 18674 52162
rect 19742 52110 19794 52162
rect 20190 52110 20242 52162
rect 21310 52110 21362 52162
rect 21870 52110 21922 52162
rect 22878 52110 22930 52162
rect 23102 52110 23154 52162
rect 23326 52110 23378 52162
rect 24222 52110 24274 52162
rect 24446 52110 24498 52162
rect 26014 52110 26066 52162
rect 27358 52110 27410 52162
rect 29822 52110 29874 52162
rect 29934 52110 29986 52162
rect 30046 52110 30098 52162
rect 30270 52110 30322 52162
rect 30942 52110 30994 52162
rect 33518 52110 33570 52162
rect 33966 52110 34018 52162
rect 35534 52110 35586 52162
rect 36094 52110 36146 52162
rect 36990 52110 37042 52162
rect 37214 52110 37266 52162
rect 37550 52110 37602 52162
rect 38334 52110 38386 52162
rect 38670 52110 38722 52162
rect 40014 52110 40066 52162
rect 41134 52110 41186 52162
rect 42478 52110 42530 52162
rect 42590 52110 42642 52162
rect 42814 52110 42866 52162
rect 43262 52110 43314 52162
rect 45726 52110 45778 52162
rect 46958 52110 47010 52162
rect 48078 52110 48130 52162
rect 48414 52110 48466 52162
rect 48862 52110 48914 52162
rect 49310 52110 49362 52162
rect 50206 52110 50258 52162
rect 8094 51998 8146 52050
rect 12238 51998 12290 52050
rect 12462 51998 12514 52050
rect 14590 51998 14642 52050
rect 17614 51998 17666 52050
rect 19294 51998 19346 52050
rect 19630 51998 19682 52050
rect 21982 51998 22034 52050
rect 26686 51998 26738 52050
rect 27022 51998 27074 52050
rect 32622 51998 32674 52050
rect 36318 51998 36370 52050
rect 36430 51998 36482 52050
rect 37438 51998 37490 52050
rect 39566 51998 39618 52050
rect 41806 51998 41858 52050
rect 47630 51998 47682 52050
rect 48190 51998 48242 52050
rect 48638 51998 48690 52050
rect 21534 51886 21586 51938
rect 30718 51886 30770 51938
rect 32734 51886 32786 51938
rect 38446 51886 38498 51938
rect 38782 51886 38834 51938
rect 50430 51886 50482 51938
rect 19838 51718 19890 51770
rect 19942 51718 19994 51770
rect 20046 51718 20098 51770
rect 50558 51718 50610 51770
rect 50662 51718 50714 51770
rect 50766 51718 50818 51770
rect 10446 51550 10498 51602
rect 10894 51550 10946 51602
rect 11118 51550 11170 51602
rect 16718 51550 16770 51602
rect 20638 51550 20690 51602
rect 21198 51550 21250 51602
rect 21646 51550 21698 51602
rect 21870 51550 21922 51602
rect 31054 51550 31106 51602
rect 34638 51550 34690 51602
rect 35646 51550 35698 51602
rect 36094 51550 36146 51602
rect 36766 51550 36818 51602
rect 39118 51550 39170 51602
rect 39454 51550 39506 51602
rect 42926 51550 42978 51602
rect 51550 51550 51602 51602
rect 8318 51438 8370 51490
rect 10222 51438 10274 51490
rect 13246 51438 13298 51490
rect 20526 51438 20578 51490
rect 20862 51438 20914 51490
rect 22542 51438 22594 51490
rect 24446 51438 24498 51490
rect 24558 51438 24610 51490
rect 24782 51438 24834 51490
rect 25566 51438 25618 51490
rect 25678 51438 25730 51490
rect 26350 51438 26402 51490
rect 27582 51438 27634 51490
rect 30382 51438 30434 51490
rect 30494 51438 30546 51490
rect 31614 51438 31666 51490
rect 32510 51438 32562 51490
rect 33070 51438 33122 51490
rect 33406 51438 33458 51490
rect 35534 51438 35586 51490
rect 37102 51438 37154 51490
rect 37438 51438 37490 51490
rect 42702 51438 42754 51490
rect 43710 51438 43762 51490
rect 45502 51438 45554 51490
rect 45614 51438 45666 51490
rect 46958 51438 47010 51490
rect 51886 51438 51938 51490
rect 6974 51326 7026 51378
rect 7758 51326 7810 51378
rect 10110 51326 10162 51378
rect 10782 51326 10834 51378
rect 11790 51326 11842 51378
rect 12014 51326 12066 51378
rect 13582 51326 13634 51378
rect 14478 51326 14530 51378
rect 16158 51326 16210 51378
rect 16382 51326 16434 51378
rect 17950 51326 18002 51378
rect 18958 51326 19010 51378
rect 19966 51326 20018 51378
rect 20302 51326 20354 51378
rect 21534 51326 21586 51378
rect 22206 51326 22258 51378
rect 27358 51326 27410 51378
rect 29934 51326 29986 51378
rect 30718 51326 30770 51378
rect 32286 51326 32338 51378
rect 34190 51326 34242 51378
rect 34414 51326 34466 51378
rect 34862 51326 34914 51378
rect 35086 51326 35138 51378
rect 35758 51326 35810 51378
rect 36318 51326 36370 51378
rect 37774 51326 37826 51378
rect 38782 51326 38834 51378
rect 40910 51326 40962 51378
rect 41358 51326 41410 51378
rect 41806 51326 41858 51378
rect 42478 51326 42530 51378
rect 43038 51326 43090 51378
rect 43486 51326 43538 51378
rect 44158 51326 44210 51378
rect 44718 51326 44770 51378
rect 45390 51326 45442 51378
rect 46286 51326 46338 51378
rect 46510 51326 46562 51378
rect 46622 51326 46674 51378
rect 47854 51326 47906 51378
rect 48750 51326 48802 51378
rect 49086 51326 49138 51378
rect 50766 51326 50818 51378
rect 50990 51326 51042 51378
rect 51326 51326 51378 51378
rect 1822 51214 1874 51266
rect 7982 51214 8034 51266
rect 12350 51214 12402 51266
rect 17502 51214 17554 51266
rect 22318 51214 22370 51266
rect 26014 51214 26066 51266
rect 34526 51214 34578 51266
rect 38558 51214 38610 51266
rect 41134 51214 41186 51266
rect 42814 51214 42866 51266
rect 47294 51214 47346 51266
rect 48974 51214 49026 51266
rect 49534 51214 49586 51266
rect 51102 51214 51154 51266
rect 12462 51102 12514 51154
rect 15822 51102 15874 51154
rect 19182 51102 19234 51154
rect 25566 51102 25618 51154
rect 29710 51102 29762 51154
rect 38222 51102 38274 51154
rect 38334 51102 38386 51154
rect 44158 51102 44210 51154
rect 46062 51102 46114 51154
rect 49758 51102 49810 51154
rect 49982 51102 50034 51154
rect 50430 51102 50482 51154
rect 4478 50934 4530 50986
rect 4582 50934 4634 50986
rect 4686 50934 4738 50986
rect 35198 50934 35250 50986
rect 35302 50934 35354 50986
rect 35406 50934 35458 50986
rect 8430 50766 8482 50818
rect 12462 50766 12514 50818
rect 17502 50766 17554 50818
rect 22542 50766 22594 50818
rect 38670 50766 38722 50818
rect 7086 50654 7138 50706
rect 8766 50654 8818 50706
rect 14254 50654 14306 50706
rect 17390 50654 17442 50706
rect 24334 50654 24386 50706
rect 27470 50654 27522 50706
rect 32622 50654 32674 50706
rect 37774 50654 37826 50706
rect 39454 50654 39506 50706
rect 41918 50654 41970 50706
rect 47854 50654 47906 50706
rect 48638 50654 48690 50706
rect 50094 50654 50146 50706
rect 6862 50542 6914 50594
rect 7198 50542 7250 50594
rect 8206 50542 8258 50594
rect 9214 50542 9266 50594
rect 11790 50542 11842 50594
rect 12014 50542 12066 50594
rect 13694 50542 13746 50594
rect 15262 50542 15314 50594
rect 16830 50542 16882 50594
rect 18174 50542 18226 50594
rect 20078 50542 20130 50594
rect 20414 50542 20466 50594
rect 22654 50542 22706 50594
rect 24222 50542 24274 50594
rect 25678 50542 25730 50594
rect 26686 50542 26738 50594
rect 27022 50542 27074 50594
rect 30494 50542 30546 50594
rect 31054 50542 31106 50594
rect 33182 50542 33234 50594
rect 34414 50542 34466 50594
rect 35086 50542 35138 50594
rect 36542 50542 36594 50594
rect 37326 50542 37378 50594
rect 38782 50542 38834 50594
rect 40350 50542 40402 50594
rect 41246 50542 41298 50594
rect 43150 50542 43202 50594
rect 43598 50542 43650 50594
rect 43934 50542 43986 50594
rect 44942 50542 44994 50594
rect 47630 50542 47682 50594
rect 48750 50542 48802 50594
rect 49534 50542 49586 50594
rect 51662 50542 51714 50594
rect 51886 50542 51938 50594
rect 1710 50430 1762 50482
rect 2942 50430 2994 50482
rect 3950 50430 4002 50482
rect 5966 50430 6018 50482
rect 7758 50430 7810 50482
rect 18398 50430 18450 50482
rect 18510 50430 18562 50482
rect 21870 50430 21922 50482
rect 21982 50430 22034 50482
rect 22542 50430 22594 50482
rect 24894 50430 24946 50482
rect 25790 50430 25842 50482
rect 27582 50430 27634 50482
rect 32958 50430 33010 50482
rect 33854 50430 33906 50482
rect 35422 50430 35474 50482
rect 36206 50430 36258 50482
rect 36318 50430 36370 50482
rect 37550 50430 37602 50482
rect 43822 50430 43874 50482
rect 45166 50430 45218 50482
rect 45614 50430 45666 50482
rect 52670 50430 52722 50482
rect 52782 50430 52834 50482
rect 53230 50430 53282 50482
rect 2046 50318 2098 50370
rect 2494 50318 2546 50370
rect 3614 50318 3666 50370
rect 5630 50318 5682 50370
rect 20190 50318 20242 50370
rect 21646 50318 21698 50370
rect 26014 50318 26066 50370
rect 42926 50318 42978 50370
rect 51438 50318 51490 50370
rect 51774 50318 51826 50370
rect 53006 50318 53058 50370
rect 53342 50318 53394 50370
rect 19838 50150 19890 50202
rect 19942 50150 19994 50202
rect 20046 50150 20098 50202
rect 50558 50150 50610 50202
rect 50662 50150 50714 50202
rect 50766 50150 50818 50202
rect 15710 49982 15762 50034
rect 20862 49982 20914 50034
rect 41806 49982 41858 50034
rect 42254 49982 42306 50034
rect 42590 49982 42642 50034
rect 44942 49982 44994 50034
rect 47406 49982 47458 50034
rect 53902 49982 53954 50034
rect 7422 49870 7474 49922
rect 11342 49870 11394 49922
rect 13582 49870 13634 49922
rect 14142 49870 14194 49922
rect 20190 49870 20242 49922
rect 21646 49870 21698 49922
rect 25790 49870 25842 49922
rect 26910 49870 26962 49922
rect 33406 49870 33458 49922
rect 37662 49870 37714 49922
rect 38894 49870 38946 49922
rect 47742 49870 47794 49922
rect 49534 49870 49586 49922
rect 53678 49870 53730 49922
rect 8430 49758 8482 49810
rect 11454 49758 11506 49810
rect 12350 49758 12402 49810
rect 13918 49758 13970 49810
rect 15374 49758 15426 49810
rect 19182 49758 19234 49810
rect 19854 49758 19906 49810
rect 20526 49758 20578 49810
rect 22990 49758 23042 49810
rect 27246 49758 27298 49810
rect 27918 49758 27970 49810
rect 29822 49758 29874 49810
rect 30158 49758 30210 49810
rect 30382 49758 30434 49810
rect 30606 49758 30658 49810
rect 32286 49758 32338 49810
rect 32510 49758 32562 49810
rect 34974 49758 35026 49810
rect 36318 49758 36370 49810
rect 36878 49758 36930 49810
rect 37550 49758 37602 49810
rect 38222 49758 38274 49810
rect 39118 49758 39170 49810
rect 41470 49758 41522 49810
rect 43038 49758 43090 49810
rect 43262 49758 43314 49810
rect 44158 49758 44210 49810
rect 44718 49758 44770 49810
rect 46622 49758 46674 49810
rect 46734 49758 46786 49810
rect 46958 49758 47010 49810
rect 50430 49758 50482 49810
rect 51774 49758 51826 49810
rect 52110 49758 52162 49810
rect 52334 49758 52386 49810
rect 52782 49758 52834 49810
rect 53006 49758 53058 49810
rect 2046 49646 2098 49698
rect 2494 49646 2546 49698
rect 2830 49646 2882 49698
rect 3390 49646 3442 49698
rect 3726 49646 3778 49698
rect 4174 49646 4226 49698
rect 4622 49646 4674 49698
rect 6862 49646 6914 49698
rect 8990 49646 9042 49698
rect 12910 49646 12962 49698
rect 14590 49646 14642 49698
rect 19630 49646 19682 49698
rect 21422 49646 21474 49698
rect 23550 49646 23602 49698
rect 25902 49646 25954 49698
rect 26014 49646 26066 49698
rect 28590 49646 28642 49698
rect 29374 49646 29426 49698
rect 33182 49646 33234 49698
rect 35758 49646 35810 49698
rect 39230 49646 39282 49698
rect 44046 49646 44098 49698
rect 48974 49646 49026 49698
rect 51998 49646 52050 49698
rect 53902 49646 53954 49698
rect 2046 49534 2098 49586
rect 2382 49534 2434 49586
rect 31054 49534 31106 49586
rect 31838 49534 31890 49586
rect 36654 49534 36706 49586
rect 47070 49534 47122 49586
rect 51214 49534 51266 49586
rect 53342 49534 53394 49586
rect 4478 49366 4530 49418
rect 4582 49366 4634 49418
rect 4686 49366 4738 49418
rect 35198 49366 35250 49418
rect 35302 49366 35354 49418
rect 35406 49366 35458 49418
rect 7310 49198 7362 49250
rect 19966 49198 20018 49250
rect 27582 49198 27634 49250
rect 34750 49198 34802 49250
rect 49534 49198 49586 49250
rect 53118 49198 53170 49250
rect 6974 49086 7026 49138
rect 7758 49086 7810 49138
rect 15486 49086 15538 49138
rect 16158 49086 16210 49138
rect 21870 49086 21922 49138
rect 24222 49086 24274 49138
rect 32734 49086 32786 49138
rect 32846 49086 32898 49138
rect 34302 49086 34354 49138
rect 34526 49086 34578 49138
rect 49086 49086 49138 49138
rect 52782 49086 52834 49138
rect 53790 49086 53842 49138
rect 2382 48974 2434 49026
rect 2942 48974 2994 49026
rect 3278 48974 3330 49026
rect 3950 48974 4002 49026
rect 4846 48974 4898 49026
rect 5182 48974 5234 49026
rect 6190 48974 6242 49026
rect 6526 48974 6578 49026
rect 6750 48974 6802 49026
rect 9214 48974 9266 49026
rect 11230 48974 11282 49026
rect 13470 48974 13522 49026
rect 13694 48974 13746 49026
rect 14030 48974 14082 49026
rect 15150 48974 15202 49026
rect 16382 48974 16434 49026
rect 18510 48974 18562 49026
rect 19294 48974 19346 49026
rect 20190 48974 20242 49026
rect 21982 48974 22034 49026
rect 22430 48974 22482 49026
rect 22654 48974 22706 49026
rect 22878 48974 22930 49026
rect 23326 48974 23378 49026
rect 23550 48974 23602 49026
rect 24110 48974 24162 49026
rect 26798 48974 26850 49026
rect 27022 48974 27074 49026
rect 28030 48974 28082 49026
rect 28254 48974 28306 49026
rect 28590 48974 28642 49026
rect 29822 48974 29874 49026
rect 31054 48974 31106 49026
rect 31502 48974 31554 49026
rect 32510 48974 32562 49026
rect 33854 48974 33906 49026
rect 35198 48974 35250 49026
rect 35534 48974 35586 49026
rect 36094 48974 36146 49026
rect 36990 48974 37042 49026
rect 37214 48974 37266 49026
rect 37662 48974 37714 49026
rect 38334 48974 38386 49026
rect 39566 48974 39618 49026
rect 40686 48974 40738 49026
rect 46734 48974 46786 49026
rect 47294 48974 47346 49026
rect 49422 48974 49474 49026
rect 50990 48974 51042 49026
rect 51550 48974 51602 49026
rect 3838 48862 3890 48914
rect 5854 48862 5906 48914
rect 6302 48862 6354 48914
rect 8206 48862 8258 48914
rect 11566 48862 11618 48914
rect 14702 48862 14754 48914
rect 17054 48862 17106 48914
rect 18846 48862 18898 48914
rect 19406 48862 19458 48914
rect 19518 48862 19570 48914
rect 20750 48862 20802 48914
rect 22542 48862 22594 48914
rect 24222 48862 24274 48914
rect 28478 48862 28530 48914
rect 30606 48862 30658 48914
rect 31166 48862 31218 48914
rect 31726 48862 31778 48914
rect 33182 48862 33234 48914
rect 33406 48862 33458 48914
rect 35646 48862 35698 48914
rect 35982 48862 36034 48914
rect 37998 48862 38050 48914
rect 39118 48862 39170 48914
rect 41358 48862 41410 48914
rect 46846 48862 46898 48914
rect 50542 48862 50594 48914
rect 52894 48862 52946 48914
rect 1710 48750 1762 48802
rect 2046 48750 2098 48802
rect 2718 48750 2770 48802
rect 3166 48750 3218 48802
rect 3614 48750 3666 48802
rect 4510 48750 4562 48802
rect 4958 48750 5010 48802
rect 5518 48750 5570 48802
rect 5742 48750 5794 48802
rect 10558 48750 10610 48802
rect 11454 48750 11506 48802
rect 20526 48750 20578 48802
rect 20862 48750 20914 48802
rect 21534 48750 21586 48802
rect 21758 48750 21810 48802
rect 30158 48750 30210 48802
rect 32062 48750 32114 48802
rect 33630 48750 33682 48802
rect 36542 48750 36594 48802
rect 37326 48750 37378 48802
rect 37438 48750 37490 48802
rect 47070 48750 47122 48802
rect 49534 48750 49586 48802
rect 51438 48750 51490 48802
rect 53678 48750 53730 48802
rect 19838 48582 19890 48634
rect 19942 48582 19994 48634
rect 20046 48582 20098 48634
rect 50558 48582 50610 48634
rect 50662 48582 50714 48634
rect 50766 48582 50818 48634
rect 16718 48414 16770 48466
rect 18734 48414 18786 48466
rect 19854 48414 19906 48466
rect 20974 48414 21026 48466
rect 21198 48414 21250 48466
rect 22654 48414 22706 48466
rect 30830 48414 30882 48466
rect 32622 48414 32674 48466
rect 35758 48414 35810 48466
rect 40238 48414 40290 48466
rect 43710 48414 43762 48466
rect 46062 48414 46114 48466
rect 50654 48414 50706 48466
rect 53118 48414 53170 48466
rect 53342 48414 53394 48466
rect 2158 48302 2210 48354
rect 2606 48302 2658 48354
rect 2718 48302 2770 48354
rect 9886 48302 9938 48354
rect 10334 48302 10386 48354
rect 11678 48302 11730 48354
rect 15038 48302 15090 48354
rect 21982 48302 22034 48354
rect 22318 48302 22370 48354
rect 25678 48302 25730 48354
rect 25790 48302 25842 48354
rect 26798 48302 26850 48354
rect 29710 48302 29762 48354
rect 31166 48302 31218 48354
rect 32286 48302 32338 48354
rect 32398 48302 32450 48354
rect 34190 48302 34242 48354
rect 36094 48302 36146 48354
rect 37774 48302 37826 48354
rect 38782 48302 38834 48354
rect 40126 48302 40178 48354
rect 41694 48302 41746 48354
rect 44494 48302 44546 48354
rect 46174 48302 46226 48354
rect 50878 48302 50930 48354
rect 50990 48302 51042 48354
rect 1934 48190 1986 48242
rect 3502 48190 3554 48242
rect 3950 48190 4002 48242
rect 4510 48190 4562 48242
rect 5070 48190 5122 48242
rect 6414 48190 6466 48242
rect 7534 48190 7586 48242
rect 7758 48190 7810 48242
rect 9774 48190 9826 48242
rect 12798 48190 12850 48242
rect 16158 48190 16210 48242
rect 18510 48190 18562 48242
rect 19294 48190 19346 48242
rect 19630 48190 19682 48242
rect 21310 48190 21362 48242
rect 21758 48190 21810 48242
rect 26238 48190 26290 48242
rect 26462 48190 26514 48242
rect 30046 48190 30098 48242
rect 33518 48190 33570 48242
rect 33742 48190 33794 48242
rect 34414 48190 34466 48242
rect 34638 48190 34690 48242
rect 34862 48190 34914 48242
rect 35086 48190 35138 48242
rect 36654 48190 36706 48242
rect 37102 48190 37154 48242
rect 38894 48190 38946 48242
rect 42030 48190 42082 48242
rect 43262 48190 43314 48242
rect 46846 48190 46898 48242
rect 47070 48190 47122 48242
rect 53678 48190 53730 48242
rect 4062 48078 4114 48130
rect 5966 48078 6018 48130
rect 8318 48078 8370 48130
rect 11006 48078 11058 48130
rect 11454 48078 11506 48130
rect 14702 48078 14754 48130
rect 26350 48078 26402 48130
rect 29822 48078 29874 48130
rect 33070 48078 33122 48130
rect 37326 48078 37378 48130
rect 44270 48078 44322 48130
rect 47742 48078 47794 48130
rect 53230 48078 53282 48130
rect 2606 47966 2658 48018
rect 14142 47966 14194 48018
rect 19518 47966 19570 48018
rect 25790 47966 25842 48018
rect 33294 47966 33346 48018
rect 4478 47798 4530 47850
rect 4582 47798 4634 47850
rect 4686 47798 4738 47850
rect 35198 47798 35250 47850
rect 35302 47798 35354 47850
rect 35406 47798 35458 47850
rect 3502 47630 3554 47682
rect 3838 47630 3890 47682
rect 4286 47630 4338 47682
rect 4622 47630 4674 47682
rect 5630 47630 5682 47682
rect 5966 47630 6018 47682
rect 32846 47630 32898 47682
rect 3726 47518 3778 47570
rect 7982 47518 8034 47570
rect 8318 47518 8370 47570
rect 11790 47518 11842 47570
rect 14590 47518 14642 47570
rect 17726 47518 17778 47570
rect 21758 47518 21810 47570
rect 23998 47518 24050 47570
rect 31390 47518 31442 47570
rect 33406 47518 33458 47570
rect 41918 47518 41970 47570
rect 47518 47518 47570 47570
rect 51214 47518 51266 47570
rect 1710 47406 1762 47458
rect 2494 47406 2546 47458
rect 2718 47406 2770 47458
rect 4062 47406 4114 47458
rect 5070 47406 5122 47458
rect 7646 47406 7698 47458
rect 9774 47406 9826 47458
rect 11006 47406 11058 47458
rect 12350 47406 12402 47458
rect 13806 47406 13858 47458
rect 14142 47406 14194 47458
rect 15934 47406 15986 47458
rect 16606 47406 16658 47458
rect 17278 47406 17330 47458
rect 17950 47406 18002 47458
rect 19630 47406 19682 47458
rect 19742 47406 19794 47458
rect 21198 47406 21250 47458
rect 21646 47406 21698 47458
rect 22766 47406 22818 47458
rect 24222 47406 24274 47458
rect 26014 47406 26066 47458
rect 27022 47406 27074 47458
rect 27358 47406 27410 47458
rect 30382 47406 30434 47458
rect 31054 47406 31106 47458
rect 32062 47406 32114 47458
rect 33182 47406 33234 47458
rect 33518 47406 33570 47458
rect 34974 47406 35026 47458
rect 35422 47406 35474 47458
rect 36318 47406 36370 47458
rect 38110 47406 38162 47458
rect 38334 47406 38386 47458
rect 39230 47406 39282 47458
rect 42142 47406 42194 47458
rect 43150 47406 43202 47458
rect 44158 47406 44210 47458
rect 49310 47406 49362 47458
rect 51102 47406 51154 47458
rect 53118 47406 53170 47458
rect 54126 47406 54178 47458
rect 54462 47406 54514 47458
rect 5854 47294 5906 47346
rect 6302 47294 6354 47346
rect 6638 47294 6690 47346
rect 9550 47294 9602 47346
rect 9662 47294 9714 47346
rect 10782 47294 10834 47346
rect 14702 47294 14754 47346
rect 15598 47294 15650 47346
rect 18622 47294 18674 47346
rect 19854 47294 19906 47346
rect 20302 47294 20354 47346
rect 24782 47294 24834 47346
rect 25566 47294 25618 47346
rect 30494 47294 30546 47346
rect 31278 47294 31330 47346
rect 35870 47294 35922 47346
rect 39006 47294 39058 47346
rect 39454 47294 39506 47346
rect 39566 47294 39618 47346
rect 42814 47294 42866 47346
rect 43822 47294 43874 47346
rect 48078 47294 48130 47346
rect 49982 47294 50034 47346
rect 51662 47294 51714 47346
rect 52894 47294 52946 47346
rect 2046 47182 2098 47234
rect 3054 47182 3106 47234
rect 3278 47182 3330 47234
rect 3390 47182 3442 47234
rect 10222 47182 10274 47234
rect 21870 47182 21922 47234
rect 22318 47182 22370 47234
rect 23102 47182 23154 47234
rect 23326 47182 23378 47234
rect 23438 47182 23490 47234
rect 30718 47182 30770 47234
rect 33294 47182 33346 47234
rect 41134 47182 41186 47234
rect 41470 47182 41522 47234
rect 43486 47182 43538 47234
rect 43934 47182 43986 47234
rect 19838 47014 19890 47066
rect 19942 47014 19994 47066
rect 20046 47014 20098 47066
rect 50558 47014 50610 47066
rect 50662 47014 50714 47066
rect 50766 47014 50818 47066
rect 3838 46846 3890 46898
rect 10894 46846 10946 46898
rect 12910 46846 12962 46898
rect 16046 46846 16098 46898
rect 18062 46846 18114 46898
rect 22430 46846 22482 46898
rect 25790 46846 25842 46898
rect 26014 46846 26066 46898
rect 26574 46846 26626 46898
rect 43150 46846 43202 46898
rect 45614 46846 45666 46898
rect 46062 46846 46114 46898
rect 47966 46846 48018 46898
rect 49086 46846 49138 46898
rect 51438 46846 51490 46898
rect 4846 46734 4898 46786
rect 5518 46734 5570 46786
rect 6750 46734 6802 46786
rect 10334 46734 10386 46786
rect 10558 46734 10610 46786
rect 13806 46734 13858 46786
rect 16270 46734 16322 46786
rect 16382 46734 16434 46786
rect 19406 46734 19458 46786
rect 19630 46734 19682 46786
rect 20302 46734 20354 46786
rect 20750 46734 20802 46786
rect 21870 46734 21922 46786
rect 22766 46734 22818 46786
rect 24222 46734 24274 46786
rect 27358 46734 27410 46786
rect 29710 46734 29762 46786
rect 30942 46734 30994 46786
rect 40014 46734 40066 46786
rect 40126 46734 40178 46786
rect 41246 46734 41298 46786
rect 42030 46734 42082 46786
rect 44158 46734 44210 46786
rect 46398 46734 46450 46786
rect 47854 46734 47906 46786
rect 48190 46734 48242 46786
rect 48974 46734 49026 46786
rect 50430 46734 50482 46786
rect 51326 46734 51378 46786
rect 54126 46734 54178 46786
rect 54238 46734 54290 46786
rect 2382 46622 2434 46674
rect 3054 46622 3106 46674
rect 3390 46622 3442 46674
rect 3726 46622 3778 46674
rect 3950 46622 4002 46674
rect 4622 46622 4674 46674
rect 6862 46622 6914 46674
rect 7982 46622 8034 46674
rect 10110 46622 10162 46674
rect 12014 46622 12066 46674
rect 12126 46622 12178 46674
rect 13358 46622 13410 46674
rect 13470 46622 13522 46674
rect 17726 46622 17778 46674
rect 20078 46622 20130 46674
rect 20526 46622 20578 46674
rect 20862 46622 20914 46674
rect 21646 46622 21698 46674
rect 22206 46622 22258 46674
rect 22542 46622 22594 46674
rect 23438 46622 23490 46674
rect 23774 46622 23826 46674
rect 25566 46622 25618 46674
rect 26126 46622 26178 46674
rect 26350 46622 26402 46674
rect 26910 46622 26962 46674
rect 29598 46622 29650 46674
rect 33070 46622 33122 46674
rect 33294 46622 33346 46674
rect 34862 46622 34914 46674
rect 36542 46622 36594 46674
rect 36990 46622 37042 46674
rect 40350 46622 40402 46674
rect 41022 46622 41074 46674
rect 41470 46622 41522 46674
rect 41806 46622 41858 46674
rect 42702 46622 42754 46674
rect 42926 46622 42978 46674
rect 45278 46622 45330 46674
rect 52670 46622 52722 46674
rect 53006 46622 53058 46674
rect 53790 46622 53842 46674
rect 2606 46510 2658 46562
rect 5854 46510 5906 46562
rect 11902 46510 11954 46562
rect 13694 46510 13746 46562
rect 19854 46510 19906 46562
rect 23662 46510 23714 46562
rect 31838 46510 31890 46562
rect 34974 46510 35026 46562
rect 37550 46510 37602 46562
rect 41918 46510 41970 46562
rect 43710 46510 43762 46562
rect 50878 46510 50930 46562
rect 53118 46510 53170 46562
rect 53454 46510 53506 46562
rect 53566 46510 53618 46562
rect 8990 46398 9042 46450
rect 39566 46398 39618 46450
rect 43262 46398 43314 46450
rect 51438 46398 51490 46450
rect 54238 46398 54290 46450
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 22654 46062 22706 46114
rect 31950 46062 32002 46114
rect 32286 46062 32338 46114
rect 33518 46062 33570 46114
rect 52782 46062 52834 46114
rect 3054 45950 3106 46002
rect 4174 45950 4226 46002
rect 15710 45950 15762 46002
rect 22094 45950 22146 46002
rect 23102 45950 23154 46002
rect 27134 45950 27186 46002
rect 29262 45950 29314 46002
rect 31390 45950 31442 46002
rect 31726 45950 31778 46002
rect 32734 45950 32786 46002
rect 48974 45950 49026 46002
rect 54126 45950 54178 46002
rect 54798 45950 54850 46002
rect 1822 45838 1874 45890
rect 3166 45838 3218 45890
rect 4510 45838 4562 45890
rect 4958 45838 5010 45890
rect 6302 45838 6354 45890
rect 7646 45838 7698 45890
rect 8430 45838 8482 45890
rect 11118 45838 11170 45890
rect 12910 45838 12962 45890
rect 13806 45838 13858 45890
rect 13918 45838 13970 45890
rect 14142 45838 14194 45890
rect 22318 45838 22370 45890
rect 24558 45838 24610 45890
rect 26014 45838 26066 45890
rect 27694 45838 27746 45890
rect 30942 45838 30994 45890
rect 33182 45838 33234 45890
rect 33518 45838 33570 45890
rect 34414 45838 34466 45890
rect 35310 45838 35362 45890
rect 35870 45838 35922 45890
rect 36094 45838 36146 45890
rect 38558 45838 38610 45890
rect 38782 45838 38834 45890
rect 40910 45838 40962 45890
rect 41358 45838 41410 45890
rect 41470 45838 41522 45890
rect 41918 45838 41970 45890
rect 42142 45838 42194 45890
rect 43486 45838 43538 45890
rect 43822 45838 43874 45890
rect 45054 45838 45106 45890
rect 45390 45838 45442 45890
rect 47406 45838 47458 45890
rect 47630 45838 47682 45890
rect 48750 45838 48802 45890
rect 49646 45838 49698 45890
rect 51774 45838 51826 45890
rect 54350 45838 54402 45890
rect 2158 45726 2210 45778
rect 5630 45726 5682 45778
rect 6414 45726 6466 45778
rect 6638 45726 6690 45778
rect 7198 45726 7250 45778
rect 11902 45726 11954 45778
rect 14254 45726 14306 45778
rect 16158 45726 16210 45778
rect 17614 45726 17666 45778
rect 17838 45726 17890 45778
rect 18734 45726 18786 45778
rect 21422 45726 21474 45778
rect 21758 45726 21810 45778
rect 23550 45726 23602 45778
rect 29710 45726 29762 45778
rect 35534 45726 35586 45778
rect 36430 45726 36482 45778
rect 39790 45726 39842 45778
rect 40798 45726 40850 45778
rect 43598 45726 43650 45778
rect 44830 45726 44882 45778
rect 46174 45726 46226 45778
rect 47518 45726 47570 45778
rect 48862 45726 48914 45778
rect 50990 45726 51042 45778
rect 51550 45726 51602 45778
rect 52670 45726 52722 45778
rect 52782 45726 52834 45778
rect 5966 45614 6018 45666
rect 9774 45614 9826 45666
rect 12798 45614 12850 45666
rect 19070 45614 19122 45666
rect 25118 45614 25170 45666
rect 26350 45614 26402 45666
rect 27022 45614 27074 45666
rect 27246 45614 27298 45666
rect 34638 45614 34690 45666
rect 37102 45614 37154 45666
rect 37438 45614 37490 45666
rect 40238 45614 40290 45666
rect 40686 45614 40738 45666
rect 41694 45614 41746 45666
rect 43038 45614 43090 45666
rect 45054 45614 45106 45666
rect 45838 45614 45890 45666
rect 46958 45614 47010 45666
rect 51326 45614 51378 45666
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 50558 45446 50610 45498
rect 50662 45446 50714 45498
rect 50766 45446 50818 45498
rect 2830 45278 2882 45330
rect 4846 45278 4898 45330
rect 9774 45278 9826 45330
rect 16382 45278 16434 45330
rect 19518 45278 19570 45330
rect 20078 45278 20130 45330
rect 23662 45278 23714 45330
rect 26350 45278 26402 45330
rect 26910 45278 26962 45330
rect 27806 45278 27858 45330
rect 32174 45278 32226 45330
rect 38894 45278 38946 45330
rect 45838 45278 45890 45330
rect 47966 45278 48018 45330
rect 48190 45278 48242 45330
rect 48302 45278 48354 45330
rect 52558 45278 52610 45330
rect 54798 45278 54850 45330
rect 2046 45166 2098 45218
rect 3950 45166 4002 45218
rect 10782 45166 10834 45218
rect 12574 45166 12626 45218
rect 15598 45166 15650 45218
rect 16606 45166 16658 45218
rect 16718 45166 16770 45218
rect 17726 45166 17778 45218
rect 20414 45166 20466 45218
rect 26574 45166 26626 45218
rect 27582 45166 27634 45218
rect 32062 45166 32114 45218
rect 34750 45166 34802 45218
rect 36206 45166 36258 45218
rect 38222 45166 38274 45218
rect 39118 45166 39170 45218
rect 45166 45166 45218 45218
rect 47742 45166 47794 45218
rect 51662 45166 51714 45218
rect 1822 45054 1874 45106
rect 2942 45054 2994 45106
rect 3166 45054 3218 45106
rect 3390 45054 3442 45106
rect 4062 45054 4114 45106
rect 4734 45054 4786 45106
rect 5294 45054 5346 45106
rect 5518 45054 5570 45106
rect 7198 45054 7250 45106
rect 8542 45054 8594 45106
rect 11006 45054 11058 45106
rect 11342 45054 11394 45106
rect 13582 45054 13634 45106
rect 15934 45054 15986 45106
rect 18958 45054 19010 45106
rect 19966 45054 20018 45106
rect 20190 45054 20242 45106
rect 23102 45054 23154 45106
rect 23326 45054 23378 45106
rect 26238 45054 26290 45106
rect 26798 45054 26850 45106
rect 27134 45054 27186 45106
rect 27470 45054 27522 45106
rect 33742 45054 33794 45106
rect 34862 45054 34914 45106
rect 37438 45054 37490 45106
rect 41694 45054 41746 45106
rect 43710 45054 43762 45106
rect 43934 45054 43986 45106
rect 44494 45054 44546 45106
rect 44942 45054 44994 45106
rect 49198 45054 49250 45106
rect 49982 45054 50034 45106
rect 51550 45054 51602 45106
rect 52446 45054 52498 45106
rect 53006 45054 53058 45106
rect 53454 45054 53506 45106
rect 53790 45054 53842 45106
rect 54238 45054 54290 45106
rect 54574 45054 54626 45106
rect 3054 44942 3106 44994
rect 7646 44942 7698 44994
rect 8990 44942 9042 44994
rect 9662 44942 9714 44994
rect 10782 44942 10834 44994
rect 12126 44942 12178 44994
rect 17502 44942 17554 44994
rect 33182 44942 33234 44994
rect 33518 44942 33570 44994
rect 34526 44942 34578 44994
rect 35758 44942 35810 44994
rect 42254 44942 42306 44994
rect 43822 44942 43874 44994
rect 45054 44942 45106 44994
rect 46286 44942 46338 44994
rect 49086 44942 49138 44994
rect 54686 44942 54738 44994
rect 9998 44830 10050 44882
rect 14926 44830 14978 44882
rect 15822 44830 15874 44882
rect 32174 44830 32226 44882
rect 38782 44830 38834 44882
rect 44046 44830 44098 44882
rect 50094 44830 50146 44882
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 4846 44494 4898 44546
rect 5630 44494 5682 44546
rect 9998 44494 10050 44546
rect 17390 44494 17442 44546
rect 21534 44494 21586 44546
rect 35758 44494 35810 44546
rect 36206 44494 36258 44546
rect 46734 44494 46786 44546
rect 2382 44382 2434 44434
rect 4286 44382 4338 44434
rect 7646 44382 7698 44434
rect 8878 44382 8930 44434
rect 12014 44382 12066 44434
rect 14366 44382 14418 44434
rect 17502 44382 17554 44434
rect 23550 44382 23602 44434
rect 34974 44382 35026 44434
rect 35422 44382 35474 44434
rect 40462 44382 40514 44434
rect 44158 44382 44210 44434
rect 45054 44382 45106 44434
rect 47070 44382 47122 44434
rect 47518 44382 47570 44434
rect 2606 44270 2658 44322
rect 2942 44270 2994 44322
rect 4622 44270 4674 44322
rect 6862 44270 6914 44322
rect 8430 44270 8482 44322
rect 9550 44270 9602 44322
rect 10894 44270 10946 44322
rect 11790 44270 11842 44322
rect 12350 44270 12402 44322
rect 13806 44270 13858 44322
rect 15822 44270 15874 44322
rect 16830 44270 16882 44322
rect 19406 44270 19458 44322
rect 19630 44270 19682 44322
rect 19854 44270 19906 44322
rect 19966 44270 20018 44322
rect 21310 44270 21362 44322
rect 21758 44270 21810 44322
rect 21870 44270 21922 44322
rect 23102 44270 23154 44322
rect 23886 44270 23938 44322
rect 25790 44270 25842 44322
rect 26798 44270 26850 44322
rect 27694 44270 27746 44322
rect 33406 44270 33458 44322
rect 36318 44270 36370 44322
rect 37326 44270 37378 44322
rect 38670 44270 38722 44322
rect 42142 44270 42194 44322
rect 43710 44270 43762 44322
rect 45166 44270 45218 44322
rect 45502 44270 45554 44322
rect 50654 44270 50706 44322
rect 51662 44270 51714 44322
rect 51774 44270 51826 44322
rect 54798 44270 54850 44322
rect 55694 44270 55746 44322
rect 2718 44158 2770 44210
rect 6302 44158 6354 44210
rect 7198 44158 7250 44210
rect 9326 44158 9378 44210
rect 9438 44158 9490 44210
rect 23774 44158 23826 44210
rect 26014 44158 26066 44210
rect 28254 44158 28306 44210
rect 32398 44158 32450 44210
rect 34414 44158 34466 44210
rect 35534 44158 35586 44210
rect 36206 44158 36258 44210
rect 36990 44158 37042 44210
rect 38446 44158 38498 44210
rect 39790 44158 39842 44210
rect 40798 44158 40850 44210
rect 42926 44158 42978 44210
rect 44270 44158 44322 44210
rect 46958 44158 47010 44210
rect 47966 44158 48018 44210
rect 49422 44158 49474 44210
rect 49646 44158 49698 44210
rect 50766 44158 50818 44210
rect 51886 44158 51938 44210
rect 53902 44158 53954 44210
rect 55806 44158 55858 44210
rect 1710 44046 1762 44098
rect 2046 44046 2098 44098
rect 3390 44046 3442 44098
rect 5742 44046 5794 44098
rect 5854 44046 5906 44098
rect 6638 44046 6690 44098
rect 7086 44046 7138 44098
rect 26574 44046 26626 44098
rect 37102 44046 37154 44098
rect 39678 44046 39730 44098
rect 46062 44046 46114 44098
rect 50990 44046 51042 44098
rect 51214 44046 51266 44098
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 50558 43878 50610 43930
rect 50662 43878 50714 43930
rect 50766 43878 50818 43930
rect 3726 43710 3778 43762
rect 9550 43710 9602 43762
rect 10782 43710 10834 43762
rect 14030 43710 14082 43762
rect 14814 43710 14866 43762
rect 20526 43710 20578 43762
rect 27918 43710 27970 43762
rect 41694 43710 41746 43762
rect 55246 43710 55298 43762
rect 4622 43598 4674 43650
rect 6078 43598 6130 43650
rect 7534 43598 7586 43650
rect 12574 43598 12626 43650
rect 15598 43598 15650 43650
rect 16606 43598 16658 43650
rect 20078 43598 20130 43650
rect 21646 43598 21698 43650
rect 23886 43598 23938 43650
rect 25342 43598 25394 43650
rect 27246 43598 27298 43650
rect 27470 43598 27522 43650
rect 28814 43598 28866 43650
rect 32174 43598 32226 43650
rect 32286 43598 32338 43650
rect 33070 43598 33122 43650
rect 33406 43598 33458 43650
rect 34078 43598 34130 43650
rect 37326 43598 37378 43650
rect 41134 43598 41186 43650
rect 41470 43598 41522 43650
rect 42590 43598 42642 43650
rect 46734 43598 46786 43650
rect 51326 43598 51378 43650
rect 55022 43598 55074 43650
rect 2718 43486 2770 43538
rect 3502 43486 3554 43538
rect 4062 43486 4114 43538
rect 5070 43486 5122 43538
rect 6862 43486 6914 43538
rect 10110 43486 10162 43538
rect 13470 43486 13522 43538
rect 14590 43486 14642 43538
rect 15710 43486 15762 43538
rect 17950 43486 18002 43538
rect 20414 43486 20466 43538
rect 20750 43486 20802 43538
rect 22542 43486 22594 43538
rect 25230 43486 25282 43538
rect 25566 43486 25618 43538
rect 27134 43486 27186 43538
rect 27582 43486 27634 43538
rect 28030 43486 28082 43538
rect 28254 43486 28306 43538
rect 31390 43486 31442 43538
rect 31614 43486 31666 43538
rect 31950 43486 32002 43538
rect 36206 43486 36258 43538
rect 43934 43486 43986 43538
rect 52446 43486 52498 43538
rect 54126 43486 54178 43538
rect 54350 43486 54402 43538
rect 2942 43374 2994 43426
rect 5518 43374 5570 43426
rect 5854 43374 5906 43426
rect 5966 43374 6018 43426
rect 6750 43374 6802 43426
rect 8094 43374 8146 43426
rect 11342 43374 11394 43426
rect 12126 43374 12178 43426
rect 16270 43374 16322 43426
rect 17726 43374 17778 43426
rect 18622 43374 18674 43426
rect 19182 43374 19234 43426
rect 19406 43374 19458 43426
rect 19742 43374 19794 43426
rect 21086 43374 21138 43426
rect 26238 43374 26290 43426
rect 28926 43374 28978 43426
rect 30718 43374 30770 43426
rect 36430 43374 36482 43426
rect 36878 43374 36930 43426
rect 41806 43374 41858 43426
rect 42254 43374 42306 43426
rect 47294 43374 47346 43426
rect 50878 43374 50930 43426
rect 53230 43374 53282 43426
rect 3054 43262 3106 43314
rect 26350 43262 26402 43314
rect 28590 43262 28642 43314
rect 39678 43262 39730 43314
rect 39790 43262 39842 43314
rect 40014 43262 40066 43314
rect 40126 43262 40178 43314
rect 40910 43262 40962 43314
rect 41134 43262 41186 43314
rect 45054 43262 45106 43314
rect 48862 43262 48914 43314
rect 48974 43262 49026 43314
rect 49198 43262 49250 43314
rect 49310 43262 49362 43314
rect 54686 43262 54738 43314
rect 55358 43262 55410 43314
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 19406 42926 19458 42978
rect 43598 42926 43650 42978
rect 46510 42926 46562 42978
rect 54350 42926 54402 42978
rect 1934 42814 1986 42866
rect 5854 42814 5906 42866
rect 12350 42814 12402 42866
rect 15710 42814 15762 42866
rect 19294 42814 19346 42866
rect 23774 42814 23826 42866
rect 26798 42814 26850 42866
rect 27246 42814 27298 42866
rect 32174 42814 32226 42866
rect 33742 42814 33794 42866
rect 34526 42814 34578 42866
rect 39006 42814 39058 42866
rect 40574 42814 40626 42866
rect 46174 42814 46226 42866
rect 48190 42814 48242 42866
rect 51214 42814 51266 42866
rect 57150 42814 57202 42866
rect 4286 42702 4338 42754
rect 4622 42702 4674 42754
rect 7310 42702 7362 42754
rect 9550 42702 9602 42754
rect 11790 42702 11842 42754
rect 11902 42702 11954 42754
rect 13806 42702 13858 42754
rect 14030 42702 14082 42754
rect 14254 42702 14306 42754
rect 20862 42702 20914 42754
rect 21870 42702 21922 42754
rect 25342 42702 25394 42754
rect 26238 42702 26290 42754
rect 26910 42702 26962 42754
rect 27470 42702 27522 42754
rect 32398 42702 32450 42754
rect 33518 42702 33570 42754
rect 35086 42702 35138 42754
rect 36094 42702 36146 42754
rect 37102 42702 37154 42754
rect 37886 42702 37938 42754
rect 38894 42702 38946 42754
rect 39790 42702 39842 42754
rect 41358 42702 41410 42754
rect 42366 42702 42418 42754
rect 42702 42702 42754 42754
rect 44942 42702 44994 42754
rect 45390 42702 45442 42754
rect 46398 42702 46450 42754
rect 46846 42702 46898 42754
rect 49870 42702 49922 42754
rect 51438 42702 51490 42754
rect 51886 42702 51938 42754
rect 54126 42702 54178 42754
rect 55246 42702 55298 42754
rect 55694 42702 55746 42754
rect 56702 42702 56754 42754
rect 6302 42590 6354 42642
rect 8542 42590 8594 42642
rect 9326 42590 9378 42642
rect 16270 42590 16322 42642
rect 17614 42590 17666 42642
rect 17838 42590 17890 42642
rect 19182 42590 19234 42642
rect 20526 42590 20578 42642
rect 20638 42590 20690 42642
rect 21310 42590 21362 42642
rect 22094 42590 22146 42642
rect 22206 42590 22258 42642
rect 24222 42590 24274 42642
rect 27806 42590 27858 42642
rect 30494 42590 30546 42642
rect 30606 42590 30658 42642
rect 35758 42590 35810 42642
rect 36990 42590 37042 42642
rect 37774 42590 37826 42642
rect 38334 42590 38386 42642
rect 48974 42590 49026 42642
rect 50318 42590 50370 42642
rect 50654 42590 50706 42642
rect 52670 42590 52722 42642
rect 4958 42478 5010 42530
rect 9774 42478 9826 42530
rect 9886 42478 9938 42530
rect 10110 42478 10162 42530
rect 10446 42478 10498 42530
rect 12686 42478 12738 42530
rect 14590 42478 14642 42530
rect 21646 42478 21698 42530
rect 22654 42478 22706 42530
rect 25790 42478 25842 42530
rect 26686 42478 26738 42530
rect 30830 42478 30882 42530
rect 35982 42478 36034 42530
rect 37550 42478 37602 42530
rect 49870 42478 49922 42530
rect 50430 42478 50482 42530
rect 51662 42478 51714 42530
rect 52782 42478 52834 42530
rect 53006 42478 53058 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 50558 42310 50610 42362
rect 50662 42310 50714 42362
rect 50766 42310 50818 42362
rect 5294 42142 5346 42194
rect 8654 42142 8706 42194
rect 10558 42142 10610 42194
rect 13358 42142 13410 42194
rect 16382 42142 16434 42194
rect 16606 42142 16658 42194
rect 22878 42142 22930 42194
rect 27134 42142 27186 42194
rect 32174 42142 32226 42194
rect 33854 42142 33906 42194
rect 36094 42142 36146 42194
rect 36990 42142 37042 42194
rect 40126 42142 40178 42194
rect 43598 42142 43650 42194
rect 2046 42030 2098 42082
rect 2494 42030 2546 42082
rect 2606 42030 2658 42082
rect 6638 42030 6690 42082
rect 8318 42030 8370 42082
rect 9886 42030 9938 42082
rect 11566 42030 11618 42082
rect 16718 42030 16770 42082
rect 18062 42030 18114 42082
rect 31614 42030 31666 42082
rect 34862 42030 34914 42082
rect 36206 42030 36258 42082
rect 37774 42030 37826 42082
rect 39230 42030 39282 42082
rect 40910 42030 40962 42082
rect 41022 42030 41074 42082
rect 42142 42030 42194 42082
rect 43374 42030 43426 42082
rect 47406 42030 47458 42082
rect 49086 42030 49138 42082
rect 54350 42030 54402 42082
rect 1710 41918 1762 41970
rect 3614 41918 3666 41970
rect 3950 41918 4002 41970
rect 4846 41918 4898 41970
rect 5406 41918 5458 41970
rect 5518 41918 5570 41970
rect 6862 41918 6914 41970
rect 7646 41918 7698 41970
rect 8878 41918 8930 41970
rect 9998 41918 10050 41970
rect 10670 41918 10722 41970
rect 12126 41918 12178 41970
rect 12798 41918 12850 41970
rect 13806 41918 13858 41970
rect 14030 41918 14082 41970
rect 14254 41918 14306 41970
rect 15374 41918 15426 41970
rect 18958 41918 19010 41970
rect 22094 41918 22146 41970
rect 22206 41918 22258 41970
rect 22542 41918 22594 41970
rect 23102 41918 23154 41970
rect 23326 41918 23378 41970
rect 23998 41918 24050 41970
rect 24670 41918 24722 41970
rect 25790 41918 25842 41970
rect 26350 41918 26402 41970
rect 28254 41918 28306 41970
rect 29262 41918 29314 41970
rect 31838 41918 31890 41970
rect 36766 41918 36818 41970
rect 37886 41918 37938 41970
rect 38558 41918 38610 41970
rect 38894 41918 38946 41970
rect 39566 41918 39618 41970
rect 40238 41918 40290 41970
rect 44046 41918 44098 41970
rect 44942 41918 44994 41970
rect 45390 41918 45442 41970
rect 47630 41918 47682 41970
rect 48862 41918 48914 41970
rect 49646 41918 49698 41970
rect 51438 41918 51490 41970
rect 52446 41918 52498 41970
rect 54238 41918 54290 41970
rect 4622 41806 4674 41858
rect 15486 41806 15538 41858
rect 17502 41806 17554 41858
rect 19630 41806 19682 41858
rect 22430 41806 22482 41858
rect 23886 41806 23938 41858
rect 25678 41806 25730 41858
rect 29150 41806 29202 41858
rect 33294 41806 33346 41858
rect 34302 41806 34354 41858
rect 41694 41806 41746 41858
rect 46174 41806 46226 41858
rect 47406 41806 47458 41858
rect 49534 41806 49586 41858
rect 52894 41806 52946 41858
rect 54910 41806 54962 41858
rect 2494 41694 2546 41746
rect 15598 41694 15650 41746
rect 23214 41694 23266 41746
rect 27582 41694 27634 41746
rect 38894 41694 38946 41746
rect 41022 41694 41074 41746
rect 50430 41694 50482 41746
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 8318 41358 8370 41410
rect 8878 41358 8930 41410
rect 14142 41358 14194 41410
rect 23662 41358 23714 41410
rect 44046 41358 44098 41410
rect 1934 41246 1986 41298
rect 7198 41246 7250 41298
rect 8094 41246 8146 41298
rect 12350 41246 12402 41298
rect 16718 41246 16770 41298
rect 20078 41246 20130 41298
rect 21534 41246 21586 41298
rect 26014 41246 26066 41298
rect 32174 41246 32226 41298
rect 33406 41246 33458 41298
rect 34078 41246 34130 41298
rect 35870 41246 35922 41298
rect 36318 41246 36370 41298
rect 4286 41134 4338 41186
rect 4734 41134 4786 41186
rect 5854 41134 5906 41186
rect 6190 41134 6242 41186
rect 7422 41134 7474 41186
rect 9326 41134 9378 41186
rect 9550 41134 9602 41186
rect 9662 41134 9714 41186
rect 10110 41134 10162 41186
rect 10894 41134 10946 41186
rect 11566 41134 11618 41186
rect 11790 41134 11842 41186
rect 14254 41134 14306 41186
rect 14590 41134 14642 41186
rect 15934 41134 15986 41186
rect 17614 41134 17666 41186
rect 17950 41134 18002 41186
rect 18510 41134 18562 41186
rect 18734 41134 18786 41186
rect 19630 41134 19682 41186
rect 21758 41134 21810 41186
rect 22542 41134 22594 41186
rect 22766 41134 22818 41186
rect 23438 41134 23490 41186
rect 31950 41134 32002 41186
rect 32286 41134 32338 41186
rect 33294 41134 33346 41186
rect 34750 41134 34802 41186
rect 35422 41134 35474 41186
rect 36542 41134 36594 41186
rect 38110 41134 38162 41186
rect 39230 41134 39282 41186
rect 41470 41134 41522 41186
rect 42590 41134 42642 41186
rect 44942 41134 44994 41186
rect 45390 41134 45442 41186
rect 47518 41134 47570 41186
rect 48638 41134 48690 41186
rect 50430 41134 50482 41186
rect 51214 41134 51266 41186
rect 51662 41134 51714 41186
rect 54238 41134 54290 41186
rect 55246 41134 55298 41186
rect 6750 41022 6802 41074
rect 8542 41022 8594 41074
rect 11678 41022 11730 41074
rect 12238 41022 12290 41074
rect 12462 41022 12514 41074
rect 13918 41022 13970 41074
rect 16494 41022 16546 41074
rect 18846 41022 18898 41074
rect 19294 41022 19346 41074
rect 19966 41022 20018 41074
rect 25118 41022 25170 41074
rect 25566 41022 25618 41074
rect 25678 41022 25730 41074
rect 25902 41022 25954 41074
rect 26238 41022 26290 41074
rect 26462 41022 26514 41074
rect 26798 41022 26850 41074
rect 26910 41022 26962 41074
rect 29486 41022 29538 41074
rect 31166 41022 31218 41074
rect 34638 41022 34690 41074
rect 37326 41022 37378 41074
rect 39342 41022 39394 41074
rect 41022 41022 41074 41074
rect 43486 41022 43538 41074
rect 44158 41022 44210 41074
rect 44830 41022 44882 41074
rect 47406 41022 47458 41074
rect 53118 41022 53170 41074
rect 55470 41022 55522 41074
rect 4958 40910 5010 40962
rect 5742 40910 5794 40962
rect 8990 40910 9042 40962
rect 18174 40910 18226 40962
rect 18286 40910 18338 40962
rect 20190 40910 20242 40962
rect 22094 40910 22146 40962
rect 25342 40910 25394 40962
rect 27134 40910 27186 40962
rect 29150 40910 29202 40962
rect 30830 40910 30882 40962
rect 31838 40910 31890 40962
rect 32510 40910 32562 40962
rect 34414 40910 34466 40962
rect 44046 40910 44098 40962
rect 48750 40910 48802 40962
rect 51998 40910 52050 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 50558 40742 50610 40794
rect 50662 40742 50714 40794
rect 50766 40742 50818 40794
rect 5182 40574 5234 40626
rect 6078 40574 6130 40626
rect 6862 40574 6914 40626
rect 7198 40574 7250 40626
rect 7422 40574 7474 40626
rect 8542 40574 8594 40626
rect 11118 40574 11170 40626
rect 19518 40574 19570 40626
rect 20526 40574 20578 40626
rect 21870 40574 21922 40626
rect 25902 40574 25954 40626
rect 33406 40574 33458 40626
rect 35310 40574 35362 40626
rect 35422 40574 35474 40626
rect 40910 40574 40962 40626
rect 47630 40574 47682 40626
rect 50654 40574 50706 40626
rect 5854 40462 5906 40514
rect 6302 40462 6354 40514
rect 9102 40462 9154 40514
rect 12014 40462 12066 40514
rect 14590 40462 14642 40514
rect 18622 40462 18674 40514
rect 19070 40462 19122 40514
rect 19294 40462 19346 40514
rect 20414 40462 20466 40514
rect 22654 40462 22706 40514
rect 25678 40462 25730 40514
rect 27134 40462 27186 40514
rect 30382 40462 30434 40514
rect 33854 40462 33906 40514
rect 35646 40462 35698 40514
rect 35870 40462 35922 40514
rect 42478 40462 42530 40514
rect 43038 40462 43090 40514
rect 44046 40462 44098 40514
rect 49198 40462 49250 40514
rect 50766 40462 50818 40514
rect 4286 40350 4338 40402
rect 5518 40350 5570 40402
rect 6414 40350 6466 40402
rect 6638 40350 6690 40402
rect 6974 40350 7026 40402
rect 7534 40350 7586 40402
rect 8318 40350 8370 40402
rect 10558 40350 10610 40402
rect 12350 40350 12402 40402
rect 13246 40350 13298 40402
rect 15598 40350 15650 40402
rect 16158 40350 16210 40402
rect 18510 40350 18562 40402
rect 18846 40350 18898 40402
rect 19742 40350 19794 40402
rect 19854 40350 19906 40402
rect 20190 40350 20242 40402
rect 21310 40350 21362 40402
rect 22878 40350 22930 40402
rect 23774 40350 23826 40402
rect 24446 40350 24498 40402
rect 25566 40350 25618 40402
rect 26014 40350 26066 40402
rect 26350 40350 26402 40402
rect 29598 40350 29650 40402
rect 33294 40350 33346 40402
rect 34078 40350 34130 40402
rect 35534 40350 35586 40402
rect 37214 40350 37266 40402
rect 38334 40350 38386 40402
rect 38894 40350 38946 40402
rect 41470 40350 41522 40402
rect 43262 40350 43314 40402
rect 43374 40350 43426 40402
rect 43598 40350 43650 40402
rect 45390 40350 45442 40402
rect 46958 40350 47010 40402
rect 48190 40350 48242 40402
rect 51550 40350 51602 40402
rect 51774 40350 51826 40402
rect 53230 40350 53282 40402
rect 54014 40350 54066 40402
rect 54238 40350 54290 40402
rect 54686 40350 54738 40402
rect 4622 40238 4674 40290
rect 4846 40238 4898 40290
rect 16270 40238 16322 40290
rect 29262 40238 29314 40290
rect 32510 40238 32562 40290
rect 34414 40238 34466 40290
rect 36318 40238 36370 40290
rect 38558 40238 38610 40290
rect 39678 40238 39730 40290
rect 45166 40238 45218 40290
rect 46286 40238 46338 40290
rect 47182 40238 47234 40290
rect 48974 40238 49026 40290
rect 51326 40238 51378 40290
rect 53342 40238 53394 40290
rect 53678 40238 53730 40290
rect 1934 40126 1986 40178
rect 21534 40126 21586 40178
rect 33406 40126 33458 40178
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 2942 39790 2994 39842
rect 4286 39790 4338 39842
rect 4622 39790 4674 39842
rect 19518 39790 19570 39842
rect 24110 39790 24162 39842
rect 29822 39790 29874 39842
rect 30158 39790 30210 39842
rect 31614 39790 31666 39842
rect 31950 39790 32002 39842
rect 37662 39790 37714 39842
rect 39790 39790 39842 39842
rect 40126 39790 40178 39842
rect 48302 39790 48354 39842
rect 2830 39678 2882 39730
rect 11118 39678 11170 39730
rect 13694 39678 13746 39730
rect 15486 39678 15538 39730
rect 28702 39678 28754 39730
rect 35870 39678 35922 39730
rect 38222 39678 38274 39730
rect 40574 39678 40626 39730
rect 44046 39678 44098 39730
rect 49086 39678 49138 39730
rect 51102 39678 51154 39730
rect 55134 39678 55186 39730
rect 1822 39566 1874 39618
rect 3054 39566 3106 39618
rect 3838 39566 3890 39618
rect 4062 39566 4114 39618
rect 6638 39566 6690 39618
rect 7422 39566 7474 39618
rect 8766 39566 8818 39618
rect 9102 39566 9154 39618
rect 10110 39566 10162 39618
rect 10894 39566 10946 39618
rect 11342 39566 11394 39618
rect 11454 39566 11506 39618
rect 16830 39566 16882 39618
rect 17502 39566 17554 39618
rect 18958 39566 19010 39618
rect 19182 39566 19234 39618
rect 23998 39566 24050 39618
rect 25006 39566 25058 39618
rect 27022 39566 27074 39618
rect 30830 39566 30882 39618
rect 32734 39566 32786 39618
rect 33854 39566 33906 39618
rect 34190 39566 34242 39618
rect 35534 39566 35586 39618
rect 37774 39566 37826 39618
rect 39454 39566 39506 39618
rect 40910 39566 40962 39618
rect 42142 39566 42194 39618
rect 42814 39566 42866 39618
rect 43598 39566 43650 39618
rect 45950 39566 46002 39618
rect 46622 39566 46674 39618
rect 47854 39566 47906 39618
rect 48078 39566 48130 39618
rect 48862 39566 48914 39618
rect 49310 39566 49362 39618
rect 49422 39566 49474 39618
rect 49982 39566 50034 39618
rect 50206 39566 50258 39618
rect 51550 39566 51602 39618
rect 52222 39566 52274 39618
rect 52670 39566 52722 39618
rect 54126 39566 54178 39618
rect 54574 39566 54626 39618
rect 55358 39566 55410 39618
rect 6414 39454 6466 39506
rect 8094 39454 8146 39506
rect 8542 39454 8594 39506
rect 15822 39454 15874 39506
rect 17838 39454 17890 39506
rect 18174 39454 18226 39506
rect 19854 39454 19906 39506
rect 20190 39454 20242 39506
rect 21646 39454 21698 39506
rect 25566 39454 25618 39506
rect 25790 39454 25842 39506
rect 27134 39454 27186 39506
rect 30942 39454 30994 39506
rect 32510 39454 32562 39506
rect 36430 39454 36482 39506
rect 37102 39454 37154 39506
rect 37214 39454 37266 39506
rect 39902 39454 39954 39506
rect 43710 39454 43762 39506
rect 46846 39454 46898 39506
rect 51886 39454 51938 39506
rect 51998 39454 52050 39506
rect 53006 39454 53058 39506
rect 54798 39454 54850 39506
rect 2046 39342 2098 39394
rect 5182 39342 5234 39394
rect 8990 39342 9042 39394
rect 9438 39342 9490 39394
rect 10446 39342 10498 39394
rect 10558 39342 10610 39394
rect 10670 39342 10722 39394
rect 14926 39342 14978 39394
rect 21310 39342 21362 39394
rect 23774 39342 23826 39394
rect 24110 39342 24162 39394
rect 25230 39342 25282 39394
rect 29486 39342 29538 39394
rect 33294 39342 33346 39394
rect 34414 39342 34466 39394
rect 34526 39342 34578 39394
rect 36878 39342 36930 39394
rect 37662 39342 37714 39394
rect 39118 39342 39170 39394
rect 42702 39342 42754 39394
rect 45390 39342 45442 39394
rect 48750 39342 48802 39394
rect 50542 39342 50594 39394
rect 55694 39342 55746 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 50558 39174 50610 39226
rect 50662 39174 50714 39226
rect 50766 39174 50818 39226
rect 4174 39006 4226 39058
rect 12126 39006 12178 39058
rect 16046 39006 16098 39058
rect 16270 39006 16322 39058
rect 16942 39006 16994 39058
rect 17390 39006 17442 39058
rect 26014 39006 26066 39058
rect 31166 39006 31218 39058
rect 45614 39006 45666 39058
rect 45838 39006 45890 39058
rect 48862 39006 48914 39058
rect 49086 39006 49138 39058
rect 52446 39006 52498 39058
rect 52782 39006 52834 39058
rect 53566 39006 53618 39058
rect 4734 38894 4786 38946
rect 6302 38894 6354 38946
rect 8318 38894 8370 38946
rect 11230 38894 11282 38946
rect 15934 38894 15986 38946
rect 16382 38894 16434 38946
rect 17726 38894 17778 38946
rect 18062 38894 18114 38946
rect 18174 38894 18226 38946
rect 23998 38894 24050 38946
rect 24222 38894 24274 38946
rect 24334 38894 24386 38946
rect 25342 38894 25394 38946
rect 33294 38894 33346 38946
rect 37102 38894 37154 38946
rect 41918 38894 41970 38946
rect 44494 38894 44546 38946
rect 45502 38894 45554 38946
rect 47742 38894 47794 38946
rect 49646 38894 49698 38946
rect 50878 38894 50930 38946
rect 51102 38894 51154 38946
rect 53118 38894 53170 38946
rect 54462 38894 54514 38946
rect 2606 38782 2658 38834
rect 3838 38782 3890 38834
rect 4622 38782 4674 38834
rect 7310 38782 7362 38834
rect 10446 38782 10498 38834
rect 10670 38782 10722 38834
rect 13806 38782 13858 38834
rect 15374 38782 15426 38834
rect 19406 38782 19458 38834
rect 19966 38782 20018 38834
rect 20414 38782 20466 38834
rect 20638 38782 20690 38834
rect 21534 38782 21586 38834
rect 22430 38782 22482 38834
rect 24558 38782 24610 38834
rect 33518 38782 33570 38834
rect 36878 38782 36930 38834
rect 37662 38782 37714 38834
rect 38558 38782 38610 38834
rect 41246 38782 41298 38834
rect 41806 38782 41858 38834
rect 43598 38782 43650 38834
rect 44382 38782 44434 38834
rect 46286 38782 46338 38834
rect 46398 38782 46450 38834
rect 46846 38782 46898 38834
rect 48750 38782 48802 38834
rect 49310 38782 49362 38834
rect 51326 38782 51378 38834
rect 53454 38782 53506 38834
rect 53790 38782 53842 38834
rect 54798 38782 54850 38834
rect 55470 38782 55522 38834
rect 2494 38670 2546 38722
rect 3054 38670 3106 38722
rect 5406 38670 5458 38722
rect 5742 38670 5794 38722
rect 14030 38670 14082 38722
rect 19182 38670 19234 38722
rect 20974 38670 21026 38722
rect 21310 38670 21362 38722
rect 22206 38670 22258 38722
rect 34078 38670 34130 38722
rect 35982 38670 36034 38722
rect 36542 38670 36594 38722
rect 37774 38670 37826 38722
rect 42590 38670 42642 38722
rect 47966 38670 48018 38722
rect 49870 38670 49922 38722
rect 50206 38670 50258 38722
rect 51886 38670 51938 38722
rect 54686 38670 54738 38722
rect 4510 38558 4562 38610
rect 14254 38558 14306 38610
rect 14366 38558 14418 38610
rect 15038 38558 15090 38610
rect 15374 38558 15426 38610
rect 18174 38558 18226 38610
rect 21870 38558 21922 38610
rect 22766 38558 22818 38610
rect 47630 38558 47682 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 2718 38222 2770 38274
rect 6526 38222 6578 38274
rect 25118 38222 25170 38274
rect 25902 38222 25954 38274
rect 41694 38222 41746 38274
rect 43710 38222 43762 38274
rect 55582 38222 55634 38274
rect 2942 38110 2994 38162
rect 8766 38110 8818 38162
rect 13582 38110 13634 38162
rect 14254 38110 14306 38162
rect 15598 38110 15650 38162
rect 17390 38110 17442 38162
rect 22206 38110 22258 38162
rect 26574 38110 26626 38162
rect 28142 38110 28194 38162
rect 33070 38110 33122 38162
rect 35310 38110 35362 38162
rect 40350 38110 40402 38162
rect 44046 38110 44098 38162
rect 48190 38110 48242 38162
rect 3054 37998 3106 38050
rect 4398 37998 4450 38050
rect 4734 37998 4786 38050
rect 5742 37998 5794 38050
rect 6302 37998 6354 38050
rect 7086 37998 7138 38050
rect 7870 37998 7922 38050
rect 8318 37998 8370 38050
rect 9326 37998 9378 38050
rect 11342 37998 11394 38050
rect 12238 37998 12290 38050
rect 15262 37998 15314 38050
rect 15934 37998 15986 38050
rect 17054 37998 17106 38050
rect 18734 37998 18786 38050
rect 19742 37998 19794 38050
rect 21422 37998 21474 38050
rect 23550 37998 23602 38050
rect 24558 37998 24610 38050
rect 24782 37998 24834 38050
rect 25454 37998 25506 38050
rect 25678 37998 25730 38050
rect 32398 37998 32450 38050
rect 36094 37998 36146 38050
rect 36430 37998 36482 38050
rect 36990 37998 37042 38050
rect 37214 37998 37266 38050
rect 37438 37998 37490 38050
rect 37886 37998 37938 38050
rect 40238 37998 40290 38050
rect 41582 37998 41634 38050
rect 45390 37998 45442 38050
rect 46398 37998 46450 38050
rect 46846 37998 46898 38050
rect 47182 37998 47234 38050
rect 47966 37998 48018 38050
rect 48750 37998 48802 38050
rect 50206 37998 50258 38050
rect 51998 37998 52050 38050
rect 53790 37998 53842 38050
rect 54462 37998 54514 38050
rect 55134 37998 55186 38050
rect 4846 37886 4898 37938
rect 9214 37886 9266 37938
rect 9438 37886 9490 37938
rect 11230 37886 11282 37938
rect 19070 37886 19122 37938
rect 20078 37886 20130 37938
rect 21646 37886 21698 37938
rect 22542 37886 22594 37938
rect 24222 37886 24274 37938
rect 26014 37886 26066 37938
rect 29822 37886 29874 37938
rect 43934 37886 43986 37938
rect 48302 37886 48354 37938
rect 50094 37886 50146 37938
rect 1822 37774 1874 37826
rect 9886 37774 9938 37826
rect 12798 37774 12850 37826
rect 18958 37774 19010 37826
rect 29934 37774 29986 37826
rect 30158 37774 30210 37826
rect 30494 37774 30546 37826
rect 35870 37774 35922 37826
rect 36318 37774 36370 37826
rect 37102 37774 37154 37826
rect 38222 37774 38274 37826
rect 45614 37774 45666 37826
rect 51886 37774 51938 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 50558 37606 50610 37658
rect 50662 37606 50714 37658
rect 50766 37606 50818 37658
rect 5518 37438 5570 37490
rect 9550 37438 9602 37490
rect 9886 37438 9938 37490
rect 10782 37438 10834 37490
rect 13470 37438 13522 37490
rect 27806 37438 27858 37490
rect 31614 37438 31666 37490
rect 33518 37438 33570 37490
rect 33966 37438 34018 37490
rect 35646 37438 35698 37490
rect 37550 37438 37602 37490
rect 40350 37438 40402 37490
rect 4734 37326 4786 37378
rect 4846 37326 4898 37378
rect 5182 37326 5234 37378
rect 6638 37326 6690 37378
rect 12014 37326 12066 37378
rect 14030 37326 14082 37378
rect 14590 37326 14642 37378
rect 15710 37326 15762 37378
rect 18062 37326 18114 37378
rect 19966 37326 20018 37378
rect 20078 37326 20130 37378
rect 21422 37326 21474 37378
rect 22542 37326 22594 37378
rect 24446 37326 24498 37378
rect 26350 37326 26402 37378
rect 26798 37326 26850 37378
rect 27918 37326 27970 37378
rect 34526 37326 34578 37378
rect 34862 37326 34914 37378
rect 38558 37326 38610 37378
rect 46846 37326 46898 37378
rect 47630 37326 47682 37378
rect 55470 37326 55522 37378
rect 57822 37326 57874 37378
rect 4174 37214 4226 37266
rect 5518 37214 5570 37266
rect 5742 37214 5794 37266
rect 6862 37214 6914 37266
rect 7870 37214 7922 37266
rect 10894 37214 10946 37266
rect 12910 37214 12962 37266
rect 13918 37214 13970 37266
rect 15150 37214 15202 37266
rect 15598 37214 15650 37266
rect 19070 37214 19122 37266
rect 21198 37214 21250 37266
rect 21534 37214 21586 37266
rect 22430 37214 22482 37266
rect 23326 37214 23378 37266
rect 23886 37214 23938 37266
rect 24110 37214 24162 37266
rect 25902 37214 25954 37266
rect 26014 37214 26066 37266
rect 26686 37214 26738 37266
rect 26910 37214 26962 37266
rect 27358 37214 27410 37266
rect 27582 37214 27634 37266
rect 28366 37214 28418 37266
rect 34302 37214 34354 37266
rect 37214 37214 37266 37266
rect 37438 37214 37490 37266
rect 37774 37214 37826 37266
rect 38110 37214 38162 37266
rect 38334 37214 38386 37266
rect 39118 37214 39170 37266
rect 42590 37214 42642 37266
rect 43486 37214 43538 37266
rect 44270 37214 44322 37266
rect 44942 37214 44994 37266
rect 46734 37214 46786 37266
rect 47518 37214 47570 37266
rect 48078 37214 48130 37266
rect 50094 37214 50146 37266
rect 50766 37214 50818 37266
rect 52670 37214 52722 37266
rect 54462 37214 54514 37266
rect 54798 37214 54850 37266
rect 55246 37214 55298 37266
rect 58158 37214 58210 37266
rect 11454 37102 11506 37154
rect 15486 37102 15538 37154
rect 17502 37102 17554 37154
rect 19630 37102 19682 37154
rect 22654 37102 22706 37154
rect 24334 37102 24386 37154
rect 25342 37102 25394 37154
rect 26238 37102 26290 37154
rect 29038 37102 29090 37154
rect 31166 37102 31218 37154
rect 38446 37102 38498 37154
rect 38894 37102 38946 37154
rect 39790 37102 39842 37154
rect 42702 37102 42754 37154
rect 43598 37102 43650 37154
rect 46174 37102 46226 37154
rect 47294 37102 47346 37154
rect 48974 37102 49026 37154
rect 52222 37102 52274 37154
rect 53902 37102 53954 37154
rect 55358 37102 55410 37154
rect 56030 37102 56082 37154
rect 57598 37102 57650 37154
rect 1934 36990 1986 37042
rect 4734 36990 4786 37042
rect 8990 36990 9042 37042
rect 11006 36990 11058 37042
rect 20078 36990 20130 37042
rect 21982 36990 22034 37042
rect 39454 36990 39506 37042
rect 40014 36990 40066 37042
rect 46846 36990 46898 37042
rect 48302 36990 48354 37042
rect 50318 36990 50370 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 2270 36654 2322 36706
rect 2606 36654 2658 36706
rect 6750 36654 6802 36706
rect 7086 36654 7138 36706
rect 10334 36654 10386 36706
rect 10782 36654 10834 36706
rect 11118 36654 11170 36706
rect 18510 36654 18562 36706
rect 18622 36654 18674 36706
rect 18958 36654 19010 36706
rect 22766 36654 22818 36706
rect 23102 36654 23154 36706
rect 24782 36654 24834 36706
rect 25118 36654 25170 36706
rect 38110 36654 38162 36706
rect 40574 36654 40626 36706
rect 43486 36654 43538 36706
rect 52670 36654 52722 36706
rect 53006 36654 53058 36706
rect 2830 36542 2882 36594
rect 3278 36542 3330 36594
rect 6526 36542 6578 36594
rect 12910 36542 12962 36594
rect 14366 36542 14418 36594
rect 14702 36542 14754 36594
rect 17166 36542 17218 36594
rect 18734 36542 18786 36594
rect 19966 36542 20018 36594
rect 26462 36542 26514 36594
rect 28590 36542 28642 36594
rect 29262 36542 29314 36594
rect 33854 36542 33906 36594
rect 34414 36542 34466 36594
rect 39902 36542 39954 36594
rect 40462 36542 40514 36594
rect 41694 36542 41746 36594
rect 44046 36542 44098 36594
rect 54126 36542 54178 36594
rect 57934 36542 57986 36594
rect 3726 36430 3778 36482
rect 4286 36430 4338 36482
rect 6190 36430 6242 36482
rect 7422 36430 7474 36482
rect 10222 36430 10274 36482
rect 11342 36430 11394 36482
rect 11678 36430 11730 36482
rect 12350 36430 12402 36482
rect 13806 36430 13858 36482
rect 15150 36430 15202 36482
rect 15598 36430 15650 36482
rect 17950 36430 18002 36482
rect 18174 36430 18226 36482
rect 19182 36430 19234 36482
rect 19854 36430 19906 36482
rect 20750 36430 20802 36482
rect 21310 36430 21362 36482
rect 22990 36430 23042 36482
rect 25678 36430 25730 36482
rect 29822 36430 29874 36482
rect 30942 36430 30994 36482
rect 37326 36430 37378 36482
rect 38222 36430 38274 36482
rect 40238 36430 40290 36482
rect 41358 36430 41410 36482
rect 43038 36430 43090 36482
rect 45614 36430 45666 36482
rect 47294 36430 47346 36482
rect 48414 36430 48466 36482
rect 50542 36430 50594 36482
rect 51214 36430 51266 36482
rect 51550 36430 51602 36482
rect 53230 36430 53282 36482
rect 54238 36430 54290 36482
rect 55246 36430 55298 36482
rect 55582 36430 55634 36482
rect 1710 36318 1762 36370
rect 2046 36318 2098 36370
rect 3614 36318 3666 36370
rect 4622 36318 4674 36370
rect 7646 36318 7698 36370
rect 7758 36318 7810 36370
rect 15822 36318 15874 36370
rect 16158 36318 16210 36370
rect 25006 36318 25058 36370
rect 31614 36318 31666 36370
rect 40910 36318 40962 36370
rect 43374 36318 43426 36370
rect 45950 36318 46002 36370
rect 46846 36318 46898 36370
rect 49086 36318 49138 36370
rect 49758 36318 49810 36370
rect 54126 36318 54178 36370
rect 1822 36206 1874 36258
rect 4734 36206 4786 36258
rect 4846 36206 4898 36258
rect 5630 36206 5682 36258
rect 8206 36206 8258 36258
rect 10334 36206 10386 36258
rect 11790 36206 11842 36258
rect 12014 36206 12066 36258
rect 16382 36206 16434 36258
rect 21646 36206 21698 36258
rect 23102 36206 23154 36258
rect 23774 36206 23826 36258
rect 29150 36206 29202 36258
rect 29374 36206 29426 36258
rect 34862 36206 34914 36258
rect 37550 36206 37602 36258
rect 38110 36206 38162 36258
rect 38670 36206 38722 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 50558 36038 50610 36090
rect 50662 36038 50714 36090
rect 50766 36038 50818 36090
rect 2606 35870 2658 35922
rect 2718 35870 2770 35922
rect 4958 35870 5010 35922
rect 5294 35870 5346 35922
rect 7310 35870 7362 35922
rect 10894 35870 10946 35922
rect 12686 35870 12738 35922
rect 13022 35870 13074 35922
rect 13582 35870 13634 35922
rect 27358 35870 27410 35922
rect 28142 35870 28194 35922
rect 28926 35870 28978 35922
rect 32174 35870 32226 35922
rect 32398 35870 32450 35922
rect 32958 35870 33010 35922
rect 33182 35870 33234 35922
rect 39678 35870 39730 35922
rect 40014 35870 40066 35922
rect 2046 35758 2098 35810
rect 2382 35758 2434 35810
rect 2942 35758 2994 35810
rect 6862 35758 6914 35810
rect 14478 35758 14530 35810
rect 17390 35758 17442 35810
rect 17614 35758 17666 35810
rect 18958 35758 19010 35810
rect 19182 35758 19234 35810
rect 23662 35758 23714 35810
rect 27694 35758 27746 35810
rect 38222 35758 38274 35810
rect 44046 35758 44098 35810
rect 45278 35758 45330 35810
rect 49870 35758 49922 35810
rect 50206 35758 50258 35810
rect 50430 35758 50482 35810
rect 51774 35758 51826 35810
rect 55470 35758 55522 35810
rect 57822 35758 57874 35810
rect 1710 35646 1762 35698
rect 2830 35646 2882 35698
rect 3726 35646 3778 35698
rect 4286 35646 4338 35698
rect 5630 35646 5682 35698
rect 6078 35646 6130 35698
rect 6526 35646 6578 35698
rect 7198 35646 7250 35698
rect 8654 35646 8706 35698
rect 10670 35646 10722 35698
rect 12910 35646 12962 35698
rect 13470 35646 13522 35698
rect 13806 35646 13858 35698
rect 14366 35646 14418 35698
rect 15038 35646 15090 35698
rect 15374 35646 15426 35698
rect 16382 35646 16434 35698
rect 17950 35646 18002 35698
rect 25230 35646 25282 35698
rect 28030 35646 28082 35698
rect 7758 35534 7810 35586
rect 9662 35534 9714 35586
rect 14254 35534 14306 35586
rect 15710 35534 15762 35586
rect 16046 35534 16098 35586
rect 17838 35534 17890 35586
rect 19294 35534 19346 35586
rect 21086 35534 21138 35586
rect 23438 35534 23490 35586
rect 24670 35534 24722 35586
rect 4398 35422 4450 35474
rect 7982 35422 8034 35474
rect 8318 35422 8370 35474
rect 8654 35422 8706 35474
rect 8990 35422 9042 35474
rect 13022 35422 13074 35474
rect 23774 35422 23826 35474
rect 28254 35646 28306 35698
rect 32510 35646 32562 35698
rect 33294 35646 33346 35698
rect 34862 35646 34914 35698
rect 38110 35646 38162 35698
rect 38446 35646 38498 35698
rect 38558 35646 38610 35698
rect 41134 35646 41186 35698
rect 41806 35646 41858 35698
rect 42590 35646 42642 35698
rect 49646 35646 49698 35698
rect 51550 35646 51602 35698
rect 54462 35646 54514 35698
rect 55246 35646 55298 35698
rect 58158 35646 58210 35698
rect 25342 35534 25394 35586
rect 25790 35534 25842 35586
rect 29374 35534 29426 35586
rect 30494 35534 30546 35586
rect 31950 35534 32002 35586
rect 33854 35534 33906 35586
rect 34190 35534 34242 35586
rect 35534 35534 35586 35586
rect 37662 35534 37714 35586
rect 38222 35534 38274 35586
rect 39118 35534 39170 35586
rect 43710 35534 43762 35586
rect 45726 35534 45778 35586
rect 57598 35534 57650 35586
rect 25790 35422 25842 35474
rect 28926 35422 28978 35474
rect 29262 35422 29314 35474
rect 42814 35422 42866 35474
rect 53118 35422 53170 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 4398 35086 4450 35138
rect 9774 35086 9826 35138
rect 10670 35086 10722 35138
rect 17726 35086 17778 35138
rect 19070 35086 19122 35138
rect 33182 35086 33234 35138
rect 34414 35086 34466 35138
rect 34638 35086 34690 35138
rect 35982 35086 36034 35138
rect 37998 35086 38050 35138
rect 39790 35086 39842 35138
rect 43150 35086 43202 35138
rect 54350 35086 54402 35138
rect 54574 35086 54626 35138
rect 4174 34974 4226 35026
rect 4734 34974 4786 35026
rect 6862 34974 6914 35026
rect 8766 34974 8818 35026
rect 9550 34974 9602 35026
rect 13582 34974 13634 35026
rect 16158 34974 16210 35026
rect 17166 34974 17218 35026
rect 18846 34974 18898 35026
rect 20190 34974 20242 35026
rect 21870 34974 21922 35026
rect 27918 34974 27970 35026
rect 30494 34974 30546 35026
rect 30942 34974 30994 35026
rect 32510 34974 32562 35026
rect 38782 34974 38834 35026
rect 39454 34974 39506 35026
rect 40350 34974 40402 35026
rect 41806 34974 41858 35026
rect 42590 34974 42642 35026
rect 52670 34974 52722 35026
rect 2606 34862 2658 34914
rect 3166 34862 3218 34914
rect 3614 34862 3666 34914
rect 5854 34862 5906 34914
rect 7310 34862 7362 34914
rect 8318 34862 8370 34914
rect 9214 34862 9266 34914
rect 10558 34862 10610 34914
rect 15150 34862 15202 34914
rect 15710 34862 15762 34914
rect 16046 34862 16098 34914
rect 16382 34862 16434 34914
rect 17502 34862 17554 34914
rect 19406 34862 19458 34914
rect 19742 34862 19794 34914
rect 19966 34862 20018 34914
rect 20414 34862 20466 34914
rect 23998 34862 24050 34914
rect 24222 34862 24274 34914
rect 24558 34862 24610 34914
rect 25006 34862 25058 34914
rect 28478 34862 28530 34914
rect 29262 34862 29314 34914
rect 29598 34862 29650 34914
rect 33518 34862 33570 34914
rect 33966 34862 34018 34914
rect 35086 34862 35138 34914
rect 38222 34862 38274 34914
rect 40798 34862 40850 34914
rect 41134 34862 41186 34914
rect 42702 34862 42754 34914
rect 43822 34862 43874 34914
rect 44158 34862 44210 34914
rect 45278 34862 45330 34914
rect 45726 34862 45778 34914
rect 47070 34862 47122 34914
rect 48526 34862 48578 34914
rect 48862 34862 48914 34914
rect 49982 34862 50034 34914
rect 51886 34862 51938 34914
rect 52222 34862 52274 34914
rect 53454 34862 53506 34914
rect 53902 34862 53954 34914
rect 54798 34862 54850 34914
rect 2046 34750 2098 34802
rect 2494 34750 2546 34802
rect 3838 34750 3890 34802
rect 7758 34750 7810 34802
rect 9102 34750 9154 34802
rect 10670 34750 10722 34802
rect 13918 34750 13970 34802
rect 25790 34750 25842 34802
rect 28366 34750 28418 34802
rect 29374 34750 29426 34802
rect 29934 34750 29986 34802
rect 30046 34750 30098 34802
rect 30830 34750 30882 34802
rect 31166 34750 31218 34802
rect 31390 34750 31442 34802
rect 32062 34750 32114 34802
rect 33854 34750 33906 34802
rect 35198 34750 35250 34802
rect 35870 34750 35922 34802
rect 37102 34750 37154 34802
rect 37214 34750 37266 34802
rect 39678 34750 39730 34802
rect 39790 34750 39842 34802
rect 44830 34750 44882 34802
rect 46174 34750 46226 34802
rect 48974 34750 49026 34802
rect 51998 34750 52050 34802
rect 52782 34750 52834 34802
rect 53006 34750 53058 34802
rect 1710 34638 1762 34690
rect 6190 34638 6242 34690
rect 10110 34638 10162 34690
rect 20526 34638 20578 34690
rect 20638 34638 20690 34690
rect 21422 34638 21474 34690
rect 24334 34638 24386 34690
rect 24446 34638 24498 34690
rect 28142 34638 28194 34690
rect 29710 34638 29762 34690
rect 32286 34638 32338 34690
rect 32510 34638 32562 34690
rect 33294 34638 33346 34690
rect 34750 34638 34802 34690
rect 35422 34638 35474 34690
rect 35982 34638 36034 34690
rect 36878 34638 36930 34690
rect 37662 34638 37714 34690
rect 40238 34638 40290 34690
rect 40462 34638 40514 34690
rect 41358 34638 41410 34690
rect 43934 34638 43986 34690
rect 46286 34638 46338 34690
rect 46510 34638 46562 34690
rect 49646 34638 49698 34690
rect 49870 34638 49922 34690
rect 53678 34638 53730 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 50558 34470 50610 34522
rect 50662 34470 50714 34522
rect 50766 34470 50818 34522
rect 4510 34302 4562 34354
rect 5854 34302 5906 34354
rect 7310 34302 7362 34354
rect 7534 34302 7586 34354
rect 8654 34302 8706 34354
rect 9662 34302 9714 34354
rect 10334 34302 10386 34354
rect 15262 34302 15314 34354
rect 15598 34302 15650 34354
rect 26014 34302 26066 34354
rect 26126 34302 26178 34354
rect 26238 34302 26290 34354
rect 27358 34302 27410 34354
rect 32958 34302 33010 34354
rect 35422 34302 35474 34354
rect 37550 34302 37602 34354
rect 41246 34302 41298 34354
rect 42926 34302 42978 34354
rect 43486 34302 43538 34354
rect 44494 34302 44546 34354
rect 45614 34302 45666 34354
rect 49310 34302 49362 34354
rect 52782 34302 52834 34354
rect 53454 34302 53506 34354
rect 5070 34190 5122 34242
rect 7086 34190 7138 34242
rect 9998 34190 10050 34242
rect 10670 34190 10722 34242
rect 12350 34190 12402 34242
rect 14254 34190 14306 34242
rect 15710 34190 15762 34242
rect 19742 34190 19794 34242
rect 20862 34190 20914 34242
rect 25342 34190 25394 34242
rect 30046 34190 30098 34242
rect 31278 34190 31330 34242
rect 31614 34190 31666 34242
rect 33742 34190 33794 34242
rect 34974 34190 35026 34242
rect 40910 34190 40962 34242
rect 41134 34190 41186 34242
rect 42142 34190 42194 34242
rect 43038 34190 43090 34242
rect 43598 34190 43650 34242
rect 44606 34190 44658 34242
rect 47518 34190 47570 34242
rect 49198 34190 49250 34242
rect 51998 34190 52050 34242
rect 53342 34190 53394 34242
rect 4286 34078 4338 34130
rect 4734 34078 4786 34130
rect 5294 34078 5346 34130
rect 5518 34078 5570 34130
rect 6750 34078 6802 34130
rect 7646 34078 7698 34130
rect 8094 34078 8146 34130
rect 8430 34078 8482 34130
rect 8542 34078 8594 34130
rect 11342 34078 11394 34130
rect 13582 34078 13634 34130
rect 14142 34078 14194 34130
rect 14926 34078 14978 34130
rect 20414 34078 20466 34130
rect 21086 34078 21138 34130
rect 24558 34078 24610 34130
rect 25118 34078 25170 34130
rect 25454 34078 25506 34130
rect 26686 34078 26738 34130
rect 27022 34078 27074 34130
rect 30718 34078 30770 34130
rect 32062 34078 32114 34130
rect 32174 34078 32226 34130
rect 32398 34078 32450 34130
rect 32622 34078 32674 34130
rect 33070 34078 33122 34130
rect 33518 34078 33570 34130
rect 33966 34078 34018 34130
rect 35198 34078 35250 34130
rect 35646 34078 35698 34130
rect 39902 34078 39954 34130
rect 41582 34078 41634 34130
rect 41806 34078 41858 34130
rect 42590 34078 42642 34130
rect 43150 34078 43202 34130
rect 43822 34078 43874 34130
rect 44158 34078 44210 34130
rect 44270 34078 44322 34130
rect 45390 34078 45442 34130
rect 45950 34078 46002 34130
rect 46622 34078 46674 34130
rect 49534 34078 49586 34130
rect 50318 34078 50370 34130
rect 50654 34078 50706 34130
rect 52446 34078 52498 34130
rect 53006 34078 53058 34130
rect 53678 34078 53730 34130
rect 6302 33966 6354 34018
rect 11566 33966 11618 34018
rect 12014 33966 12066 34018
rect 17614 33966 17666 34018
rect 21758 33966 21810 34018
rect 23886 33966 23938 34018
rect 27918 33966 27970 34018
rect 33294 33966 33346 34018
rect 35310 33966 35362 34018
rect 36654 33966 36706 34018
rect 39230 33966 39282 34018
rect 40126 33966 40178 34018
rect 41918 33966 41970 34018
rect 48078 33966 48130 34018
rect 49758 33966 49810 34018
rect 1934 33854 1986 33906
rect 12462 33854 12514 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 19518 33518 19570 33570
rect 19854 33518 19906 33570
rect 30606 33518 30658 33570
rect 40350 33518 40402 33570
rect 41022 33518 41074 33570
rect 41806 33518 41858 33570
rect 42142 33518 42194 33570
rect 43822 33518 43874 33570
rect 3614 33406 3666 33458
rect 8430 33406 8482 33458
rect 9326 33406 9378 33458
rect 9998 33406 10050 33458
rect 12798 33406 12850 33458
rect 14478 33406 14530 33458
rect 19182 33406 19234 33458
rect 23550 33406 23602 33458
rect 27806 33406 27858 33458
rect 29262 33406 29314 33458
rect 31950 33406 32002 33458
rect 34414 33406 34466 33458
rect 37102 33406 37154 33458
rect 40126 33406 40178 33458
rect 41134 33406 41186 33458
rect 46174 33406 46226 33458
rect 48414 33406 48466 33458
rect 51326 33406 51378 33458
rect 54910 33406 54962 33458
rect 57822 33406 57874 33458
rect 3502 33294 3554 33346
rect 3838 33294 3890 33346
rect 4062 33294 4114 33346
rect 5966 33294 6018 33346
rect 7086 33294 7138 33346
rect 11566 33294 11618 33346
rect 14366 33294 14418 33346
rect 15262 33294 15314 33346
rect 20638 33294 20690 33346
rect 21758 33294 21810 33346
rect 26798 33294 26850 33346
rect 31390 33294 31442 33346
rect 31614 33294 31666 33346
rect 34526 33294 34578 33346
rect 35534 33294 35586 33346
rect 37886 33294 37938 33346
rect 38558 33294 38610 33346
rect 41918 33294 41970 33346
rect 42702 33294 42754 33346
rect 42926 33294 42978 33346
rect 43934 33294 43986 33346
rect 45166 33294 45218 33346
rect 46286 33294 46338 33346
rect 47182 33294 47234 33346
rect 47518 33294 47570 33346
rect 48078 33294 48130 33346
rect 49870 33294 49922 33346
rect 53790 33294 53842 33346
rect 54574 33294 54626 33346
rect 55582 33294 55634 33346
rect 2046 33182 2098 33234
rect 2718 33182 2770 33234
rect 4958 33182 5010 33234
rect 6190 33182 6242 33234
rect 7758 33182 7810 33234
rect 10446 33182 10498 33234
rect 20526 33182 20578 33234
rect 21422 33182 21474 33234
rect 28142 33182 28194 33234
rect 30158 33182 30210 33234
rect 30494 33182 30546 33234
rect 30606 33182 30658 33234
rect 31054 33182 31106 33234
rect 31166 33182 31218 33234
rect 34862 33182 34914 33234
rect 35870 33182 35922 33234
rect 36094 33182 36146 33234
rect 37326 33182 37378 33234
rect 38334 33182 38386 33234
rect 42254 33182 42306 33234
rect 44830 33182 44882 33234
rect 46062 33182 46114 33234
rect 50766 33182 50818 33234
rect 53118 33182 53170 33234
rect 53566 33182 53618 33234
rect 54126 33182 54178 33234
rect 1710 33070 1762 33122
rect 2382 33070 2434 33122
rect 6526 33070 6578 33122
rect 7310 33070 7362 33122
rect 7870 33070 7922 33122
rect 8094 33070 8146 33122
rect 8878 33070 8930 33122
rect 28478 33070 28530 33122
rect 29710 33070 29762 33122
rect 31950 33070 32002 33122
rect 32174 33070 32226 33122
rect 32734 33070 32786 33122
rect 34974 33070 35026 33122
rect 35198 33070 35250 33122
rect 35758 33070 35810 33122
rect 37102 33070 37154 33122
rect 38222 33070 38274 33122
rect 40686 33070 40738 33122
rect 49310 33070 49362 33122
rect 53230 33070 53282 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 50558 32902 50610 32954
rect 50662 32902 50714 32954
rect 50766 32902 50818 32954
rect 3278 32734 3330 32786
rect 5518 32734 5570 32786
rect 7086 32734 7138 32786
rect 9662 32734 9714 32786
rect 17838 32734 17890 32786
rect 18734 32734 18786 32786
rect 20526 32734 20578 32786
rect 25454 32734 25506 32786
rect 26574 32734 26626 32786
rect 29822 32734 29874 32786
rect 42142 32734 42194 32786
rect 49646 32734 49698 32786
rect 51662 32734 51714 32786
rect 52222 32734 52274 32786
rect 56702 32734 56754 32786
rect 2494 32622 2546 32674
rect 5966 32622 6018 32674
rect 6190 32622 6242 32674
rect 9550 32622 9602 32674
rect 10110 32622 10162 32674
rect 20862 32622 20914 32674
rect 31054 32622 31106 32674
rect 42814 32622 42866 32674
rect 42926 32622 42978 32674
rect 43710 32622 43762 32674
rect 45166 32622 45218 32674
rect 49758 32622 49810 32674
rect 51550 32622 51602 32674
rect 52670 32622 52722 32674
rect 53006 32622 53058 32674
rect 53230 32622 53282 32674
rect 57262 32622 57314 32674
rect 2270 32510 2322 32562
rect 3950 32510 4002 32562
rect 4958 32510 5010 32562
rect 5854 32510 5906 32562
rect 6638 32510 6690 32562
rect 7422 32510 7474 32562
rect 7646 32510 7698 32562
rect 8094 32510 8146 32562
rect 8542 32510 8594 32562
rect 10222 32510 10274 32562
rect 11902 32510 11954 32562
rect 13470 32510 13522 32562
rect 14478 32510 14530 32562
rect 15262 32510 15314 32562
rect 17390 32510 17442 32562
rect 17726 32510 17778 32562
rect 18062 32510 18114 32562
rect 21310 32510 21362 32562
rect 24558 32510 24610 32562
rect 25118 32510 25170 32562
rect 25454 32510 25506 32562
rect 25790 32510 25842 32562
rect 26350 32510 26402 32562
rect 28702 32510 28754 32562
rect 29038 32510 29090 32562
rect 30718 32510 30770 32562
rect 34750 32510 34802 32562
rect 42366 32510 42418 32562
rect 42590 32510 42642 32562
rect 43822 32510 43874 32562
rect 44718 32510 44770 32562
rect 45278 32510 45330 32562
rect 45838 32510 45890 32562
rect 46622 32510 46674 32562
rect 51886 32510 51938 32562
rect 52110 32510 52162 32562
rect 52446 32510 52498 32562
rect 54462 32510 54514 32562
rect 54686 32510 54738 32562
rect 54910 32510 54962 32562
rect 56590 32510 56642 32562
rect 57150 32510 57202 32562
rect 12350 32398 12402 32450
rect 13582 32398 13634 32450
rect 15150 32398 15202 32450
rect 17950 32398 18002 32450
rect 21758 32398 21810 32450
rect 23886 32398 23938 32450
rect 27022 32398 27074 32450
rect 27470 32398 27522 32450
rect 27918 32398 27970 32450
rect 28254 32398 28306 32450
rect 29486 32398 29538 32450
rect 30382 32398 30434 32450
rect 31502 32398 31554 32450
rect 33182 32398 33234 32450
rect 38334 32398 38386 32450
rect 43934 32398 43986 32450
rect 52782 32398 52834 32450
rect 6862 32286 6914 32338
rect 8094 32286 8146 32338
rect 9662 32286 9714 32338
rect 27470 32286 27522 32338
rect 27918 32286 27970 32338
rect 28366 32286 28418 32338
rect 30158 32286 30210 32338
rect 42030 32286 42082 32338
rect 49646 32286 49698 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 17502 31950 17554 32002
rect 23886 31950 23938 32002
rect 26574 31950 26626 32002
rect 27694 31950 27746 32002
rect 34974 31950 35026 32002
rect 45278 31950 45330 32002
rect 1934 31838 1986 31890
rect 5630 31838 5682 31890
rect 7982 31838 8034 31890
rect 8654 31838 8706 31890
rect 12014 31838 12066 31890
rect 13694 31838 13746 31890
rect 16382 31838 16434 31890
rect 16830 31838 16882 31890
rect 19182 31838 19234 31890
rect 22206 31838 22258 31890
rect 22766 31838 22818 31890
rect 23662 31838 23714 31890
rect 23998 31838 24050 31890
rect 26126 31838 26178 31890
rect 28030 31838 28082 31890
rect 29598 31838 29650 31890
rect 32398 31838 32450 31890
rect 34638 31838 34690 31890
rect 35086 31838 35138 31890
rect 35982 31838 36034 31890
rect 39902 31838 39954 31890
rect 45054 31838 45106 31890
rect 47966 31838 48018 31890
rect 49198 31838 49250 31890
rect 51550 31838 51602 31890
rect 52110 31838 52162 31890
rect 57934 31838 57986 31890
rect 4286 31726 4338 31778
rect 4622 31726 4674 31778
rect 6190 31726 6242 31778
rect 7422 31726 7474 31778
rect 8542 31726 8594 31778
rect 8878 31726 8930 31778
rect 9662 31726 9714 31778
rect 10110 31726 10162 31778
rect 10334 31726 10386 31778
rect 11790 31726 11842 31778
rect 13918 31726 13970 31778
rect 14254 31726 14306 31778
rect 14590 31726 14642 31778
rect 14926 31726 14978 31778
rect 16158 31726 16210 31778
rect 16606 31726 16658 31778
rect 17726 31726 17778 31778
rect 25118 31726 25170 31778
rect 25454 31726 25506 31778
rect 26014 31726 26066 31778
rect 26350 31726 26402 31778
rect 26574 31726 26626 31778
rect 27694 31726 27746 31778
rect 28254 31726 28306 31778
rect 29374 31726 29426 31778
rect 29822 31726 29874 31778
rect 31054 31726 31106 31778
rect 31950 31726 32002 31778
rect 33182 31726 33234 31778
rect 33854 31726 33906 31778
rect 36430 31726 36482 31778
rect 37102 31726 37154 31778
rect 40350 31726 40402 31778
rect 45502 31726 45554 31778
rect 46622 31726 46674 31778
rect 48190 31726 48242 31778
rect 48750 31726 48802 31778
rect 49086 31726 49138 31778
rect 51886 31726 51938 31778
rect 53454 31726 53506 31778
rect 54126 31726 54178 31778
rect 55582 31726 55634 31778
rect 4958 31614 5010 31666
rect 11678 31614 11730 31666
rect 16830 31614 16882 31666
rect 18174 31614 18226 31666
rect 18734 31614 18786 31666
rect 24446 31614 24498 31666
rect 25230 31614 25282 31666
rect 27358 31614 27410 31666
rect 31166 31614 31218 31666
rect 31502 31614 31554 31666
rect 33518 31614 33570 31666
rect 34190 31614 34242 31666
rect 34302 31614 34354 31666
rect 35310 31614 35362 31666
rect 35646 31614 35698 31666
rect 35870 31614 35922 31666
rect 37774 31614 37826 31666
rect 44942 31614 44994 31666
rect 45950 31614 46002 31666
rect 46062 31614 46114 31666
rect 46510 31614 46562 31666
rect 47070 31614 47122 31666
rect 47182 31614 47234 31666
rect 49646 31614 49698 31666
rect 54350 31614 54402 31666
rect 6526 31502 6578 31554
rect 6862 31502 6914 31554
rect 7086 31502 7138 31554
rect 7310 31502 7362 31554
rect 9326 31502 9378 31554
rect 10222 31502 10274 31554
rect 14814 31502 14866 31554
rect 17054 31502 17106 31554
rect 17950 31502 18002 31554
rect 18062 31502 18114 31554
rect 20302 31502 20354 31554
rect 20750 31502 20802 31554
rect 21310 31502 21362 31554
rect 21646 31502 21698 31554
rect 23102 31502 23154 31554
rect 24782 31502 24834 31554
rect 28590 31502 28642 31554
rect 29598 31502 29650 31554
rect 32846 31502 32898 31554
rect 33406 31502 33458 31554
rect 34078 31502 34130 31554
rect 45726 31502 45778 31554
rect 46286 31502 46338 31554
rect 47406 31502 47458 31554
rect 47630 31502 47682 31554
rect 52894 31502 52946 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 50558 31334 50610 31386
rect 50662 31334 50714 31386
rect 50766 31334 50818 31386
rect 8094 31166 8146 31218
rect 8878 31166 8930 31218
rect 9774 31166 9826 31218
rect 21198 31166 21250 31218
rect 21310 31166 21362 31218
rect 22094 31166 22146 31218
rect 22318 31166 22370 31218
rect 26574 31166 26626 31218
rect 26910 31166 26962 31218
rect 32958 31166 33010 31218
rect 35982 31166 36034 31218
rect 36430 31166 36482 31218
rect 37550 31166 37602 31218
rect 38558 31166 38610 31218
rect 38670 31166 38722 31218
rect 48974 31166 49026 31218
rect 49310 31166 49362 31218
rect 54798 31166 54850 31218
rect 2382 31054 2434 31106
rect 2606 31054 2658 31106
rect 6750 31054 6802 31106
rect 10222 31054 10274 31106
rect 12462 31054 12514 31106
rect 21086 31054 21138 31106
rect 23662 31054 23714 31106
rect 23998 31054 24050 31106
rect 24558 31054 24610 31106
rect 25230 31054 25282 31106
rect 25342 31054 25394 31106
rect 25454 31054 25506 31106
rect 34190 31054 34242 31106
rect 35198 31054 35250 31106
rect 35646 31054 35698 31106
rect 39230 31054 39282 31106
rect 42478 31054 42530 31106
rect 43150 31054 43202 31106
rect 44494 31054 44546 31106
rect 45838 31054 45890 31106
rect 46846 31054 46898 31106
rect 48750 31054 48802 31106
rect 49198 31054 49250 31106
rect 49534 31054 49586 31106
rect 51102 31054 51154 31106
rect 3054 30942 3106 30994
rect 3502 30942 3554 30994
rect 4510 30942 4562 30994
rect 5630 30942 5682 30994
rect 5854 30942 5906 30994
rect 6078 30942 6130 30994
rect 6526 30942 6578 30994
rect 7086 30942 7138 30994
rect 7646 30942 7698 30994
rect 7870 30942 7922 30994
rect 8542 30942 8594 30994
rect 8766 30942 8818 30994
rect 8990 30942 9042 30994
rect 9550 30942 9602 30994
rect 10670 30942 10722 30994
rect 11790 30942 11842 30994
rect 16158 30942 16210 30994
rect 16606 30942 16658 30994
rect 20190 30942 20242 30994
rect 20638 30942 20690 30994
rect 21422 30942 21474 30994
rect 21646 30942 21698 30994
rect 22990 30942 23042 30994
rect 23326 30942 23378 30994
rect 24334 30942 24386 30994
rect 26014 30942 26066 30994
rect 27246 30942 27298 30994
rect 33070 30942 33122 30994
rect 34078 30942 34130 30994
rect 35086 30942 35138 30994
rect 37326 30942 37378 30994
rect 38222 30942 38274 30994
rect 38446 30942 38498 30994
rect 39118 30942 39170 30994
rect 41358 30942 41410 30994
rect 42254 30942 42306 30994
rect 42814 30942 42866 30994
rect 44382 30942 44434 30994
rect 44606 30942 44658 30994
rect 45054 30942 45106 30994
rect 46286 30942 46338 30994
rect 46622 30942 46674 30994
rect 47630 30942 47682 30994
rect 48078 30942 48130 30994
rect 50206 30942 50258 30994
rect 52670 30942 52722 30994
rect 53006 30942 53058 30994
rect 53790 30942 53842 30994
rect 54126 30942 54178 30994
rect 54350 30942 54402 30994
rect 2270 30830 2322 30882
rect 3278 30830 3330 30882
rect 3726 30830 3778 30882
rect 4062 30830 4114 30882
rect 5406 30830 5458 30882
rect 12126 30830 12178 30882
rect 13246 30830 13298 30882
rect 15374 30830 15426 30882
rect 17390 30830 17442 30882
rect 19518 30830 19570 30882
rect 22206 30830 22258 30882
rect 24110 30830 24162 30882
rect 31838 30830 31890 30882
rect 36318 30830 36370 30882
rect 39678 30830 39730 30882
rect 41022 30830 41074 30882
rect 42366 30830 42418 30882
rect 46398 30830 46450 30882
rect 47182 30830 47234 30882
rect 51662 30830 51714 30882
rect 54686 30830 54738 30882
rect 7086 30718 7138 30770
rect 8206 30718 8258 30770
rect 25790 30718 25842 30770
rect 36654 30718 36706 30770
rect 37662 30718 37714 30770
rect 37998 30718 38050 30770
rect 45278 30718 45330 30770
rect 45614 30718 45666 30770
rect 52558 30718 52610 30770
rect 55022 30718 55074 30770
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 9998 30382 10050 30434
rect 16046 30382 16098 30434
rect 19406 30382 19458 30434
rect 28254 30382 28306 30434
rect 31502 30382 31554 30434
rect 45166 30382 45218 30434
rect 57934 30382 57986 30434
rect 5966 30270 6018 30322
rect 9662 30270 9714 30322
rect 12462 30270 12514 30322
rect 26350 30270 26402 30322
rect 28478 30270 28530 30322
rect 29598 30270 29650 30322
rect 31838 30270 31890 30322
rect 37662 30270 37714 30322
rect 37998 30270 38050 30322
rect 42702 30270 42754 30322
rect 43374 30270 43426 30322
rect 43598 30270 43650 30322
rect 43934 30270 43986 30322
rect 45614 30270 45666 30322
rect 51214 30270 51266 30322
rect 52670 30270 52722 30322
rect 54798 30270 54850 30322
rect 4286 30158 4338 30210
rect 4622 30158 4674 30210
rect 7422 30158 7474 30210
rect 8990 30158 9042 30210
rect 10110 30158 10162 30210
rect 10894 30158 10946 30210
rect 11454 30158 11506 30210
rect 14478 30158 14530 30210
rect 15710 30158 15762 30210
rect 16830 30158 16882 30210
rect 18286 30158 18338 30210
rect 20190 30158 20242 30210
rect 24558 30158 24610 30210
rect 26798 30158 26850 30210
rect 27358 30158 27410 30210
rect 28030 30158 28082 30210
rect 29486 30158 29538 30210
rect 30494 30158 30546 30210
rect 32286 30158 32338 30210
rect 33294 30158 33346 30210
rect 34526 30158 34578 30210
rect 35310 30158 35362 30210
rect 36318 30158 36370 30210
rect 37214 30158 37266 30210
rect 39566 30158 39618 30210
rect 39790 30158 39842 30210
rect 40574 30158 40626 30210
rect 44270 30158 44322 30210
rect 45726 30158 45778 30210
rect 46286 30158 46338 30210
rect 47182 30158 47234 30210
rect 47742 30158 47794 30210
rect 48974 30158 49026 30210
rect 49982 30158 50034 30210
rect 50318 30158 50370 30210
rect 50990 30158 51042 30210
rect 53342 30158 53394 30210
rect 55582 30158 55634 30210
rect 2494 30046 2546 30098
rect 4958 30046 5010 30098
rect 6526 30046 6578 30098
rect 8094 30046 8146 30098
rect 14702 30046 14754 30098
rect 15374 30046 15426 30098
rect 16606 30046 16658 30098
rect 18510 30046 18562 30098
rect 19070 30046 19122 30098
rect 20078 30046 20130 30098
rect 23886 30046 23938 30098
rect 27582 30046 27634 30098
rect 30830 30046 30882 30098
rect 31278 30046 31330 30098
rect 32510 30046 32562 30098
rect 34414 30046 34466 30098
rect 34974 30046 35026 30098
rect 37774 30046 37826 30098
rect 38558 30046 38610 30098
rect 47070 30046 47122 30098
rect 49870 30046 49922 30098
rect 54238 30046 54290 30098
rect 20750 29934 20802 29986
rect 21646 29934 21698 29986
rect 25230 29934 25282 29986
rect 25566 29934 25618 29986
rect 27022 29934 27074 29986
rect 29822 29934 29874 29986
rect 34302 29934 34354 29986
rect 35758 29934 35810 29986
rect 36990 29934 37042 29986
rect 38894 29934 38946 29986
rect 43038 29934 43090 29986
rect 44046 29934 44098 29986
rect 46398 29934 46450 29986
rect 46622 29934 46674 29986
rect 48974 29934 49026 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 50558 29766 50610 29818
rect 50662 29766 50714 29818
rect 50766 29766 50818 29818
rect 7758 29598 7810 29650
rect 8990 29598 9042 29650
rect 20078 29598 20130 29650
rect 23214 29598 23266 29650
rect 23662 29598 23714 29650
rect 24222 29598 24274 29650
rect 24782 29598 24834 29650
rect 25454 29598 25506 29650
rect 28590 29598 28642 29650
rect 28702 29598 28754 29650
rect 29150 29598 29202 29650
rect 30046 29598 30098 29650
rect 31950 29598 32002 29650
rect 32286 29598 32338 29650
rect 34638 29598 34690 29650
rect 37998 29598 38050 29650
rect 40350 29598 40402 29650
rect 40798 29598 40850 29650
rect 45838 29598 45890 29650
rect 46062 29598 46114 29650
rect 7534 29486 7586 29538
rect 8318 29486 8370 29538
rect 14590 29486 14642 29538
rect 16718 29486 16770 29538
rect 20302 29486 20354 29538
rect 20862 29486 20914 29538
rect 22206 29486 22258 29538
rect 23550 29486 23602 29538
rect 26014 29486 26066 29538
rect 26798 29486 26850 29538
rect 30382 29486 30434 29538
rect 34750 29486 34802 29538
rect 35534 29486 35586 29538
rect 35982 29486 36034 29538
rect 37326 29486 37378 29538
rect 37550 29486 37602 29538
rect 42030 29486 42082 29538
rect 42702 29486 42754 29538
rect 44606 29486 44658 29538
rect 46174 29486 46226 29538
rect 4286 29374 4338 29426
rect 5294 29374 5346 29426
rect 5518 29374 5570 29426
rect 6414 29374 6466 29426
rect 6638 29374 6690 29426
rect 7422 29374 7474 29426
rect 7870 29374 7922 29426
rect 8430 29374 8482 29426
rect 8542 29374 8594 29426
rect 14366 29374 14418 29426
rect 15598 29374 15650 29426
rect 16606 29374 16658 29426
rect 21310 29374 21362 29426
rect 21534 29374 21586 29426
rect 22542 29374 22594 29426
rect 22878 29374 22930 29426
rect 25790 29374 25842 29426
rect 26350 29374 26402 29426
rect 26574 29374 26626 29426
rect 27134 29374 27186 29426
rect 27582 29374 27634 29426
rect 27806 29374 27858 29426
rect 28030 29374 28082 29426
rect 28478 29374 28530 29426
rect 29374 29374 29426 29426
rect 30606 29374 30658 29426
rect 31614 29374 31666 29426
rect 33406 29374 33458 29426
rect 34638 29374 34690 29426
rect 35310 29374 35362 29426
rect 36206 29374 36258 29426
rect 36766 29374 36818 29426
rect 37102 29374 37154 29426
rect 37886 29374 37938 29426
rect 38110 29374 38162 29426
rect 38558 29374 38610 29426
rect 40910 29374 40962 29426
rect 41918 29374 41970 29426
rect 42814 29374 42866 29426
rect 45278 29374 45330 29426
rect 45502 29374 45554 29426
rect 15934 29262 15986 29314
rect 18174 29262 18226 29314
rect 19630 29262 19682 29314
rect 26462 29262 26514 29314
rect 27694 29262 27746 29314
rect 31166 29262 31218 29314
rect 37438 29262 37490 29314
rect 39902 29262 39954 29314
rect 1934 29150 1986 29202
rect 6638 29150 6690 29202
rect 21758 29150 21810 29202
rect 21870 29150 21922 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 5630 28814 5682 28866
rect 5966 28814 6018 28866
rect 17390 28814 17442 28866
rect 28478 28814 28530 28866
rect 41246 28814 41298 28866
rect 2270 28702 2322 28754
rect 13470 28702 13522 28754
rect 15598 28702 15650 28754
rect 19070 28702 19122 28754
rect 19630 28702 19682 28754
rect 20750 28702 20802 28754
rect 29262 28702 29314 28754
rect 31166 28702 31218 28754
rect 36430 28702 36482 28754
rect 49758 28702 49810 28754
rect 57934 28702 57986 28754
rect 1934 28590 1986 28642
rect 2718 28590 2770 28642
rect 3054 28590 3106 28642
rect 16382 28590 16434 28642
rect 17054 28590 17106 28642
rect 17950 28590 18002 28642
rect 26686 28590 26738 28642
rect 27694 28590 27746 28642
rect 28030 28590 28082 28642
rect 29598 28590 29650 28642
rect 30046 28590 30098 28642
rect 30830 28590 30882 28642
rect 31614 28590 31666 28642
rect 32174 28590 32226 28642
rect 32510 28590 32562 28642
rect 33294 28590 33346 28642
rect 34526 28590 34578 28642
rect 35086 28590 35138 28642
rect 35310 28590 35362 28642
rect 35982 28590 36034 28642
rect 36990 28590 37042 28642
rect 37662 28590 37714 28642
rect 38670 28590 38722 28642
rect 40350 28590 40402 28642
rect 41022 28590 41074 28642
rect 41582 28590 41634 28642
rect 42254 28590 42306 28642
rect 42702 28590 42754 28642
rect 42926 28590 42978 28642
rect 43710 28590 43762 28642
rect 50318 28590 50370 28642
rect 50654 28590 50706 28642
rect 51102 28590 51154 28642
rect 51774 28590 51826 28642
rect 51998 28590 52050 28642
rect 55582 28590 55634 28642
rect 5854 28478 5906 28530
rect 18062 28478 18114 28530
rect 19294 28478 19346 28530
rect 19518 28478 19570 28530
rect 22094 28478 22146 28530
rect 27470 28478 27522 28530
rect 28366 28478 28418 28530
rect 33630 28478 33682 28530
rect 34974 28478 35026 28530
rect 37326 28478 37378 28530
rect 37998 28478 38050 28530
rect 39342 28478 39394 28530
rect 41806 28478 41858 28530
rect 43150 28478 43202 28530
rect 43262 28478 43314 28530
rect 3390 28366 3442 28418
rect 20190 28366 20242 28418
rect 27582 28366 27634 28418
rect 28478 28366 28530 28418
rect 30382 28366 30434 28418
rect 32846 28366 32898 28418
rect 33966 28366 34018 28418
rect 34750 28366 34802 28418
rect 35758 28366 35810 28418
rect 35870 28366 35922 28418
rect 38558 28366 38610 28418
rect 39118 28366 39170 28418
rect 39230 28366 39282 28418
rect 39902 28366 39954 28418
rect 40798 28366 40850 28418
rect 41694 28366 41746 28418
rect 42142 28366 42194 28418
rect 42366 28366 42418 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 50558 28198 50610 28250
rect 50662 28198 50714 28250
rect 50766 28198 50818 28250
rect 2046 28030 2098 28082
rect 2718 28030 2770 28082
rect 3614 28030 3666 28082
rect 18062 28030 18114 28082
rect 18510 28030 18562 28082
rect 18734 28030 18786 28082
rect 21646 28030 21698 28082
rect 22430 28030 22482 28082
rect 23326 28030 23378 28082
rect 25566 28030 25618 28082
rect 33294 28030 33346 28082
rect 33630 28030 33682 28082
rect 35422 28030 35474 28082
rect 36654 28030 36706 28082
rect 37102 28030 37154 28082
rect 37326 28030 37378 28082
rect 39230 28030 39282 28082
rect 39342 28030 39394 28082
rect 39790 28030 39842 28082
rect 40014 28030 40066 28082
rect 52670 28030 52722 28082
rect 16270 27918 16322 27970
rect 16606 27918 16658 27970
rect 17614 27918 17666 27970
rect 19070 27918 19122 27970
rect 20302 27918 20354 27970
rect 21758 27918 21810 27970
rect 22206 27918 22258 27970
rect 22654 27918 22706 27970
rect 23662 27918 23714 27970
rect 24110 27918 24162 27970
rect 29374 27918 29426 27970
rect 35198 27918 35250 27970
rect 35870 27918 35922 27970
rect 38446 27918 38498 27970
rect 41694 27918 41746 27970
rect 44494 27918 44546 27970
rect 48750 27918 48802 27970
rect 53230 27918 53282 27970
rect 1822 27806 1874 27858
rect 2382 27806 2434 27858
rect 18398 27806 18450 27858
rect 19294 27806 19346 27858
rect 19630 27806 19682 27858
rect 20190 27806 20242 27858
rect 21198 27806 21250 27858
rect 23886 27806 23938 27858
rect 24222 27806 24274 27858
rect 25678 27806 25730 27858
rect 26126 27806 26178 27858
rect 29598 27806 29650 27858
rect 30046 27806 30098 27858
rect 30942 27806 30994 27858
rect 33966 27806 34018 27858
rect 34974 27806 35026 27858
rect 35982 27806 36034 27858
rect 37774 27806 37826 27858
rect 38222 27806 38274 27858
rect 38558 27806 38610 27858
rect 38782 27806 38834 27858
rect 39454 27806 39506 27858
rect 40462 27806 40514 27858
rect 40910 27806 40962 27858
rect 45166 27806 45218 27858
rect 46286 27806 46338 27858
rect 47966 27806 48018 27858
rect 49198 27806 49250 27858
rect 50990 27806 51042 27858
rect 51214 27806 51266 27858
rect 51886 27806 51938 27858
rect 52558 27806 52610 27858
rect 53118 27806 53170 27858
rect 3166 27694 3218 27746
rect 18958 27694 19010 27746
rect 22542 27694 22594 27746
rect 24670 27694 24722 27746
rect 26798 27694 26850 27746
rect 28926 27694 28978 27746
rect 30606 27694 30658 27746
rect 31390 27694 31442 27746
rect 32510 27694 32562 27746
rect 37214 27694 37266 27746
rect 39902 27694 39954 27746
rect 43822 27694 43874 27746
rect 45390 27694 45442 27746
rect 47630 27694 47682 27746
rect 49086 27694 49138 27746
rect 52110 27694 52162 27746
rect 57598 27694 57650 27746
rect 19966 27582 20018 27634
rect 25566 27582 25618 27634
rect 45950 27582 46002 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 18958 27246 19010 27298
rect 22094 27246 22146 27298
rect 57934 27246 57986 27298
rect 15150 27134 15202 27186
rect 17278 27134 17330 27186
rect 20078 27134 20130 27186
rect 20526 27134 20578 27186
rect 22654 27134 22706 27186
rect 22878 27134 22930 27186
rect 25006 27134 25058 27186
rect 26574 27134 26626 27186
rect 27134 27134 27186 27186
rect 27694 27134 27746 27186
rect 28590 27134 28642 27186
rect 29262 27134 29314 27186
rect 30382 27134 30434 27186
rect 32174 27134 32226 27186
rect 32510 27134 32562 27186
rect 37774 27134 37826 27186
rect 39902 27134 39954 27186
rect 41022 27134 41074 27186
rect 43150 27134 43202 27186
rect 47966 27134 48018 27186
rect 51774 27134 51826 27186
rect 52670 27134 52722 27186
rect 1710 27022 1762 27074
rect 2494 27022 2546 27074
rect 3166 27022 3218 27074
rect 3614 27022 3666 27074
rect 6862 27022 6914 27074
rect 7758 27022 7810 27074
rect 17950 27022 18002 27074
rect 19070 27022 19122 27074
rect 19294 27022 19346 27074
rect 19406 27022 19458 27074
rect 21310 27022 21362 27074
rect 21534 27022 21586 27074
rect 21646 27022 21698 27074
rect 25678 27022 25730 27074
rect 26014 27022 26066 27074
rect 27582 27022 27634 27074
rect 28254 27022 28306 27074
rect 29710 27022 29762 27074
rect 30830 27022 30882 27074
rect 32622 27022 32674 27074
rect 32846 27022 32898 27074
rect 33966 27022 34018 27074
rect 35310 27022 35362 27074
rect 35982 27022 36034 27074
rect 36990 27022 37042 27074
rect 40350 27022 40402 27074
rect 45502 27022 45554 27074
rect 46622 27022 46674 27074
rect 47406 27022 47458 27074
rect 48078 27022 48130 27074
rect 49086 27022 49138 27074
rect 50206 27022 50258 27074
rect 50990 27022 51042 27074
rect 51886 27022 51938 27074
rect 53118 27022 53170 27074
rect 53566 27022 53618 27074
rect 55582 27022 55634 27074
rect 2046 26910 2098 26962
rect 2718 26910 2770 26962
rect 6526 26910 6578 26962
rect 9102 26910 9154 26962
rect 18622 26910 18674 26962
rect 26462 26910 26514 26962
rect 33070 26910 33122 26962
rect 33294 26910 33346 26962
rect 35198 26910 35250 26962
rect 36094 26910 36146 26962
rect 45614 26910 45666 26962
rect 48750 26910 48802 26962
rect 49198 26910 49250 26962
rect 54350 26910 54402 26962
rect 54462 26910 54514 26962
rect 54686 26910 54738 26962
rect 54910 26910 54962 26962
rect 26686 26798 26738 26850
rect 27806 26798 27858 26850
rect 31614 26798 31666 26850
rect 33854 26798 33906 26850
rect 46510 26798 46562 26850
rect 49982 26798 50034 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 50558 26630 50610 26682
rect 50662 26630 50714 26682
rect 50766 26630 50818 26682
rect 2046 26462 2098 26514
rect 2718 26462 2770 26514
rect 3390 26462 3442 26514
rect 12686 26462 12738 26514
rect 14926 26462 14978 26514
rect 15486 26462 15538 26514
rect 25566 26462 25618 26514
rect 26462 26462 26514 26514
rect 26686 26462 26738 26514
rect 28142 26462 28194 26514
rect 28926 26462 28978 26514
rect 29934 26462 29986 26514
rect 31726 26462 31778 26514
rect 41806 26462 41858 26514
rect 42478 26462 42530 26514
rect 47518 26462 47570 26514
rect 51662 26462 51714 26514
rect 52558 26462 52610 26514
rect 55582 26462 55634 26514
rect 4734 26350 4786 26402
rect 5406 26350 5458 26402
rect 6302 26350 6354 26402
rect 12462 26350 12514 26402
rect 13806 26350 13858 26402
rect 14030 26350 14082 26402
rect 18398 26350 18450 26402
rect 26126 26350 26178 26402
rect 27694 26350 27746 26402
rect 29710 26350 29762 26402
rect 30606 26350 30658 26402
rect 30942 26350 30994 26402
rect 31166 26350 31218 26402
rect 32174 26350 32226 26402
rect 33518 26350 33570 26402
rect 41918 26350 41970 26402
rect 42814 26350 42866 26402
rect 45950 26350 46002 26402
rect 50318 26350 50370 26402
rect 51886 26350 51938 26402
rect 51998 26350 52050 26402
rect 52446 26350 52498 26402
rect 52670 26350 52722 26402
rect 53118 26350 53170 26402
rect 54126 26350 54178 26402
rect 57822 26350 57874 26402
rect 1822 26238 1874 26290
rect 2382 26238 2434 26290
rect 3054 26238 3106 26290
rect 5182 26238 5234 26290
rect 6862 26238 6914 26290
rect 7758 26238 7810 26290
rect 8206 26238 8258 26290
rect 9550 26238 9602 26290
rect 9886 26238 9938 26290
rect 10110 26238 10162 26290
rect 11118 26238 11170 26290
rect 11454 26238 11506 26290
rect 11566 26238 11618 26290
rect 12350 26238 12402 26290
rect 13134 26238 13186 26290
rect 14366 26238 14418 26290
rect 14702 26238 14754 26290
rect 16494 26238 16546 26290
rect 18286 26238 18338 26290
rect 18622 26238 18674 26290
rect 23662 26238 23714 26290
rect 25118 26238 25170 26290
rect 25454 26238 25506 26290
rect 25678 26238 25730 26290
rect 27134 26238 27186 26290
rect 27470 26238 27522 26290
rect 30158 26238 30210 26290
rect 30382 26238 30434 26290
rect 30718 26238 30770 26290
rect 31278 26238 31330 26290
rect 31502 26238 31554 26290
rect 31838 26238 31890 26290
rect 32510 26238 32562 26290
rect 33742 26238 33794 26290
rect 34078 26238 34130 26290
rect 34974 26238 35026 26290
rect 41582 26238 41634 26290
rect 43262 26238 43314 26290
rect 44494 26238 44546 26290
rect 45166 26238 45218 26290
rect 46062 26238 46114 26290
rect 47742 26238 47794 26290
rect 49646 26238 49698 26290
rect 50094 26238 50146 26290
rect 50430 26238 50482 26290
rect 52894 26238 52946 26290
rect 53230 26238 53282 26290
rect 54798 26238 54850 26290
rect 55358 26238 55410 26290
rect 55694 26238 55746 26290
rect 55918 26238 55970 26290
rect 56590 26238 56642 26290
rect 58158 26238 58210 26290
rect 3838 26126 3890 26178
rect 4286 26126 4338 26178
rect 9998 26126 10050 26178
rect 12910 26126 12962 26178
rect 18958 26126 19010 26178
rect 19406 26126 19458 26178
rect 20750 26126 20802 26178
rect 22990 26126 23042 26178
rect 24222 26126 24274 26178
rect 25902 26126 25954 26178
rect 26574 26126 26626 26178
rect 29262 26126 29314 26178
rect 30046 26126 30098 26178
rect 33182 26126 33234 26178
rect 33966 26126 34018 26178
rect 34526 26126 34578 26178
rect 37102 26126 37154 26178
rect 41022 26126 41074 26178
rect 43710 26126 43762 26178
rect 44382 26126 44434 26178
rect 45278 26126 45330 26178
rect 49422 26126 49474 26178
rect 53790 26126 53842 26178
rect 54574 26126 54626 26178
rect 57374 26126 57426 26178
rect 13470 26014 13522 26066
rect 14142 26014 14194 26066
rect 15038 26014 15090 26066
rect 16606 26014 16658 26066
rect 18734 26014 18786 26066
rect 19518 26014 19570 26066
rect 40798 26014 40850 26066
rect 41470 26014 41522 26066
rect 45950 26014 46002 26066
rect 47406 26014 47458 26066
rect 49086 26014 49138 26066
rect 56590 26014 56642 26066
rect 56926 26014 56978 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 5966 25678 6018 25730
rect 22990 25678 23042 25730
rect 23214 25678 23266 25730
rect 23774 25678 23826 25730
rect 37774 25678 37826 25730
rect 38222 25678 38274 25730
rect 38446 25678 38498 25730
rect 45502 25678 45554 25730
rect 52782 25678 52834 25730
rect 54686 25678 54738 25730
rect 57486 25678 57538 25730
rect 1934 25566 1986 25618
rect 6750 25566 6802 25618
rect 13918 25566 13970 25618
rect 20526 25566 20578 25618
rect 24894 25566 24946 25618
rect 27022 25566 27074 25618
rect 27470 25566 27522 25618
rect 29934 25566 29986 25618
rect 33070 25566 33122 25618
rect 35758 25566 35810 25618
rect 38446 25566 38498 25618
rect 46286 25566 46338 25618
rect 46958 25566 47010 25618
rect 49982 25566 50034 25618
rect 55022 25566 55074 25618
rect 4286 25454 4338 25506
rect 4846 25454 4898 25506
rect 5966 25454 6018 25506
rect 6638 25454 6690 25506
rect 7534 25454 7586 25506
rect 7870 25454 7922 25506
rect 8878 25454 8930 25506
rect 9438 25454 9490 25506
rect 9774 25454 9826 25506
rect 9998 25454 10050 25506
rect 11454 25454 11506 25506
rect 11678 25454 11730 25506
rect 14030 25454 14082 25506
rect 14702 25454 14754 25506
rect 15038 25454 15090 25506
rect 16606 25454 16658 25506
rect 18174 25454 18226 25506
rect 18734 25454 18786 25506
rect 19518 25454 19570 25506
rect 23662 25454 23714 25506
rect 24222 25454 24274 25506
rect 27806 25454 27858 25506
rect 29262 25454 29314 25506
rect 32622 25454 32674 25506
rect 33406 25454 33458 25506
rect 34190 25454 34242 25506
rect 35086 25454 35138 25506
rect 35982 25454 36034 25506
rect 37550 25454 37602 25506
rect 37998 25454 38050 25506
rect 40238 25454 40290 25506
rect 40686 25454 40738 25506
rect 41134 25454 41186 25506
rect 41582 25454 41634 25506
rect 44830 25454 44882 25506
rect 45166 25454 45218 25506
rect 45950 25454 46002 25506
rect 46734 25454 46786 25506
rect 47182 25454 47234 25506
rect 47630 25454 47682 25506
rect 47966 25454 48018 25506
rect 48638 25454 48690 25506
rect 49534 25454 49586 25506
rect 50206 25454 50258 25506
rect 50318 25454 50370 25506
rect 50654 25454 50706 25506
rect 53566 25454 53618 25506
rect 53902 25454 53954 25506
rect 54574 25454 54626 25506
rect 55582 25454 55634 25506
rect 5630 25342 5682 25394
rect 7198 25342 7250 25394
rect 7646 25342 7698 25394
rect 8430 25342 8482 25394
rect 10670 25342 10722 25394
rect 12350 25342 12402 25394
rect 16270 25342 16322 25394
rect 18510 25342 18562 25394
rect 20078 25342 20130 25394
rect 28142 25342 28194 25394
rect 33070 25342 33122 25394
rect 33182 25342 33234 25394
rect 35198 25342 35250 25394
rect 36206 25342 36258 25394
rect 37438 25342 37490 25394
rect 47406 25342 47458 25394
rect 47854 25342 47906 25394
rect 49758 25342 49810 25394
rect 52782 25342 52834 25394
rect 52894 25342 52946 25394
rect 53678 25342 53730 25394
rect 5070 25230 5122 25282
rect 9326 25230 9378 25282
rect 10334 25230 10386 25282
rect 10782 25230 10834 25282
rect 11006 25230 11058 25282
rect 12014 25230 12066 25282
rect 12462 25230 12514 25282
rect 12574 25230 12626 25282
rect 15150 25230 15202 25282
rect 15374 25230 15426 25282
rect 17614 25230 17666 25282
rect 19070 25230 19122 25282
rect 19854 25230 19906 25282
rect 20190 25230 20242 25282
rect 22878 25230 22930 25282
rect 32174 25230 32226 25282
rect 37214 25230 37266 25282
rect 39006 25230 39058 25282
rect 39454 25230 39506 25282
rect 39902 25230 39954 25282
rect 41694 25230 41746 25282
rect 42142 25230 42194 25282
rect 44942 25230 44994 25282
rect 48862 25230 48914 25282
rect 50542 25230 50594 25282
rect 52110 25230 52162 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 50558 25062 50610 25114
rect 50662 25062 50714 25114
rect 50766 25062 50818 25114
rect 4286 24894 4338 24946
rect 5406 24894 5458 24946
rect 16718 24894 16770 24946
rect 20862 24894 20914 24946
rect 21646 24894 21698 24946
rect 22206 24894 22258 24946
rect 24110 24894 24162 24946
rect 26462 24894 26514 24946
rect 3278 24782 3330 24834
rect 16270 24782 16322 24834
rect 16606 24782 16658 24834
rect 26910 24838 26962 24890
rect 27246 24894 27298 24946
rect 32174 24894 32226 24946
rect 32510 24894 32562 24946
rect 35422 24894 35474 24946
rect 42590 24894 42642 24946
rect 45614 24894 45666 24946
rect 46062 24894 46114 24946
rect 27022 24782 27074 24834
rect 27694 24782 27746 24834
rect 27806 24782 27858 24834
rect 30270 24782 30322 24834
rect 30382 24782 30434 24834
rect 33518 24782 33570 24834
rect 34302 24782 34354 24834
rect 34638 24782 34690 24834
rect 35758 24782 35810 24834
rect 39902 24782 39954 24834
rect 41022 24782 41074 24834
rect 41694 24782 41746 24834
rect 43822 24782 43874 24834
rect 2046 24670 2098 24722
rect 3054 24670 3106 24722
rect 3390 24670 3442 24722
rect 3838 24670 3890 24722
rect 4734 24670 4786 24722
rect 6302 24670 6354 24722
rect 7870 24670 7922 24722
rect 8094 24670 8146 24722
rect 8318 24670 8370 24722
rect 9102 24670 9154 24722
rect 9774 24670 9826 24722
rect 11790 24670 11842 24722
rect 12686 24670 12738 24722
rect 13582 24670 13634 24722
rect 15598 24670 15650 24722
rect 16942 24670 16994 24722
rect 17278 24670 17330 24722
rect 18062 24670 18114 24722
rect 19294 24670 19346 24722
rect 20190 24670 20242 24722
rect 20526 24670 20578 24722
rect 20862 24670 20914 24722
rect 21198 24670 21250 24722
rect 21422 24670 21474 24722
rect 21758 24670 21810 24722
rect 30046 24670 30098 24722
rect 30830 24670 30882 24722
rect 32958 24670 33010 24722
rect 33294 24670 33346 24722
rect 34414 24670 34466 24722
rect 34862 24670 34914 24722
rect 35198 24670 35250 24722
rect 35646 24670 35698 24722
rect 36318 24670 36370 24722
rect 40014 24670 40066 24722
rect 41134 24670 41186 24722
rect 41582 24670 41634 24722
rect 42478 24670 42530 24722
rect 44270 24670 44322 24722
rect 45390 24670 45442 24722
rect 49086 24670 49138 24722
rect 49422 24670 49474 24722
rect 49982 24670 50034 24722
rect 50318 24670 50370 24722
rect 50654 24670 50706 24722
rect 52110 24670 52162 24722
rect 52558 24670 52610 24722
rect 53454 24670 53506 24722
rect 57150 24670 57202 24722
rect 2494 24558 2546 24610
rect 2830 24558 2882 24610
rect 4510 24558 4562 24610
rect 5742 24558 5794 24610
rect 6078 24558 6130 24610
rect 10558 24558 10610 24610
rect 11566 24558 11618 24610
rect 13470 24558 13522 24610
rect 15374 24558 15426 24610
rect 18510 24558 18562 24610
rect 19742 24558 19794 24610
rect 23662 24558 23714 24610
rect 28366 24558 28418 24610
rect 30382 24558 30434 24610
rect 33182 24558 33234 24610
rect 34750 24558 34802 24610
rect 35982 24558 36034 24610
rect 37102 24558 37154 24610
rect 39230 24558 39282 24610
rect 44158 24558 44210 24610
rect 49646 24558 49698 24610
rect 50430 24558 50482 24610
rect 53006 24558 53058 24610
rect 56702 24558 56754 24610
rect 57374 24558 57426 24610
rect 4958 24446 5010 24498
rect 6526 24446 6578 24498
rect 6750 24446 6802 24498
rect 7198 24446 7250 24498
rect 18286 24446 18338 24498
rect 27806 24446 27858 24498
rect 39902 24446 39954 24498
rect 41246 24446 41298 24498
rect 55358 24446 55410 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 3838 24110 3890 24162
rect 17838 24110 17890 24162
rect 18174 24110 18226 24162
rect 18622 24110 18674 24162
rect 20190 24110 20242 24162
rect 24222 24110 24274 24162
rect 34974 24110 35026 24162
rect 35198 24110 35250 24162
rect 37102 24110 37154 24162
rect 57934 24110 57986 24162
rect 2382 23998 2434 24050
rect 9214 23998 9266 24050
rect 10782 23998 10834 24050
rect 12910 23998 12962 24050
rect 17166 23998 17218 24050
rect 24446 23998 24498 24050
rect 25118 23998 25170 24050
rect 28366 23998 28418 24050
rect 30046 23998 30098 24050
rect 31726 23998 31778 24050
rect 33742 23998 33794 24050
rect 38222 23998 38274 24050
rect 39790 23998 39842 24050
rect 44942 23998 44994 24050
rect 45838 23998 45890 24050
rect 48414 23998 48466 24050
rect 2046 23886 2098 23938
rect 2830 23886 2882 23938
rect 3390 23886 3442 23938
rect 4622 23886 4674 23938
rect 5854 23886 5906 23938
rect 6526 23886 6578 23938
rect 6862 23886 6914 23938
rect 7086 23886 7138 23938
rect 7534 23886 7586 23938
rect 7870 23886 7922 23938
rect 8206 23886 8258 23938
rect 8542 23886 8594 23938
rect 12238 23886 12290 23938
rect 13694 23886 13746 23938
rect 14142 23886 14194 23938
rect 15598 23886 15650 23938
rect 16494 23886 16546 23938
rect 19742 23886 19794 23938
rect 19966 23886 20018 23938
rect 23998 23886 24050 23938
rect 25454 23886 25506 23938
rect 29598 23886 29650 23938
rect 30494 23886 30546 23938
rect 31614 23886 31666 23938
rect 34638 23886 34690 23938
rect 35870 23886 35922 23938
rect 36990 23886 37042 23938
rect 37774 23886 37826 23938
rect 39902 23886 39954 23938
rect 41022 23886 41074 23938
rect 41470 23886 41522 23938
rect 41918 23886 41970 23938
rect 44270 23886 44322 23938
rect 46286 23886 46338 23938
rect 46734 23886 46786 23938
rect 47518 23886 47570 23938
rect 49086 23886 49138 23938
rect 49870 23886 49922 23938
rect 52110 23886 52162 23938
rect 53678 23886 53730 23938
rect 55582 23886 55634 23938
rect 2942 23774 2994 23826
rect 3166 23774 3218 23826
rect 8878 23774 8930 23826
rect 11230 23774 11282 23826
rect 14366 23774 14418 23826
rect 14478 23774 14530 23826
rect 15486 23774 15538 23826
rect 18062 23774 18114 23826
rect 18510 23774 18562 23826
rect 19406 23774 19458 23826
rect 23326 23774 23378 23826
rect 23438 23774 23490 23826
rect 24558 23774 24610 23826
rect 26238 23774 26290 23826
rect 29262 23774 29314 23826
rect 30158 23774 30210 23826
rect 31278 23774 31330 23826
rect 34414 23774 34466 23826
rect 37102 23774 37154 23826
rect 37662 23774 37714 23826
rect 39342 23774 39394 23826
rect 43934 23774 43986 23826
rect 44046 23774 44098 23826
rect 49982 23774 50034 23826
rect 50990 23774 51042 23826
rect 51214 23774 51266 23826
rect 51438 23774 51490 23826
rect 53454 23774 53506 23826
rect 55022 23774 55074 23826
rect 55246 23774 55298 23826
rect 4062 23662 4114 23714
rect 5182 23662 5234 23714
rect 6190 23662 6242 23714
rect 6974 23662 7026 23714
rect 7198 23662 7250 23714
rect 7870 23662 7922 23714
rect 10446 23662 10498 23714
rect 13918 23662 13970 23714
rect 18622 23662 18674 23714
rect 19518 23662 19570 23714
rect 20526 23662 20578 23714
rect 22542 23662 22594 23714
rect 22878 23662 22930 23714
rect 23102 23662 23154 23714
rect 29374 23662 29426 23714
rect 29822 23662 29874 23714
rect 30046 23662 30098 23714
rect 30942 23662 30994 23714
rect 31166 23662 31218 23714
rect 33294 23662 33346 23714
rect 35198 23662 35250 23714
rect 35982 23662 36034 23714
rect 36206 23662 36258 23714
rect 37438 23662 37490 23714
rect 47742 23662 47794 23714
rect 50878 23662 50930 23714
rect 51774 23662 51826 23714
rect 51998 23662 52050 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 50558 23494 50610 23546
rect 50662 23494 50714 23546
rect 50766 23494 50818 23546
rect 7310 23326 7362 23378
rect 11678 23326 11730 23378
rect 15486 23326 15538 23378
rect 22318 23326 22370 23378
rect 24110 23326 24162 23378
rect 27358 23326 27410 23378
rect 27470 23326 27522 23378
rect 27806 23326 27858 23378
rect 30046 23326 30098 23378
rect 30830 23326 30882 23378
rect 31054 23326 31106 23378
rect 38558 23326 38610 23378
rect 40238 23326 40290 23378
rect 40462 23326 40514 23378
rect 41022 23326 41074 23378
rect 41470 23326 41522 23378
rect 42142 23326 42194 23378
rect 44046 23326 44098 23378
rect 46734 23326 46786 23378
rect 48078 23326 48130 23378
rect 53902 23326 53954 23378
rect 56142 23326 56194 23378
rect 58158 23326 58210 23378
rect 3726 23214 3778 23266
rect 4734 23214 4786 23266
rect 6862 23214 6914 23266
rect 8766 23214 8818 23266
rect 10670 23214 10722 23266
rect 13470 23214 13522 23266
rect 14926 23214 14978 23266
rect 15710 23214 15762 23266
rect 29822 23214 29874 23266
rect 35982 23214 36034 23266
rect 40126 23214 40178 23266
rect 47070 23214 47122 23266
rect 52334 23214 52386 23266
rect 55022 23214 55074 23266
rect 55806 23214 55858 23266
rect 55918 23214 55970 23266
rect 2270 23102 2322 23154
rect 4174 23102 4226 23154
rect 4846 23102 4898 23154
rect 7086 23102 7138 23154
rect 7758 23102 7810 23154
rect 8206 23102 8258 23154
rect 8654 23102 8706 23154
rect 9550 23102 9602 23154
rect 10110 23102 10162 23154
rect 11342 23102 11394 23154
rect 12462 23102 12514 23154
rect 12686 23102 12738 23154
rect 13806 23102 13858 23154
rect 14814 23102 14866 23154
rect 15822 23102 15874 23154
rect 16158 23102 16210 23154
rect 16718 23102 16770 23154
rect 18174 23102 18226 23154
rect 20862 23102 20914 23154
rect 21310 23102 21362 23154
rect 21982 23102 22034 23154
rect 22542 23102 22594 23154
rect 22878 23102 22930 23154
rect 23102 23102 23154 23154
rect 27582 23102 27634 23154
rect 29710 23102 29762 23154
rect 30718 23102 30770 23154
rect 33966 23102 34018 23154
rect 34414 23102 34466 23154
rect 34638 23102 34690 23154
rect 35310 23102 35362 23154
rect 40910 23102 40962 23154
rect 41246 23102 41298 23154
rect 41582 23102 41634 23154
rect 43038 23102 43090 23154
rect 43710 23102 43762 23154
rect 43934 23102 43986 23154
rect 44270 23102 44322 23154
rect 46398 23102 46450 23154
rect 47406 23102 47458 23154
rect 48190 23102 48242 23154
rect 50430 23102 50482 23154
rect 50878 23102 50930 23154
rect 53566 23102 53618 23154
rect 54686 23102 54738 23154
rect 55246 23102 55298 23154
rect 55470 23102 55522 23154
rect 57038 23102 57090 23154
rect 1822 22990 1874 23042
rect 2830 22990 2882 23042
rect 4286 22990 4338 23042
rect 10558 22990 10610 23042
rect 12350 22990 12402 23042
rect 14030 22990 14082 23042
rect 18734 22990 18786 23042
rect 20526 22990 20578 23042
rect 21758 22990 21810 23042
rect 22766 22990 22818 23042
rect 23550 22990 23602 23042
rect 23774 22990 23826 23042
rect 24670 22990 24722 23042
rect 34526 22990 34578 23042
rect 38110 22990 38162 23042
rect 42814 22990 42866 23042
rect 50542 22990 50594 23042
rect 52110 22990 52162 23042
rect 56702 22990 56754 23042
rect 57262 22990 57314 23042
rect 8766 22878 8818 22930
rect 14926 22878 14978 22930
rect 17838 22878 17890 22930
rect 18174 22878 18226 22930
rect 43374 22878 43426 22930
rect 51102 22878 51154 22930
rect 54462 22878 54514 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 8990 22542 9042 22594
rect 12910 22542 12962 22594
rect 13806 22542 13858 22594
rect 22542 22542 22594 22594
rect 28030 22542 28082 22594
rect 47854 22542 47906 22594
rect 49982 22542 50034 22594
rect 56814 22542 56866 22594
rect 4510 22430 4562 22482
rect 5854 22430 5906 22482
rect 14030 22430 14082 22482
rect 23662 22430 23714 22482
rect 25118 22430 25170 22482
rect 26462 22430 26514 22482
rect 29262 22430 29314 22482
rect 37886 22430 37938 22482
rect 39566 22430 39618 22482
rect 41134 22430 41186 22482
rect 42030 22430 42082 22482
rect 45166 22430 45218 22482
rect 47742 22430 47794 22482
rect 50542 22430 50594 22482
rect 56590 22430 56642 22482
rect 2494 22318 2546 22370
rect 5070 22318 5122 22370
rect 6750 22318 6802 22370
rect 7646 22318 7698 22370
rect 10670 22318 10722 22370
rect 11678 22318 11730 22370
rect 18174 22318 18226 22370
rect 19070 22318 19122 22370
rect 21870 22318 21922 22370
rect 22094 22318 22146 22370
rect 22654 22318 22706 22370
rect 23214 22318 23266 22370
rect 25566 22318 25618 22370
rect 26350 22318 26402 22370
rect 27918 22318 27970 22370
rect 28254 22318 28306 22370
rect 30942 22318 30994 22370
rect 31502 22318 31554 22370
rect 31726 22318 31778 22370
rect 32062 22318 32114 22370
rect 34078 22318 34130 22370
rect 34526 22318 34578 22370
rect 35198 22318 35250 22370
rect 35982 22318 36034 22370
rect 36206 22318 36258 22370
rect 36542 22318 36594 22370
rect 37438 22318 37490 22370
rect 40014 22318 40066 22370
rect 40462 22318 40514 22370
rect 40910 22318 40962 22370
rect 42590 22318 42642 22370
rect 43598 22318 43650 22370
rect 44830 22318 44882 22370
rect 45390 22318 45442 22370
rect 46286 22318 46338 22370
rect 47518 22318 47570 22370
rect 50318 22318 50370 22370
rect 51662 22318 51714 22370
rect 51886 22318 51938 22370
rect 52222 22318 52274 22370
rect 53902 22318 53954 22370
rect 54462 22318 54514 22370
rect 54910 22318 54962 22370
rect 55134 22318 55186 22370
rect 56254 22318 56306 22370
rect 56814 22318 56866 22370
rect 57150 22318 57202 22370
rect 57374 22318 57426 22370
rect 2718 22206 2770 22258
rect 3614 22206 3666 22258
rect 6638 22206 6690 22258
rect 10558 22206 10610 22258
rect 17950 22206 18002 22258
rect 20414 22206 20466 22258
rect 22542 22206 22594 22258
rect 23550 22206 23602 22258
rect 24334 22206 24386 22258
rect 24558 22206 24610 22258
rect 26014 22206 26066 22258
rect 26574 22206 26626 22258
rect 28590 22206 28642 22258
rect 33854 22206 33906 22258
rect 34190 22206 34242 22258
rect 34974 22206 35026 22258
rect 36318 22206 36370 22258
rect 36990 22206 37042 22258
rect 41246 22206 41298 22258
rect 43934 22206 43986 22258
rect 45950 22206 46002 22258
rect 46062 22206 46114 22258
rect 51326 22206 51378 22258
rect 51998 22206 52050 22258
rect 52670 22206 52722 22258
rect 53006 22206 53058 22258
rect 53454 22206 53506 22258
rect 55470 22206 55522 22258
rect 13470 22094 13522 22146
rect 21534 22094 21586 22146
rect 23326 22094 23378 22146
rect 23662 22094 23714 22146
rect 24446 22094 24498 22146
rect 27806 22094 27858 22146
rect 31054 22094 31106 22146
rect 31166 22094 31218 22146
rect 31950 22094 32002 22146
rect 34302 22094 34354 22146
rect 35086 22094 35138 22146
rect 47854 22094 47906 22146
rect 51438 22094 51490 22146
rect 54350 22094 54402 22146
rect 55134 22094 55186 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 50558 21926 50610 21978
rect 50662 21926 50714 21978
rect 50766 21926 50818 21978
rect 1822 21758 1874 21810
rect 9102 21758 9154 21810
rect 11230 21758 11282 21810
rect 11566 21758 11618 21810
rect 11790 21758 11842 21810
rect 12014 21758 12066 21810
rect 33182 21758 33234 21810
rect 33742 21758 33794 21810
rect 34862 21758 34914 21810
rect 38670 21758 38722 21810
rect 39342 21758 39394 21810
rect 39566 21758 39618 21810
rect 39678 21758 39730 21810
rect 41918 21758 41970 21810
rect 47742 21758 47794 21810
rect 49758 21758 49810 21810
rect 50990 21758 51042 21810
rect 51998 21758 52050 21810
rect 53230 21758 53282 21810
rect 54350 21758 54402 21810
rect 54686 21758 54738 21810
rect 2046 21646 2098 21698
rect 4286 21646 4338 21698
rect 8206 21646 8258 21698
rect 14478 21646 14530 21698
rect 16158 21646 16210 21698
rect 1710 21310 1762 21362
rect 25678 21646 25730 21698
rect 27022 21646 27074 21698
rect 28590 21646 28642 21698
rect 30270 21646 30322 21698
rect 35646 21646 35698 21698
rect 35870 21646 35922 21698
rect 35982 21646 36034 21698
rect 39902 21646 39954 21698
rect 41022 21646 41074 21698
rect 45054 21646 45106 21698
rect 46286 21646 46338 21698
rect 50766 21646 50818 21698
rect 51886 21646 51938 21698
rect 53006 21646 53058 21698
rect 55918 21646 55970 21698
rect 56702 21646 56754 21698
rect 2270 21534 2322 21586
rect 2494 21534 2546 21586
rect 2718 21534 2770 21586
rect 2830 21534 2882 21586
rect 4510 21534 4562 21586
rect 5630 21534 5682 21586
rect 6862 21534 6914 21586
rect 8430 21534 8482 21586
rect 8654 21534 8706 21586
rect 9438 21534 9490 21586
rect 10334 21534 10386 21586
rect 12126 21534 12178 21586
rect 15486 21534 15538 21586
rect 17614 21534 17666 21586
rect 18734 21534 18786 21586
rect 20302 21534 20354 21586
rect 21310 21534 21362 21586
rect 21758 21534 21810 21586
rect 23550 21534 23602 21586
rect 26350 21534 26402 21586
rect 27134 21534 27186 21586
rect 27470 21534 27522 21586
rect 29486 21534 29538 21586
rect 33966 21534 34018 21586
rect 34414 21534 34466 21586
rect 35086 21534 35138 21586
rect 35534 21534 35586 21586
rect 38558 21534 38610 21586
rect 38894 21534 38946 21586
rect 39006 21534 39058 21586
rect 40238 21534 40290 21586
rect 40910 21534 40962 21586
rect 41806 21534 41858 21586
rect 43710 21534 43762 21586
rect 44382 21534 44434 21586
rect 45278 21534 45330 21586
rect 47294 21534 47346 21586
rect 49534 21534 49586 21586
rect 51214 21534 51266 21586
rect 52110 21534 52162 21586
rect 52558 21534 52610 21586
rect 53566 21534 53618 21586
rect 54910 21534 54962 21586
rect 55582 21534 55634 21586
rect 56590 21534 56642 21586
rect 57486 21534 57538 21586
rect 3278 21422 3330 21474
rect 5182 21422 5234 21474
rect 8094 21422 8146 21474
rect 10110 21422 10162 21474
rect 12574 21422 12626 21474
rect 14030 21422 14082 21474
rect 17726 21422 17778 21474
rect 18174 21422 18226 21474
rect 19182 21422 19234 21474
rect 23662 21422 23714 21474
rect 24334 21422 24386 21474
rect 26014 21422 26066 21474
rect 28702 21422 28754 21474
rect 29150 21422 29202 21474
rect 32398 21422 32450 21474
rect 33854 21422 33906 21474
rect 34974 21422 35026 21474
rect 36430 21422 36482 21474
rect 38334 21422 38386 21474
rect 42478 21422 42530 21474
rect 43934 21422 43986 21474
rect 44606 21422 44658 21474
rect 45950 21422 46002 21474
rect 53342 21422 53394 21474
rect 55694 21422 55746 21474
rect 56814 21422 56866 21474
rect 10446 21310 10498 21362
rect 21758 21310 21810 21362
rect 27694 21310 27746 21362
rect 28030 21310 28082 21362
rect 28366 21310 28418 21362
rect 50654 21310 50706 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 7198 20974 7250 21026
rect 15374 20974 15426 21026
rect 15934 20974 15986 21026
rect 22878 20974 22930 21026
rect 23438 20974 23490 21026
rect 27470 20974 27522 21026
rect 36206 20974 36258 21026
rect 44046 20974 44098 21026
rect 46062 20974 46114 21026
rect 51662 20974 51714 21026
rect 55806 20974 55858 21026
rect 2494 20862 2546 20914
rect 3278 20862 3330 20914
rect 4846 20862 4898 20914
rect 9102 20862 9154 20914
rect 9886 20862 9938 20914
rect 13582 20862 13634 20914
rect 15374 20862 15426 20914
rect 17278 20862 17330 20914
rect 18622 20862 18674 20914
rect 22878 20862 22930 20914
rect 26014 20862 26066 20914
rect 27694 20862 27746 20914
rect 28030 20862 28082 20914
rect 32510 20862 32562 20914
rect 33630 20862 33682 20914
rect 35758 20862 35810 20914
rect 41358 20862 41410 20914
rect 50430 20862 50482 20914
rect 57262 20862 57314 20914
rect 1710 20750 1762 20802
rect 3726 20750 3778 20802
rect 4286 20750 4338 20802
rect 6190 20750 6242 20802
rect 6414 20750 6466 20802
rect 6974 20750 7026 20802
rect 7422 20750 7474 20802
rect 7870 20750 7922 20802
rect 8430 20750 8482 20802
rect 9326 20750 9378 20802
rect 10894 20750 10946 20802
rect 16830 20750 16882 20802
rect 18062 20750 18114 20802
rect 19070 20750 19122 20802
rect 19406 20750 19458 20802
rect 21758 20750 21810 20802
rect 22206 20750 22258 20802
rect 24222 20750 24274 20802
rect 24558 20750 24610 20802
rect 25230 20750 25282 20802
rect 26910 20750 26962 20802
rect 30718 20750 30770 20802
rect 31278 20750 31330 20802
rect 32398 20750 32450 20802
rect 32846 20750 32898 20802
rect 36094 20750 36146 20802
rect 40014 20750 40066 20802
rect 43374 20750 43426 20802
rect 43710 20750 43762 20802
rect 46958 20750 47010 20802
rect 49086 20750 49138 20802
rect 51102 20750 51154 20802
rect 56814 20750 56866 20802
rect 57038 20750 57090 20802
rect 58158 20750 58210 20802
rect 2046 20638 2098 20690
rect 3838 20638 3890 20690
rect 8990 20638 9042 20690
rect 9774 20638 9826 20690
rect 10334 20638 10386 20690
rect 10670 20638 10722 20690
rect 11118 20638 11170 20690
rect 11230 20638 11282 20690
rect 11678 20638 11730 20690
rect 12798 20638 12850 20690
rect 12910 20638 12962 20690
rect 21310 20638 21362 20690
rect 27358 20638 27410 20690
rect 27918 20638 27970 20690
rect 29262 20638 29314 20690
rect 29934 20638 29986 20690
rect 31726 20638 31778 20690
rect 32062 20638 32114 20690
rect 39454 20638 39506 20690
rect 41134 20638 41186 20690
rect 43934 20638 43986 20690
rect 45950 20638 46002 20690
rect 46062 20638 46114 20690
rect 46734 20638 46786 20690
rect 47294 20638 47346 20690
rect 49310 20638 49362 20690
rect 49646 20638 49698 20690
rect 50094 20638 50146 20690
rect 50542 20638 50594 20690
rect 50990 20638 51042 20690
rect 51214 20638 51266 20690
rect 55694 20638 55746 20690
rect 55806 20638 55858 20690
rect 57822 20638 57874 20690
rect 2830 20526 2882 20578
rect 4062 20526 4114 20578
rect 4510 20526 4562 20578
rect 4734 20526 4786 20578
rect 4846 20526 4898 20578
rect 5966 20526 6018 20578
rect 6302 20526 6354 20578
rect 8542 20526 8594 20578
rect 8766 20526 8818 20578
rect 9550 20526 9602 20578
rect 9886 20526 9938 20578
rect 12014 20526 12066 20578
rect 12686 20526 12738 20578
rect 15934 20526 15986 20578
rect 23326 20526 23378 20578
rect 27134 20526 27186 20578
rect 29710 20526 29762 20578
rect 29822 20526 29874 20578
rect 36206 20526 36258 20578
rect 37102 20526 37154 20578
rect 46958 20526 47010 20578
rect 48414 20526 48466 20578
rect 48526 20526 48578 20578
rect 48638 20526 48690 20578
rect 50318 20526 50370 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 50558 20358 50610 20410
rect 50662 20358 50714 20410
rect 50766 20358 50818 20410
rect 6750 20190 6802 20242
rect 24222 20190 24274 20242
rect 31054 20190 31106 20242
rect 33854 20190 33906 20242
rect 40350 20190 40402 20242
rect 56478 20190 56530 20242
rect 58270 20190 58322 20242
rect 3278 20078 3330 20130
rect 4958 20078 5010 20130
rect 5854 20078 5906 20130
rect 7198 20078 7250 20130
rect 7534 20078 7586 20130
rect 10446 20078 10498 20130
rect 12462 20078 12514 20130
rect 12574 20078 12626 20130
rect 13134 20078 13186 20130
rect 14478 20078 14530 20130
rect 16494 20078 16546 20130
rect 18174 20078 18226 20130
rect 19294 20078 19346 20130
rect 19630 20078 19682 20130
rect 20078 20078 20130 20130
rect 20414 20078 20466 20130
rect 21198 20078 21250 20130
rect 22878 20078 22930 20130
rect 23550 20078 23602 20130
rect 24446 20078 24498 20130
rect 25566 20078 25618 20130
rect 28254 20078 28306 20130
rect 29374 20078 29426 20130
rect 29822 20078 29874 20130
rect 30270 20078 30322 20130
rect 31502 20078 31554 20130
rect 31614 20078 31666 20130
rect 32622 20078 32674 20130
rect 35198 20078 35250 20130
rect 37774 20078 37826 20130
rect 39790 20078 39842 20130
rect 40126 20078 40178 20130
rect 40910 20078 40962 20130
rect 42478 20078 42530 20130
rect 42926 20078 42978 20130
rect 43822 20078 43874 20130
rect 48750 20078 48802 20130
rect 51326 20078 51378 20130
rect 52894 20078 52946 20130
rect 56702 20078 56754 20130
rect 2158 19966 2210 20018
rect 2606 19966 2658 20018
rect 3726 19966 3778 20018
rect 5070 19966 5122 20018
rect 6526 19966 6578 20018
rect 6862 19966 6914 20018
rect 9550 19966 9602 20018
rect 10334 19966 10386 20018
rect 11342 19966 11394 20018
rect 12238 19966 12290 20018
rect 12910 19966 12962 20018
rect 13470 19966 13522 20018
rect 15374 19966 15426 20018
rect 17390 19966 17442 20018
rect 18398 19966 18450 20018
rect 18958 19966 19010 20018
rect 21646 19966 21698 20018
rect 23102 19966 23154 20018
rect 24558 19966 24610 20018
rect 25230 19966 25282 20018
rect 27470 19966 27522 20018
rect 28142 19966 28194 20018
rect 29710 19966 29762 20018
rect 30046 19966 30098 20018
rect 30494 19966 30546 20018
rect 30718 19966 30770 20018
rect 30830 19966 30882 20018
rect 33070 19966 33122 20018
rect 33294 19966 33346 20018
rect 33854 19966 33906 20018
rect 34414 19966 34466 20018
rect 40238 19966 40290 20018
rect 41358 19966 41410 20018
rect 42366 19966 42418 20018
rect 42702 19966 42754 20018
rect 43150 19966 43202 20018
rect 43486 19966 43538 20018
rect 43598 19966 43650 20018
rect 43934 19966 43986 20018
rect 44158 19966 44210 20018
rect 49086 19966 49138 20018
rect 49310 19966 49362 20018
rect 50878 19966 50930 20018
rect 51102 19966 51154 20018
rect 51550 19966 51602 20018
rect 53118 19966 53170 20018
rect 54238 19966 54290 20018
rect 55022 19966 55074 20018
rect 56814 19966 56866 20018
rect 9998 19854 10050 19906
rect 11566 19854 11618 19906
rect 12014 19854 12066 19906
rect 13022 19854 13074 19906
rect 14030 19854 14082 19906
rect 17838 19854 17890 19906
rect 28030 19854 28082 19906
rect 37326 19854 37378 19906
rect 41694 19854 41746 19906
rect 43262 19854 43314 19906
rect 53790 19854 53842 19906
rect 54798 19854 54850 19906
rect 28926 19742 28978 19794
rect 29486 19742 29538 19794
rect 31726 19742 31778 19794
rect 33630 19742 33682 19794
rect 48862 19742 48914 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 4622 19406 4674 19458
rect 27806 19406 27858 19458
rect 33070 19406 33122 19458
rect 42366 19406 42418 19458
rect 42814 19406 42866 19458
rect 46286 19406 46338 19458
rect 47518 19406 47570 19458
rect 53006 19406 53058 19458
rect 54126 19406 54178 19458
rect 55806 19406 55858 19458
rect 4958 19294 5010 19346
rect 10558 19294 10610 19346
rect 11342 19294 11394 19346
rect 14254 19294 14306 19346
rect 17054 19294 17106 19346
rect 17950 19294 18002 19346
rect 19630 19294 19682 19346
rect 21422 19294 21474 19346
rect 23662 19294 23714 19346
rect 29598 19294 29650 19346
rect 33630 19294 33682 19346
rect 36990 19294 37042 19346
rect 37438 19294 37490 19346
rect 38334 19294 38386 19346
rect 40574 19294 40626 19346
rect 41022 19294 41074 19346
rect 45278 19294 45330 19346
rect 46622 19294 46674 19346
rect 47182 19294 47234 19346
rect 50430 19294 50482 19346
rect 51214 19294 51266 19346
rect 54462 19294 54514 19346
rect 54910 19294 54962 19346
rect 1822 19182 1874 19234
rect 3614 19182 3666 19234
rect 3950 19182 4002 19234
rect 4398 19182 4450 19234
rect 6078 19182 6130 19234
rect 6302 19182 6354 19234
rect 6862 19182 6914 19234
rect 8318 19182 8370 19234
rect 8878 19182 8930 19234
rect 10110 19182 10162 19234
rect 11230 19182 11282 19234
rect 14478 19182 14530 19234
rect 16494 19182 16546 19234
rect 18510 19182 18562 19234
rect 19518 19182 19570 19234
rect 20526 19182 20578 19234
rect 21646 19182 21698 19234
rect 22878 19182 22930 19234
rect 24782 19182 24834 19234
rect 25006 19182 25058 19234
rect 26014 19182 26066 19234
rect 26126 19182 26178 19234
rect 27582 19182 27634 19234
rect 28030 19182 28082 19234
rect 29150 19182 29202 19234
rect 30046 19182 30098 19234
rect 31614 19182 31666 19234
rect 32174 19182 32226 19234
rect 32734 19182 32786 19234
rect 37662 19182 37714 19234
rect 38782 19182 38834 19234
rect 39230 19182 39282 19234
rect 42030 19182 42082 19234
rect 42590 19182 42642 19234
rect 43486 19182 43538 19234
rect 43710 19182 43762 19234
rect 45166 19182 45218 19234
rect 48414 19182 48466 19234
rect 49646 19182 49698 19234
rect 50766 19182 50818 19234
rect 53342 19182 53394 19234
rect 53902 19182 53954 19234
rect 56142 19182 56194 19234
rect 57150 19182 57202 19234
rect 57486 19182 57538 19234
rect 2046 19070 2098 19122
rect 2382 19070 2434 19122
rect 2718 19070 2770 19122
rect 4062 19070 4114 19122
rect 5742 19070 5794 19122
rect 6414 19070 6466 19122
rect 15038 19070 15090 19122
rect 16606 19070 16658 19122
rect 18734 19070 18786 19122
rect 19742 19070 19794 19122
rect 20414 19070 20466 19122
rect 20750 19070 20802 19122
rect 25230 19070 25282 19122
rect 25566 19070 25618 19122
rect 25790 19070 25842 19122
rect 26686 19070 26738 19122
rect 29262 19070 29314 19122
rect 31502 19070 31554 19122
rect 32510 19070 32562 19122
rect 41806 19070 41858 19122
rect 43822 19070 43874 19122
rect 44270 19070 44322 19122
rect 46846 19070 46898 19122
rect 49422 19070 49474 19122
rect 53566 19070 53618 19122
rect 54798 19070 54850 19122
rect 55022 19070 55074 19122
rect 15934 18958 15986 19010
rect 17502 18958 17554 19010
rect 26798 18958 26850 19010
rect 27022 18958 27074 19010
rect 27694 18958 27746 19010
rect 32062 18958 32114 19010
rect 39678 18958 39730 19010
rect 40014 18958 40066 19010
rect 42254 18958 42306 19010
rect 43150 18958 43202 19010
rect 44942 18958 44994 19010
rect 45390 18958 45442 19010
rect 47406 18958 47458 19010
rect 48526 18958 48578 19010
rect 48750 18958 48802 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 50558 18790 50610 18842
rect 50662 18790 50714 18842
rect 50766 18790 50818 18842
rect 3390 18622 3442 18674
rect 3726 18622 3778 18674
rect 4062 18622 4114 18674
rect 14254 18622 14306 18674
rect 15822 18622 15874 18674
rect 24558 18622 24610 18674
rect 26574 18622 26626 18674
rect 28590 18622 28642 18674
rect 28814 18622 28866 18674
rect 31390 18622 31442 18674
rect 31502 18622 31554 18674
rect 32398 18622 32450 18674
rect 33294 18622 33346 18674
rect 35422 18622 35474 18674
rect 35870 18622 35922 18674
rect 37214 18622 37266 18674
rect 39118 18622 39170 18674
rect 42366 18622 42418 18674
rect 44942 18622 44994 18674
rect 2046 18510 2098 18562
rect 2718 18510 2770 18562
rect 3054 18510 3106 18562
rect 6974 18510 7026 18562
rect 10894 18510 10946 18562
rect 13134 18510 13186 18562
rect 15150 18510 15202 18562
rect 15710 18510 15762 18562
rect 16830 18510 16882 18562
rect 18062 18510 18114 18562
rect 21086 18510 21138 18562
rect 23214 18510 23266 18562
rect 23662 18510 23714 18562
rect 24446 18510 24498 18562
rect 26910 18510 26962 18562
rect 27694 18510 27746 18562
rect 30494 18510 30546 18562
rect 31278 18510 31330 18562
rect 35086 18510 35138 18562
rect 36990 18510 37042 18562
rect 37886 18510 37938 18562
rect 39902 18510 39954 18562
rect 44158 18510 44210 18562
rect 44270 18510 44322 18562
rect 46174 18510 46226 18562
rect 47182 18510 47234 18562
rect 51550 18510 51602 18562
rect 54126 18510 54178 18562
rect 56590 18510 56642 18562
rect 1822 18398 1874 18450
rect 2494 18398 2546 18450
rect 4510 18398 4562 18450
rect 4734 18398 4786 18450
rect 5070 18398 5122 18450
rect 5294 18398 5346 18450
rect 5518 18398 5570 18450
rect 5854 18398 5906 18450
rect 7758 18398 7810 18450
rect 9102 18398 9154 18450
rect 11902 18398 11954 18450
rect 13470 18398 13522 18450
rect 13694 18398 13746 18450
rect 13806 18398 13858 18450
rect 14590 18398 14642 18450
rect 14814 18398 14866 18450
rect 16046 18398 16098 18450
rect 16270 18398 16322 18450
rect 16494 18398 16546 18450
rect 16718 18398 16770 18450
rect 19294 18398 19346 18450
rect 20974 18398 21026 18450
rect 22766 18398 22818 18450
rect 23886 18398 23938 18450
rect 24782 18398 24834 18450
rect 25678 18398 25730 18450
rect 26014 18398 26066 18450
rect 26238 18398 26290 18450
rect 27470 18398 27522 18450
rect 28254 18398 28306 18450
rect 28926 18398 28978 18450
rect 30606 18398 30658 18450
rect 30830 18398 30882 18450
rect 35982 18398 36034 18450
rect 37438 18398 37490 18450
rect 38334 18398 38386 18450
rect 38894 18398 38946 18450
rect 40238 18398 40290 18450
rect 41134 18398 41186 18450
rect 42142 18398 42194 18450
rect 43150 18398 43202 18450
rect 45278 18398 45330 18450
rect 47406 18398 47458 18450
rect 47742 18398 47794 18450
rect 48974 18398 49026 18450
rect 50318 18398 50370 18450
rect 52222 18398 52274 18450
rect 53566 18398 53618 18450
rect 54574 18398 54626 18450
rect 57150 18398 57202 18450
rect 4846 18286 4898 18338
rect 6302 18286 6354 18338
rect 10334 18286 10386 18338
rect 15038 18286 15090 18338
rect 17838 18286 17890 18338
rect 20638 18286 20690 18338
rect 31838 18286 31890 18338
rect 36430 18286 36482 18338
rect 37326 18286 37378 18338
rect 37886 18286 37938 18338
rect 40350 18286 40402 18338
rect 41470 18286 41522 18338
rect 41694 18286 41746 18338
rect 42702 18286 42754 18338
rect 43038 18286 43090 18338
rect 46622 18286 46674 18338
rect 49086 18286 49138 18338
rect 53454 18286 53506 18338
rect 55022 18286 55074 18338
rect 57486 18286 57538 18338
rect 30494 18174 30546 18226
rect 32062 18174 32114 18226
rect 35870 18174 35922 18226
rect 44158 18174 44210 18226
rect 50542 18174 50594 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 9438 17838 9490 17890
rect 9550 17838 9602 17890
rect 14030 17838 14082 17890
rect 26126 17838 26178 17890
rect 29262 17838 29314 17890
rect 31502 17838 31554 17890
rect 34862 17838 34914 17890
rect 37550 17838 37602 17890
rect 5742 17726 5794 17778
rect 6526 17726 6578 17778
rect 8654 17726 8706 17778
rect 10558 17726 10610 17778
rect 12574 17726 12626 17778
rect 15150 17726 15202 17778
rect 15934 17726 15986 17778
rect 20862 17726 20914 17778
rect 23326 17726 23378 17778
rect 29710 17726 29762 17778
rect 31166 17726 31218 17778
rect 32734 17726 32786 17778
rect 34302 17726 34354 17778
rect 40798 17726 40850 17778
rect 42254 17726 42306 17778
rect 45166 17726 45218 17778
rect 47294 17726 47346 17778
rect 48526 17726 48578 17778
rect 55582 17726 55634 17778
rect 1710 17614 1762 17666
rect 3054 17614 3106 17666
rect 3950 17614 4002 17666
rect 7982 17614 8034 17666
rect 8990 17614 9042 17666
rect 9214 17614 9266 17666
rect 11902 17614 11954 17666
rect 13470 17614 13522 17666
rect 13694 17614 13746 17666
rect 14478 17614 14530 17666
rect 15486 17614 15538 17666
rect 17166 17614 17218 17666
rect 18622 17614 18674 17666
rect 19182 17614 19234 17666
rect 19294 17614 19346 17666
rect 19630 17614 19682 17666
rect 21646 17614 21698 17666
rect 21982 17614 22034 17666
rect 22206 17614 22258 17666
rect 22878 17614 22930 17666
rect 24446 17614 24498 17666
rect 25454 17614 25506 17666
rect 25790 17614 25842 17666
rect 29262 17614 29314 17666
rect 29822 17614 29874 17666
rect 31054 17614 31106 17666
rect 33070 17614 33122 17666
rect 33518 17614 33570 17666
rect 34526 17614 34578 17666
rect 35310 17614 35362 17666
rect 35646 17614 35698 17666
rect 35982 17614 36034 17666
rect 38558 17614 38610 17666
rect 38782 17614 38834 17666
rect 40350 17614 40402 17666
rect 41358 17614 41410 17666
rect 42478 17614 42530 17666
rect 45838 17614 45890 17666
rect 50878 17614 50930 17666
rect 56142 17614 56194 17666
rect 57150 17614 57202 17666
rect 2046 17502 2098 17554
rect 2382 17502 2434 17554
rect 2718 17502 2770 17554
rect 3390 17502 3442 17554
rect 4510 17502 4562 17554
rect 4846 17502 4898 17554
rect 6974 17502 7026 17554
rect 10894 17502 10946 17554
rect 14254 17502 14306 17554
rect 17278 17502 17330 17554
rect 19742 17502 19794 17554
rect 20526 17502 20578 17554
rect 21310 17502 21362 17554
rect 22318 17502 22370 17554
rect 37438 17502 37490 17554
rect 46846 17502 46898 17554
rect 48750 17502 48802 17554
rect 50318 17502 50370 17554
rect 50990 17502 51042 17554
rect 57374 17502 57426 17554
rect 4174 17390 4226 17442
rect 13918 17390 13970 17442
rect 16046 17390 16098 17442
rect 16158 17390 16210 17442
rect 17054 17390 17106 17442
rect 21422 17390 21474 17442
rect 35534 17390 35586 17442
rect 35758 17390 35810 17442
rect 36542 17390 36594 17442
rect 37102 17390 37154 17442
rect 50430 17390 50482 17442
rect 51214 17390 51266 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 50558 17222 50610 17274
rect 50662 17222 50714 17274
rect 50766 17222 50818 17274
rect 2046 17054 2098 17106
rect 2382 17054 2434 17106
rect 3054 17054 3106 17106
rect 3838 17054 3890 17106
rect 4510 17054 4562 17106
rect 4734 17054 4786 17106
rect 6302 17054 6354 17106
rect 6750 17054 6802 17106
rect 7646 17054 7698 17106
rect 11790 17054 11842 17106
rect 12462 17054 12514 17106
rect 14366 17054 14418 17106
rect 14590 17054 14642 17106
rect 20974 17054 21026 17106
rect 28142 17054 28194 17106
rect 28366 17054 28418 17106
rect 28702 17054 28754 17106
rect 28926 17054 28978 17106
rect 34974 17054 35026 17106
rect 35310 17054 35362 17106
rect 38334 17054 38386 17106
rect 43598 17054 43650 17106
rect 47854 17054 47906 17106
rect 53342 17054 53394 17106
rect 56926 17054 56978 17106
rect 5294 16942 5346 16994
rect 7758 16942 7810 16994
rect 12126 16942 12178 16994
rect 12798 16942 12850 16994
rect 14142 16942 14194 16994
rect 19518 16942 19570 16994
rect 21758 16942 21810 16994
rect 24334 16942 24386 16994
rect 25566 16942 25618 16994
rect 27470 16942 27522 16994
rect 37550 16942 37602 16994
rect 39566 16942 39618 16994
rect 41582 16942 41634 16994
rect 43038 16942 43090 16994
rect 46622 16942 46674 16994
rect 47966 16942 48018 16994
rect 52110 16942 52162 16994
rect 55022 16942 55074 16994
rect 57374 16942 57426 16994
rect 1822 16830 1874 16882
rect 2606 16830 2658 16882
rect 3278 16830 3330 16882
rect 3726 16830 3778 16882
rect 4286 16830 4338 16882
rect 4958 16830 5010 16882
rect 5854 16830 5906 16882
rect 7534 16830 7586 16882
rect 13022 16830 13074 16882
rect 13358 16830 13410 16882
rect 13582 16830 13634 16882
rect 15038 16830 15090 16882
rect 15374 16830 15426 16882
rect 15486 16830 15538 16882
rect 16270 16830 16322 16882
rect 18174 16830 18226 16882
rect 18846 16830 18898 16882
rect 19182 16830 19234 16882
rect 22094 16830 22146 16882
rect 22990 16830 23042 16882
rect 26126 16830 26178 16882
rect 26798 16830 26850 16882
rect 28030 16830 28082 16882
rect 28590 16830 28642 16882
rect 29262 16830 29314 16882
rect 29486 16830 29538 16882
rect 31390 16830 31442 16882
rect 34526 16830 34578 16882
rect 35758 16830 35810 16882
rect 36206 16830 36258 16882
rect 36766 16830 36818 16882
rect 39790 16830 39842 16882
rect 40462 16830 40514 16882
rect 46846 16830 46898 16882
rect 53230 16830 53282 16882
rect 54574 16830 54626 16882
rect 54910 16830 54962 16882
rect 55246 16830 55298 16882
rect 55470 16830 55522 16882
rect 56030 16830 56082 16882
rect 56702 16830 56754 16882
rect 57822 16830 57874 16882
rect 4622 16718 4674 16770
rect 13246 16718 13298 16770
rect 14478 16718 14530 16770
rect 31502 16718 31554 16770
rect 31838 16718 31890 16770
rect 38894 16718 38946 16770
rect 39902 16718 39954 16770
rect 41694 16718 41746 16770
rect 51662 16718 51714 16770
rect 3838 16606 3890 16658
rect 29710 16606 29762 16658
rect 29822 16606 29874 16658
rect 34638 16606 34690 16658
rect 37326 16606 37378 16658
rect 37662 16606 37714 16658
rect 38670 16606 38722 16658
rect 55694 16606 55746 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 5854 16270 5906 16322
rect 6190 16270 6242 16322
rect 6974 16270 7026 16322
rect 14478 16270 14530 16322
rect 18286 16270 18338 16322
rect 19182 16270 19234 16322
rect 22990 16270 23042 16322
rect 33294 16270 33346 16322
rect 43486 16270 43538 16322
rect 46510 16270 46562 16322
rect 55582 16270 55634 16322
rect 2494 16158 2546 16210
rect 3502 16158 3554 16210
rect 18958 16158 19010 16210
rect 22318 16158 22370 16210
rect 22654 16158 22706 16210
rect 28030 16158 28082 16210
rect 37998 16158 38050 16210
rect 38782 16158 38834 16210
rect 41134 16158 41186 16210
rect 49198 16158 49250 16210
rect 53230 16158 53282 16210
rect 55358 16158 55410 16210
rect 57934 16158 57986 16210
rect 4286 16046 4338 16098
rect 4510 16046 4562 16098
rect 5630 16046 5682 16098
rect 6638 16046 6690 16098
rect 7982 16046 8034 16098
rect 8654 16046 8706 16098
rect 10782 16046 10834 16098
rect 11006 16046 11058 16098
rect 13694 16046 13746 16098
rect 13918 16046 13970 16098
rect 16046 16046 16098 16098
rect 16942 16046 16994 16098
rect 18846 16046 18898 16098
rect 19182 16046 19234 16098
rect 20078 16046 20130 16098
rect 21422 16046 21474 16098
rect 21646 16046 21698 16098
rect 24222 16046 24274 16098
rect 25118 16046 25170 16098
rect 25790 16046 25842 16098
rect 26014 16046 26066 16098
rect 26686 16046 26738 16098
rect 27022 16046 27074 16098
rect 27582 16046 27634 16098
rect 29822 16046 29874 16098
rect 30046 16046 30098 16098
rect 35534 16046 35586 16098
rect 36206 16046 36258 16098
rect 37102 16046 37154 16098
rect 37326 16046 37378 16098
rect 39790 16046 39842 16098
rect 41582 16046 41634 16098
rect 41918 16046 41970 16098
rect 44046 16046 44098 16098
rect 45278 16046 45330 16098
rect 47854 16046 47906 16098
rect 50766 16046 50818 16098
rect 51102 16046 51154 16098
rect 55134 16046 55186 16098
rect 56142 16046 56194 16098
rect 56478 16046 56530 16098
rect 56814 16046 56866 16098
rect 1710 15934 1762 15986
rect 2046 15934 2098 15986
rect 3166 15934 3218 15986
rect 3614 15934 3666 15986
rect 3950 15934 4002 15986
rect 4734 15934 4786 15986
rect 5070 15934 5122 15986
rect 7534 15934 7586 15986
rect 11678 15934 11730 15986
rect 14030 15934 14082 15986
rect 15934 15934 15986 15986
rect 20302 15934 20354 15986
rect 20414 15934 20466 15986
rect 23326 15934 23378 15986
rect 23662 15934 23714 15986
rect 24110 15934 24162 15986
rect 25230 15934 25282 15986
rect 28142 15934 28194 15986
rect 33406 15934 33458 15986
rect 34414 15934 34466 15986
rect 34974 15934 35026 15986
rect 35310 15934 35362 15986
rect 35870 15934 35922 15986
rect 36094 15934 36146 15986
rect 41022 15934 41074 15986
rect 41806 15934 41858 15986
rect 43374 15934 43426 15986
rect 44270 15934 44322 15986
rect 44942 15934 44994 15986
rect 45502 15934 45554 15986
rect 48974 15934 49026 15986
rect 50094 15934 50146 15986
rect 50990 15934 51042 15986
rect 53566 15934 53618 15986
rect 53678 15934 53730 15986
rect 53902 15934 53954 15986
rect 54238 15934 54290 15986
rect 2830 15822 2882 15874
rect 6862 15822 6914 15874
rect 7198 15822 7250 15874
rect 7422 15822 7474 15874
rect 8318 15822 8370 15874
rect 8990 15822 9042 15874
rect 22766 15822 22818 15874
rect 23886 15822 23938 15874
rect 25454 15822 25506 15874
rect 30382 15822 30434 15874
rect 33294 15822 33346 15874
rect 34078 15822 34130 15874
rect 43486 15822 43538 15874
rect 51550 15822 51602 15874
rect 54350 15822 54402 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 50558 15654 50610 15706
rect 50662 15654 50714 15706
rect 50766 15654 50818 15706
rect 4958 15486 5010 15538
rect 13246 15486 13298 15538
rect 13582 15486 13634 15538
rect 14926 15486 14978 15538
rect 20638 15486 20690 15538
rect 31502 15486 31554 15538
rect 34638 15486 34690 15538
rect 35646 15486 35698 15538
rect 39902 15486 39954 15538
rect 49982 15486 50034 15538
rect 50542 15486 50594 15538
rect 56478 15486 56530 15538
rect 56590 15486 56642 15538
rect 6526 15374 6578 15426
rect 11006 15374 11058 15426
rect 11678 15374 11730 15426
rect 11790 15374 11842 15426
rect 13358 15374 13410 15426
rect 16494 15374 16546 15426
rect 19406 15374 19458 15426
rect 22430 15374 22482 15426
rect 26014 15374 26066 15426
rect 27918 15374 27970 15426
rect 31054 15374 31106 15426
rect 34862 15374 34914 15426
rect 37774 15374 37826 15426
rect 45950 15374 46002 15426
rect 49870 15374 49922 15426
rect 50430 15374 50482 15426
rect 54014 15374 54066 15426
rect 55918 15374 55970 15426
rect 4286 15262 4338 15314
rect 7758 15262 7810 15314
rect 10222 15262 10274 15314
rect 10558 15262 10610 15314
rect 11454 15262 11506 15314
rect 13918 15262 13970 15314
rect 15150 15262 15202 15314
rect 16046 15262 16098 15314
rect 20302 15262 20354 15314
rect 22542 15262 22594 15314
rect 23438 15262 23490 15314
rect 26350 15262 26402 15314
rect 27246 15262 27298 15314
rect 29262 15262 29314 15314
rect 29598 15262 29650 15314
rect 29710 15262 29762 15314
rect 30382 15262 30434 15314
rect 30942 15262 30994 15314
rect 31278 15262 31330 15314
rect 31614 15262 31666 15314
rect 31838 15262 31890 15314
rect 33742 15262 33794 15314
rect 34974 15262 35026 15314
rect 35982 15262 36034 15314
rect 36878 15262 36930 15314
rect 37326 15262 37378 15314
rect 37662 15262 37714 15314
rect 39454 15262 39506 15314
rect 41470 15262 41522 15314
rect 42926 15262 42978 15314
rect 43934 15262 43986 15314
rect 45726 15262 45778 15314
rect 47518 15262 47570 15314
rect 48750 15262 48802 15314
rect 49086 15262 49138 15314
rect 50206 15262 50258 15314
rect 50766 15262 50818 15314
rect 50990 15262 51042 15314
rect 52222 15262 52274 15314
rect 52782 15262 52834 15314
rect 55246 15262 55298 15314
rect 56814 15262 56866 15314
rect 57038 15262 57090 15314
rect 5518 15150 5570 15202
rect 6078 15150 6130 15202
rect 8766 15150 8818 15202
rect 11006 15150 11058 15202
rect 18846 15150 18898 15202
rect 24670 15150 24722 15202
rect 34078 15150 34130 15202
rect 34414 15150 34466 15202
rect 36542 15150 36594 15202
rect 41134 15150 41186 15202
rect 43598 15150 43650 15202
rect 44382 15150 44434 15202
rect 47294 15150 47346 15202
rect 51662 15150 51714 15202
rect 53790 15150 53842 15202
rect 1934 15038 1986 15090
rect 49422 15038 49474 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 6638 14702 6690 14754
rect 6862 14702 6914 14754
rect 17950 14702 18002 14754
rect 21310 14702 21362 14754
rect 29822 14702 29874 14754
rect 33070 14702 33122 14754
rect 39790 14702 39842 14754
rect 43822 14702 43874 14754
rect 48526 14702 48578 14754
rect 52782 14702 52834 14754
rect 55134 14702 55186 14754
rect 2270 14590 2322 14642
rect 3390 14590 3442 14642
rect 3838 14590 3890 14642
rect 4622 14590 4674 14642
rect 4958 14590 5010 14642
rect 6414 14590 6466 14642
rect 9550 14590 9602 14642
rect 10782 14590 10834 14642
rect 12910 14590 12962 14642
rect 15598 14590 15650 14642
rect 16270 14590 16322 14642
rect 17838 14590 17890 14642
rect 19294 14590 19346 14642
rect 20078 14590 20130 14642
rect 22654 14590 22706 14642
rect 23550 14590 23602 14642
rect 26910 14590 26962 14642
rect 30830 14590 30882 14642
rect 36990 14590 37042 14642
rect 42478 14590 42530 14642
rect 47406 14590 47458 14642
rect 50766 14590 50818 14642
rect 52894 14590 52946 14642
rect 55470 14590 55522 14642
rect 1822 14478 1874 14530
rect 2606 14478 2658 14530
rect 8094 14478 8146 14530
rect 8430 14478 8482 14530
rect 8766 14478 8818 14530
rect 8990 14478 9042 14530
rect 9998 14478 10050 14530
rect 15262 14478 15314 14530
rect 16382 14478 16434 14530
rect 16606 14478 16658 14530
rect 17726 14478 17778 14530
rect 19518 14478 19570 14530
rect 21646 14478 21698 14530
rect 23102 14478 23154 14530
rect 23438 14478 23490 14530
rect 25006 14478 25058 14530
rect 25902 14478 25954 14530
rect 26350 14478 26402 14530
rect 28366 14478 28418 14530
rect 28702 14478 28754 14530
rect 29710 14478 29762 14530
rect 30046 14478 30098 14530
rect 30270 14478 30322 14530
rect 31278 14478 31330 14530
rect 32398 14478 32450 14530
rect 33630 14478 33682 14530
rect 34526 14478 34578 14530
rect 34750 14478 34802 14530
rect 38334 14478 38386 14530
rect 41134 14478 41186 14530
rect 43374 14478 43426 14530
rect 43710 14478 43762 14530
rect 44046 14478 44098 14530
rect 44270 14478 44322 14530
rect 44942 14478 44994 14530
rect 45390 14478 45442 14530
rect 45726 14478 45778 14530
rect 46174 14478 46226 14530
rect 47518 14478 47570 14530
rect 49310 14478 49362 14530
rect 50430 14478 50482 14530
rect 53006 14478 53058 14530
rect 53230 14478 53282 14530
rect 54238 14478 54290 14530
rect 54462 14478 54514 14530
rect 54686 14478 54738 14530
rect 55246 14478 55298 14530
rect 55806 14478 55858 14530
rect 56142 14478 56194 14530
rect 2942 14366 2994 14418
rect 8654 14366 8706 14418
rect 10334 14366 10386 14418
rect 11230 14366 11282 14418
rect 12574 14366 12626 14418
rect 30382 14366 30434 14418
rect 33518 14366 33570 14418
rect 35422 14366 35474 14418
rect 36206 14366 36258 14418
rect 37214 14366 37266 14418
rect 38670 14366 38722 14418
rect 42030 14366 42082 14418
rect 43038 14366 43090 14418
rect 55694 14366 55746 14418
rect 56478 14366 56530 14418
rect 7310 14254 7362 14306
rect 8206 14254 8258 14306
rect 21422 14254 21474 14306
rect 28478 14254 28530 14306
rect 29486 14254 29538 14306
rect 32734 14254 32786 14306
rect 32958 14254 33010 14306
rect 33854 14254 33906 14306
rect 35086 14254 35138 14306
rect 35534 14254 35586 14306
rect 35646 14254 35698 14306
rect 36318 14254 36370 14306
rect 36542 14254 36594 14306
rect 43150 14254 43202 14306
rect 56366 14254 56418 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 50558 14086 50610 14138
rect 50662 14086 50714 14138
rect 50766 14086 50818 14138
rect 2046 13918 2098 13970
rect 2718 13918 2770 13970
rect 3166 13918 3218 13970
rect 3614 13918 3666 13970
rect 5966 13918 6018 13970
rect 6190 13918 6242 13970
rect 8766 13918 8818 13970
rect 10558 13918 10610 13970
rect 17614 13918 17666 13970
rect 24558 13918 24610 13970
rect 26350 13918 26402 13970
rect 28478 13918 28530 13970
rect 31278 13918 31330 13970
rect 32510 13918 32562 13970
rect 48302 13918 48354 13970
rect 53454 13918 53506 13970
rect 54462 13918 54514 13970
rect 55582 13918 55634 13970
rect 1710 13806 1762 13858
rect 8318 13806 8370 13858
rect 11342 13806 11394 13858
rect 13918 13806 13970 13858
rect 15262 13806 15314 13858
rect 15486 13806 15538 13858
rect 23662 13806 23714 13858
rect 23886 13806 23938 13858
rect 26574 13806 26626 13858
rect 28254 13806 28306 13858
rect 30270 13806 30322 13858
rect 43598 13806 43650 13858
rect 45838 13806 45890 13858
rect 48750 13806 48802 13858
rect 50766 13806 50818 13858
rect 52670 13806 52722 13858
rect 55358 13806 55410 13858
rect 2382 13694 2434 13746
rect 6526 13694 6578 13746
rect 8542 13694 8594 13746
rect 8878 13694 8930 13746
rect 9774 13694 9826 13746
rect 9886 13694 9938 13746
rect 10110 13694 10162 13746
rect 11678 13694 11730 13746
rect 12574 13694 12626 13746
rect 22430 13694 22482 13746
rect 22654 13694 22706 13746
rect 23326 13694 23378 13746
rect 24110 13694 24162 13746
rect 26238 13694 26290 13746
rect 27246 13694 27298 13746
rect 27694 13694 27746 13746
rect 27806 13694 27858 13746
rect 28142 13694 28194 13746
rect 30718 13694 30770 13746
rect 31166 13694 31218 13746
rect 32398 13694 32450 13746
rect 33854 13694 33906 13746
rect 34974 13694 35026 13746
rect 35646 13694 35698 13746
rect 36654 13694 36706 13746
rect 37550 13694 37602 13746
rect 37774 13694 37826 13746
rect 39566 13694 39618 13746
rect 41246 13694 41298 13746
rect 41582 13694 41634 13746
rect 44718 13694 44770 13746
rect 47294 13694 47346 13746
rect 47630 13694 47682 13746
rect 48974 13694 49026 13746
rect 49086 13694 49138 13746
rect 51998 13694 52050 13746
rect 53678 13694 53730 13746
rect 54350 13694 54402 13746
rect 54574 13694 54626 13746
rect 55022 13694 55074 13746
rect 55246 13694 55298 13746
rect 4062 13582 4114 13634
rect 6078 13582 6130 13634
rect 8766 13582 8818 13634
rect 9550 13582 9602 13634
rect 18062 13582 18114 13634
rect 22878 13582 22930 13634
rect 23550 13582 23602 13634
rect 36878 13582 36930 13634
rect 40126 13582 40178 13634
rect 41470 13582 41522 13634
rect 43150 13582 43202 13634
rect 47966 13582 48018 13634
rect 50206 13582 50258 13634
rect 15598 13470 15650 13522
rect 39790 13470 39842 13522
rect 41918 13470 41970 13522
rect 53342 13470 53394 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 42366 13134 42418 13186
rect 43486 13134 43538 13186
rect 53678 13134 53730 13186
rect 3166 13022 3218 13074
rect 6302 13022 6354 13074
rect 15038 13022 15090 13074
rect 15934 13022 15986 13074
rect 28590 13022 28642 13074
rect 29262 13022 29314 13074
rect 31390 13022 31442 13074
rect 33182 13022 33234 13074
rect 39342 13022 39394 13074
rect 41134 13022 41186 13074
rect 42478 13022 42530 13074
rect 45726 13022 45778 13074
rect 48974 13022 49026 13074
rect 51662 13022 51714 13074
rect 55470 13022 55522 13074
rect 2494 12910 2546 12962
rect 5742 12910 5794 12962
rect 6750 12910 6802 12962
rect 8990 12910 9042 12962
rect 13694 12910 13746 12962
rect 14590 12910 14642 12962
rect 15262 12910 15314 12962
rect 17390 12910 17442 12962
rect 18958 12910 19010 12962
rect 20414 12910 20466 12962
rect 21758 12910 21810 12962
rect 23326 12910 23378 12962
rect 23998 12910 24050 12962
rect 27246 12910 27298 12962
rect 27918 12910 27970 12962
rect 34190 12910 34242 12962
rect 35086 12910 35138 12962
rect 38222 12910 38274 12962
rect 40126 12910 40178 12962
rect 41694 12910 41746 12962
rect 44158 12910 44210 12962
rect 45054 12910 45106 12962
rect 46622 12910 46674 12962
rect 47518 12910 47570 12962
rect 48414 12910 48466 12962
rect 48750 12910 48802 12962
rect 50990 12910 51042 12962
rect 52110 12910 52162 12962
rect 54574 12910 54626 12962
rect 54798 12910 54850 12962
rect 1710 12798 1762 12850
rect 2046 12798 2098 12850
rect 2718 12798 2770 12850
rect 3614 12798 3666 12850
rect 9326 12798 9378 12850
rect 9998 12798 10050 12850
rect 12574 12798 12626 12850
rect 14366 12798 14418 12850
rect 16494 12798 16546 12850
rect 18062 12798 18114 12850
rect 18734 12798 18786 12850
rect 19294 12798 19346 12850
rect 19966 12798 20018 12850
rect 20078 12798 20130 12850
rect 20750 12798 20802 12850
rect 21646 12798 21698 12850
rect 22094 12798 22146 12850
rect 23102 12798 23154 12850
rect 24670 12798 24722 12850
rect 25790 12798 25842 12850
rect 25902 12798 25954 12850
rect 26126 12798 26178 12850
rect 26686 12798 26738 12850
rect 29486 12798 29538 12850
rect 31166 12798 31218 12850
rect 35310 12798 35362 12850
rect 38334 12798 38386 12850
rect 38558 12798 38610 12850
rect 39678 12798 39730 12850
rect 43934 12798 43986 12850
rect 44046 12798 44098 12850
rect 44830 12798 44882 12850
rect 49422 12798 49474 12850
rect 51102 12798 51154 12850
rect 53006 12798 53058 12850
rect 53342 12798 53394 12850
rect 7086 12686 7138 12738
rect 9662 12686 9714 12738
rect 12910 12686 12962 12738
rect 14030 12686 14082 12738
rect 19182 12686 19234 12738
rect 19742 12686 19794 12738
rect 37102 12686 37154 12738
rect 38782 12686 38834 12738
rect 42590 12686 42642 12738
rect 47630 12686 47682 12738
rect 47854 12686 47906 12738
rect 52670 12686 52722 12738
rect 53566 12686 53618 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 50558 12518 50610 12570
rect 50662 12518 50714 12570
rect 50766 12518 50818 12570
rect 2046 12350 2098 12402
rect 4958 12350 5010 12402
rect 20638 12350 20690 12402
rect 37662 12350 37714 12402
rect 40126 12350 40178 12402
rect 41806 12350 41858 12402
rect 42702 12350 42754 12402
rect 43374 12350 43426 12402
rect 43710 12350 43762 12402
rect 45054 12350 45106 12402
rect 50766 12350 50818 12402
rect 51886 12350 51938 12402
rect 6414 12238 6466 12290
rect 8430 12238 8482 12290
rect 16494 12238 16546 12290
rect 18174 12238 18226 12290
rect 18958 12238 19010 12290
rect 23326 12238 23378 12290
rect 31054 12238 31106 12290
rect 36206 12238 36258 12290
rect 36766 12238 36818 12290
rect 38334 12238 38386 12290
rect 38894 12238 38946 12290
rect 39342 12238 39394 12290
rect 39790 12238 39842 12290
rect 44382 12238 44434 12290
rect 44606 12238 44658 12290
rect 48190 12238 48242 12290
rect 51662 12238 51714 12290
rect 52110 12238 52162 12290
rect 54798 12238 54850 12290
rect 54910 12238 54962 12290
rect 1710 12126 1762 12178
rect 2494 12126 2546 12178
rect 4846 12126 4898 12178
rect 5182 12126 5234 12178
rect 5966 12126 6018 12178
rect 6190 12126 6242 12178
rect 6974 12126 7026 12178
rect 8766 12126 8818 12178
rect 9774 12126 9826 12178
rect 11342 12126 11394 12178
rect 12350 12126 12402 12178
rect 12798 12126 12850 12178
rect 15262 12126 15314 12178
rect 15934 12126 15986 12178
rect 19182 12126 19234 12178
rect 20190 12126 20242 12178
rect 22094 12126 22146 12178
rect 22542 12126 22594 12178
rect 22990 12126 23042 12178
rect 23774 12126 23826 12178
rect 24334 12126 24386 12178
rect 25454 12126 25506 12178
rect 27022 12126 27074 12178
rect 28030 12126 28082 12178
rect 28590 12126 28642 12178
rect 30382 12126 30434 12178
rect 36430 12126 36482 12178
rect 37102 12126 37154 12178
rect 37550 12126 37602 12178
rect 37886 12126 37938 12178
rect 38110 12126 38162 12178
rect 38446 12126 38498 12178
rect 40238 12126 40290 12178
rect 41358 12126 41410 12178
rect 41470 12126 41522 12178
rect 42926 12126 42978 12178
rect 44046 12126 44098 12178
rect 47070 12126 47122 12178
rect 47406 12126 47458 12178
rect 47966 12126 48018 12178
rect 49646 12126 49698 12178
rect 50206 12126 50258 12178
rect 51550 12126 51602 12178
rect 52894 12126 52946 12178
rect 53902 12126 53954 12178
rect 2942 12014 2994 12066
rect 6750 12014 6802 12066
rect 8990 12014 9042 12066
rect 10222 12014 10274 12066
rect 14590 12014 14642 12066
rect 23998 12014 24050 12066
rect 25902 12014 25954 12066
rect 27246 12014 27298 12066
rect 30606 12014 30658 12066
rect 36318 12014 36370 12066
rect 41918 12014 41970 12066
rect 47518 12014 47570 12066
rect 49534 12014 49586 12066
rect 50430 12014 50482 12066
rect 53790 12014 53842 12066
rect 7310 11902 7362 11954
rect 13022 11902 13074 11954
rect 17726 11902 17778 11954
rect 17838 11902 17890 11954
rect 18062 11902 18114 11954
rect 49086 11902 49138 11954
rect 54910 11902 54962 11954
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 6526 11566 6578 11618
rect 11454 11566 11506 11618
rect 25566 11566 25618 11618
rect 39902 11566 39954 11618
rect 48078 11566 48130 11618
rect 48638 11566 48690 11618
rect 6862 11454 6914 11506
rect 8654 11454 8706 11506
rect 14254 11454 14306 11506
rect 15374 11454 15426 11506
rect 18286 11454 18338 11506
rect 19294 11454 19346 11506
rect 23886 11454 23938 11506
rect 28030 11454 28082 11506
rect 33182 11454 33234 11506
rect 34078 11454 34130 11506
rect 34862 11454 34914 11506
rect 40238 11454 40290 11506
rect 44830 11454 44882 11506
rect 47518 11454 47570 11506
rect 52894 11454 52946 11506
rect 53678 11454 53730 11506
rect 5182 11342 5234 11394
rect 5630 11342 5682 11394
rect 5966 11342 6018 11394
rect 6302 11342 6354 11394
rect 7310 11342 7362 11394
rect 7422 11342 7474 11394
rect 7534 11342 7586 11394
rect 10222 11342 10274 11394
rect 12238 11342 12290 11394
rect 12686 11342 12738 11394
rect 13470 11342 13522 11394
rect 15710 11342 15762 11394
rect 17950 11342 18002 11394
rect 19854 11342 19906 11394
rect 20302 11342 20354 11394
rect 20750 11342 20802 11394
rect 21534 11342 21586 11394
rect 24334 11342 24386 11394
rect 25342 11342 25394 11394
rect 27022 11342 27074 11394
rect 27582 11342 27634 11394
rect 32398 11342 32450 11394
rect 32958 11342 33010 11394
rect 34414 11342 34466 11394
rect 36206 11342 36258 11394
rect 37774 11342 37826 11394
rect 38894 11342 38946 11394
rect 40350 11342 40402 11394
rect 40910 11342 40962 11394
rect 43822 11342 43874 11394
rect 44158 11342 44210 11394
rect 45502 11342 45554 11394
rect 46398 11342 46450 11394
rect 47630 11342 47682 11394
rect 49982 11342 50034 11394
rect 50766 11342 50818 11394
rect 53230 11342 53282 11394
rect 1710 11230 1762 11282
rect 2046 11230 2098 11282
rect 5742 11230 5794 11282
rect 7982 11230 8034 11282
rect 8990 11230 9042 11282
rect 12910 11230 12962 11282
rect 13694 11230 13746 11282
rect 13806 11230 13858 11282
rect 16606 11230 16658 11282
rect 18062 11230 18114 11282
rect 18734 11230 18786 11282
rect 21870 11230 21922 11282
rect 22430 11230 22482 11282
rect 28030 11230 28082 11282
rect 36542 11230 36594 11282
rect 37326 11230 37378 11282
rect 43934 11230 43986 11282
rect 46734 11230 46786 11282
rect 50878 11230 50930 11282
rect 54014 11230 54066 11282
rect 2494 11118 2546 11170
rect 17054 11118 17106 11170
rect 22094 11118 22146 11170
rect 36318 11118 36370 11170
rect 54126 11118 54178 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 50558 10950 50610 11002
rect 50662 10950 50714 11002
rect 50766 10950 50818 11002
rect 2046 10782 2098 10834
rect 5742 10782 5794 10834
rect 6862 10782 6914 10834
rect 7646 10782 7698 10834
rect 10446 10782 10498 10834
rect 23214 10782 23266 10834
rect 6078 10670 6130 10722
rect 6190 10670 6242 10722
rect 6974 10670 7026 10722
rect 28030 10726 28082 10778
rect 28142 10782 28194 10834
rect 41246 10782 41298 10834
rect 47294 10782 47346 10834
rect 47854 10782 47906 10834
rect 53230 10782 53282 10834
rect 53342 10782 53394 10834
rect 53902 10782 53954 10834
rect 54238 10782 54290 10834
rect 55022 10782 55074 10834
rect 7198 10670 7250 10722
rect 10782 10670 10834 10722
rect 11342 10670 11394 10722
rect 12462 10670 12514 10722
rect 14926 10670 14978 10722
rect 15374 10670 15426 10722
rect 30158 10670 30210 10722
rect 32510 10670 32562 10722
rect 38222 10670 38274 10722
rect 39566 10670 39618 10722
rect 42478 10670 42530 10722
rect 44718 10670 44770 10722
rect 46062 10670 46114 10722
rect 46286 10670 46338 10722
rect 49198 10670 49250 10722
rect 53790 10670 53842 10722
rect 1710 10558 1762 10610
rect 6414 10558 6466 10610
rect 6526 10558 6578 10610
rect 9662 10558 9714 10610
rect 10110 10558 10162 10610
rect 11118 10558 11170 10610
rect 11790 10558 11842 10610
rect 13582 10558 13634 10610
rect 15598 10558 15650 10610
rect 16606 10558 16658 10610
rect 17838 10558 17890 10610
rect 18510 10558 18562 10610
rect 19406 10558 19458 10610
rect 20414 10558 20466 10610
rect 20974 10558 21026 10610
rect 22654 10558 22706 10610
rect 22878 10558 22930 10610
rect 28926 10558 28978 10610
rect 29374 10558 29426 10610
rect 29822 10558 29874 10610
rect 30606 10558 30658 10610
rect 33518 10558 33570 10610
rect 34078 10558 34130 10610
rect 35086 10558 35138 10610
rect 36430 10558 36482 10610
rect 38110 10558 38162 10610
rect 39006 10558 39058 10610
rect 39790 10558 39842 10610
rect 40014 10558 40066 10610
rect 41582 10558 41634 10610
rect 44942 10558 44994 10610
rect 47070 10558 47122 10610
rect 47518 10558 47570 10610
rect 47854 10558 47906 10610
rect 48190 10558 48242 10610
rect 49870 10558 49922 10610
rect 54014 10558 54066 10610
rect 54686 10558 54738 10610
rect 2494 10446 2546 10498
rect 11566 10446 11618 10498
rect 12126 10446 12178 10498
rect 15710 10446 15762 10498
rect 30382 10446 30434 10498
rect 31950 10446 32002 10498
rect 36542 10446 36594 10498
rect 38446 10446 38498 10498
rect 43038 10446 43090 10498
rect 50094 10446 50146 10498
rect 9774 10334 9826 10386
rect 9998 10334 10050 10386
rect 20526 10334 20578 10386
rect 28142 10334 28194 10386
rect 32174 10334 32226 10386
rect 37438 10334 37490 10386
rect 39454 10334 39506 10386
rect 53454 10334 53506 10386
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 14366 9998 14418 10050
rect 23998 9998 24050 10050
rect 26910 9998 26962 10050
rect 54462 9998 54514 10050
rect 6638 9886 6690 9938
rect 7086 9886 7138 9938
rect 8430 9886 8482 9938
rect 10446 9886 10498 9938
rect 20190 9886 20242 9938
rect 28478 9886 28530 9938
rect 29262 9886 29314 9938
rect 31390 9886 31442 9938
rect 32286 9886 32338 9938
rect 32958 9886 33010 9938
rect 34862 9886 34914 9938
rect 37102 9886 37154 9938
rect 38894 9886 38946 9938
rect 43150 9886 43202 9938
rect 43934 9886 43986 9938
rect 44830 9886 44882 9938
rect 53454 9886 53506 9938
rect 6414 9774 6466 9826
rect 9998 9774 10050 9826
rect 12798 9774 12850 9826
rect 14142 9774 14194 9826
rect 15374 9774 15426 9826
rect 16270 9774 16322 9826
rect 17054 9774 17106 9826
rect 18734 9774 18786 9826
rect 19294 9774 19346 9826
rect 20526 9774 20578 9826
rect 23438 9774 23490 9826
rect 25902 9774 25954 9826
rect 26462 9774 26514 9826
rect 30718 9774 30770 9826
rect 32622 9774 32674 9826
rect 32734 9774 32786 9826
rect 33070 9774 33122 9826
rect 33406 9774 33458 9826
rect 34750 9774 34802 9826
rect 35086 9774 35138 9826
rect 35422 9774 35474 9826
rect 37550 9774 37602 9826
rect 38222 9774 38274 9826
rect 38446 9774 38498 9826
rect 39454 9774 39506 9826
rect 40798 9774 40850 9826
rect 41582 9774 41634 9826
rect 43486 9774 43538 9826
rect 45278 9774 45330 9826
rect 53118 9774 53170 9826
rect 53678 9774 53730 9826
rect 53902 9774 53954 9826
rect 54126 9774 54178 9826
rect 7646 9662 7698 9714
rect 7758 9662 7810 9714
rect 8878 9662 8930 9714
rect 12686 9662 12738 9714
rect 14478 9662 14530 9714
rect 14702 9662 14754 9714
rect 15822 9662 15874 9714
rect 16942 9662 16994 9714
rect 17838 9662 17890 9714
rect 17950 9662 18002 9714
rect 21422 9662 21474 9714
rect 21534 9662 21586 9714
rect 23662 9662 23714 9714
rect 24782 9662 24834 9714
rect 24894 9662 24946 9714
rect 26014 9662 26066 9714
rect 26238 9662 26290 9714
rect 28366 9662 28418 9714
rect 28590 9662 28642 9714
rect 29486 9662 29538 9714
rect 34526 9662 34578 9714
rect 35758 9662 35810 9714
rect 37886 9662 37938 9714
rect 40574 9662 40626 9714
rect 51998 9662 52050 9714
rect 53230 9662 53282 9714
rect 7982 9550 8034 9602
rect 12462 9550 12514 9602
rect 16382 9550 16434 9602
rect 16718 9550 16770 9602
rect 18174 9550 18226 9602
rect 21198 9550 21250 9602
rect 24110 9550 24162 9602
rect 24222 9550 24274 9602
rect 24558 9550 24610 9602
rect 32062 9550 32114 9602
rect 32286 9550 32338 9602
rect 35422 9550 35474 9602
rect 38782 9550 38834 9602
rect 39006 9550 39058 9602
rect 42030 9550 42082 9602
rect 51662 9550 51714 9602
rect 51886 9550 51938 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 50558 9382 50610 9434
rect 50662 9382 50714 9434
rect 50766 9382 50818 9434
rect 5630 9214 5682 9266
rect 7422 9214 7474 9266
rect 14254 9214 14306 9266
rect 15822 9214 15874 9266
rect 18734 9214 18786 9266
rect 19182 9214 19234 9266
rect 19518 9214 19570 9266
rect 26126 9214 26178 9266
rect 27694 9214 27746 9266
rect 30606 9214 30658 9266
rect 30830 9214 30882 9266
rect 34302 9214 34354 9266
rect 35198 9214 35250 9266
rect 36094 9214 36146 9266
rect 38334 9214 38386 9266
rect 38782 9214 38834 9266
rect 43374 9214 43426 9266
rect 44830 9214 44882 9266
rect 47070 9214 47122 9266
rect 48862 9214 48914 9266
rect 52894 9214 52946 9266
rect 2046 9102 2098 9154
rect 6190 9102 6242 9154
rect 6526 9102 6578 9154
rect 6750 9102 6802 9154
rect 7086 9102 7138 9154
rect 8654 9102 8706 9154
rect 8990 9102 9042 9154
rect 12574 9102 12626 9154
rect 15150 9102 15202 9154
rect 15486 9102 15538 9154
rect 20638 9102 20690 9154
rect 22878 9102 22930 9154
rect 27470 9102 27522 9154
rect 28254 9102 28306 9154
rect 30158 9102 30210 9154
rect 31166 9102 31218 9154
rect 31838 9102 31890 9154
rect 33182 9102 33234 9154
rect 35310 9102 35362 9154
rect 36542 9102 36594 9154
rect 37214 9102 37266 9154
rect 37662 9102 37714 9154
rect 37774 9102 37826 9154
rect 38670 9102 38722 9154
rect 39006 9102 39058 9154
rect 39230 9102 39282 9154
rect 40350 9102 40402 9154
rect 42254 9102 42306 9154
rect 43934 9102 43986 9154
rect 46062 9102 46114 9154
rect 47182 9102 47234 9154
rect 49758 9102 49810 9154
rect 50654 9102 50706 9154
rect 52110 9102 52162 9154
rect 1710 8990 1762 9042
rect 5966 8990 6018 9042
rect 7982 8990 8034 9042
rect 9550 8990 9602 9042
rect 9886 8990 9938 9042
rect 10110 8990 10162 9042
rect 13022 8990 13074 9042
rect 13806 8990 13858 9042
rect 14814 8990 14866 9042
rect 17726 8990 17778 9042
rect 17950 8990 18002 9042
rect 21646 8990 21698 9042
rect 23662 8990 23714 9042
rect 24446 8990 24498 9042
rect 25230 8990 25282 9042
rect 25454 8990 25506 9042
rect 27358 8990 27410 9042
rect 28590 8990 28642 9042
rect 29486 8990 29538 9042
rect 30494 8990 30546 9042
rect 32174 8990 32226 9042
rect 33742 8990 33794 9042
rect 33966 8990 34018 9042
rect 35646 8990 35698 9042
rect 35870 8990 35922 9042
rect 36206 8990 36258 9042
rect 36990 8990 37042 9042
rect 37886 8990 37938 9042
rect 40910 8990 40962 9042
rect 41022 8990 41074 9042
rect 41134 8990 41186 9042
rect 41358 8990 41410 9042
rect 41806 8990 41858 9042
rect 42030 8990 42082 9042
rect 42366 8990 42418 9042
rect 42814 8990 42866 9042
rect 43262 8990 43314 9042
rect 43486 8990 43538 9042
rect 44158 8990 44210 9042
rect 44718 8990 44770 9042
rect 45726 8990 45778 9042
rect 46846 8990 46898 9042
rect 48750 8990 48802 9042
rect 49982 8990 50034 9042
rect 51214 8990 51266 9042
rect 51438 8990 51490 9042
rect 51550 8990 51602 9042
rect 51774 8990 51826 9042
rect 52558 8990 52610 9042
rect 52894 8990 52946 9042
rect 2494 8878 2546 8930
rect 6974 8878 7026 8930
rect 9998 8878 10050 8930
rect 17502 8878 17554 8930
rect 20078 8878 20130 8930
rect 23998 8878 24050 8930
rect 24334 8878 24386 8930
rect 31166 8878 31218 8930
rect 25678 8766 25730 8818
rect 31390 8766 31442 8818
rect 33070 8766 33122 8818
rect 33406 8766 33458 8818
rect 39902 8766 39954 8818
rect 40014 8766 40066 8818
rect 40238 8766 40290 8818
rect 48974 8766 49026 8818
rect 49198 8766 49250 8818
rect 50430 8766 50482 8818
rect 50766 8766 50818 8818
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 7422 8430 7474 8482
rect 19182 8430 19234 8482
rect 26910 8430 26962 8482
rect 34414 8430 34466 8482
rect 39454 8430 39506 8482
rect 42590 8430 42642 8482
rect 44270 8430 44322 8482
rect 6526 8318 6578 8370
rect 7758 8318 7810 8370
rect 8206 8318 8258 8370
rect 11678 8318 11730 8370
rect 14478 8318 14530 8370
rect 15934 8318 15986 8370
rect 22094 8318 22146 8370
rect 22878 8318 22930 8370
rect 24110 8318 24162 8370
rect 29374 8318 29426 8370
rect 29710 8318 29762 8370
rect 31054 8318 31106 8370
rect 33518 8318 33570 8370
rect 36430 8318 36482 8370
rect 37102 8318 37154 8370
rect 42926 8318 42978 8370
rect 43150 8318 43202 8370
rect 44942 8318 44994 8370
rect 46174 8318 46226 8370
rect 48862 8318 48914 8370
rect 49422 8318 49474 8370
rect 52558 8318 52610 8370
rect 6750 8206 6802 8258
rect 7086 8206 7138 8258
rect 9662 8206 9714 8258
rect 11006 8206 11058 8258
rect 11230 8206 11282 8258
rect 11790 8206 11842 8258
rect 13582 8206 13634 8258
rect 13806 8206 13858 8258
rect 15262 8206 15314 8258
rect 15374 8206 15426 8258
rect 16942 8206 16994 8258
rect 17838 8206 17890 8258
rect 20078 8206 20130 8258
rect 20526 8206 20578 8258
rect 20750 8206 20802 8258
rect 21310 8206 21362 8258
rect 21534 8206 21586 8258
rect 22430 8206 22482 8258
rect 25566 8206 25618 8258
rect 27470 8206 27522 8258
rect 28366 8206 28418 8258
rect 34078 8206 34130 8258
rect 34302 8206 34354 8258
rect 35534 8206 35586 8258
rect 35758 8206 35810 8258
rect 38558 8206 38610 8258
rect 40798 8206 40850 8258
rect 41134 8206 41186 8258
rect 43486 8206 43538 8258
rect 44718 8206 44770 8258
rect 45054 8206 45106 8258
rect 45278 8206 45330 8258
rect 47294 8206 47346 8258
rect 49758 8206 49810 8258
rect 50878 8206 50930 8258
rect 53006 8206 53058 8258
rect 53230 8206 53282 8258
rect 53454 8206 53506 8258
rect 53902 8206 53954 8258
rect 54014 8206 54066 8258
rect 7646 8094 7698 8146
rect 8654 8094 8706 8146
rect 12350 8094 12402 8146
rect 12686 8094 12738 8146
rect 12798 8094 12850 8146
rect 15486 8094 15538 8146
rect 16718 8094 16770 8146
rect 23438 8094 23490 8146
rect 23550 8094 23602 8146
rect 24558 8094 24610 8146
rect 27582 8094 27634 8146
rect 29150 8094 29202 8146
rect 31166 8094 31218 8146
rect 32846 8094 32898 8146
rect 36094 8094 36146 8146
rect 37662 8094 37714 8146
rect 40462 8094 40514 8146
rect 43710 8094 43762 8146
rect 43822 8094 43874 8146
rect 48302 8094 48354 8146
rect 51438 8094 51490 8146
rect 54238 8094 54290 8146
rect 6974 7982 7026 8034
rect 13022 7982 13074 8034
rect 23214 7982 23266 8034
rect 28478 7982 28530 8034
rect 36318 7982 36370 8034
rect 40238 7982 40290 8034
rect 41694 7982 41746 8034
rect 53790 7982 53842 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 50558 7814 50610 7866
rect 50662 7814 50714 7866
rect 50766 7814 50818 7866
rect 8766 7646 8818 7698
rect 8878 7646 8930 7698
rect 8990 7646 9042 7698
rect 10446 7646 10498 7698
rect 12798 7646 12850 7698
rect 14142 7646 14194 7698
rect 14926 7646 14978 7698
rect 15374 7646 15426 7698
rect 25342 7646 25394 7698
rect 25678 7646 25730 7698
rect 26798 7646 26850 7698
rect 27582 7646 27634 7698
rect 32622 7646 32674 7698
rect 34190 7646 34242 7698
rect 34862 7646 34914 7698
rect 45726 7646 45778 7698
rect 47630 7646 47682 7698
rect 48302 7646 48354 7698
rect 49534 7646 49586 7698
rect 53342 7646 53394 7698
rect 11790 7534 11842 7586
rect 11902 7534 11954 7586
rect 12350 7534 12402 7586
rect 19406 7534 19458 7586
rect 20526 7534 20578 7586
rect 24446 7534 24498 7586
rect 26014 7534 26066 7586
rect 26574 7534 26626 7586
rect 27806 7534 27858 7586
rect 28030 7534 28082 7586
rect 30158 7534 30210 7586
rect 33070 7534 33122 7586
rect 37102 7534 37154 7586
rect 39342 7534 39394 7586
rect 47070 7534 47122 7586
rect 47182 7534 47234 7586
rect 48078 7534 48130 7586
rect 50206 7534 50258 7586
rect 50430 7534 50482 7586
rect 50542 7534 50594 7586
rect 51214 7534 51266 7586
rect 8430 7422 8482 7474
rect 9550 7422 9602 7474
rect 9998 7422 10050 7474
rect 10782 7422 10834 7474
rect 11006 7422 11058 7474
rect 11566 7422 11618 7474
rect 15262 7422 15314 7474
rect 15598 7422 15650 7474
rect 16046 7422 16098 7474
rect 16382 7422 16434 7474
rect 16606 7422 16658 7474
rect 18174 7422 18226 7474
rect 18622 7422 18674 7474
rect 19966 7422 20018 7474
rect 20302 7422 20354 7474
rect 22766 7422 22818 7474
rect 24110 7422 24162 7474
rect 26350 7422 26402 7474
rect 27022 7422 27074 7474
rect 27246 7422 27298 7474
rect 29150 7422 29202 7474
rect 30270 7422 30322 7474
rect 30606 7422 30658 7474
rect 31726 7422 31778 7474
rect 31950 7422 32002 7474
rect 33294 7422 33346 7474
rect 33742 7422 33794 7474
rect 34638 7422 34690 7474
rect 35646 7422 35698 7474
rect 35870 7422 35922 7474
rect 36206 7422 36258 7474
rect 36318 7422 36370 7474
rect 37214 7422 37266 7474
rect 37550 7422 37602 7474
rect 38558 7422 38610 7474
rect 39230 7422 39282 7474
rect 39454 7422 39506 7474
rect 39902 7422 39954 7474
rect 41134 7422 41186 7474
rect 42926 7422 42978 7474
rect 43934 7422 43986 7474
rect 46062 7422 46114 7474
rect 46846 7422 46898 7474
rect 47966 7422 48018 7474
rect 48750 7422 48802 7474
rect 48974 7422 49026 7474
rect 49310 7422 49362 7474
rect 49422 7422 49474 7474
rect 49646 7422 49698 7474
rect 52446 7422 52498 7474
rect 14254 7310 14306 7362
rect 18734 7310 18786 7362
rect 20862 7310 20914 7362
rect 22430 7310 22482 7362
rect 28926 7310 28978 7362
rect 41246 7310 41298 7362
rect 43598 7310 43650 7362
rect 44382 7310 44434 7362
rect 50990 7310 51042 7362
rect 9774 7198 9826 7250
rect 11342 7198 11394 7250
rect 12238 7198 12290 7250
rect 13918 7198 13970 7250
rect 29262 7198 29314 7250
rect 32174 7198 32226 7250
rect 33518 7198 33570 7250
rect 35310 7198 35362 7250
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 10670 6862 10722 6914
rect 15486 6862 15538 6914
rect 37438 6862 37490 6914
rect 37886 6862 37938 6914
rect 44830 6862 44882 6914
rect 52782 6862 52834 6914
rect 52894 6862 52946 6914
rect 53230 6862 53282 6914
rect 11006 6750 11058 6802
rect 11342 6750 11394 6802
rect 11678 6750 11730 6802
rect 13582 6750 13634 6802
rect 16494 6750 16546 6802
rect 18062 6750 18114 6802
rect 22206 6750 22258 6802
rect 23998 6750 24050 6802
rect 36990 6750 37042 6802
rect 37214 6750 37266 6802
rect 40350 6750 40402 6802
rect 41582 6750 41634 6802
rect 44158 6750 44210 6802
rect 44942 6750 44994 6802
rect 50766 6750 50818 6802
rect 9326 6638 9378 6690
rect 9662 6638 9714 6690
rect 12462 6638 12514 6690
rect 14030 6638 14082 6690
rect 15150 6638 15202 6690
rect 16382 6638 16434 6690
rect 17278 6638 17330 6690
rect 17950 6638 18002 6690
rect 18510 6638 18562 6690
rect 18734 6638 18786 6690
rect 22094 6638 22146 6690
rect 22542 6638 22594 6690
rect 22990 6638 23042 6690
rect 24110 6638 24162 6690
rect 24558 6638 24610 6690
rect 24782 6638 24834 6690
rect 25454 6638 25506 6690
rect 28142 6638 28194 6690
rect 31390 6638 31442 6690
rect 31838 6638 31890 6690
rect 32398 6638 32450 6690
rect 32734 6638 32786 6690
rect 34302 6638 34354 6690
rect 39006 6638 39058 6690
rect 42702 6638 42754 6690
rect 46398 6638 46450 6690
rect 47294 6638 47346 6690
rect 50654 6638 50706 6690
rect 51438 6638 51490 6690
rect 53118 6638 53170 6690
rect 9438 6526 9490 6578
rect 10894 6526 10946 6578
rect 11566 6526 11618 6578
rect 12350 6526 12402 6578
rect 19854 6526 19906 6578
rect 20190 6526 20242 6578
rect 20302 6526 20354 6578
rect 23662 6526 23714 6578
rect 27806 6526 27858 6578
rect 27918 6526 27970 6578
rect 30494 6526 30546 6578
rect 33630 6526 33682 6578
rect 34526 6526 34578 6578
rect 36094 6526 36146 6578
rect 38558 6526 38610 6578
rect 40126 6526 40178 6578
rect 40686 6526 40738 6578
rect 41022 6526 41074 6578
rect 43486 6526 43538 6578
rect 46846 6526 46898 6578
rect 49534 6526 49586 6578
rect 50318 6526 50370 6578
rect 12126 6414 12178 6466
rect 12574 6414 12626 6466
rect 17726 6414 17778 6466
rect 18174 6414 18226 6466
rect 19070 6414 19122 6466
rect 20526 6414 20578 6466
rect 31054 6414 31106 6466
rect 36430 6414 36482 6466
rect 45054 6414 45106 6466
rect 45614 6414 45666 6466
rect 47406 6414 47458 6466
rect 49982 6414 50034 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 50558 6246 50610 6298
rect 50662 6246 50714 6298
rect 50766 6246 50818 6298
rect 12238 6078 12290 6130
rect 16270 6078 16322 6130
rect 16494 6078 16546 6130
rect 35870 6078 35922 6130
rect 40014 6078 40066 6130
rect 41918 6078 41970 6130
rect 42702 6078 42754 6130
rect 46062 6078 46114 6130
rect 48862 6078 48914 6130
rect 51662 6078 51714 6130
rect 51886 6078 51938 6130
rect 52670 6078 52722 6130
rect 12350 5966 12402 6018
rect 13806 5966 13858 6018
rect 16158 5966 16210 6018
rect 34190 5966 34242 6018
rect 34974 5966 35026 6018
rect 38670 5966 38722 6018
rect 41022 5966 41074 6018
rect 49310 5966 49362 6018
rect 52110 5966 52162 6018
rect 52222 5966 52274 6018
rect 12910 5854 12962 5906
rect 13134 5854 13186 5906
rect 19070 5854 19122 5906
rect 20862 5854 20914 5906
rect 21646 5854 21698 5906
rect 29486 5854 29538 5906
rect 30046 5854 30098 5906
rect 30494 5854 30546 5906
rect 30942 5854 30994 5906
rect 31390 5854 31442 5906
rect 33070 5854 33122 5906
rect 34078 5854 34130 5906
rect 34414 5854 34466 5906
rect 36094 5854 36146 5906
rect 36542 5854 36594 5906
rect 37774 5854 37826 5906
rect 39342 5854 39394 5906
rect 40238 5854 40290 5906
rect 41358 5854 41410 5906
rect 41806 5854 41858 5906
rect 43150 5854 43202 5906
rect 43374 5854 43426 5906
rect 43598 5854 43650 5906
rect 44046 5854 44098 5906
rect 44606 5854 44658 5906
rect 45390 5854 45442 5906
rect 45950 5854 46002 5906
rect 48974 5854 49026 5906
rect 49982 5854 50034 5906
rect 50430 5854 50482 5906
rect 51326 5854 51378 5906
rect 19182 5742 19234 5794
rect 21870 5742 21922 5794
rect 29262 5742 29314 5794
rect 31838 5742 31890 5794
rect 32622 5742 32674 5794
rect 33518 5742 33570 5794
rect 39566 5742 39618 5794
rect 42478 5742 42530 5794
rect 45166 5742 45218 5794
rect 46622 5742 46674 5794
rect 47070 5742 47122 5794
rect 22318 5630 22370 5682
rect 46062 5630 46114 5682
rect 48862 5630 48914 5682
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 20750 5294 20802 5346
rect 22094 5294 22146 5346
rect 22430 5294 22482 5346
rect 31166 5294 31218 5346
rect 47518 5294 47570 5346
rect 17950 5182 18002 5234
rect 21870 5182 21922 5234
rect 30942 5182 30994 5234
rect 33518 5182 33570 5234
rect 35870 5182 35922 5234
rect 37438 5182 37490 5234
rect 40126 5182 40178 5234
rect 41806 5182 41858 5234
rect 45614 5182 45666 5234
rect 45950 5182 46002 5234
rect 46958 5182 47010 5234
rect 49534 5182 49586 5234
rect 19406 5070 19458 5122
rect 28366 5070 28418 5122
rect 29710 5070 29762 5122
rect 31614 5070 31666 5122
rect 31950 5070 32002 5122
rect 32174 5070 32226 5122
rect 32510 5070 32562 5122
rect 35758 5070 35810 5122
rect 36430 5070 36482 5122
rect 39454 5070 39506 5122
rect 40574 5070 40626 5122
rect 42254 5070 42306 5122
rect 43038 5070 43090 5122
rect 43486 5070 43538 5122
rect 43598 5070 43650 5122
rect 43934 5070 43986 5122
rect 44830 5070 44882 5122
rect 46062 5070 46114 5122
rect 47182 5070 47234 5122
rect 47742 5070 47794 5122
rect 49086 5070 49138 5122
rect 49982 5070 50034 5122
rect 18398 4958 18450 5010
rect 28590 4958 28642 5010
rect 30046 4958 30098 5010
rect 31726 4958 31778 5010
rect 44158 4958 44210 5010
rect 44270 4958 44322 5010
rect 45166 4958 45218 5010
rect 47966 4958 48018 5010
rect 48078 4958 48130 5010
rect 50318 4958 50370 5010
rect 29374 4846 29426 4898
rect 30382 4846 30434 4898
rect 35982 4846 36034 4898
rect 36206 4846 36258 4898
rect 43262 4846 43314 4898
rect 43374 4846 43426 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 50558 4678 50610 4730
rect 50662 4678 50714 4730
rect 50766 4678 50818 4730
rect 27694 4510 27746 4562
rect 32622 4510 32674 4562
rect 37774 4510 37826 4562
rect 40350 4510 40402 4562
rect 41694 4510 41746 4562
rect 43822 4510 43874 4562
rect 44718 4510 44770 4562
rect 45390 4510 45442 4562
rect 46062 4510 46114 4562
rect 31726 4398 31778 4450
rect 31950 4398 32002 4450
rect 33966 4398 34018 4450
rect 34862 4398 34914 4450
rect 36654 4398 36706 4450
rect 39006 4398 39058 4450
rect 40910 4398 40962 4450
rect 46398 4398 46450 4450
rect 28814 4286 28866 4338
rect 31614 4286 31666 4338
rect 32174 4286 32226 4338
rect 34414 4286 34466 4338
rect 36318 4286 36370 4338
rect 36990 4286 37042 4338
rect 39230 4286 39282 4338
rect 41134 4286 41186 4338
rect 42254 4286 42306 4338
rect 42478 4286 42530 4338
rect 42702 4286 42754 4338
rect 43150 4286 43202 4338
rect 43262 4286 43314 4338
rect 43486 4286 43538 4338
rect 44382 4286 44434 4338
rect 44942 4286 44994 4338
rect 45614 4286 45666 4338
rect 25342 4174 25394 4226
rect 28254 4174 28306 4226
rect 34974 4174 35026 4226
rect 42030 4174 42082 4226
rect 46846 4174 46898 4226
rect 47294 4174 47346 4226
rect 47742 4174 47794 4226
rect 48190 4174 48242 4226
rect 48862 4174 48914 4226
rect 49758 4174 49810 4226
rect 29486 4062 29538 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 40014 3726 40066 3778
rect 41134 3726 41186 3778
rect 41470 3726 41522 3778
rect 26798 3614 26850 3666
rect 29262 3614 29314 3666
rect 32398 3614 32450 3666
rect 36990 3614 37042 3666
rect 40350 3614 40402 3666
rect 40910 3614 40962 3666
rect 41806 3614 41858 3666
rect 49310 3614 49362 3666
rect 24894 3502 24946 3554
rect 27694 3502 27746 3554
rect 31166 3502 31218 3554
rect 34638 3502 34690 3554
rect 35310 3502 35362 3554
rect 36430 3502 36482 3554
rect 39118 3502 39170 3554
rect 39790 3502 39842 3554
rect 42254 3502 42306 3554
rect 43934 3502 43986 3554
rect 44494 3502 44546 3554
rect 45166 3502 45218 3554
rect 45950 3502 46002 3554
rect 46622 3502 46674 3554
rect 47630 3502 47682 3554
rect 48190 3502 48242 3554
rect 49982 3502 50034 3554
rect 22206 3390 22258 3442
rect 22430 3390 22482 3442
rect 22766 3390 22818 3442
rect 24558 3390 24610 3442
rect 28366 3390 28418 3442
rect 28702 3390 28754 3442
rect 35086 3390 35138 3442
rect 38894 3390 38946 3442
rect 42702 3390 42754 3442
rect 43038 3390 43090 3442
rect 43598 3390 43650 3442
rect 44270 3390 44322 3442
rect 44942 3390 44994 3442
rect 45614 3390 45666 3442
rect 46286 3390 46338 3442
rect 47406 3390 47458 3442
rect 48414 3390 48466 3442
rect 50318 3390 50370 3442
rect 19742 3278 19794 3330
rect 48862 3278 48914 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
rect 50558 3110 50610 3162
rect 50662 3110 50714 3162
rect 50766 3110 50818 3162
<< metal2 >>
rect 23520 59200 23632 60000
rect 24192 59200 24304 60000
rect 24864 59200 24976 60000
rect 25536 59200 25648 60000
rect 26208 59200 26320 60000
rect 26880 59200 26992 60000
rect 27552 59200 27664 60000
rect 28224 59200 28336 60000
rect 28896 59200 29008 60000
rect 29568 59200 29680 60000
rect 30240 59200 30352 60000
rect 30912 59200 31024 60000
rect 31584 59200 31696 60000
rect 32256 59200 32368 60000
rect 32928 59200 33040 60000
rect 33600 59200 33712 60000
rect 34272 59200 34384 60000
rect 34944 59200 35056 60000
rect 35616 59200 35728 60000
rect 36288 59200 36400 60000
rect 36960 59200 37072 60000
rect 37632 59200 37744 60000
rect 38304 59200 38416 60000
rect 40320 59200 40432 60000
rect 40572 59276 40964 59332
rect 19836 56476 20100 56486
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 19836 56410 20100 56420
rect 23436 56308 23492 56318
rect 23548 56308 23604 59200
rect 24220 57428 24276 59200
rect 24220 57372 24724 57428
rect 24220 56754 24276 56766
rect 24220 56702 24222 56754
rect 24274 56702 24276 56754
rect 23996 56642 24052 56654
rect 23996 56590 23998 56642
rect 24050 56590 24052 56642
rect 23436 56306 23716 56308
rect 23436 56254 23438 56306
rect 23490 56254 23716 56306
rect 23436 56252 23716 56254
rect 23436 56242 23492 56252
rect 23660 56194 23716 56252
rect 23660 56142 23662 56194
rect 23714 56142 23716 56194
rect 23660 56130 23716 56142
rect 23996 56194 24052 56590
rect 23996 56142 23998 56194
rect 24050 56142 24052 56194
rect 23996 56130 24052 56142
rect 4476 55692 4740 55702
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4476 55626 4740 55636
rect 24220 55410 24276 56702
rect 24220 55358 24222 55410
rect 24274 55358 24276 55410
rect 24220 55346 24276 55358
rect 24556 56194 24612 56206
rect 24556 56142 24558 56194
rect 24610 56142 24612 56194
rect 19836 54908 20100 54918
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 19836 54842 20100 54852
rect 4476 54124 4740 54134
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4476 54058 4740 54068
rect 22652 53842 22708 53854
rect 22652 53790 22654 53842
rect 22706 53790 22708 53842
rect 13468 53730 13524 53742
rect 13692 53732 13748 53742
rect 13468 53678 13470 53730
rect 13522 53678 13524 53730
rect 12572 53058 12628 53070
rect 12572 53006 12574 53058
rect 12626 53006 12628 53058
rect 10444 52946 10500 52958
rect 10444 52894 10446 52946
rect 10498 52894 10500 52946
rect 10332 52834 10388 52846
rect 10332 52782 10334 52834
rect 10386 52782 10388 52834
rect 4476 52556 4740 52566
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4476 52490 4740 52500
rect 10332 52274 10388 52782
rect 10332 52222 10334 52274
rect 10386 52222 10388 52274
rect 7644 52164 7700 52174
rect 7644 52162 7812 52164
rect 7644 52110 7646 52162
rect 7698 52110 7812 52162
rect 7644 52108 7812 52110
rect 7644 52098 7700 52108
rect 6972 51380 7028 51390
rect 6860 51378 7028 51380
rect 6860 51326 6974 51378
rect 7026 51326 7028 51378
rect 6860 51324 7028 51326
rect 1820 51268 1876 51278
rect 1820 51266 1988 51268
rect 1820 51214 1822 51266
rect 1874 51214 1988 51266
rect 1820 51212 1988 51214
rect 1820 51202 1876 51212
rect 1708 50484 1764 50494
rect 1932 50428 1988 51212
rect 5964 51044 6020 51054
rect 4476 50988 4740 50998
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4476 50922 4740 50932
rect 1708 50390 1764 50428
rect 1820 50372 1988 50428
rect 2940 50484 2996 50494
rect 2940 50390 2996 50428
rect 3948 50482 4004 50494
rect 3948 50430 3950 50482
rect 4002 50430 4004 50482
rect 2044 50372 2100 50382
rect 2492 50372 2548 50382
rect 1708 49364 1764 49374
rect 1484 48804 1540 48814
rect 1708 48804 1764 49308
rect 1372 44436 1428 44446
rect 1260 39396 1316 39406
rect 1260 31780 1316 39340
rect 1372 34804 1428 44380
rect 1372 34738 1428 34748
rect 1484 34468 1540 48748
rect 1596 48802 1764 48804
rect 1596 48750 1710 48802
rect 1762 48750 1764 48802
rect 1596 48748 1764 48750
rect 1596 44324 1652 48748
rect 1708 48738 1764 48748
rect 1708 48580 1764 48590
rect 1708 47458 1764 48524
rect 1708 47406 1710 47458
rect 1762 47406 1764 47458
rect 1708 47394 1764 47406
rect 1820 47012 1876 50372
rect 2044 50278 2100 50316
rect 2268 50370 2548 50372
rect 2268 50318 2494 50370
rect 2546 50318 2548 50370
rect 2268 50316 2548 50318
rect 2268 49812 2324 50316
rect 2492 50306 2548 50316
rect 3612 50372 3668 50382
rect 3612 50370 3892 50372
rect 3612 50318 3614 50370
rect 3666 50318 3892 50370
rect 3612 50316 3892 50318
rect 3612 50306 3668 50316
rect 2156 49756 2324 49812
rect 2044 49698 2100 49710
rect 2044 49646 2046 49698
rect 2098 49646 2100 49698
rect 2044 49586 2100 49646
rect 2044 49534 2046 49586
rect 2098 49534 2100 49586
rect 2044 49522 2100 49534
rect 2044 48804 2100 48814
rect 2044 48710 2100 48748
rect 2156 48580 2212 49756
rect 2492 49698 2548 49710
rect 2492 49646 2494 49698
rect 2546 49646 2548 49698
rect 2380 49586 2436 49598
rect 2380 49534 2382 49586
rect 2434 49534 2436 49586
rect 2380 49028 2436 49534
rect 2492 49252 2548 49646
rect 2828 49700 2884 49710
rect 3388 49700 3444 49710
rect 2828 49606 2884 49644
rect 3052 49698 3444 49700
rect 3052 49646 3390 49698
rect 3442 49646 3444 49698
rect 3052 49644 3444 49646
rect 2492 49186 2548 49196
rect 2940 49028 2996 49038
rect 2380 48934 2436 48972
rect 2492 49026 2996 49028
rect 2492 48974 2942 49026
rect 2994 48974 2996 49026
rect 2492 48972 2996 48974
rect 2156 48524 2324 48580
rect 2156 48356 2212 48366
rect 2156 48262 2212 48300
rect 1708 46956 1876 47012
rect 1932 48242 1988 48254
rect 1932 48190 1934 48242
rect 1986 48190 1988 48242
rect 1708 45108 1764 46956
rect 1820 46788 1876 46798
rect 1820 45890 1876 46732
rect 1820 45838 1822 45890
rect 1874 45838 1876 45890
rect 1820 45444 1876 45838
rect 1932 45780 1988 48190
rect 2044 47236 2100 47246
rect 2044 47142 2100 47180
rect 2268 46788 2324 48524
rect 2492 47684 2548 48972
rect 2940 48962 2996 48972
rect 2716 48804 2772 48814
rect 2716 48802 2996 48804
rect 2716 48750 2718 48802
rect 2770 48750 2996 48802
rect 2716 48748 2996 48750
rect 2716 48738 2772 48748
rect 2716 48468 2772 48478
rect 2604 48354 2660 48366
rect 2604 48302 2606 48354
rect 2658 48302 2660 48354
rect 2604 48244 2660 48302
rect 2716 48354 2772 48412
rect 2716 48302 2718 48354
rect 2770 48302 2772 48354
rect 2716 48290 2772 48302
rect 2604 48178 2660 48188
rect 2268 46722 2324 46732
rect 2380 47628 2548 47684
rect 2604 48018 2660 48030
rect 2604 47966 2606 48018
rect 2658 47966 2660 48018
rect 2380 46674 2436 47628
rect 2380 46622 2382 46674
rect 2434 46622 2436 46674
rect 2380 46610 2436 46622
rect 2492 47460 2548 47470
rect 2156 45780 2212 45790
rect 1932 45778 2324 45780
rect 1932 45726 2158 45778
rect 2210 45726 2324 45778
rect 1932 45724 2324 45726
rect 2156 45714 2212 45724
rect 1820 45388 1988 45444
rect 1820 45108 1876 45118
rect 1708 45106 1876 45108
rect 1708 45054 1822 45106
rect 1874 45054 1876 45106
rect 1708 45052 1876 45054
rect 1596 44258 1652 44268
rect 1708 44100 1764 44110
rect 1708 44006 1764 44044
rect 1708 41972 1764 41982
rect 1708 41300 1764 41916
rect 1596 41244 1764 41300
rect 1596 36484 1652 41244
rect 1708 41076 1764 41086
rect 1820 41076 1876 45052
rect 1932 44548 1988 45388
rect 2156 45332 2212 45342
rect 1932 44482 1988 44492
rect 2044 45218 2100 45230
rect 2044 45166 2046 45218
rect 2098 45166 2100 45218
rect 2044 44324 2100 45166
rect 1932 44268 2100 44324
rect 2156 44324 2212 45276
rect 1932 43092 1988 44268
rect 2044 44098 2100 44110
rect 2044 44046 2046 44098
rect 2098 44046 2100 44098
rect 2044 43764 2100 44046
rect 2044 43698 2100 43708
rect 1932 43036 2100 43092
rect 1932 42866 1988 42878
rect 1932 42814 1934 42866
rect 1986 42814 1988 42866
rect 1932 42420 1988 42814
rect 2044 42868 2100 43036
rect 2044 42802 2100 42812
rect 1932 42354 1988 42364
rect 2044 42082 2100 42094
rect 2044 42030 2046 42082
rect 2098 42030 2100 42082
rect 1764 41020 1876 41076
rect 1932 41298 1988 41310
rect 1932 41246 1934 41298
rect 1986 41246 1988 41298
rect 1708 41010 1764 41020
rect 1932 40404 1988 41246
rect 1932 40338 1988 40348
rect 1932 40178 1988 40190
rect 1932 40126 1934 40178
rect 1986 40126 1988 40178
rect 1932 39732 1988 40126
rect 1932 39666 1988 39676
rect 1820 39618 1876 39630
rect 1820 39566 1822 39618
rect 1874 39566 1876 39618
rect 1708 38612 1764 38622
rect 1708 36596 1764 38556
rect 1820 37826 1876 39566
rect 2044 39620 2100 42030
rect 2044 39554 2100 39564
rect 2044 39396 2100 39406
rect 2044 39302 2100 39340
rect 2156 39172 2212 44268
rect 2268 44100 2324 45724
rect 2380 44436 2436 44446
rect 2492 44436 2548 47404
rect 2604 47460 2660 47966
rect 2716 47460 2772 47470
rect 2604 47458 2772 47460
rect 2604 47406 2718 47458
rect 2770 47406 2772 47458
rect 2604 47404 2772 47406
rect 2604 46562 2660 47404
rect 2716 47394 2772 47404
rect 2604 46510 2606 46562
rect 2658 46510 2660 46562
rect 2604 46498 2660 46510
rect 2940 45556 2996 48748
rect 3052 48244 3108 49644
rect 3388 49634 3444 49644
rect 3724 49698 3780 49710
rect 3724 49646 3726 49698
rect 3778 49646 3780 49698
rect 3388 49140 3444 49150
rect 3276 49028 3332 49038
rect 3276 48934 3332 48972
rect 3164 48804 3220 48814
rect 3164 48802 3332 48804
rect 3164 48750 3166 48802
rect 3218 48750 3332 48802
rect 3164 48748 3332 48750
rect 3164 48738 3220 48748
rect 3052 47460 3108 48188
rect 3052 47394 3108 47404
rect 3276 48356 3332 48748
rect 3388 48468 3444 49084
rect 3612 48802 3668 48814
rect 3612 48750 3614 48802
rect 3666 48750 3668 48802
rect 3612 48692 3668 48750
rect 3612 48626 3668 48636
rect 3724 48468 3780 49646
rect 3836 48916 3892 50316
rect 3948 49364 4004 50430
rect 5964 50482 6020 50988
rect 6860 50596 6916 51324
rect 6972 51314 7028 51324
rect 7756 51378 7812 52108
rect 7756 51326 7758 51378
rect 7810 51326 7812 51378
rect 5964 50430 5966 50482
rect 6018 50430 6020 50482
rect 5964 50418 6020 50430
rect 6524 50594 6916 50596
rect 6524 50542 6862 50594
rect 6914 50542 6916 50594
rect 6524 50540 6916 50542
rect 4844 50372 4900 50382
rect 3948 49298 4004 49308
rect 4172 49700 4228 49710
rect 4620 49700 4676 49710
rect 4172 49698 4676 49700
rect 4172 49646 4174 49698
rect 4226 49646 4622 49698
rect 4674 49646 4676 49698
rect 4172 49644 4676 49646
rect 3948 49140 4004 49150
rect 3948 49026 4004 49084
rect 3948 48974 3950 49026
rect 4002 48974 4004 49026
rect 3948 48962 4004 48974
rect 4172 49028 4228 49644
rect 4620 49634 4676 49644
rect 4476 49420 4740 49430
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4476 49354 4740 49364
rect 4844 49140 4900 50316
rect 5628 50372 5684 50382
rect 5628 50278 5684 50316
rect 4172 48962 4228 48972
rect 4732 49028 4788 49038
rect 3836 48822 3892 48860
rect 4508 48802 4564 48814
rect 4508 48750 4510 48802
rect 4562 48750 4564 48802
rect 3388 48402 3444 48412
rect 3612 48412 3780 48468
rect 3948 48692 4004 48702
rect 3276 47348 3332 48300
rect 3500 48242 3556 48254
rect 3500 48190 3502 48242
rect 3554 48190 3556 48242
rect 3388 48132 3444 48142
rect 3388 47460 3444 48076
rect 3500 47682 3556 48190
rect 3500 47630 3502 47682
rect 3554 47630 3556 47682
rect 3500 47618 3556 47630
rect 3388 47404 3556 47460
rect 3052 47234 3108 47246
rect 3052 47182 3054 47234
rect 3106 47182 3108 47234
rect 3052 47124 3108 47182
rect 3052 47058 3108 47068
rect 3276 47234 3332 47292
rect 3276 47182 3278 47234
rect 3330 47182 3332 47234
rect 3052 46676 3108 46686
rect 3052 46002 3108 46620
rect 3052 45950 3054 46002
rect 3106 45950 3108 46002
rect 3052 45938 3108 45950
rect 3164 45892 3220 45902
rect 3164 45798 3220 45836
rect 2716 45500 2996 45556
rect 2716 44660 2772 45500
rect 2828 45332 2884 45342
rect 3276 45332 3332 47182
rect 3388 47234 3444 47246
rect 3388 47182 3390 47234
rect 3442 47182 3444 47234
rect 3388 46674 3444 47182
rect 3388 46622 3390 46674
rect 3442 46622 3444 46674
rect 3388 46610 3444 46622
rect 2828 45330 3332 45332
rect 2828 45278 2830 45330
rect 2882 45278 3332 45330
rect 2828 45276 3332 45278
rect 2828 45266 2884 45276
rect 2940 45108 2996 45118
rect 2436 44380 2548 44436
rect 2604 44604 2716 44660
rect 2380 44342 2436 44380
rect 2604 44322 2660 44604
rect 2716 44594 2772 44604
rect 2828 45106 2996 45108
rect 2828 45054 2942 45106
rect 2994 45054 2996 45106
rect 2828 45052 2996 45054
rect 2716 44436 2772 44446
rect 2828 44436 2884 45052
rect 2940 45042 2996 45052
rect 3164 45106 3220 45118
rect 3164 45054 3166 45106
rect 3218 45054 3220 45106
rect 3052 44996 3108 45006
rect 3052 44902 3108 44940
rect 2772 44380 2884 44436
rect 2716 44370 2772 44380
rect 2604 44270 2606 44322
rect 2658 44270 2660 44322
rect 2604 44258 2660 44270
rect 2940 44324 2996 44334
rect 3164 44324 3220 45054
rect 3388 45106 3444 45118
rect 3388 45054 3390 45106
rect 3442 45054 3444 45106
rect 3388 44884 3444 45054
rect 3500 45108 3556 47404
rect 3500 45042 3556 45052
rect 3388 44818 3444 44828
rect 2996 44268 3220 44324
rect 2940 44230 2996 44268
rect 2716 44210 2772 44222
rect 2716 44158 2718 44210
rect 2770 44158 2772 44210
rect 2716 44100 2772 44158
rect 2268 44044 2772 44100
rect 2828 44212 2884 44222
rect 2828 43988 2884 44156
rect 3388 44100 3444 44110
rect 3444 44044 3556 44100
rect 3388 44006 3444 44044
rect 2604 43932 2884 43988
rect 2492 42084 2548 42094
rect 2268 42082 2548 42084
rect 2268 42030 2494 42082
rect 2546 42030 2548 42082
rect 2268 42028 2548 42030
rect 2268 39284 2324 42028
rect 2492 42018 2548 42028
rect 2604 42082 2660 43932
rect 2716 43652 2772 43662
rect 2716 43538 2772 43596
rect 2716 43486 2718 43538
rect 2770 43486 2772 43538
rect 2716 43474 2772 43486
rect 3500 43538 3556 44044
rect 3500 43486 3502 43538
rect 3554 43486 3556 43538
rect 3500 43474 3556 43486
rect 3612 43876 3668 48412
rect 3948 48242 4004 48636
rect 4508 48580 4564 48750
rect 4732 48580 4788 48972
rect 4844 49026 4900 49084
rect 5740 49084 6244 49140
rect 4844 48974 4846 49026
rect 4898 48974 4900 49026
rect 4844 48962 4900 48974
rect 5180 49028 5236 49038
rect 5740 49028 5796 49084
rect 5180 49026 5796 49028
rect 5180 48974 5182 49026
rect 5234 48974 5796 49026
rect 5180 48972 5796 48974
rect 6188 49026 6244 49084
rect 6188 48974 6190 49026
rect 6242 48974 6244 49026
rect 5180 48962 5236 48972
rect 6188 48962 6244 48974
rect 6300 49028 6356 49038
rect 4956 48916 5012 48926
rect 4956 48802 5012 48860
rect 5852 48916 5908 48926
rect 6076 48916 6132 48926
rect 5852 48914 6076 48916
rect 5852 48862 5854 48914
rect 5906 48862 6076 48914
rect 5852 48860 6076 48862
rect 5852 48850 5908 48860
rect 6076 48850 6132 48860
rect 6300 48914 6356 48972
rect 6524 49026 6580 50540
rect 6860 50530 6916 50540
rect 7084 50706 7140 50718
rect 7084 50654 7086 50706
rect 7138 50654 7140 50706
rect 7084 50428 7140 50654
rect 6524 48974 6526 49026
rect 6578 48974 6580 49026
rect 6524 48962 6580 48974
rect 6636 50372 7140 50428
rect 7196 50596 7252 50606
rect 6636 49028 6692 50372
rect 6860 49700 6916 49710
rect 6860 49606 6916 49644
rect 6972 49140 7028 49150
rect 6972 49046 7028 49084
rect 6636 48962 6692 48972
rect 6748 49026 6804 49038
rect 6748 48974 6750 49026
rect 6802 48974 6804 49026
rect 6300 48862 6302 48914
rect 6354 48862 6356 48914
rect 6300 48850 6356 48862
rect 5516 48804 5572 48814
rect 4956 48750 4958 48802
rect 5010 48750 5012 48802
rect 4732 48524 4900 48580
rect 4508 48514 4564 48524
rect 3948 48190 3950 48242
rect 4002 48190 4004 48242
rect 3948 47908 4004 48190
rect 4508 48242 4564 48254
rect 4508 48190 4510 48242
rect 4562 48190 4564 48242
rect 4060 48132 4116 48142
rect 4060 48038 4116 48076
rect 4508 48132 4564 48190
rect 4508 48066 4564 48076
rect 3948 47852 4340 47908
rect 3836 47682 3892 47694
rect 3836 47630 3838 47682
rect 3890 47630 3892 47682
rect 3724 47572 3780 47582
rect 3724 47478 3780 47516
rect 3836 47460 3892 47630
rect 4284 47682 4340 47852
rect 4476 47852 4740 47862
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4476 47786 4740 47796
rect 4284 47630 4286 47682
rect 4338 47630 4340 47682
rect 4284 47618 4340 47630
rect 4620 47684 4676 47694
rect 4844 47684 4900 48524
rect 4620 47682 4900 47684
rect 4620 47630 4622 47682
rect 4674 47630 4900 47682
rect 4620 47628 4900 47630
rect 4620 47618 4676 47628
rect 4172 47572 4228 47582
rect 4060 47460 4116 47470
rect 3836 47458 4116 47460
rect 3836 47406 4062 47458
rect 4114 47406 4116 47458
rect 3836 47404 4116 47406
rect 3836 46898 3892 47404
rect 4060 47394 4116 47404
rect 4172 47236 4228 47516
rect 3836 46846 3838 46898
rect 3890 46846 3892 46898
rect 3836 46834 3892 46846
rect 4060 47180 4228 47236
rect 2940 43428 2996 43438
rect 2604 42030 2606 42082
rect 2658 42030 2660 42082
rect 2604 42018 2660 42030
rect 2716 42868 2772 42878
rect 2492 41748 2548 41758
rect 2492 41746 2660 41748
rect 2492 41694 2494 41746
rect 2546 41694 2660 41746
rect 2492 41692 2660 41694
rect 2492 41682 2548 41692
rect 2268 39228 2436 39284
rect 2156 39116 2324 39172
rect 2156 38948 2212 38958
rect 2156 38612 2212 38892
rect 2156 38546 2212 38556
rect 2268 38276 2324 39116
rect 1820 37774 1822 37826
rect 1874 37774 1876 37826
rect 1820 36708 1876 37774
rect 2156 38220 2324 38276
rect 1932 37044 1988 37054
rect 1932 36950 1988 36988
rect 1820 36652 1988 36708
rect 1708 36540 1876 36596
rect 1596 36418 1652 36428
rect 1708 36370 1764 36382
rect 1708 36318 1710 36370
rect 1762 36318 1764 36370
rect 1708 35924 1764 36318
rect 1820 36260 1876 36540
rect 1820 36166 1876 36204
rect 1932 36036 1988 36652
rect 2156 36596 2212 38220
rect 2268 38052 2324 38062
rect 2268 36706 2324 37996
rect 2380 37604 2436 39228
rect 2604 38834 2660 41692
rect 2716 38948 2772 42812
rect 2940 39842 2996 43372
rect 3052 43316 3108 43326
rect 3612 43316 3668 43820
rect 3724 46674 3780 46686
rect 3724 46622 3726 46674
rect 3778 46622 3780 46674
rect 3724 45892 3780 46622
rect 3948 46676 4004 46686
rect 3948 46582 4004 46620
rect 4060 46340 4116 47180
rect 4844 46788 4900 46798
rect 4956 46788 5012 48750
rect 5068 48802 5572 48804
rect 5068 48750 5518 48802
rect 5570 48750 5572 48802
rect 5068 48748 5572 48750
rect 5068 48242 5124 48748
rect 5516 48468 5572 48748
rect 5740 48804 5796 48814
rect 5740 48710 5796 48748
rect 6636 48804 6692 48814
rect 5516 48412 5908 48468
rect 5068 48190 5070 48242
rect 5122 48190 5124 48242
rect 5068 48178 5124 48190
rect 5628 48132 5684 48142
rect 5628 47682 5684 48076
rect 5628 47630 5630 47682
rect 5682 47630 5684 47682
rect 5628 47618 5684 47630
rect 5068 47460 5124 47470
rect 5068 47366 5124 47404
rect 5852 47346 5908 48412
rect 6412 48244 6468 48254
rect 6076 48242 6468 48244
rect 6076 48190 6414 48242
rect 6466 48190 6468 48242
rect 6076 48188 6468 48190
rect 5964 48132 6020 48142
rect 5964 48038 6020 48076
rect 5964 47684 6020 47694
rect 6076 47684 6132 48188
rect 6412 48178 6468 48188
rect 5964 47682 6132 47684
rect 5964 47630 5966 47682
rect 6018 47630 6132 47682
rect 5964 47628 6132 47630
rect 5964 47618 6020 47628
rect 5852 47294 5854 47346
rect 5906 47294 5908 47346
rect 5852 47282 5908 47294
rect 6300 47348 6356 47358
rect 6300 47254 6356 47292
rect 6636 47346 6692 48748
rect 6636 47294 6638 47346
rect 6690 47294 6692 47346
rect 6636 47282 6692 47294
rect 4844 46786 5012 46788
rect 4844 46734 4846 46786
rect 4898 46734 5012 46786
rect 4844 46732 5012 46734
rect 5404 47124 5460 47134
rect 4620 46676 4676 46686
rect 3724 43762 3780 45836
rect 3724 43710 3726 43762
rect 3778 43710 3780 43762
rect 3724 43698 3780 43710
rect 3836 46284 4116 46340
rect 4172 46674 4676 46676
rect 4172 46622 4622 46674
rect 4674 46622 4676 46674
rect 4172 46620 4676 46622
rect 3052 43222 3108 43260
rect 3388 43260 3668 43316
rect 2940 39790 2942 39842
rect 2994 39790 2996 39842
rect 2940 39778 2996 39790
rect 2716 38882 2772 38892
rect 2828 39730 2884 39742
rect 2828 39678 2830 39730
rect 2882 39678 2884 39730
rect 2604 38782 2606 38834
rect 2658 38782 2660 38834
rect 2380 37538 2436 37548
rect 2492 38722 2548 38734
rect 2492 38670 2494 38722
rect 2546 38670 2548 38722
rect 2268 36654 2270 36706
rect 2322 36654 2324 36706
rect 2268 36642 2324 36654
rect 2380 37380 2436 37390
rect 2156 36530 2212 36540
rect 2044 36372 2100 36382
rect 2268 36372 2324 36382
rect 2044 36370 2212 36372
rect 2044 36318 2046 36370
rect 2098 36318 2212 36370
rect 2044 36316 2212 36318
rect 2044 36306 2100 36316
rect 2156 36148 2212 36316
rect 2156 36082 2212 36092
rect 1708 35858 1764 35868
rect 1820 35980 1988 36036
rect 1708 35698 1764 35710
rect 1708 35646 1710 35698
rect 1762 35646 1764 35698
rect 1708 35364 1764 35646
rect 1708 35298 1764 35308
rect 1484 34402 1540 34412
rect 1708 34690 1764 34702
rect 1708 34638 1710 34690
rect 1762 34638 1764 34690
rect 1708 34132 1764 34638
rect 1708 34066 1764 34076
rect 1708 33124 1764 33134
rect 1708 33030 1764 33068
rect 1820 33012 1876 35980
rect 2044 35812 2100 35822
rect 2268 35812 2324 36316
rect 2044 35810 2324 35812
rect 2044 35758 2046 35810
rect 2098 35758 2324 35810
rect 2044 35756 2324 35758
rect 2380 35810 2436 37324
rect 2380 35758 2382 35810
rect 2434 35758 2436 35810
rect 1932 35252 1988 35262
rect 1932 34804 1988 35196
rect 2044 35140 2100 35756
rect 2380 35588 2436 35758
rect 2044 35074 2100 35084
rect 2156 35532 2436 35588
rect 2044 34804 2100 34814
rect 1932 34802 2100 34804
rect 1932 34750 2046 34802
rect 2098 34750 2100 34802
rect 1932 34748 2100 34750
rect 2044 34020 2100 34748
rect 2044 33954 2100 33964
rect 1932 33908 1988 33918
rect 1932 33814 1988 33852
rect 2044 33236 2100 33246
rect 2156 33236 2212 35532
rect 2044 33234 2212 33236
rect 2044 33182 2046 33234
rect 2098 33182 2212 33234
rect 2044 33180 2212 33182
rect 2268 35364 2324 35374
rect 2044 33170 2100 33180
rect 1820 32946 1876 32956
rect 2268 32562 2324 35308
rect 2380 35252 2436 35532
rect 2492 36148 2548 38670
rect 2604 38500 2660 38782
rect 2828 38668 2884 39678
rect 3052 39618 3108 39630
rect 3052 39566 3054 39618
rect 3106 39566 3108 39618
rect 3052 38722 3108 39566
rect 3052 38670 3054 38722
rect 3106 38670 3108 38722
rect 2828 38612 2996 38668
rect 2604 38434 2660 38444
rect 2716 38274 2772 38286
rect 2716 38222 2718 38274
rect 2770 38222 2772 38274
rect 2716 38052 2772 38222
rect 2604 37996 2716 38052
rect 2604 36706 2660 37996
rect 2716 37986 2772 37996
rect 2940 38162 2996 38612
rect 2940 38110 2942 38162
rect 2994 38110 2996 38162
rect 2604 36654 2606 36706
rect 2658 36654 2660 36706
rect 2604 36642 2660 36654
rect 2716 37604 2772 37614
rect 2716 36372 2772 37548
rect 2828 37044 2884 37054
rect 2828 36594 2884 36988
rect 2828 36542 2830 36594
rect 2882 36542 2884 36594
rect 2828 36530 2884 36542
rect 2940 36596 2996 38110
rect 3052 38050 3108 38670
rect 3388 38388 3444 43260
rect 3612 41970 3668 41982
rect 3612 41918 3614 41970
rect 3666 41918 3668 41970
rect 3612 40404 3668 41918
rect 3836 41748 3892 46284
rect 4172 46004 4228 46620
rect 4620 46610 4676 46620
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 4172 45910 4228 45948
rect 4508 45892 4564 45902
rect 4844 45892 4900 46732
rect 4508 45890 4900 45892
rect 4508 45838 4510 45890
rect 4562 45838 4900 45890
rect 4508 45836 4900 45838
rect 4956 45890 5012 45902
rect 4956 45838 4958 45890
rect 5010 45838 5012 45890
rect 4508 45780 4564 45836
rect 4956 45780 5012 45838
rect 4060 45724 4564 45780
rect 4732 45724 5012 45780
rect 3948 45218 4004 45230
rect 3948 45166 3950 45218
rect 4002 45166 4004 45218
rect 3948 44884 4004 45166
rect 4060 45106 4116 45724
rect 4620 45668 4676 45678
rect 4620 45108 4676 45612
rect 4732 45332 4788 45724
rect 4732 45266 4788 45276
rect 4844 45332 4900 45342
rect 4844 45330 5348 45332
rect 4844 45278 4846 45330
rect 4898 45278 5348 45330
rect 4844 45276 5348 45278
rect 4844 45266 4900 45276
rect 4732 45108 4788 45118
rect 4060 45054 4062 45106
rect 4114 45054 4116 45106
rect 4060 45042 4116 45054
rect 4284 45106 4788 45108
rect 4284 45054 4734 45106
rect 4786 45054 4788 45106
rect 4284 45052 4788 45054
rect 3948 44818 4004 44828
rect 4284 44434 4340 45052
rect 4732 45042 4788 45052
rect 5068 45108 5124 45118
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 4284 44382 4286 44434
rect 4338 44382 4340 44434
rect 4284 44370 4340 44382
rect 4844 44546 4900 44558
rect 4844 44494 4846 44546
rect 4898 44494 4900 44546
rect 4620 44324 4676 44334
rect 4620 44230 4676 44268
rect 4620 43652 4676 43662
rect 4620 43558 4676 43596
rect 4060 43540 4116 43550
rect 4060 43446 4116 43484
rect 4844 43540 4900 44494
rect 4844 43474 4900 43484
rect 5068 44436 5124 45052
rect 5292 45106 5348 45276
rect 5292 45054 5294 45106
rect 5346 45054 5348 45106
rect 5292 45042 5348 45054
rect 5068 43538 5124 44380
rect 5068 43486 5070 43538
rect 5122 43486 5124 43538
rect 5068 43474 5124 43486
rect 3836 41682 3892 41692
rect 3948 43428 4004 43438
rect 5404 43428 5460 47068
rect 6748 47012 6804 48974
rect 7196 48356 7252 50540
rect 7756 50482 7812 51326
rect 7980 52162 8036 52174
rect 7980 52110 7982 52162
rect 8034 52110 8036 52162
rect 7980 51268 8036 52110
rect 8092 52052 8148 52062
rect 8092 52050 8484 52052
rect 8092 51998 8094 52050
rect 8146 51998 8484 52050
rect 8092 51996 8484 51998
rect 8092 51986 8148 51996
rect 8316 51492 8372 51502
rect 8316 51398 8372 51436
rect 7980 51266 8372 51268
rect 7980 51214 7982 51266
rect 8034 51214 8372 51266
rect 7980 51212 8372 51214
rect 7980 51202 8036 51212
rect 7756 50430 7758 50482
rect 7810 50430 7812 50482
rect 7420 49924 7476 49934
rect 7644 49924 7700 49934
rect 7308 49922 7644 49924
rect 7308 49870 7422 49922
rect 7474 49870 7644 49922
rect 7308 49868 7644 49870
rect 7308 49250 7364 49868
rect 7420 49858 7476 49868
rect 7644 49858 7700 49868
rect 7308 49198 7310 49250
rect 7362 49198 7364 49250
rect 7308 49186 7364 49198
rect 7756 49700 7812 50430
rect 7756 49138 7812 49644
rect 7756 49086 7758 49138
rect 7810 49086 7812 49138
rect 7756 49074 7812 49086
rect 8204 50594 8260 50606
rect 8204 50542 8206 50594
rect 8258 50542 8260 50594
rect 8204 49924 8260 50542
rect 8204 48914 8260 49868
rect 8204 48862 8206 48914
rect 8258 48862 8260 48914
rect 8204 48850 8260 48862
rect 8316 49812 8372 51212
rect 8428 50818 8484 51996
rect 10220 51490 10276 51502
rect 10220 51438 10222 51490
rect 10274 51438 10276 51490
rect 10108 51378 10164 51390
rect 10108 51326 10110 51378
rect 10162 51326 10164 51378
rect 10108 51044 10164 51326
rect 10108 50978 10164 50988
rect 8428 50766 8430 50818
rect 8482 50766 8484 50818
rect 8428 50754 8484 50766
rect 8764 50708 8820 50718
rect 8764 50614 8820 50652
rect 9212 50596 9268 50606
rect 9212 50502 9268 50540
rect 8428 49812 8484 49822
rect 8316 49810 8484 49812
rect 8316 49758 8430 49810
rect 8482 49758 8484 49810
rect 8316 49756 8484 49758
rect 8316 48916 8372 49756
rect 8428 49746 8484 49756
rect 7196 48300 7364 48356
rect 6412 46956 6804 47012
rect 5516 46786 5572 46798
rect 5516 46734 5518 46786
rect 5570 46734 5572 46786
rect 5516 46116 5572 46734
rect 5852 46562 5908 46574
rect 5852 46510 5854 46562
rect 5906 46510 5908 46562
rect 5628 46116 5684 46126
rect 5516 46060 5628 46116
rect 5628 45778 5684 46060
rect 5628 45726 5630 45778
rect 5682 45726 5684 45778
rect 5628 45714 5684 45726
rect 5516 45106 5572 45118
rect 5516 45054 5518 45106
rect 5570 45054 5572 45106
rect 5516 43652 5572 45054
rect 5852 45108 5908 46510
rect 6300 46116 6356 46126
rect 6300 45890 6356 46060
rect 6300 45838 6302 45890
rect 6354 45838 6356 45890
rect 6300 45826 6356 45838
rect 6412 45780 6468 46956
rect 6748 46786 6804 46798
rect 6748 46734 6750 46786
rect 6802 46734 6804 46786
rect 6412 45686 6468 45724
rect 6636 45780 6692 45790
rect 6748 45780 6804 46734
rect 6860 46676 6916 46686
rect 6860 46582 6916 46620
rect 7196 45780 7252 45790
rect 6636 45778 7252 45780
rect 6636 45726 6638 45778
rect 6690 45726 7198 45778
rect 7250 45726 7252 45778
rect 6636 45724 7252 45726
rect 6636 45714 6692 45724
rect 7196 45714 7252 45724
rect 5852 45042 5908 45052
rect 5964 45666 6020 45678
rect 5964 45614 5966 45666
rect 6018 45614 6020 45666
rect 5628 44996 5684 45006
rect 5628 44546 5684 44940
rect 5964 44884 6020 45614
rect 5964 44818 6020 44828
rect 6412 45332 6468 45342
rect 5628 44494 5630 44546
rect 5682 44494 5684 44546
rect 5628 44482 5684 44494
rect 6300 44212 6356 44222
rect 6300 44118 6356 44156
rect 5740 44098 5796 44110
rect 5740 44046 5742 44098
rect 5794 44046 5796 44098
rect 5740 43652 5796 44046
rect 5852 44100 5908 44110
rect 5852 44006 5908 44044
rect 6412 44100 6468 45276
rect 7196 45108 7252 45118
rect 7196 45014 7252 45052
rect 5516 43596 5684 43652
rect 5516 43428 5572 43438
rect 5404 43426 5572 43428
rect 5404 43374 5518 43426
rect 5570 43374 5572 43426
rect 5404 43372 5572 43374
rect 3948 41970 4004 43372
rect 4284 43316 4340 43326
rect 4284 42754 4340 43260
rect 5516 43204 5572 43372
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 5516 43138 5572 43148
rect 4476 43082 4740 43092
rect 5628 42980 5684 43596
rect 5740 43586 5796 43596
rect 6076 43650 6132 43662
rect 6076 43598 6078 43650
rect 6130 43598 6132 43650
rect 5852 43428 5908 43438
rect 5852 43334 5908 43372
rect 5964 43426 6020 43438
rect 5964 43374 5966 43426
rect 6018 43374 6020 43426
rect 5628 42924 5908 42980
rect 4284 42702 4286 42754
rect 4338 42702 4340 42754
rect 4284 42690 4340 42702
rect 4620 42868 4676 42878
rect 4620 42754 4676 42812
rect 4620 42702 4622 42754
rect 4674 42702 4676 42754
rect 4620 42690 4676 42702
rect 4956 42530 5012 42542
rect 4956 42478 4958 42530
rect 5010 42478 5012 42530
rect 3948 41918 3950 41970
rect 4002 41918 4004 41970
rect 3612 40338 3668 40348
rect 3724 41076 3780 41086
rect 3388 38322 3444 38332
rect 3052 37998 3054 38050
rect 3106 37998 3108 38050
rect 3052 37986 3108 37998
rect 3724 37716 3780 41020
rect 3948 40180 4004 41918
rect 4844 41970 4900 41982
rect 4844 41918 4846 41970
rect 4898 41918 4900 41970
rect 4620 41860 4676 41870
rect 4620 41766 4676 41804
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 4284 41412 4340 41422
rect 4284 41186 4340 41356
rect 4284 41134 4286 41186
rect 4338 41134 4340 41186
rect 4284 41122 4340 41134
rect 4732 41186 4788 41198
rect 4732 41134 4734 41186
rect 4786 41134 4788 41186
rect 4732 41076 4788 41134
rect 4732 41010 4788 41020
rect 4284 40852 4340 40862
rect 4172 40740 4228 40750
rect 3948 40114 4004 40124
rect 4060 40404 4116 40414
rect 3836 39620 3892 39630
rect 3836 39618 4004 39620
rect 3836 39566 3838 39618
rect 3890 39566 4004 39618
rect 3836 39564 4004 39566
rect 3836 39554 3892 39564
rect 3724 37650 3780 37660
rect 3836 38834 3892 38846
rect 3836 38782 3838 38834
rect 3890 38782 3892 38834
rect 3836 37492 3892 38782
rect 3724 37436 3892 37492
rect 3724 37380 3780 37436
rect 3724 37314 3780 37324
rect 3276 36596 3332 36606
rect 2940 36594 3332 36596
rect 2940 36542 3278 36594
rect 3330 36542 3332 36594
rect 2940 36540 3332 36542
rect 3276 36530 3332 36540
rect 3724 36482 3780 36494
rect 3724 36430 3726 36482
rect 3778 36430 3780 36482
rect 2716 36306 2772 36316
rect 3612 36370 3668 36382
rect 3612 36318 3614 36370
rect 3666 36318 3668 36370
rect 2940 36260 2996 36270
rect 2492 35364 2548 36092
rect 2716 36148 2772 36158
rect 2604 35924 2660 35934
rect 2604 35588 2660 35868
rect 2716 35922 2772 36092
rect 2716 35870 2718 35922
rect 2770 35870 2772 35922
rect 2716 35858 2772 35870
rect 2940 35812 2996 36204
rect 2940 35810 3332 35812
rect 2940 35758 2942 35810
rect 2994 35758 3332 35810
rect 2940 35756 3332 35758
rect 2940 35746 2996 35756
rect 2828 35698 2884 35710
rect 2828 35646 2830 35698
rect 2882 35646 2884 35698
rect 2604 35532 2772 35588
rect 2604 35364 2660 35374
rect 2492 35308 2604 35364
rect 2604 35298 2660 35308
rect 2380 35196 2548 35252
rect 2492 34802 2548 35196
rect 2492 34750 2494 34802
rect 2546 34750 2548 34802
rect 2492 34738 2548 34750
rect 2604 35140 2660 35150
rect 2716 35140 2772 35532
rect 2828 35476 2884 35646
rect 3276 35476 3332 35756
rect 3612 35700 3668 36318
rect 3724 36148 3780 36430
rect 3836 36148 3892 36158
rect 3724 36092 3836 36148
rect 3836 36082 3892 36092
rect 3724 35700 3780 35710
rect 3948 35700 4004 39564
rect 4060 39618 4116 40348
rect 4060 39566 4062 39618
rect 4114 39566 4116 39618
rect 4060 39554 4116 39566
rect 4172 39058 4228 40684
rect 4284 40402 4340 40796
rect 4844 40516 4900 41918
rect 4956 41972 5012 42478
rect 5292 42196 5348 42206
rect 5292 42194 5684 42196
rect 5292 42142 5294 42194
rect 5346 42142 5684 42194
rect 5292 42140 5684 42142
rect 5292 42130 5348 42140
rect 5404 41972 5460 41982
rect 4956 41916 5124 41972
rect 4956 40964 5012 40974
rect 4956 40870 5012 40908
rect 5068 40516 5124 41916
rect 5404 41878 5460 41916
rect 5516 41970 5572 41982
rect 5516 41918 5518 41970
rect 5570 41918 5572 41970
rect 5516 41076 5572 41918
rect 5180 41020 5572 41076
rect 5180 40626 5236 41020
rect 5180 40574 5182 40626
rect 5234 40574 5236 40626
rect 5180 40562 5236 40574
rect 4844 40460 5012 40516
rect 4284 40350 4286 40402
rect 4338 40350 4340 40402
rect 4284 40338 4340 40350
rect 4620 40292 4676 40302
rect 4620 40198 4676 40236
rect 4844 40290 4900 40302
rect 4844 40238 4846 40290
rect 4898 40238 4900 40290
rect 4284 40180 4340 40190
rect 4284 39842 4340 40124
rect 4732 40180 4788 40190
rect 4844 40180 4900 40238
rect 4788 40124 4900 40180
rect 4732 40114 4788 40124
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4956 39956 5012 40460
rect 5068 40450 5124 40460
rect 4476 39946 4740 39956
rect 4844 39900 5012 39956
rect 5516 40402 5572 40414
rect 5516 40350 5518 40402
rect 5570 40350 5572 40402
rect 4284 39790 4286 39842
rect 4338 39790 4340 39842
rect 4284 39778 4340 39790
rect 4620 39844 4676 39854
rect 4844 39844 4900 39900
rect 4620 39842 4900 39844
rect 4620 39790 4622 39842
rect 4674 39790 4900 39842
rect 4620 39788 4900 39790
rect 4620 39778 4676 39788
rect 5180 39396 5236 39406
rect 5180 39394 5348 39396
rect 5180 39342 5182 39394
rect 5234 39342 5348 39394
rect 5180 39340 5348 39342
rect 5180 39330 5236 39340
rect 4172 39006 4174 39058
rect 4226 39006 4228 39058
rect 4172 38994 4228 39006
rect 4732 38946 4788 38958
rect 4732 38894 4734 38946
rect 4786 38894 4788 38946
rect 4620 38836 4676 38846
rect 4620 38742 4676 38780
rect 4508 38612 4564 38622
rect 4284 38610 4564 38612
rect 4284 38558 4510 38610
rect 4562 38558 4564 38610
rect 4284 38556 4564 38558
rect 4732 38612 4788 38894
rect 5180 38836 5236 38846
rect 4732 38556 4900 38612
rect 3612 35698 3780 35700
rect 3612 35646 3726 35698
rect 3778 35646 3780 35698
rect 3612 35644 3780 35646
rect 2828 35420 3220 35476
rect 3164 35308 3220 35420
rect 3276 35410 3332 35420
rect 3164 35252 3556 35308
rect 3500 35186 3556 35196
rect 2716 35084 3444 35140
rect 2604 34914 2660 35084
rect 3164 34916 3220 34926
rect 2604 34862 2606 34914
rect 2658 34862 2660 34914
rect 2268 32510 2270 32562
rect 2322 32510 2324 32562
rect 2268 32498 2324 32510
rect 2380 33122 2436 33134
rect 2380 33070 2382 33122
rect 2434 33070 2436 33122
rect 1260 31714 1316 31724
rect 1932 31890 1988 31902
rect 1932 31838 1934 31890
rect 1986 31838 1988 31890
rect 1932 30996 1988 31838
rect 2380 31892 2436 33070
rect 2492 33124 2548 33134
rect 2492 32676 2548 33068
rect 2604 32788 2660 34862
rect 2716 34914 3220 34916
rect 2716 34862 3166 34914
rect 3218 34862 3220 34914
rect 2716 34860 3220 34862
rect 2716 33348 2772 34860
rect 3164 34850 3220 34860
rect 2716 33234 2772 33292
rect 2716 33182 2718 33234
rect 2770 33182 2772 33234
rect 2716 33170 2772 33182
rect 3388 34804 3444 35084
rect 3612 34914 3668 34926
rect 3612 34862 3614 34914
rect 3666 34862 3668 34914
rect 3612 34804 3668 34862
rect 3388 34748 3668 34804
rect 3276 32788 3332 32798
rect 2604 32732 2772 32788
rect 2548 32620 2660 32676
rect 2492 32582 2548 32620
rect 2380 31106 2436 31836
rect 2380 31054 2382 31106
rect 2434 31054 2436 31106
rect 2380 31042 2436 31054
rect 2604 31106 2660 32620
rect 2604 31054 2606 31106
rect 2658 31054 2660 31106
rect 2604 31042 2660 31054
rect 2716 31332 2772 32732
rect 3276 32694 3332 32732
rect 1932 30930 1988 30940
rect 2268 30884 2324 30894
rect 2716 30884 2772 31276
rect 3052 31556 3108 31566
rect 3388 31556 3444 34748
rect 3724 34244 3780 35644
rect 3836 35644 4004 35700
rect 4060 38500 4116 38510
rect 4060 35700 4116 38444
rect 4172 38276 4228 38286
rect 4172 37266 4228 38220
rect 4284 38052 4340 38556
rect 4508 38546 4564 38556
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 4844 38276 4900 38556
rect 4620 38220 4900 38276
rect 4956 38500 5012 38510
rect 4284 37986 4340 37996
rect 4396 38052 4452 38062
rect 4620 38052 4676 38220
rect 4396 38050 4676 38052
rect 4396 37998 4398 38050
rect 4450 37998 4676 38050
rect 4396 37996 4676 37998
rect 4732 38052 4788 38062
rect 4172 37214 4174 37266
rect 4226 37214 4228 37266
rect 4172 37202 4228 37214
rect 4396 37044 4452 37996
rect 4732 37958 4788 37996
rect 4844 37938 4900 37950
rect 4844 37886 4846 37938
rect 4898 37886 4900 37938
rect 4844 37604 4900 37886
rect 4844 37538 4900 37548
rect 4732 37380 4788 37390
rect 4732 37286 4788 37324
rect 4844 37380 4900 37390
rect 4956 37380 5012 38444
rect 4844 37378 5012 37380
rect 4844 37326 4846 37378
rect 4898 37326 5012 37378
rect 4844 37324 5012 37326
rect 4844 37314 4900 37324
rect 4732 37044 4788 37054
rect 4452 37042 4900 37044
rect 4452 36990 4734 37042
rect 4786 36990 4900 37042
rect 4452 36988 4900 36990
rect 4396 36978 4452 36988
rect 4732 36978 4788 36988
rect 4844 36932 4900 36988
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4844 36866 4900 36876
rect 4476 36810 4740 36820
rect 4284 36540 4900 36596
rect 4284 36482 4340 36540
rect 4284 36430 4286 36482
rect 4338 36430 4340 36482
rect 4284 36418 4340 36430
rect 4620 36372 4676 36382
rect 4620 36278 4676 36316
rect 4732 36258 4788 36270
rect 4732 36206 4734 36258
rect 4786 36206 4788 36258
rect 4284 36148 4340 36158
rect 4284 35700 4340 36092
rect 4732 35700 4788 36206
rect 4060 35644 4228 35700
rect 3836 35028 3892 35644
rect 3836 34962 3892 34972
rect 4060 35252 4116 35262
rect 3724 34178 3780 34188
rect 3836 34802 3892 34814
rect 3836 34750 3838 34802
rect 3890 34750 3892 34802
rect 3500 33908 3556 33918
rect 3500 33346 3556 33852
rect 3836 33908 3892 34750
rect 4060 34692 4116 35196
rect 4172 35026 4228 35644
rect 4284 35698 4788 35700
rect 4284 35646 4286 35698
rect 4338 35646 4788 35698
rect 4284 35644 4788 35646
rect 4844 36258 4900 36540
rect 4844 36206 4846 36258
rect 4898 36206 4900 36258
rect 4284 35634 4340 35644
rect 4396 35476 4452 35514
rect 4396 35410 4452 35420
rect 4284 35364 4340 35374
rect 4284 35140 4340 35308
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4396 35140 4452 35150
rect 4284 35138 4452 35140
rect 4284 35086 4398 35138
rect 4450 35086 4452 35138
rect 4284 35084 4452 35086
rect 4396 35074 4452 35084
rect 4172 34974 4174 35026
rect 4226 34974 4228 35026
rect 4172 34962 4228 34974
rect 4508 35028 4564 35038
rect 4732 35028 4788 35038
rect 4564 35026 4788 35028
rect 4564 34974 4734 35026
rect 4786 34974 4788 35026
rect 4564 34972 4788 34974
rect 4508 34962 4564 34972
rect 4732 34962 4788 34972
rect 4060 34626 4116 34636
rect 4508 34356 4564 34366
rect 4844 34356 4900 36206
rect 4956 35922 5012 37324
rect 5180 37378 5236 38780
rect 5180 37326 5182 37378
rect 5234 37326 5236 37378
rect 5180 37314 5236 37326
rect 5292 36260 5348 39340
rect 5516 39060 5572 40350
rect 5516 38994 5572 39004
rect 5404 38722 5460 38734
rect 5404 38670 5406 38722
rect 5458 38670 5460 38722
rect 5404 38276 5460 38670
rect 5628 38724 5684 42140
rect 5740 40962 5796 42924
rect 5852 42866 5908 42924
rect 5852 42814 5854 42866
rect 5906 42814 5908 42866
rect 5852 42802 5908 42814
rect 5852 41188 5908 41198
rect 5964 41188 6020 43374
rect 5852 41186 6020 41188
rect 5852 41134 5854 41186
rect 5906 41134 6020 41186
rect 5852 41132 6020 41134
rect 5852 41122 5908 41132
rect 5740 40910 5742 40962
rect 5794 40910 5796 40962
rect 5740 40898 5796 40910
rect 6076 40626 6132 43598
rect 6300 42642 6356 42654
rect 6300 42590 6302 42642
rect 6354 42590 6356 42642
rect 6300 41972 6356 42590
rect 6300 41906 6356 41916
rect 6188 41860 6244 41870
rect 6188 41300 6244 41804
rect 6188 41186 6244 41244
rect 6188 41134 6190 41186
rect 6242 41134 6244 41186
rect 6188 41122 6244 41134
rect 6076 40574 6078 40626
rect 6130 40574 6132 40626
rect 5852 40514 5908 40526
rect 5852 40462 5854 40514
rect 5906 40462 5908 40514
rect 5852 40068 5908 40462
rect 6076 40404 6132 40574
rect 6300 40516 6356 40526
rect 6300 40422 6356 40460
rect 6076 40338 6132 40348
rect 6412 40402 6468 44044
rect 6636 44884 6692 44894
rect 6636 44100 6692 44828
rect 6860 44324 6916 44334
rect 6860 44230 6916 44268
rect 7196 44210 7252 44222
rect 7196 44158 7198 44210
rect 7250 44158 7252 44210
rect 7084 44100 7140 44110
rect 6636 44098 7140 44100
rect 6636 44046 6638 44098
rect 6690 44046 7086 44098
rect 7138 44046 7140 44098
rect 6636 44044 7140 44046
rect 6636 44034 6692 44044
rect 7084 44034 7140 44044
rect 7196 44100 7252 44158
rect 7196 44034 7252 44044
rect 7308 43876 7364 48300
rect 7532 48242 7588 48254
rect 7756 48244 7812 48254
rect 7532 48190 7534 48242
rect 7586 48190 7588 48242
rect 7532 48132 7588 48190
rect 7532 47572 7588 48076
rect 7532 47506 7588 47516
rect 7644 48242 7812 48244
rect 7644 48190 7758 48242
rect 7810 48190 7812 48242
rect 7644 48188 7812 48190
rect 7644 47458 7700 48188
rect 7756 48178 7812 48188
rect 8316 48130 8372 48860
rect 8988 49698 9044 49710
rect 8988 49646 8990 49698
rect 9042 49646 9044 49698
rect 8988 48244 9044 49646
rect 9212 49026 9268 49038
rect 9212 48974 9214 49026
rect 9266 48974 9268 49026
rect 9212 48916 9268 48974
rect 9212 48850 9268 48860
rect 8988 48178 9044 48188
rect 9100 48356 9156 48366
rect 8316 48078 8318 48130
rect 8370 48078 8372 48130
rect 8316 48066 8372 48078
rect 7644 47406 7646 47458
rect 7698 47406 7700 47458
rect 7644 46676 7700 47406
rect 7644 45890 7700 46620
rect 7644 45838 7646 45890
rect 7698 45838 7700 45890
rect 7644 44994 7700 45838
rect 7980 47572 8036 47582
rect 7980 46674 8036 47516
rect 8316 47572 8372 47582
rect 8316 47478 8372 47516
rect 7980 46622 7982 46674
rect 8034 46622 8036 46674
rect 7980 45892 8036 46622
rect 8876 47348 8932 47358
rect 8540 46116 8596 46126
rect 8428 45892 8484 45902
rect 7980 45890 8484 45892
rect 7980 45838 8430 45890
rect 8482 45838 8484 45890
rect 7980 45836 8484 45838
rect 8428 45826 8484 45836
rect 8540 45106 8596 46060
rect 8652 45780 8708 45790
rect 8708 45724 8820 45780
rect 8652 45714 8708 45724
rect 8540 45054 8542 45106
rect 8594 45054 8596 45106
rect 8540 45042 8596 45054
rect 7644 44942 7646 44994
rect 7698 44942 7700 44994
rect 7644 44930 7700 44942
rect 7644 44436 7700 44446
rect 7644 44342 7700 44380
rect 7084 43820 7364 43876
rect 7532 44324 7588 44334
rect 6748 43540 6804 43550
rect 6748 43426 6804 43484
rect 6748 43374 6750 43426
rect 6802 43374 6804 43426
rect 6748 43362 6804 43374
rect 6860 43538 6916 43550
rect 6860 43486 6862 43538
rect 6914 43486 6916 43538
rect 6636 42082 6692 42094
rect 6636 42030 6638 42082
rect 6690 42030 6692 42082
rect 6636 41972 6692 42030
rect 6636 40628 6692 41916
rect 6860 42084 6916 43486
rect 6860 41970 6916 42028
rect 6860 41918 6862 41970
rect 6914 41918 6916 41970
rect 6860 41906 6916 41918
rect 6636 40562 6692 40572
rect 6748 41188 6804 41198
rect 6748 41074 6804 41132
rect 6748 41022 6750 41074
rect 6802 41022 6804 41074
rect 6412 40350 6414 40402
rect 6466 40350 6468 40402
rect 6412 40292 6468 40350
rect 5852 40002 5908 40012
rect 6188 40236 6468 40292
rect 6636 40402 6692 40414
rect 6636 40350 6638 40402
rect 6690 40350 6692 40402
rect 5964 39620 6020 39630
rect 5740 38724 5796 38762
rect 5628 38722 5796 38724
rect 5628 38670 5742 38722
rect 5794 38670 5796 38722
rect 5628 38668 5796 38670
rect 5404 38210 5460 38220
rect 5516 38612 5796 38668
rect 5516 37490 5572 38612
rect 5740 38164 5796 38174
rect 5740 38050 5796 38108
rect 5740 37998 5742 38050
rect 5794 37998 5796 38050
rect 5740 37986 5796 37998
rect 5516 37438 5518 37490
rect 5570 37438 5572 37490
rect 5516 37426 5572 37438
rect 5740 37604 5796 37614
rect 5516 37266 5572 37278
rect 5516 37214 5518 37266
rect 5570 37214 5572 37266
rect 5516 37044 5572 37214
rect 5740 37268 5796 37548
rect 5740 37174 5796 37212
rect 5516 36978 5572 36988
rect 5628 36260 5684 36270
rect 5292 36258 5684 36260
rect 5292 36206 5630 36258
rect 5682 36206 5684 36258
rect 5292 36204 5684 36206
rect 4956 35870 4958 35922
rect 5010 35870 5012 35922
rect 4956 35858 5012 35870
rect 5292 35924 5348 35934
rect 5292 35830 5348 35868
rect 5404 35812 5460 35822
rect 5516 35812 5572 36204
rect 5628 36194 5684 36204
rect 5964 35924 6020 39564
rect 6076 38724 6132 38734
rect 6188 38724 6244 40236
rect 6636 39844 6692 40350
rect 6412 39788 6692 39844
rect 6412 39508 6468 39788
rect 6748 39732 6804 41022
rect 6860 40740 6916 40750
rect 6860 40626 6916 40684
rect 6860 40574 6862 40626
rect 6914 40574 6916 40626
rect 6860 40562 6916 40574
rect 6636 39676 6804 39732
rect 6972 40402 7028 40414
rect 6972 40350 6974 40402
rect 7026 40350 7028 40402
rect 6636 39620 6692 39676
rect 6300 39506 6468 39508
rect 6300 39454 6414 39506
rect 6466 39454 6468 39506
rect 6300 39452 6468 39454
rect 6300 38946 6356 39452
rect 6412 39442 6468 39452
rect 6524 39618 6692 39620
rect 6524 39566 6638 39618
rect 6690 39566 6692 39618
rect 6524 39564 6692 39566
rect 6300 38894 6302 38946
rect 6354 38894 6356 38946
rect 6300 38882 6356 38894
rect 6132 38668 6244 38724
rect 6076 38658 6132 38668
rect 6524 38274 6580 39564
rect 6636 39554 6692 39564
rect 6524 38222 6526 38274
rect 6578 38222 6580 38274
rect 6524 38210 6580 38222
rect 6300 38050 6356 38062
rect 6300 37998 6302 38050
rect 6354 37998 6356 38050
rect 6300 37156 6356 37998
rect 6748 38052 6804 38062
rect 6300 37090 6356 37100
rect 6636 37378 6692 37390
rect 6636 37326 6638 37378
rect 6690 37326 6692 37378
rect 6524 36932 6580 36942
rect 6524 36594 6580 36876
rect 6636 36708 6692 37326
rect 6636 36642 6692 36652
rect 6748 36706 6804 37996
rect 6860 37266 6916 37278
rect 6860 37214 6862 37266
rect 6914 37214 6916 37266
rect 6860 37156 6916 37214
rect 6860 37090 6916 37100
rect 6748 36654 6750 36706
rect 6802 36654 6804 36706
rect 6748 36642 6804 36654
rect 6524 36542 6526 36594
rect 6578 36542 6580 36594
rect 6524 36530 6580 36542
rect 5964 35858 6020 35868
rect 6188 36482 6244 36494
rect 6188 36430 6190 36482
rect 6242 36430 6244 36482
rect 5460 35756 5572 35812
rect 5404 35746 5460 35756
rect 5628 35700 5684 35710
rect 5684 35644 5908 35700
rect 5628 35606 5684 35644
rect 4508 34354 4900 34356
rect 4508 34302 4510 34354
rect 4562 34302 4900 34354
rect 4508 34300 4900 34302
rect 4956 35588 5012 35598
rect 4956 34356 5012 35532
rect 4508 34290 4564 34300
rect 4956 34290 5012 34300
rect 5068 34916 5124 34926
rect 5852 34916 5908 35644
rect 6076 35698 6132 35710
rect 6076 35646 6078 35698
rect 6130 35646 6132 35698
rect 6076 35364 6132 35646
rect 6076 35298 6132 35308
rect 6188 34916 6244 36430
rect 6524 36260 6580 36270
rect 6524 35698 6580 36204
rect 6972 36148 7028 40350
rect 7084 38668 7140 43820
rect 7532 43650 7588 44268
rect 8428 44322 8484 44334
rect 8428 44270 8430 44322
rect 8482 44270 8484 44322
rect 8428 44212 8484 44270
rect 8484 44156 8708 44212
rect 8428 44146 8484 44156
rect 7532 43598 7534 43650
rect 7586 43598 7588 43650
rect 7532 43586 7588 43598
rect 7308 43540 7364 43550
rect 7308 42756 7364 43484
rect 8092 43426 8148 43438
rect 8092 43374 8094 43426
rect 8146 43374 8148 43426
rect 8092 43316 8148 43374
rect 8092 43250 8148 43260
rect 7308 42754 7700 42756
rect 7308 42702 7310 42754
rect 7362 42702 7700 42754
rect 7308 42700 7700 42702
rect 7308 42690 7364 42700
rect 7644 41970 7700 42700
rect 8540 42642 8596 42654
rect 8540 42590 8542 42642
rect 8594 42590 8596 42642
rect 7644 41918 7646 41970
rect 7698 41918 7700 41970
rect 7644 41906 7700 41918
rect 8316 42082 8372 42094
rect 8316 42030 8318 42082
rect 8370 42030 8372 42082
rect 8316 41972 8372 42030
rect 8316 41906 8372 41916
rect 8540 41748 8596 42590
rect 8652 42194 8708 44156
rect 8652 42142 8654 42194
rect 8706 42142 8708 42194
rect 8652 42130 8708 42142
rect 8652 41748 8708 41758
rect 8540 41692 8652 41748
rect 8652 41682 8708 41692
rect 8092 41636 8148 41646
rect 7196 41300 7252 41310
rect 7252 41244 7364 41300
rect 7196 41206 7252 41244
rect 7196 40628 7252 40638
rect 7196 40534 7252 40572
rect 7308 39620 7364 41244
rect 8092 41298 8148 41580
rect 8092 41246 8094 41298
rect 8146 41246 8148 41298
rect 8092 41234 8148 41246
rect 8316 41410 8372 41422
rect 8316 41358 8318 41410
rect 8370 41358 8372 41410
rect 7420 41188 7476 41198
rect 7420 41094 7476 41132
rect 7420 40628 7476 40638
rect 7420 40534 7476 40572
rect 7532 40404 7588 40414
rect 7532 40310 7588 40348
rect 8316 40404 8372 41358
rect 8540 41076 8596 41086
rect 8540 40982 8596 41020
rect 8764 40852 8820 45724
rect 8876 44434 8932 47292
rect 8988 46450 9044 46462
rect 8988 46398 8990 46450
rect 9042 46398 9044 46450
rect 8988 45220 9044 46398
rect 8988 45154 9044 45164
rect 8988 44996 9044 45006
rect 9100 44996 9156 48300
rect 9884 48356 9940 48366
rect 10220 48356 10276 51438
rect 10332 51492 10388 52222
rect 10444 52162 10500 52894
rect 12460 52948 12516 52958
rect 11116 52836 11172 52846
rect 11116 52834 11284 52836
rect 11116 52782 11118 52834
rect 11170 52782 11284 52834
rect 11116 52780 11284 52782
rect 11116 52770 11172 52780
rect 11004 52388 11060 52398
rect 11004 52294 11060 52332
rect 10444 52110 10446 52162
rect 10498 52110 10500 52162
rect 10444 51604 10500 52110
rect 11116 52164 11172 52174
rect 10892 51604 10948 51614
rect 10444 51602 10948 51604
rect 10444 51550 10446 51602
rect 10498 51550 10894 51602
rect 10946 51550 10948 51602
rect 10444 51548 10948 51550
rect 10444 51538 10500 51548
rect 10892 51538 10948 51548
rect 11116 51602 11172 52108
rect 11116 51550 11118 51602
rect 11170 51550 11172 51602
rect 11116 51538 11172 51550
rect 10332 51426 10388 51436
rect 10780 51380 10836 51390
rect 10780 51286 10836 51324
rect 11228 51380 11284 52780
rect 12460 52388 12516 52892
rect 11788 52164 11844 52174
rect 11788 52070 11844 52108
rect 12348 52164 12404 52174
rect 12348 52070 12404 52108
rect 12236 52052 12292 52062
rect 11228 51314 11284 51324
rect 11788 51378 11844 51390
rect 11788 51326 11790 51378
rect 11842 51326 11844 51378
rect 11788 50594 11844 51326
rect 11788 50542 11790 50594
rect 11842 50542 11844 50594
rect 11340 49980 11732 50036
rect 11340 49922 11396 49980
rect 11340 49870 11342 49922
rect 11394 49870 11396 49922
rect 11340 49858 11396 49870
rect 11676 49924 11732 49980
rect 11452 49810 11508 49822
rect 11452 49758 11454 49810
rect 11506 49758 11508 49810
rect 11228 49026 11284 49038
rect 11228 48974 11230 49026
rect 11282 48974 11284 49026
rect 10556 48804 10612 48814
rect 10556 48710 10612 48748
rect 10332 48356 10388 48366
rect 10220 48354 10388 48356
rect 10220 48302 10334 48354
rect 10386 48302 10388 48354
rect 10220 48300 10388 48302
rect 9884 48262 9940 48300
rect 9772 48242 9828 48254
rect 9772 48190 9774 48242
rect 9826 48190 9828 48242
rect 9772 47572 9828 48190
rect 9772 47458 9828 47516
rect 9772 47406 9774 47458
rect 9826 47406 9828 47458
rect 9772 47394 9828 47406
rect 9548 47348 9604 47358
rect 9548 47254 9604 47292
rect 9660 47346 9716 47358
rect 9660 47294 9662 47346
rect 9714 47294 9716 47346
rect 9212 47236 9268 47246
rect 9212 45108 9268 47180
rect 9660 46116 9716 47294
rect 10332 47348 10388 48300
rect 11004 48130 11060 48142
rect 11004 48078 11006 48130
rect 11058 48078 11060 48130
rect 11004 47458 11060 48078
rect 11004 47406 11006 47458
rect 11058 47406 11060 47458
rect 11004 47394 11060 47406
rect 10220 47234 10276 47246
rect 10220 47182 10222 47234
rect 10274 47182 10276 47234
rect 9660 46050 9716 46060
rect 10108 46674 10164 46686
rect 10108 46622 10110 46674
rect 10162 46622 10164 46674
rect 9772 45668 9828 45678
rect 9772 45574 9828 45612
rect 9772 45332 9828 45342
rect 9828 45276 9940 45332
rect 9772 45238 9828 45276
rect 9212 45042 9268 45052
rect 8988 44994 9156 44996
rect 8988 44942 8990 44994
rect 9042 44942 9156 44994
rect 8988 44940 9156 44942
rect 9660 44996 9716 45006
rect 8988 44930 9044 44940
rect 9660 44902 9716 44940
rect 9884 44548 9940 45276
rect 9996 44884 10052 44894
rect 9996 44790 10052 44828
rect 9996 44548 10052 44558
rect 9884 44546 10052 44548
rect 9884 44494 9998 44546
rect 10050 44494 10052 44546
rect 9884 44492 10052 44494
rect 9996 44482 10052 44492
rect 8876 44382 8878 44434
rect 8930 44382 8932 44434
rect 8876 44370 8932 44382
rect 9548 44324 9604 44334
rect 10108 44324 10164 46622
rect 10220 46676 10276 47182
rect 10332 46786 10388 47292
rect 10780 47346 10836 47358
rect 10780 47294 10782 47346
rect 10834 47294 10836 47346
rect 10556 46788 10612 46798
rect 10332 46734 10334 46786
rect 10386 46734 10388 46786
rect 10332 46722 10388 46734
rect 10444 46786 10612 46788
rect 10444 46734 10558 46786
rect 10610 46734 10612 46786
rect 10444 46732 10612 46734
rect 10220 46610 10276 46620
rect 9604 44268 10164 44324
rect 10444 45444 10500 46732
rect 10556 46722 10612 46732
rect 9548 44230 9604 44268
rect 9324 44210 9380 44222
rect 9324 44158 9326 44210
rect 9378 44158 9380 44210
rect 9324 43876 9380 44158
rect 9436 44212 9492 44222
rect 9436 43988 9492 44156
rect 9436 43932 9716 43988
rect 9212 43820 9604 43876
rect 8876 41970 8932 41982
rect 8876 41918 8878 41970
rect 8930 41918 8932 41970
rect 8876 41410 8932 41918
rect 8876 41358 8878 41410
rect 8930 41358 8932 41410
rect 8876 41346 8932 41358
rect 8988 41412 9044 41422
rect 8540 40796 8820 40852
rect 8540 40626 8596 40796
rect 8540 40574 8542 40626
rect 8594 40574 8596 40626
rect 8540 40562 8596 40574
rect 8372 40348 8484 40404
rect 8316 40310 8372 40348
rect 7420 39620 7476 39630
rect 7308 39618 7476 39620
rect 7308 39566 7422 39618
rect 7474 39566 7476 39618
rect 7308 39564 7476 39566
rect 7308 38834 7364 39564
rect 7420 39554 7476 39564
rect 8092 39508 8148 39518
rect 8092 39414 8148 39452
rect 8316 38948 8372 38958
rect 8316 38854 8372 38892
rect 7308 38782 7310 38834
rect 7362 38782 7364 38834
rect 7308 38770 7364 38782
rect 7084 38612 7364 38668
rect 7084 38050 7140 38062
rect 7084 37998 7086 38050
rect 7138 37998 7140 38050
rect 7084 36706 7140 37998
rect 7084 36654 7086 36706
rect 7138 36654 7140 36706
rect 7084 36642 7140 36654
rect 6972 36082 7028 36092
rect 7196 35924 7252 35934
rect 6860 35812 6916 35822
rect 6860 35810 7028 35812
rect 6860 35758 6862 35810
rect 6914 35758 7028 35810
rect 6860 35756 7028 35758
rect 6860 35746 6916 35756
rect 6524 35646 6526 35698
rect 6578 35646 6580 35698
rect 6524 35588 6580 35646
rect 6524 35522 6580 35532
rect 6860 35476 6916 35486
rect 6860 35026 6916 35420
rect 6860 34974 6862 35026
rect 6914 34974 6916 35026
rect 6860 34962 6916 34974
rect 5068 34242 5124 34860
rect 5068 34190 5070 34242
rect 5122 34190 5124 34242
rect 5068 34178 5124 34190
rect 5516 34914 5908 34916
rect 5516 34862 5854 34914
rect 5906 34862 5908 34914
rect 5516 34860 5908 34862
rect 3836 33842 3892 33852
rect 3948 34132 4004 34142
rect 3724 33572 3780 33582
rect 3612 33516 3724 33572
rect 3612 33458 3668 33516
rect 3724 33506 3780 33516
rect 3612 33406 3614 33458
rect 3666 33406 3668 33458
rect 3612 33394 3668 33406
rect 3836 33348 3892 33358
rect 3500 33294 3502 33346
rect 3554 33294 3556 33346
rect 3500 33282 3556 33294
rect 3724 33346 3892 33348
rect 3724 33294 3838 33346
rect 3890 33294 3892 33346
rect 3724 33292 3892 33294
rect 3612 31668 3668 31678
rect 3500 31556 3556 31566
rect 3388 31500 3500 31556
rect 3052 30994 3108 31500
rect 3500 31490 3556 31500
rect 3500 30996 3556 31006
rect 3052 30942 3054 30994
rect 3106 30942 3108 30994
rect 3052 30930 3108 30942
rect 3388 30994 3556 30996
rect 3388 30942 3502 30994
rect 3554 30942 3556 30994
rect 3388 30940 3556 30942
rect 2268 30882 2772 30884
rect 2268 30830 2270 30882
rect 2322 30830 2772 30882
rect 2268 30828 2772 30830
rect 3276 30884 3332 30894
rect 2268 30818 2324 30828
rect 3276 30790 3332 30828
rect 2268 30660 2324 30670
rect 1708 30324 1764 30334
rect 1596 28868 1652 28878
rect 1260 28196 1316 28206
rect 1260 11284 1316 28140
rect 1484 22820 1540 22830
rect 1372 22764 1484 22820
rect 1372 18228 1428 22764
rect 1484 22754 1540 22764
rect 1484 22372 1540 22382
rect 1484 18452 1540 22316
rect 1484 18386 1540 18396
rect 1372 18162 1428 18172
rect 1596 12628 1652 28812
rect 1708 27076 1764 30268
rect 1932 29204 1988 29214
rect 1932 29110 1988 29148
rect 2268 28754 2324 30604
rect 3388 30660 3444 30940
rect 3500 30930 3556 30940
rect 3388 30594 3444 30604
rect 2492 30098 2548 30110
rect 2492 30046 2494 30098
rect 2546 30046 2548 30098
rect 2492 29652 2548 30046
rect 2492 29586 2548 29596
rect 2828 29764 2884 29774
rect 2268 28702 2270 28754
rect 2322 28702 2324 28754
rect 2268 28690 2324 28702
rect 2716 29428 2772 29438
rect 1932 28642 1988 28654
rect 1932 28590 1934 28642
rect 1986 28590 1988 28642
rect 1932 28308 1988 28590
rect 1932 28242 1988 28252
rect 2044 28644 2100 28654
rect 2044 28082 2100 28588
rect 2716 28644 2772 29372
rect 2716 28550 2772 28588
rect 2044 28030 2046 28082
rect 2098 28030 2100 28082
rect 2044 28018 2100 28030
rect 2716 28084 2772 28094
rect 2828 28084 2884 29708
rect 3052 28642 3108 28654
rect 3052 28590 3054 28642
rect 3106 28590 3108 28642
rect 2716 28082 2884 28084
rect 2716 28030 2718 28082
rect 2770 28030 2884 28082
rect 2716 28028 2884 28030
rect 2940 28420 2996 28430
rect 2716 28018 2772 28028
rect 1820 27860 1876 27870
rect 1820 27766 1876 27804
rect 2380 27858 2436 27870
rect 2380 27806 2382 27858
rect 2434 27806 2436 27858
rect 2380 27636 2436 27806
rect 2380 27570 2436 27580
rect 1708 26982 1764 27020
rect 2044 27188 2100 27198
rect 2044 26962 2100 27132
rect 2044 26910 2046 26962
rect 2098 26910 2100 26962
rect 2044 26898 2100 26910
rect 2492 27074 2548 27086
rect 2492 27022 2494 27074
rect 2546 27022 2548 27074
rect 2492 26852 2548 27022
rect 2716 26964 2772 26974
rect 2940 26964 2996 28364
rect 3052 28308 3108 28590
rect 3388 28644 3444 28654
rect 3388 28418 3444 28588
rect 3388 28366 3390 28418
rect 3442 28366 3444 28418
rect 3388 28354 3444 28366
rect 3052 28242 3108 28252
rect 3612 28082 3668 31612
rect 3724 31108 3780 33292
rect 3836 33282 3892 33292
rect 3724 30882 3780 31052
rect 3724 30830 3726 30882
rect 3778 30830 3780 30882
rect 3724 30818 3780 30830
rect 3948 32562 4004 34076
rect 4284 34130 4340 34142
rect 4284 34078 4286 34130
rect 4338 34078 4340 34130
rect 4284 33908 4340 34078
rect 4732 34132 4788 34142
rect 4732 34038 4788 34076
rect 5292 34130 5348 34142
rect 5292 34078 5294 34130
rect 5346 34078 5348 34130
rect 4284 33842 4340 33852
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 5292 33572 5348 34078
rect 5516 34130 5572 34860
rect 5852 34850 5908 34860
rect 6076 34860 6244 34916
rect 6972 34916 7028 35756
rect 5516 34078 5518 34130
rect 5570 34078 5572 34130
rect 5516 34066 5572 34078
rect 5852 34692 5908 34702
rect 5852 34354 5908 34636
rect 5852 34302 5854 34354
rect 5906 34302 5908 34354
rect 4060 33348 4116 33358
rect 4060 33346 4228 33348
rect 4060 33294 4062 33346
rect 4114 33294 4228 33346
rect 4060 33292 4228 33294
rect 4060 33282 4116 33292
rect 3948 32510 3950 32562
rect 4002 32510 4004 32562
rect 3948 30660 4004 32510
rect 4060 31892 4116 31902
rect 4060 30882 4116 31836
rect 4060 30830 4062 30882
rect 4114 30830 4116 30882
rect 4060 30818 4116 30830
rect 4172 31444 4228 33292
rect 4956 33234 5012 33246
rect 4956 33182 4958 33234
rect 5010 33182 5012 33234
rect 4956 32788 5012 33182
rect 5012 32732 5124 32788
rect 4956 32722 5012 32732
rect 4956 32562 5012 32574
rect 4956 32510 4958 32562
rect 5010 32510 5012 32562
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4732 32004 4788 32014
rect 4284 31778 4340 31790
rect 4620 31780 4676 31790
rect 4284 31726 4286 31778
rect 4338 31726 4340 31778
rect 4284 31668 4340 31726
rect 4284 31602 4340 31612
rect 4508 31724 4620 31780
rect 3948 30594 4004 30604
rect 4172 30436 4228 31388
rect 4508 30994 4564 31724
rect 4620 31686 4676 31724
rect 4732 31668 4788 31948
rect 4956 31892 5012 32510
rect 4956 31826 5012 31836
rect 4956 31668 5012 31678
rect 4732 31666 5012 31668
rect 4732 31614 4958 31666
rect 5010 31614 5012 31666
rect 4732 31612 5012 31614
rect 4956 31602 5012 31612
rect 4508 30942 4510 30994
rect 4562 30942 4564 30994
rect 4508 30930 4564 30942
rect 4956 31220 5012 31230
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4172 30380 4676 30436
rect 4284 30210 4340 30222
rect 4284 30158 4286 30210
rect 4338 30158 4340 30210
rect 4284 29988 4340 30158
rect 4620 30210 4676 30380
rect 4620 30158 4622 30210
rect 4674 30158 4676 30210
rect 4620 30146 4676 30158
rect 4956 30098 5012 31164
rect 5068 31108 5124 32732
rect 5292 32676 5348 33516
rect 5404 34020 5460 34030
rect 5404 32788 5460 33964
rect 5852 33236 5908 34302
rect 6076 33572 6132 34860
rect 6972 34850 7028 34860
rect 7196 35698 7252 35868
rect 7196 35646 7198 35698
rect 7250 35646 7252 35698
rect 6300 34804 6356 34814
rect 6188 34692 6244 34702
rect 6188 34598 6244 34636
rect 6300 34020 6356 34748
rect 7196 34356 7252 35646
rect 7308 35922 7364 38612
rect 7868 38050 7924 38062
rect 7868 37998 7870 38050
rect 7922 37998 7924 38050
rect 7644 37940 7700 37950
rect 7420 36708 7476 36718
rect 7420 36482 7476 36652
rect 7420 36430 7422 36482
rect 7474 36430 7476 36482
rect 7420 36418 7476 36430
rect 7308 35870 7310 35922
rect 7362 35870 7364 35922
rect 7308 35140 7364 35870
rect 7644 36370 7700 37884
rect 7868 37268 7924 37998
rect 7868 37174 7924 37212
rect 8316 38050 8372 38062
rect 8316 37998 8318 38050
rect 8370 37998 8372 38050
rect 8316 37044 8372 37998
rect 8428 37156 8484 40348
rect 8764 39618 8820 40796
rect 8988 40962 9044 41356
rect 8988 40910 8990 40962
rect 9042 40910 9044 40962
rect 8988 40180 9044 40910
rect 9100 40852 9156 40862
rect 9100 40516 9156 40796
rect 9212 40628 9268 43820
rect 9548 43762 9604 43820
rect 9548 43710 9550 43762
rect 9602 43710 9604 43762
rect 9548 43698 9604 43710
rect 9548 42756 9604 42766
rect 9660 42756 9716 43932
rect 10108 43540 10164 43550
rect 10444 43540 10500 45388
rect 10780 45218 10836 47294
rect 10780 45166 10782 45218
rect 10834 45166 10836 45218
rect 10780 45154 10836 45166
rect 10892 46898 10948 46910
rect 10892 46846 10894 46898
rect 10946 46846 10948 46898
rect 10780 44994 10836 45006
rect 10780 44942 10782 44994
rect 10834 44942 10836 44994
rect 10780 43764 10836 44942
rect 10892 44322 10948 46846
rect 11228 46676 11284 48974
rect 11452 48802 11508 49758
rect 11452 48750 11454 48802
rect 11506 48750 11508 48802
rect 11452 48130 11508 48750
rect 11564 48914 11620 48926
rect 11564 48862 11566 48914
rect 11618 48862 11620 48914
rect 11564 48468 11620 48862
rect 11564 48402 11620 48412
rect 11676 48354 11732 49868
rect 11676 48302 11678 48354
rect 11730 48302 11732 48354
rect 11676 48290 11732 48302
rect 11788 48692 11844 50542
rect 12012 51378 12068 51390
rect 12012 51326 12014 51378
rect 12066 51326 12068 51378
rect 12012 50708 12068 51326
rect 12236 50820 12292 51996
rect 12460 52050 12516 52332
rect 12572 52276 12628 53006
rect 12572 52210 12628 52220
rect 12796 52946 12852 52958
rect 12796 52894 12798 52946
rect 12850 52894 12852 52946
rect 12796 52724 12852 52894
rect 13468 52948 13524 53678
rect 13468 52854 13524 52892
rect 13580 53730 13748 53732
rect 13580 53678 13694 53730
rect 13746 53678 13748 53730
rect 13580 53676 13748 53678
rect 13580 52724 13636 53676
rect 13692 53666 13748 53676
rect 21980 53730 22036 53742
rect 21980 53678 21982 53730
rect 22034 53678 22036 53730
rect 14252 53618 14308 53630
rect 14252 53566 14254 53618
rect 14306 53566 14308 53618
rect 12796 52668 13636 52724
rect 12460 51998 12462 52050
rect 12514 51998 12516 52050
rect 12460 51986 12516 51998
rect 12796 52052 12852 52668
rect 12796 51986 12852 51996
rect 13244 52276 13300 52286
rect 13244 51490 13300 52220
rect 13244 51438 13246 51490
rect 13298 51438 13300 51490
rect 13244 51426 13300 51438
rect 12348 51380 12404 51390
rect 12348 51266 12404 51324
rect 13580 51378 13636 52668
rect 13580 51326 13582 51378
rect 13634 51326 13636 51378
rect 13580 51314 13636 51326
rect 13916 53170 13972 53182
rect 13916 53118 13918 53170
rect 13970 53118 13972 53170
rect 12348 51214 12350 51266
rect 12402 51214 12404 51266
rect 12348 51202 12404 51214
rect 12460 51156 12516 51166
rect 12460 51062 12516 51100
rect 13692 51156 13748 51166
rect 12460 50820 12516 50830
rect 12236 50818 12516 50820
rect 12236 50766 12462 50818
rect 12514 50766 12516 50818
rect 12236 50764 12516 50766
rect 12460 50754 12516 50764
rect 12012 50594 12068 50652
rect 12012 50542 12014 50594
rect 12066 50542 12068 50594
rect 12012 50530 12068 50542
rect 13692 50594 13748 51100
rect 13692 50542 13694 50594
rect 13746 50542 13748 50594
rect 13692 50530 13748 50542
rect 13916 50596 13972 53118
rect 13916 50530 13972 50540
rect 14140 52162 14196 52174
rect 14140 52110 14142 52162
rect 14194 52110 14196 52162
rect 14140 50148 14196 52110
rect 14252 50706 14308 53566
rect 21308 53618 21364 53630
rect 21532 53620 21588 53630
rect 21308 53566 21310 53618
rect 21362 53566 21364 53618
rect 19836 53340 20100 53350
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 19836 53274 20100 53284
rect 14924 53060 14980 53070
rect 14924 52834 14980 53004
rect 15596 53060 15652 53070
rect 15596 52966 15652 53004
rect 16156 53060 16212 53070
rect 16156 52966 16212 53004
rect 18060 53058 18116 53070
rect 18060 53006 18062 53058
rect 18114 53006 18116 53058
rect 14924 52782 14926 52834
rect 14978 52782 14980 52834
rect 14588 52276 14644 52286
rect 14588 52182 14644 52220
rect 14588 52052 14644 52062
rect 14924 52052 14980 52782
rect 15484 52946 15540 52958
rect 17388 52948 17444 52958
rect 15484 52894 15486 52946
rect 15538 52894 15540 52946
rect 15260 52276 15316 52286
rect 15148 52164 15204 52174
rect 15148 52070 15204 52108
rect 14588 52050 14980 52052
rect 14588 51998 14590 52050
rect 14642 51998 14980 52050
rect 14588 51996 14980 51998
rect 14476 51380 14532 51390
rect 14476 51286 14532 51324
rect 14252 50654 14254 50706
rect 14306 50654 14308 50706
rect 14252 50642 14308 50654
rect 14140 50082 14196 50092
rect 13580 49924 13636 49934
rect 13580 49830 13636 49868
rect 14028 49924 14084 49934
rect 11452 48078 11454 48130
rect 11506 48078 11508 48130
rect 11452 48066 11508 48078
rect 11788 47570 11844 48636
rect 12348 49810 12404 49822
rect 12348 49758 12350 49810
rect 12402 49758 12404 49810
rect 12348 48804 12404 49758
rect 13916 49810 13972 49822
rect 13916 49758 13918 49810
rect 13970 49758 13972 49810
rect 12908 49700 12964 49710
rect 12908 49606 12964 49644
rect 11900 48468 11956 48478
rect 11956 48412 12068 48468
rect 11900 48402 11956 48412
rect 11788 47518 11790 47570
rect 11842 47518 11844 47570
rect 11788 47506 11844 47518
rect 11900 48244 11956 48254
rect 11228 46610 11284 46620
rect 11900 46562 11956 48188
rect 11900 46510 11902 46562
rect 11954 46510 11956 46562
rect 11900 46498 11956 46510
rect 12012 46674 12068 48412
rect 12348 47458 12404 48748
rect 13468 49026 13524 49038
rect 13468 48974 13470 49026
rect 13522 48974 13524 49026
rect 12796 48244 12852 48254
rect 12796 48150 12852 48188
rect 12348 47406 12350 47458
rect 12402 47406 12404 47458
rect 12348 47394 12404 47406
rect 13468 47348 13524 48974
rect 13692 49026 13748 49038
rect 13692 48974 13694 49026
rect 13746 48974 13748 49026
rect 13692 48692 13748 48974
rect 13356 47292 13524 47348
rect 13580 48636 13692 48692
rect 12908 46900 12964 46910
rect 13356 46900 13412 47292
rect 12908 46898 13412 46900
rect 12908 46846 12910 46898
rect 12962 46846 13412 46898
rect 12908 46844 13412 46846
rect 12908 46834 12964 46844
rect 12012 46622 12014 46674
rect 12066 46622 12068 46674
rect 11116 45890 11172 45902
rect 11116 45838 11118 45890
rect 11170 45838 11172 45890
rect 11116 45332 11172 45838
rect 11900 45778 11956 45790
rect 11900 45726 11902 45778
rect 11954 45726 11956 45778
rect 11004 45108 11060 45118
rect 11116 45108 11172 45276
rect 11004 45106 11172 45108
rect 11004 45054 11006 45106
rect 11058 45054 11172 45106
rect 11004 45052 11172 45054
rect 11340 45668 11396 45678
rect 11340 45106 11396 45612
rect 11900 45668 11956 45726
rect 11900 45602 11956 45612
rect 11340 45054 11342 45106
rect 11394 45054 11396 45106
rect 11004 45042 11060 45052
rect 11340 45042 11396 45054
rect 12012 45332 12068 46622
rect 12124 46676 12180 46686
rect 12124 46582 12180 46620
rect 13356 46674 13412 46844
rect 13356 46622 13358 46674
rect 13410 46622 13412 46674
rect 13356 46610 13412 46622
rect 13468 46676 13524 46686
rect 13580 46676 13636 48636
rect 13692 48626 13748 48636
rect 13916 48356 13972 49758
rect 13916 47796 13972 48300
rect 13916 47730 13972 47740
rect 14028 49026 14084 49868
rect 14140 49922 14196 49934
rect 14140 49870 14142 49922
rect 14194 49870 14196 49922
rect 14140 49700 14196 49870
rect 14588 49700 14644 51996
rect 15260 50594 15316 52220
rect 15484 51492 15540 52894
rect 16716 52946 17444 52948
rect 16716 52894 17390 52946
rect 17442 52894 17444 52946
rect 16716 52892 17444 52894
rect 15596 52724 15652 52734
rect 15596 52722 15764 52724
rect 15596 52670 15598 52722
rect 15650 52670 15764 52722
rect 15596 52668 15764 52670
rect 15596 52658 15652 52668
rect 15484 51044 15540 51436
rect 15708 52162 15764 52668
rect 16604 52276 16660 52286
rect 16604 52182 16660 52220
rect 15708 52110 15710 52162
rect 15762 52110 15764 52162
rect 15708 51380 15764 52110
rect 16380 52164 16436 52174
rect 16156 51380 16212 51390
rect 15708 51378 16212 51380
rect 15708 51326 16158 51378
rect 16210 51326 16212 51378
rect 15708 51324 16212 51326
rect 16156 51314 16212 51324
rect 16380 51378 16436 52108
rect 16716 51602 16772 52892
rect 17388 52882 17444 52892
rect 17948 52946 18004 52958
rect 17948 52894 17950 52946
rect 18002 52894 18004 52946
rect 16716 51550 16718 51602
rect 16770 51550 16772 51602
rect 16716 51538 16772 51550
rect 17276 52388 17332 52398
rect 17276 52274 17332 52332
rect 17276 52222 17278 52274
rect 17330 52222 17332 52274
rect 16380 51326 16382 51378
rect 16434 51326 16436 51378
rect 16380 51314 16436 51326
rect 17276 51268 17332 52222
rect 17948 52276 18004 52894
rect 18060 52388 18116 53006
rect 19628 52948 19684 52958
rect 19628 52854 19684 52892
rect 20636 52948 20692 52958
rect 18396 52836 18452 52846
rect 18396 52742 18452 52780
rect 19180 52836 19236 52846
rect 19180 52742 19236 52780
rect 20076 52834 20132 52846
rect 20076 52782 20078 52834
rect 20130 52782 20132 52834
rect 20076 52500 20132 52782
rect 20076 52434 20132 52444
rect 18060 52322 18116 52332
rect 17948 52210 18004 52220
rect 18620 52276 18676 52286
rect 18620 52164 18676 52220
rect 19740 52276 19796 52286
rect 18620 52162 19012 52164
rect 18620 52110 18622 52162
rect 18674 52110 19012 52162
rect 18620 52108 19012 52110
rect 18620 52098 18676 52108
rect 17612 52050 17668 52062
rect 17612 51998 17614 52050
rect 17666 51998 17668 52050
rect 17612 51380 17668 51998
rect 17948 51380 18004 51390
rect 17612 51378 18004 51380
rect 17612 51326 17950 51378
rect 18002 51326 18004 51378
rect 17612 51324 18004 51326
rect 17500 51268 17556 51278
rect 17276 51266 17556 51268
rect 17276 51214 17502 51266
rect 17554 51214 17556 51266
rect 17276 51212 17556 51214
rect 15820 51156 15876 51166
rect 15820 51154 16100 51156
rect 15820 51102 15822 51154
rect 15874 51102 16100 51154
rect 15820 51100 16100 51102
rect 15820 51090 15876 51100
rect 15484 50978 15540 50988
rect 15260 50542 15262 50594
rect 15314 50542 15316 50594
rect 15260 50530 15316 50542
rect 15708 50484 15764 50494
rect 14140 49698 14644 49700
rect 14140 49646 14590 49698
rect 14642 49646 14644 49698
rect 14140 49644 14644 49646
rect 14028 48974 14030 49026
rect 14082 48974 14084 49026
rect 13804 47458 13860 47470
rect 13804 47406 13806 47458
rect 13858 47406 13860 47458
rect 13804 46786 13860 47406
rect 13804 46734 13806 46786
rect 13858 46734 13860 46786
rect 13804 46722 13860 46734
rect 13468 46674 13636 46676
rect 13468 46622 13470 46674
rect 13522 46622 13636 46674
rect 13468 46620 13636 46622
rect 13468 46610 13524 46620
rect 13692 46564 13748 46574
rect 14028 46564 14084 48974
rect 14140 48018 14196 48030
rect 14140 47966 14142 48018
rect 14194 47966 14196 48018
rect 14140 47684 14196 47966
rect 14140 47458 14196 47628
rect 14140 47406 14142 47458
rect 14194 47406 14196 47458
rect 14140 47394 14196 47406
rect 14476 47124 14532 49644
rect 14588 49634 14644 49644
rect 14700 50148 14756 50158
rect 14700 49140 14756 50092
rect 15708 50034 15764 50428
rect 15708 49982 15710 50034
rect 15762 49982 15764 50034
rect 15708 49970 15764 49982
rect 15372 49810 15428 49822
rect 15372 49758 15374 49810
rect 15426 49758 15428 49810
rect 14700 49074 14756 49084
rect 15148 49700 15204 49710
rect 15148 49026 15204 49644
rect 15372 49140 15428 49758
rect 15372 49074 15428 49084
rect 15484 49138 15540 49150
rect 15484 49086 15486 49138
rect 15538 49086 15540 49138
rect 15148 48974 15150 49026
rect 15202 48974 15204 49026
rect 15148 48962 15204 48974
rect 14700 48916 14756 48926
rect 14700 48130 14756 48860
rect 14700 48078 14702 48130
rect 14754 48078 14756 48130
rect 14700 48066 14756 48078
rect 15036 48354 15092 48366
rect 15036 48302 15038 48354
rect 15090 48302 15092 48354
rect 14588 47572 14644 47582
rect 14588 47478 14644 47516
rect 14700 47348 14756 47358
rect 14700 47254 14756 47292
rect 15036 47236 15092 48302
rect 15036 47170 15092 47180
rect 14476 47068 14756 47124
rect 13692 46562 14084 46564
rect 13692 46510 13694 46562
rect 13746 46510 14084 46562
rect 13692 46508 14084 46510
rect 13692 46498 13748 46508
rect 12908 45890 12964 45902
rect 12908 45838 12910 45890
rect 12962 45838 12964 45890
rect 12796 45780 12852 45790
rect 12796 45666 12852 45724
rect 12796 45614 12798 45666
rect 12850 45614 12852 45666
rect 12796 45602 12852 45614
rect 10892 44270 10894 44322
rect 10946 44270 10948 44322
rect 10892 44258 10948 44270
rect 11340 44884 11396 44894
rect 10108 43538 10500 43540
rect 10108 43486 10110 43538
rect 10162 43486 10500 43538
rect 10108 43484 10500 43486
rect 10556 43762 10836 43764
rect 10556 43710 10782 43762
rect 10834 43710 10836 43762
rect 10556 43708 10836 43710
rect 10108 43474 10164 43484
rect 9548 42754 9716 42756
rect 9548 42702 9550 42754
rect 9602 42702 9716 42754
rect 9548 42700 9716 42702
rect 9324 42642 9380 42654
rect 9324 42590 9326 42642
rect 9378 42590 9380 42642
rect 9324 41636 9380 42590
rect 9324 41570 9380 41580
rect 9324 41186 9380 41198
rect 9324 41134 9326 41186
rect 9378 41134 9380 41186
rect 9324 40964 9380 41134
rect 9548 41186 9604 42700
rect 9772 42532 9828 42542
rect 9548 41134 9550 41186
rect 9602 41134 9604 41186
rect 9548 41122 9604 41134
rect 9660 41636 9716 41646
rect 9660 41186 9716 41580
rect 9660 41134 9662 41186
rect 9714 41134 9716 41186
rect 9660 41122 9716 41134
rect 9772 40964 9828 42476
rect 9884 42530 9940 42542
rect 9884 42478 9886 42530
rect 9938 42478 9940 42530
rect 9884 42082 9940 42478
rect 10108 42532 10164 42542
rect 10108 42438 10164 42476
rect 10444 42530 10500 42542
rect 10444 42478 10446 42530
rect 10498 42478 10500 42530
rect 9884 42030 9886 42082
rect 9938 42030 9940 42082
rect 9884 42018 9940 42030
rect 10444 42084 10500 42478
rect 10556 42194 10612 43708
rect 10780 43698 10836 43708
rect 11340 43428 11396 44828
rect 12012 44434 12068 45276
rect 12348 45220 12404 45230
rect 12012 44382 12014 44434
rect 12066 44382 12068 44434
rect 12012 44370 12068 44382
rect 12124 44996 12180 45006
rect 11340 43334 11396 43372
rect 11788 44322 11844 44334
rect 11788 44270 11790 44322
rect 11842 44270 11844 44322
rect 10556 42142 10558 42194
rect 10610 42142 10612 42194
rect 10556 42130 10612 42142
rect 11228 43204 11284 43214
rect 10444 42018 10500 42028
rect 9996 41970 10052 41982
rect 9996 41918 9998 41970
rect 10050 41918 10052 41970
rect 9324 40908 9828 40964
rect 9884 40964 9940 40974
rect 9324 40740 9380 40908
rect 9324 40674 9380 40684
rect 9212 40562 9268 40572
rect 9100 40422 9156 40460
rect 8988 40114 9044 40124
rect 8764 39566 8766 39618
rect 8818 39566 8820 39618
rect 8540 39508 8596 39518
rect 8540 39506 8708 39508
rect 8540 39454 8542 39506
rect 8594 39454 8708 39506
rect 8540 39452 8708 39454
rect 8540 39442 8596 39452
rect 8652 38164 8708 39452
rect 8764 38668 8820 39566
rect 9100 39620 9156 39630
rect 9100 39526 9156 39564
rect 8988 39394 9044 39406
rect 8988 39342 8990 39394
rect 9042 39342 9044 39394
rect 8764 38612 8932 38668
rect 8876 38276 8932 38612
rect 8988 38500 9044 39342
rect 9436 39394 9492 39406
rect 9436 39342 9438 39394
rect 9490 39342 9492 39394
rect 9436 39060 9492 39342
rect 9436 38994 9492 39004
rect 9884 38668 9940 40908
rect 9996 39396 10052 41918
rect 10668 41972 10724 41982
rect 10668 41878 10724 41916
rect 10892 41748 10948 41758
rect 10108 41188 10164 41198
rect 10108 41094 10164 41132
rect 10892 41186 10948 41692
rect 10892 41134 10894 41186
rect 10946 41134 10948 41186
rect 10668 40516 10724 40526
rect 10556 40404 10612 40414
rect 10668 40404 10724 40460
rect 10556 40402 10724 40404
rect 10556 40350 10558 40402
rect 10610 40350 10724 40402
rect 10556 40348 10724 40350
rect 10892 40404 10948 41134
rect 10556 40338 10612 40348
rect 10892 40338 10948 40348
rect 11116 41076 11172 41086
rect 11116 40626 11172 41020
rect 11116 40574 11118 40626
rect 11170 40574 11172 40626
rect 11116 39730 11172 40574
rect 11116 39678 11118 39730
rect 11170 39678 11172 39730
rect 11116 39666 11172 39678
rect 9996 39330 10052 39340
rect 10108 39618 10164 39630
rect 10892 39620 10948 39630
rect 10108 39566 10110 39618
rect 10162 39566 10164 39618
rect 10108 38948 10164 39566
rect 10108 38882 10164 38892
rect 10332 39618 10948 39620
rect 10332 39566 10894 39618
rect 10946 39566 10948 39618
rect 10332 39564 10948 39566
rect 9884 38612 10052 38668
rect 8988 38434 9044 38444
rect 9772 38500 9828 38510
rect 8876 38220 9380 38276
rect 8764 38164 8820 38174
rect 8652 38162 8820 38164
rect 8652 38110 8766 38162
rect 8818 38110 8820 38162
rect 8652 38108 8820 38110
rect 8764 37716 8820 38108
rect 9324 38050 9380 38220
rect 9324 37998 9326 38050
rect 9378 37998 9380 38050
rect 9324 37986 9380 37998
rect 9212 37940 9268 37950
rect 9212 37846 9268 37884
rect 9436 37938 9492 37950
rect 9436 37886 9438 37938
rect 9490 37886 9492 37938
rect 9436 37716 9492 37886
rect 8764 37660 9492 37716
rect 9548 37940 9604 37950
rect 9548 37490 9604 37884
rect 9548 37438 9550 37490
rect 9602 37438 9604 37490
rect 9548 37426 9604 37438
rect 9772 37492 9828 38444
rect 9884 37828 9940 37838
rect 9884 37734 9940 37772
rect 9884 37492 9940 37502
rect 9772 37490 9940 37492
rect 9772 37438 9886 37490
rect 9938 37438 9940 37490
rect 9772 37436 9940 37438
rect 9884 37380 9940 37436
rect 9884 37314 9940 37324
rect 8764 37156 8820 37166
rect 8428 37100 8708 37156
rect 8316 36978 8372 36988
rect 7644 36318 7646 36370
rect 7698 36318 7700 36370
rect 7644 35924 7700 36318
rect 7756 36370 7812 36382
rect 7756 36318 7758 36370
rect 7810 36318 7812 36370
rect 7756 36148 7812 36318
rect 8204 36260 8260 36270
rect 8204 36166 8260 36204
rect 7756 36082 7812 36092
rect 8652 35924 8708 37100
rect 7644 35868 7924 35924
rect 7756 35700 7812 35710
rect 7756 35588 7812 35644
rect 7308 35074 7364 35084
rect 7644 35586 7812 35588
rect 7644 35534 7758 35586
rect 7810 35534 7812 35586
rect 7644 35532 7812 35534
rect 7196 34290 7252 34300
rect 7308 34916 7364 34926
rect 7644 34916 7700 35532
rect 7756 35522 7812 35532
rect 7308 34914 7700 34916
rect 7308 34862 7310 34914
rect 7362 34862 7700 34914
rect 7308 34860 7700 34862
rect 7308 34354 7364 34860
rect 7756 34804 7812 34814
rect 7756 34710 7812 34748
rect 7868 34580 7924 35868
rect 8652 35858 8708 35868
rect 8652 35700 8708 35738
rect 8652 35634 8708 35644
rect 7980 35476 8036 35486
rect 8316 35476 8372 35486
rect 7980 35382 8036 35420
rect 8092 35474 8372 35476
rect 8092 35422 8318 35474
rect 8370 35422 8372 35474
rect 8092 35420 8372 35422
rect 7308 34302 7310 34354
rect 7362 34302 7364 34354
rect 7308 34290 7364 34302
rect 7532 34524 7924 34580
rect 7980 35140 8036 35150
rect 7532 34354 7588 34524
rect 7532 34302 7534 34354
rect 7586 34302 7588 34354
rect 7084 34242 7140 34254
rect 7084 34190 7086 34242
rect 7138 34190 7140 34242
rect 6076 33506 6132 33516
rect 6188 34018 6356 34020
rect 6188 33966 6302 34018
rect 6354 33966 6356 34018
rect 6188 33964 6356 33966
rect 6188 33460 6244 33964
rect 6300 33954 6356 33964
rect 6748 34130 6804 34142
rect 6748 34078 6750 34130
rect 6802 34078 6804 34130
rect 5516 32788 5572 32798
rect 5404 32732 5516 32788
rect 5516 32694 5572 32732
rect 5292 32610 5348 32620
rect 5852 32562 5908 33180
rect 5964 33348 6020 33358
rect 5964 32674 6020 33292
rect 6188 33234 6244 33404
rect 6748 33348 6804 34078
rect 7084 34132 7140 34190
rect 7532 34132 7588 34302
rect 7084 34076 7588 34132
rect 7644 34356 7700 34366
rect 7644 34130 7700 34300
rect 7644 34078 7646 34130
rect 7698 34078 7700 34130
rect 6748 33282 6804 33292
rect 7084 33346 7140 33358
rect 7084 33294 7086 33346
rect 7138 33294 7140 33346
rect 6188 33182 6190 33234
rect 6242 33182 6244 33234
rect 6188 33170 6244 33182
rect 6524 33122 6580 33134
rect 6524 33070 6526 33122
rect 6578 33070 6580 33122
rect 5964 32622 5966 32674
rect 6018 32622 6020 32674
rect 5964 32610 6020 32622
rect 6188 33012 6244 33022
rect 6188 32674 6244 32956
rect 6188 32622 6190 32674
rect 6242 32622 6244 32674
rect 6188 32610 6244 32622
rect 5852 32510 5854 32562
rect 5906 32510 5908 32562
rect 5852 32498 5908 32510
rect 6188 32340 6244 32350
rect 5628 31892 5684 31902
rect 5628 31798 5684 31836
rect 6188 31778 6244 32284
rect 6188 31726 6190 31778
rect 6242 31726 6244 31778
rect 6188 31714 6244 31726
rect 6524 31780 6580 33070
rect 7084 32788 7140 33294
rect 7644 33348 7700 34078
rect 7644 33282 7700 33292
rect 7756 33236 7812 33246
rect 7756 33142 7812 33180
rect 7308 33122 7364 33134
rect 7308 33070 7310 33122
rect 7362 33070 7364 33122
rect 7308 33012 7364 33070
rect 7308 32946 7364 32956
rect 7868 33122 7924 33134
rect 7868 33070 7870 33122
rect 7922 33070 7924 33122
rect 6636 32786 7140 32788
rect 6636 32734 7086 32786
rect 7138 32734 7140 32786
rect 6636 32732 7140 32734
rect 6636 32562 6692 32732
rect 7084 32722 7140 32732
rect 7420 32788 7476 32798
rect 6636 32510 6638 32562
rect 6690 32510 6692 32562
rect 6636 32498 6692 32510
rect 7420 32562 7476 32732
rect 7868 32788 7924 33070
rect 7644 32676 7700 32686
rect 7644 32564 7700 32620
rect 7420 32510 7422 32562
rect 7474 32510 7476 32562
rect 7420 32498 7476 32510
rect 7532 32562 7700 32564
rect 7532 32510 7646 32562
rect 7698 32510 7700 32562
rect 7532 32508 7700 32510
rect 6860 32338 6916 32350
rect 6860 32286 6862 32338
rect 6914 32286 6916 32338
rect 6860 31892 6916 32286
rect 6860 31826 6916 31836
rect 6524 31714 6580 31724
rect 7420 31780 7476 31790
rect 7532 31780 7588 32508
rect 7644 32498 7700 32508
rect 7868 32004 7924 32732
rect 7868 31938 7924 31948
rect 7980 32564 8036 35084
rect 8092 34130 8148 35420
rect 8316 35410 8372 35420
rect 8652 35474 8708 35486
rect 8652 35422 8654 35474
rect 8706 35422 8708 35474
rect 8652 35364 8708 35422
rect 8428 35308 8708 35364
rect 8428 35252 8484 35308
rect 8316 35196 8484 35252
rect 8316 34914 8372 35196
rect 8764 35026 8820 37100
rect 8764 34974 8766 35026
rect 8818 34974 8820 35026
rect 8764 34962 8820 34974
rect 8876 37044 8932 37054
rect 8316 34862 8318 34914
rect 8370 34862 8372 34914
rect 8316 34850 8372 34862
rect 8652 34692 8708 34702
rect 8652 34354 8708 34636
rect 8652 34302 8654 34354
rect 8706 34302 8708 34354
rect 8652 34290 8708 34302
rect 8092 34078 8094 34130
rect 8146 34078 8148 34130
rect 8092 34066 8148 34078
rect 8428 34132 8484 34142
rect 8428 34038 8484 34076
rect 8540 34132 8596 34142
rect 8876 34132 8932 36988
rect 8988 37042 9044 37054
rect 8988 36990 8990 37042
rect 9042 36990 9044 37042
rect 8988 36484 9044 36990
rect 8988 36418 9044 36428
rect 9548 35700 9604 35710
rect 8988 35476 9044 35486
rect 8988 35382 9044 35420
rect 9548 35026 9604 35644
rect 9660 35586 9716 35598
rect 9660 35534 9662 35586
rect 9714 35534 9716 35586
rect 9660 35364 9716 35534
rect 9660 35298 9716 35308
rect 9772 35476 9828 35486
rect 9772 35138 9828 35420
rect 9772 35086 9774 35138
rect 9826 35086 9828 35138
rect 9772 35074 9828 35086
rect 9548 34974 9550 35026
rect 9602 34974 9604 35026
rect 9548 34962 9604 34974
rect 9212 34914 9268 34926
rect 9212 34862 9214 34914
rect 9266 34862 9268 34914
rect 8540 34130 8932 34132
rect 8540 34078 8542 34130
rect 8594 34078 8932 34130
rect 8540 34076 8932 34078
rect 9100 34802 9156 34814
rect 9100 34750 9102 34802
rect 9154 34750 9156 34802
rect 8540 34066 8596 34076
rect 8428 33460 8484 33470
rect 8428 33366 8484 33404
rect 9100 33460 9156 34750
rect 9212 34804 9268 34862
rect 9212 34020 9268 34748
rect 9996 34468 10052 38612
rect 10332 36706 10388 39564
rect 10892 39554 10948 39564
rect 10444 39394 10500 39406
rect 10444 39342 10446 39394
rect 10498 39342 10500 39394
rect 10444 38834 10500 39342
rect 10556 39396 10612 39406
rect 10556 39302 10612 39340
rect 10668 39394 10724 39406
rect 10668 39342 10670 39394
rect 10722 39342 10724 39394
rect 10444 38782 10446 38834
rect 10498 38782 10500 38834
rect 10444 37828 10500 38782
rect 10444 37762 10500 37772
rect 10668 38834 10724 39342
rect 11228 39396 11284 43148
rect 11788 42980 11844 44270
rect 12124 43426 12180 44940
rect 12348 44324 12404 45164
rect 12348 44230 12404 44268
rect 12572 45220 12628 45230
rect 12572 43650 12628 45164
rect 12572 43598 12574 43650
rect 12626 43598 12628 43650
rect 12572 43586 12628 43598
rect 12124 43374 12126 43426
rect 12178 43374 12180 43426
rect 12124 43362 12180 43374
rect 12908 43428 12964 45838
rect 13804 45890 13860 45902
rect 13804 45838 13806 45890
rect 13858 45838 13860 45890
rect 13804 45780 13860 45838
rect 13580 45668 13636 45678
rect 13580 45106 13636 45612
rect 13580 45054 13582 45106
rect 13634 45054 13636 45106
rect 13580 45042 13636 45054
rect 13468 44324 13524 44334
rect 13468 43538 13524 44268
rect 13804 44322 13860 45724
rect 13916 45890 13972 45902
rect 13916 45838 13918 45890
rect 13970 45838 13972 45890
rect 13916 45332 13972 45838
rect 13916 45266 13972 45276
rect 14140 45890 14196 45902
rect 14140 45838 14142 45890
rect 14194 45838 14196 45890
rect 14140 45220 14196 45838
rect 14140 45154 14196 45164
rect 14252 45778 14308 45790
rect 14252 45726 14254 45778
rect 14306 45726 14308 45778
rect 13804 44270 13806 44322
rect 13858 44270 13860 44322
rect 13804 44258 13860 44270
rect 14028 43764 14084 43774
rect 14028 43670 14084 43708
rect 13468 43486 13470 43538
rect 13522 43486 13524 43538
rect 13468 43474 13524 43486
rect 14252 43540 14308 45726
rect 14364 45332 14420 45342
rect 14364 44434 14420 45276
rect 14364 44382 14366 44434
rect 14418 44382 14420 44434
rect 14364 44370 14420 44382
rect 14588 43540 14644 43550
rect 14252 43538 14644 43540
rect 14252 43486 14590 43538
rect 14642 43486 14644 43538
rect 14252 43484 14644 43486
rect 14588 43474 14644 43484
rect 12908 43362 12964 43372
rect 14028 43428 14084 43438
rect 11676 42924 11844 42980
rect 11564 42082 11620 42094
rect 11564 42030 11566 42082
rect 11618 42030 11620 42082
rect 11564 41860 11620 42030
rect 11564 41794 11620 41804
rect 11564 41188 11620 41198
rect 11564 41094 11620 41132
rect 11676 41074 11732 42924
rect 12348 42866 12404 42878
rect 12348 42814 12350 42866
rect 12402 42814 12404 42866
rect 11676 41022 11678 41074
rect 11730 41022 11732 41074
rect 11676 41010 11732 41022
rect 11788 42754 11844 42766
rect 11788 42702 11790 42754
rect 11842 42702 11844 42754
rect 11788 41186 11844 42702
rect 11788 41134 11790 41186
rect 11842 41134 11844 41186
rect 11788 40516 11844 41134
rect 11900 42754 11956 42766
rect 11900 42702 11902 42754
rect 11954 42702 11956 42754
rect 11900 41188 11956 42702
rect 12348 42084 12404 42814
rect 13804 42754 13860 42766
rect 13804 42702 13806 42754
rect 13858 42702 13860 42754
rect 12684 42532 12740 42542
rect 12684 42438 12740 42476
rect 13804 42532 13860 42702
rect 13356 42194 13412 42206
rect 13356 42142 13358 42194
rect 13410 42142 13412 42194
rect 12348 42028 12628 42084
rect 12124 41972 12180 41982
rect 12124 41970 12404 41972
rect 12124 41918 12126 41970
rect 12178 41918 12404 41970
rect 12124 41916 12404 41918
rect 12124 41906 12180 41916
rect 11900 41122 11956 41132
rect 12012 41860 12068 41870
rect 11788 40450 11844 40460
rect 12012 40514 12068 41804
rect 12348 41298 12404 41916
rect 12348 41246 12350 41298
rect 12402 41246 12404 41298
rect 12236 41076 12292 41086
rect 12236 40982 12292 41020
rect 12012 40462 12014 40514
rect 12066 40462 12068 40514
rect 12012 40450 12068 40462
rect 12348 40402 12404 41246
rect 12460 41188 12516 41198
rect 12460 41074 12516 41132
rect 12460 41022 12462 41074
rect 12514 41022 12516 41074
rect 12460 41010 12516 41022
rect 12348 40350 12350 40402
rect 12402 40350 12404 40402
rect 12348 40338 12404 40350
rect 12460 40404 12516 40414
rect 12572 40404 12628 42028
rect 12796 41972 12852 41982
rect 12796 41878 12852 41916
rect 13356 41972 13412 42142
rect 13356 41906 13412 41916
rect 13804 41970 13860 42476
rect 14028 42754 14084 43372
rect 14028 42702 14030 42754
rect 14082 42702 14084 42754
rect 13804 41918 13806 41970
rect 13858 41918 13860 41970
rect 13804 41906 13860 41918
rect 13916 42084 13972 42094
rect 13916 41076 13972 42028
rect 14028 41970 14084 42702
rect 14028 41918 14030 41970
rect 14082 41918 14084 41970
rect 14028 41906 14084 41918
rect 14252 42754 14308 42766
rect 14252 42702 14254 42754
rect 14306 42702 14308 42754
rect 14252 41970 14308 42702
rect 14588 42530 14644 42542
rect 14588 42478 14590 42530
rect 14642 42478 14644 42530
rect 14252 41918 14254 41970
rect 14306 41918 14308 41970
rect 14252 41860 14308 41918
rect 14140 41412 14196 41422
rect 14252 41412 14308 41804
rect 14140 41410 14308 41412
rect 14140 41358 14142 41410
rect 14194 41358 14308 41410
rect 14140 41356 14308 41358
rect 14364 42084 14420 42094
rect 14140 41346 14196 41356
rect 14252 41188 14308 41198
rect 14364 41188 14420 42028
rect 14252 41186 14532 41188
rect 14252 41134 14254 41186
rect 14306 41134 14532 41186
rect 14252 41132 14532 41134
rect 14252 41122 14308 41132
rect 13692 41074 13972 41076
rect 13692 41022 13918 41074
rect 13970 41022 13972 41074
rect 13692 41020 13972 41022
rect 13356 40628 13412 40638
rect 12516 40348 12628 40404
rect 13244 40404 13300 40414
rect 12460 40338 12516 40348
rect 13244 40310 13300 40348
rect 13244 40180 13300 40190
rect 11340 39620 11396 39630
rect 11340 39526 11396 39564
rect 11452 39618 11508 39630
rect 11452 39566 11454 39618
rect 11506 39566 11508 39618
rect 11452 39508 11508 39566
rect 11452 39442 11508 39452
rect 12908 39508 12964 39518
rect 11228 39340 11396 39396
rect 11228 38948 11284 38958
rect 11228 38854 11284 38892
rect 10668 38782 10670 38834
rect 10722 38782 10724 38834
rect 10668 37044 10724 38782
rect 11340 38668 11396 39340
rect 12124 39060 12180 39070
rect 12124 38966 12180 39004
rect 11788 38948 11844 38958
rect 11788 38668 11844 38892
rect 11340 38612 11620 38668
rect 11788 38612 12292 38668
rect 11340 38050 11396 38062
rect 11340 37998 11342 38050
rect 11394 37998 11396 38050
rect 11228 37938 11284 37950
rect 11228 37886 11230 37938
rect 11282 37886 11284 37938
rect 10780 37828 10836 37838
rect 10780 37490 10836 37772
rect 10780 37438 10782 37490
rect 10834 37438 10836 37490
rect 10780 37426 10836 37438
rect 11228 37492 11284 37886
rect 11228 37426 11284 37436
rect 10892 37268 10948 37278
rect 10892 37266 11172 37268
rect 10892 37214 10894 37266
rect 10946 37214 11172 37266
rect 10892 37212 11172 37214
rect 10892 37202 10948 37212
rect 11116 37156 11172 37212
rect 11340 37156 11396 37998
rect 11452 37156 11508 37166
rect 11116 37154 11508 37156
rect 11116 37102 11454 37154
rect 11506 37102 11508 37154
rect 11116 37100 11508 37102
rect 11452 37090 11508 37100
rect 11004 37044 11060 37054
rect 10668 37042 11060 37044
rect 10668 36990 11006 37042
rect 11058 36990 11060 37042
rect 10668 36988 11060 36990
rect 10332 36654 10334 36706
rect 10386 36654 10388 36706
rect 10332 36642 10388 36654
rect 10780 36706 10836 36988
rect 11004 36978 11060 36988
rect 10780 36654 10782 36706
rect 10834 36654 10836 36706
rect 10780 36642 10836 36654
rect 11116 36708 11172 36718
rect 11116 36706 11508 36708
rect 11116 36654 11118 36706
rect 11170 36654 11508 36706
rect 11116 36652 11508 36654
rect 10220 36484 10276 36494
rect 10220 36390 10276 36428
rect 11116 36484 11172 36652
rect 11116 36418 11172 36428
rect 11340 36482 11396 36494
rect 11340 36430 11342 36482
rect 11394 36430 11396 36482
rect 10332 36260 10388 36270
rect 11340 36260 11396 36430
rect 10332 36258 11396 36260
rect 10332 36206 10334 36258
rect 10386 36206 11396 36258
rect 10332 36204 11396 36206
rect 10332 36194 10388 36204
rect 10668 36036 10724 36046
rect 10668 35700 10724 35980
rect 10892 35924 10948 35934
rect 10892 35830 10948 35868
rect 10668 35698 10836 35700
rect 10668 35646 10670 35698
rect 10722 35646 10836 35698
rect 10668 35644 10836 35646
rect 10668 35634 10724 35644
rect 10668 35140 10724 35150
rect 10444 35138 10724 35140
rect 10444 35086 10670 35138
rect 10722 35086 10724 35138
rect 10444 35084 10724 35086
rect 10332 34916 10388 34926
rect 10108 34692 10164 34702
rect 10108 34598 10164 34636
rect 9660 34412 10164 34468
rect 9660 34354 9716 34412
rect 9660 34302 9662 34354
rect 9714 34302 9716 34354
rect 9660 34290 9716 34302
rect 9996 34244 10052 34254
rect 9996 34150 10052 34188
rect 9884 34132 9940 34142
rect 9212 33954 9268 33964
rect 9772 34076 9884 34132
rect 9100 33394 9156 33404
rect 9324 33908 9380 33918
rect 9324 33572 9380 33852
rect 9324 33458 9380 33516
rect 9324 33406 9326 33458
rect 9378 33406 9380 33458
rect 9324 33394 9380 33406
rect 9548 33348 9604 33358
rect 8092 33122 8148 33134
rect 8092 33070 8094 33122
rect 8146 33070 8148 33122
rect 8092 33012 8148 33070
rect 8092 32946 8148 32956
rect 8876 33122 8932 33134
rect 8876 33070 8878 33122
rect 8930 33070 8932 33122
rect 8092 32564 8148 32574
rect 7980 32562 8148 32564
rect 7980 32510 8094 32562
rect 8146 32510 8148 32562
rect 7980 32508 8148 32510
rect 7980 31890 8036 32508
rect 8092 32498 8148 32508
rect 8540 32564 8596 32574
rect 8540 32470 8596 32508
rect 7980 31838 7982 31890
rect 8034 31838 8036 31890
rect 7980 31826 8036 31838
rect 8092 32338 8148 32350
rect 8092 32286 8094 32338
rect 8146 32286 8148 32338
rect 7420 31778 7588 31780
rect 7420 31726 7422 31778
rect 7474 31726 7588 31778
rect 7420 31724 7588 31726
rect 7420 31714 7476 31724
rect 6524 31556 6580 31566
rect 6524 31462 6580 31500
rect 6860 31554 6916 31566
rect 6860 31502 6862 31554
rect 6914 31502 6916 31554
rect 5852 31220 5908 31230
rect 5068 31052 5684 31108
rect 4956 30046 4958 30098
rect 5010 30046 5012 30098
rect 4956 30034 5012 30046
rect 4284 29922 4340 29932
rect 4284 29540 4340 29550
rect 4284 29426 4340 29484
rect 4284 29374 4286 29426
rect 4338 29374 4340 29426
rect 4284 29362 4340 29374
rect 5292 29426 5348 31052
rect 5628 30994 5684 31052
rect 5628 30942 5630 30994
rect 5682 30942 5684 30994
rect 5628 30930 5684 30942
rect 5852 30994 5908 31164
rect 6636 31220 6692 31230
rect 5852 30942 5854 30994
rect 5906 30942 5908 30994
rect 5852 30930 5908 30942
rect 6076 31108 6132 31118
rect 6076 30994 6132 31052
rect 6076 30942 6078 30994
rect 6130 30942 6132 30994
rect 6076 30930 6132 30942
rect 6412 31108 6468 31118
rect 5292 29374 5294 29426
rect 5346 29374 5348 29426
rect 5292 29204 5348 29374
rect 5404 30884 5460 30894
rect 5404 29428 5460 30828
rect 5964 30322 6020 30334
rect 5964 30270 5966 30322
rect 6018 30270 6020 30322
rect 5516 29428 5572 29438
rect 5404 29426 5908 29428
rect 5404 29374 5518 29426
rect 5570 29374 5908 29426
rect 5404 29372 5908 29374
rect 5516 29362 5572 29372
rect 5292 29148 5684 29204
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 5628 28866 5684 29148
rect 5628 28814 5630 28866
rect 5682 28814 5684 28866
rect 5628 28802 5684 28814
rect 5852 28530 5908 29372
rect 5964 28866 6020 30270
rect 6412 29426 6468 31052
rect 6524 30996 6580 31006
rect 6524 30902 6580 30940
rect 6524 30098 6580 30110
rect 6524 30046 6526 30098
rect 6578 30046 6580 30098
rect 6524 29876 6580 30046
rect 6524 29810 6580 29820
rect 6412 29374 6414 29426
rect 6466 29374 6468 29426
rect 6412 29362 6468 29374
rect 6636 29426 6692 31164
rect 6748 31108 6804 31118
rect 6748 31014 6804 31052
rect 6636 29374 6638 29426
rect 6690 29374 6692 29426
rect 6636 29362 6692 29374
rect 6860 29428 6916 31502
rect 7084 31554 7140 31566
rect 7084 31502 7086 31554
rect 7138 31502 7140 31554
rect 7084 31444 7140 31502
rect 7308 31556 7364 31566
rect 7308 31462 7364 31500
rect 7084 31378 7140 31388
rect 8092 31220 8148 32286
rect 8876 32340 8932 33070
rect 9548 32674 9604 33292
rect 9660 32788 9716 32798
rect 9660 32694 9716 32732
rect 9548 32622 9550 32674
rect 9602 32622 9604 32674
rect 9548 32610 9604 32622
rect 8876 32274 8932 32284
rect 9660 32338 9716 32350
rect 9660 32286 9662 32338
rect 9714 32286 9716 32338
rect 8652 31892 8708 31902
rect 8708 31836 8820 31892
rect 8652 31798 8708 31836
rect 8540 31780 8596 31790
rect 8092 31218 8372 31220
rect 8092 31166 8094 31218
rect 8146 31166 8372 31218
rect 8092 31164 8372 31166
rect 8092 31154 8148 31164
rect 7084 31108 7140 31118
rect 7084 30994 7140 31052
rect 7084 30942 7086 30994
rect 7138 30942 7140 30994
rect 7084 30930 7140 30942
rect 7532 30996 7588 31006
rect 7084 30772 7140 30782
rect 7084 30770 7476 30772
rect 7084 30718 7086 30770
rect 7138 30718 7476 30770
rect 7084 30716 7476 30718
rect 7084 30706 7140 30716
rect 7420 30210 7476 30716
rect 7420 30158 7422 30210
rect 7474 30158 7476 30210
rect 7420 30146 7476 30158
rect 6860 29362 6916 29372
rect 7420 29876 7476 29886
rect 7420 29426 7476 29820
rect 7420 29374 7422 29426
rect 7474 29374 7476 29426
rect 7420 29362 7476 29374
rect 7532 29538 7588 30940
rect 7532 29486 7534 29538
rect 7586 29486 7588 29538
rect 7532 29428 7588 29486
rect 7644 30994 7700 31006
rect 7644 30942 7646 30994
rect 7698 30942 7700 30994
rect 7644 29428 7700 30942
rect 7868 30996 7924 31006
rect 7868 30902 7924 30940
rect 8204 30770 8260 30782
rect 8204 30718 8206 30770
rect 8258 30718 8260 30770
rect 8204 30212 8260 30718
rect 8204 30146 8260 30156
rect 8092 30100 8148 30110
rect 8092 30006 8148 30044
rect 8316 29876 8372 31164
rect 8540 30994 8596 31724
rect 8540 30942 8542 30994
rect 8594 30942 8596 30994
rect 8540 30930 8596 30942
rect 8764 30994 8820 31836
rect 8876 31780 8932 31790
rect 9660 31780 9716 32286
rect 8876 31778 9716 31780
rect 8876 31726 8878 31778
rect 8930 31726 9662 31778
rect 9714 31726 9716 31778
rect 8876 31724 9716 31726
rect 8876 31714 8932 31724
rect 8876 31218 8932 31230
rect 8876 31166 8878 31218
rect 8930 31166 8932 31218
rect 8876 31108 8932 31166
rect 8876 31042 8932 31052
rect 8764 30942 8766 30994
rect 8818 30942 8820 30994
rect 8764 30930 8820 30942
rect 8988 30994 9044 31724
rect 9660 31714 9716 31724
rect 9324 31554 9380 31566
rect 9324 31502 9326 31554
rect 9378 31502 9380 31554
rect 9324 31220 9380 31502
rect 9436 31220 9492 31230
rect 9324 31164 9436 31220
rect 9436 31154 9492 31164
rect 9772 31218 9828 34076
rect 9884 34066 9940 34076
rect 9772 31166 9774 31218
rect 9826 31166 9828 31218
rect 9772 31154 9828 31166
rect 9996 33460 10052 33470
rect 9548 30996 9604 31006
rect 8988 30942 8990 30994
rect 9042 30942 9044 30994
rect 8988 30930 9044 30942
rect 9100 30994 9604 30996
rect 9100 30942 9550 30994
rect 9602 30942 9604 30994
rect 9100 30940 9604 30942
rect 8988 30212 9044 30222
rect 8988 30118 9044 30156
rect 7756 29764 7812 29774
rect 7756 29650 7812 29708
rect 7756 29598 7758 29650
rect 7810 29598 7812 29650
rect 7756 29586 7812 29598
rect 8316 29538 8372 29820
rect 8988 29652 9044 29662
rect 9100 29652 9156 30940
rect 9548 30930 9604 30940
rect 9996 30434 10052 33404
rect 10108 32676 10164 34412
rect 10332 34354 10388 34860
rect 10332 34302 10334 34354
rect 10386 34302 10388 34354
rect 10332 34290 10388 34302
rect 10444 33234 10500 35084
rect 10668 35074 10724 35084
rect 10556 34916 10612 34926
rect 10556 34822 10612 34860
rect 10668 34804 10724 34814
rect 10668 34468 10724 34748
rect 10556 34412 10724 34468
rect 10556 34244 10612 34412
rect 10556 34178 10612 34188
rect 10668 34244 10724 34254
rect 10780 34244 10836 35644
rect 11340 35028 11396 36204
rect 11340 34962 11396 34972
rect 11452 34916 11508 36652
rect 11564 36484 11620 38612
rect 12236 38050 12292 38612
rect 12236 37998 12238 38050
rect 12290 37998 12292 38050
rect 12236 37986 12292 37998
rect 12796 37828 12852 37838
rect 12796 37734 12852 37772
rect 12012 37492 12068 37502
rect 12012 37378 12068 37436
rect 12012 37326 12014 37378
rect 12066 37326 12068 37378
rect 12012 37314 12068 37326
rect 12908 37266 12964 39452
rect 12908 37214 12910 37266
rect 12962 37214 12964 37266
rect 12908 37202 12964 37214
rect 13020 38052 13076 38062
rect 12908 36596 12964 36606
rect 12684 36540 12908 36596
rect 11676 36484 11732 36494
rect 11564 36428 11676 36484
rect 11676 36390 11732 36428
rect 12348 36484 12404 36494
rect 12348 36390 12404 36428
rect 11788 36260 11844 36270
rect 11788 36166 11844 36204
rect 12012 36260 12068 36270
rect 12012 36258 12180 36260
rect 12012 36206 12014 36258
rect 12066 36206 12180 36258
rect 12012 36204 12180 36206
rect 12012 36194 12068 36204
rect 11452 34850 11508 34860
rect 10668 34242 10836 34244
rect 10668 34190 10670 34242
rect 10722 34190 10836 34242
rect 10668 34188 10836 34190
rect 10668 33460 10724 34188
rect 11340 34132 11396 34142
rect 11340 34038 11396 34076
rect 10668 33394 10724 33404
rect 11564 34020 11620 34030
rect 12012 34020 12068 34030
rect 11564 33346 11620 33964
rect 11900 34018 12068 34020
rect 11900 33966 12014 34018
rect 12066 33966 12068 34018
rect 11900 33964 12068 33966
rect 11564 33294 11566 33346
rect 11618 33294 11620 33346
rect 11564 33282 11620 33294
rect 11788 33460 11844 33470
rect 10444 33182 10446 33234
rect 10498 33182 10500 33234
rect 10444 33170 10500 33182
rect 10108 32582 10164 32620
rect 11676 32676 11732 32686
rect 10220 32564 10276 32574
rect 10220 32470 10276 32508
rect 10332 31892 10388 31902
rect 10108 31780 10164 31790
rect 10108 31686 10164 31724
rect 10332 31778 10388 31836
rect 10332 31726 10334 31778
rect 10386 31726 10388 31778
rect 10332 31714 10388 31726
rect 11676 31666 11732 32620
rect 11788 31778 11844 33404
rect 11900 32562 11956 33964
rect 12012 33954 12068 33964
rect 11900 32510 11902 32562
rect 11954 32510 11956 32562
rect 11900 32498 11956 32510
rect 12012 31892 12068 31902
rect 12012 31798 12068 31836
rect 11788 31726 11790 31778
rect 11842 31726 11844 31778
rect 11788 31714 11844 31726
rect 11676 31614 11678 31666
rect 11730 31614 11732 31666
rect 11676 31602 11732 31614
rect 10220 31556 10276 31566
rect 10220 31462 10276 31500
rect 11452 31220 11508 31230
rect 10220 31108 10276 31118
rect 10220 31014 10276 31052
rect 9996 30382 9998 30434
rect 10050 30382 10052 30434
rect 9996 30370 10052 30382
rect 10668 30994 10724 31006
rect 10668 30942 10670 30994
rect 10722 30942 10724 30994
rect 9660 30322 9716 30334
rect 9660 30270 9662 30322
rect 9714 30270 9716 30322
rect 9660 29764 9716 30270
rect 10108 30212 10164 30222
rect 10108 30118 10164 30156
rect 10668 30212 10724 30942
rect 10892 30212 10948 30222
rect 10668 30210 10948 30212
rect 10668 30158 10894 30210
rect 10946 30158 10948 30210
rect 10668 30156 10948 30158
rect 10668 30100 10724 30156
rect 10892 30146 10948 30156
rect 11452 30212 11508 31164
rect 11788 30996 11844 31006
rect 11788 30902 11844 30940
rect 12124 30882 12180 36204
rect 12348 35924 12404 35934
rect 12348 34242 12404 35868
rect 12684 35922 12740 36540
rect 12908 36502 12964 36540
rect 13020 35924 13076 37996
rect 12684 35870 12686 35922
rect 12738 35870 12740 35922
rect 12684 35700 12740 35870
rect 12684 35634 12740 35644
rect 12796 35922 13076 35924
rect 12796 35870 13022 35922
rect 13074 35870 13076 35922
rect 12796 35868 13076 35870
rect 12796 34804 12852 35868
rect 13020 35858 13076 35868
rect 12908 35700 12964 35710
rect 12908 35606 12964 35644
rect 12796 34738 12852 34748
rect 13020 35474 13076 35486
rect 13020 35422 13022 35474
rect 13074 35422 13076 35474
rect 13020 34804 13076 35422
rect 13020 34738 13076 34748
rect 12348 34190 12350 34242
rect 12402 34190 12404 34242
rect 12348 34178 12404 34190
rect 12460 33906 12516 33918
rect 12460 33854 12462 33906
rect 12514 33854 12516 33906
rect 12460 33460 12516 33854
rect 12348 33404 12516 33460
rect 12796 33460 12852 33470
rect 12348 32450 12404 33404
rect 12796 33366 12852 33404
rect 12348 32398 12350 32450
rect 12402 32398 12404 32450
rect 12348 32386 12404 32398
rect 12460 31108 12516 31118
rect 12460 31014 12516 31052
rect 12124 30830 12126 30882
rect 12178 30830 12180 30882
rect 12124 30818 12180 30830
rect 13244 30884 13300 40124
rect 13356 37716 13412 40572
rect 13692 39730 13748 41020
rect 13916 41010 13972 41020
rect 13692 39678 13694 39730
rect 13746 39678 13748 39730
rect 13692 39666 13748 39678
rect 14028 40516 14084 40526
rect 13804 39060 13860 39070
rect 13804 38834 13860 39004
rect 13804 38782 13806 38834
rect 13858 38782 13860 38834
rect 13804 38770 13860 38782
rect 14028 38722 14084 40460
rect 14028 38670 14030 38722
rect 14082 38670 14084 38722
rect 13356 37650 13412 37660
rect 13468 38612 13524 38622
rect 13468 37490 13524 38556
rect 13916 38388 13972 38398
rect 13580 38164 13636 38174
rect 13636 38108 13860 38164
rect 13580 38070 13636 38108
rect 13468 37438 13470 37490
rect 13522 37438 13524 37490
rect 13468 37426 13524 37438
rect 13804 37268 13860 38108
rect 13916 37492 13972 38332
rect 14028 38164 14084 38670
rect 14140 38836 14196 38846
rect 14140 38164 14196 38780
rect 14252 38610 14308 38622
rect 14252 38558 14254 38610
rect 14306 38558 14308 38610
rect 14252 38388 14308 38558
rect 14252 38322 14308 38332
rect 14364 38610 14420 38622
rect 14364 38558 14366 38610
rect 14418 38558 14420 38610
rect 14252 38164 14308 38174
rect 14140 38162 14308 38164
rect 14140 38110 14254 38162
rect 14306 38110 14308 38162
rect 14140 38108 14308 38110
rect 14028 38098 14084 38108
rect 13916 37426 13972 37436
rect 14028 37380 14084 37390
rect 14028 37286 14084 37324
rect 13916 37268 13972 37278
rect 13804 37266 13972 37268
rect 13804 37214 13918 37266
rect 13970 37214 13972 37266
rect 13804 37212 13972 37214
rect 13804 36596 13860 37212
rect 13916 37202 13972 37212
rect 13804 36482 13860 36540
rect 13804 36430 13806 36482
rect 13858 36430 13860 36482
rect 13804 36418 13860 36430
rect 13580 35922 13636 35934
rect 13580 35870 13582 35922
rect 13634 35870 13636 35922
rect 13580 35812 13636 35870
rect 13692 35812 13748 35822
rect 13580 35756 13692 35812
rect 13692 35746 13748 35756
rect 13468 35698 13524 35710
rect 13468 35646 13470 35698
rect 13522 35646 13524 35698
rect 13468 35364 13524 35646
rect 13804 35700 13860 35710
rect 13804 35606 13860 35644
rect 14252 35586 14308 38108
rect 14364 37940 14420 38558
rect 14364 37874 14420 37884
rect 14364 36596 14420 36606
rect 14476 36596 14532 41132
rect 14588 41186 14644 42478
rect 14588 41134 14590 41186
rect 14642 41134 14644 41186
rect 14588 41122 14644 41134
rect 14588 40516 14644 40526
rect 14588 40422 14644 40460
rect 14588 37492 14644 37502
rect 14588 37378 14644 37436
rect 14588 37326 14590 37378
rect 14642 37326 14644 37378
rect 14588 37314 14644 37326
rect 14364 36594 14476 36596
rect 14364 36542 14366 36594
rect 14418 36542 14476 36594
rect 14364 36540 14476 36542
rect 14364 36530 14420 36540
rect 14476 36502 14532 36540
rect 14700 36708 14756 47068
rect 14812 46004 14868 46014
rect 14812 43762 14868 45948
rect 15484 46004 15540 49086
rect 16044 49140 16100 51100
rect 17500 50818 17556 51212
rect 17500 50766 17502 50818
rect 17554 50766 17556 50818
rect 17500 50754 17556 50766
rect 17388 50706 17444 50718
rect 17388 50654 17390 50706
rect 17442 50654 17444 50706
rect 16828 50596 16884 50606
rect 16828 50502 16884 50540
rect 16156 49140 16212 49150
rect 16044 49138 16212 49140
rect 16044 49086 16158 49138
rect 16210 49086 16212 49138
rect 16044 49084 16212 49086
rect 15932 48468 15988 48478
rect 15932 47572 15988 48412
rect 16156 48244 16212 49084
rect 16380 49028 16436 49038
rect 16380 48934 16436 48972
rect 17052 48916 17108 48926
rect 17052 48822 17108 48860
rect 16716 48466 16772 48478
rect 16716 48414 16718 48466
rect 16770 48414 16772 48466
rect 16156 48242 16660 48244
rect 16156 48190 16158 48242
rect 16210 48190 16660 48242
rect 16156 48188 16660 48190
rect 16156 48178 16212 48188
rect 15932 47458 15988 47516
rect 15932 47406 15934 47458
rect 15986 47406 15988 47458
rect 15932 47394 15988 47406
rect 16380 47796 16436 47806
rect 16380 47572 16436 47740
rect 15596 47346 15652 47358
rect 15596 47294 15598 47346
rect 15650 47294 15652 47346
rect 15596 47236 15652 47294
rect 15596 46900 15652 47180
rect 16044 46900 16100 46910
rect 15596 46898 16100 46900
rect 15596 46846 16046 46898
rect 16098 46846 16100 46898
rect 15596 46844 16100 46846
rect 16044 46834 16100 46844
rect 16268 46786 16324 46798
rect 16268 46734 16270 46786
rect 16322 46734 16324 46786
rect 16268 46564 16324 46734
rect 16380 46786 16436 47516
rect 16604 47458 16660 48188
rect 16604 47406 16606 47458
rect 16658 47406 16660 47458
rect 16604 47394 16660 47406
rect 16380 46734 16382 46786
rect 16434 46734 16436 46786
rect 16380 46722 16436 46734
rect 16716 46788 16772 48414
rect 17388 48468 17444 50654
rect 17948 50596 18004 51324
rect 18956 51378 19012 52108
rect 19740 52162 19796 52220
rect 19740 52110 19742 52162
rect 19794 52110 19796 52162
rect 19740 52098 19796 52110
rect 20188 52164 20244 52174
rect 20188 52070 20244 52108
rect 18956 51326 18958 51378
rect 19010 51326 19012 51378
rect 18956 51314 19012 51326
rect 19292 52050 19348 52062
rect 19292 51998 19294 52050
rect 19346 51998 19348 52050
rect 19180 51154 19236 51166
rect 19180 51102 19182 51154
rect 19234 51102 19236 51154
rect 18172 50596 18228 50606
rect 17948 50594 18228 50596
rect 17948 50542 18174 50594
rect 18226 50542 18228 50594
rect 17948 50540 18228 50542
rect 18172 50530 18228 50540
rect 18396 50482 18452 50494
rect 18396 50430 18398 50482
rect 18450 50430 18452 50482
rect 18396 49028 18452 50430
rect 18508 50484 18564 50494
rect 18508 50390 18564 50428
rect 19180 49810 19236 51102
rect 19292 50428 19348 51998
rect 19628 52050 19684 52062
rect 20636 52052 20692 52892
rect 20748 52836 20804 52846
rect 20748 52742 20804 52780
rect 21308 52836 21364 53566
rect 21308 52770 21364 52780
rect 21420 53618 21588 53620
rect 21420 53566 21534 53618
rect 21586 53566 21588 53618
rect 21420 53564 21588 53566
rect 21308 52500 21364 52510
rect 21308 52162 21364 52444
rect 21308 52110 21310 52162
rect 21362 52110 21364 52162
rect 21308 52098 21364 52110
rect 19628 51998 19630 52050
rect 19682 51998 19684 52050
rect 19628 51604 19684 51998
rect 20412 51996 20692 52052
rect 21196 52052 21252 52062
rect 19836 51772 20100 51782
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 19836 51706 20100 51716
rect 19628 51548 20020 51604
rect 19964 51378 20020 51548
rect 19964 51326 19966 51378
rect 20018 51326 20020 51378
rect 19964 51314 20020 51326
rect 20076 51492 20132 51502
rect 20076 50594 20132 51436
rect 20076 50542 20078 50594
rect 20130 50542 20132 50594
rect 20076 50530 20132 50542
rect 20300 51378 20356 51390
rect 20300 51326 20302 51378
rect 20354 51326 20356 51378
rect 20300 50596 20356 51326
rect 20300 50530 20356 50540
rect 20412 50594 20468 51996
rect 20636 51604 20692 51614
rect 20636 51510 20692 51548
rect 21196 51602 21252 51996
rect 21420 51716 21476 53564
rect 21532 53554 21588 53564
rect 21756 53506 21812 53518
rect 21756 53454 21758 53506
rect 21810 53454 21812 53506
rect 21532 53060 21588 53070
rect 21532 52966 21588 53004
rect 21644 52052 21700 52062
rect 21532 51940 21588 51950
rect 21532 51846 21588 51884
rect 21196 51550 21198 51602
rect 21250 51550 21252 51602
rect 21196 51538 21252 51550
rect 21308 51660 21476 51716
rect 21532 51716 21588 51726
rect 20412 50542 20414 50594
rect 20466 50542 20468 50594
rect 20412 50530 20468 50542
rect 20524 51490 20580 51502
rect 20524 51438 20526 51490
rect 20578 51438 20580 51490
rect 20524 51268 20580 51438
rect 20860 51492 20916 51502
rect 20860 51398 20916 51436
rect 21308 51380 21364 51660
rect 20972 51324 21364 51380
rect 21532 51378 21588 51660
rect 21644 51604 21700 51996
rect 21644 51510 21700 51548
rect 21532 51326 21534 51378
rect 21586 51326 21588 51378
rect 20972 51268 21028 51324
rect 20524 51212 21028 51268
rect 20524 50428 20580 51212
rect 19292 50372 19460 50428
rect 19180 49758 19182 49810
rect 19234 49758 19236 49810
rect 19180 49746 19236 49758
rect 19292 49812 19348 49822
rect 18508 49028 18564 49038
rect 19292 49028 19348 49756
rect 19404 49140 19460 50372
rect 20188 50372 20580 50428
rect 20188 50370 20244 50372
rect 20188 50318 20190 50370
rect 20242 50318 20244 50370
rect 20188 50306 20244 50318
rect 19836 50204 20100 50214
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 19836 50138 20100 50148
rect 20860 50036 20916 51212
rect 20748 50034 20916 50036
rect 20748 49982 20862 50034
rect 20914 49982 20916 50034
rect 20748 49980 20916 49982
rect 20188 49924 20244 49934
rect 20188 49830 20244 49868
rect 19852 49812 19908 49822
rect 20524 49812 20580 49822
rect 19852 49810 20020 49812
rect 19852 49758 19854 49810
rect 19906 49758 20020 49810
rect 19852 49756 20020 49758
rect 19852 49746 19908 49756
rect 19404 49074 19460 49084
rect 19628 49698 19684 49710
rect 19628 49646 19630 49698
rect 19682 49646 19684 49698
rect 17388 48402 17444 48412
rect 18060 49026 18564 49028
rect 18060 48974 18510 49026
rect 18562 48974 18564 49026
rect 18060 48972 18564 48974
rect 17724 47684 17780 47694
rect 17724 47572 17780 47628
rect 17612 47570 17780 47572
rect 17612 47518 17726 47570
rect 17778 47518 17780 47570
rect 17612 47516 17780 47518
rect 17276 47460 17332 47470
rect 17276 47366 17332 47404
rect 16716 46722 16772 46732
rect 17500 47348 17556 47358
rect 16604 46676 16660 46686
rect 16604 46564 16660 46620
rect 16268 46508 16660 46564
rect 15708 46004 15764 46014
rect 15540 46002 15764 46004
rect 15540 45950 15710 46002
rect 15762 45950 15764 46002
rect 15540 45948 15764 45950
rect 15484 45910 15540 45948
rect 15708 45938 15764 45948
rect 15932 45780 15988 45790
rect 15932 45444 15988 45724
rect 15596 45220 15652 45230
rect 15484 45218 15652 45220
rect 15484 45166 15598 45218
rect 15650 45166 15652 45218
rect 15484 45164 15652 45166
rect 14812 43710 14814 43762
rect 14866 43710 14868 43762
rect 14812 43698 14868 43710
rect 14924 44882 14980 44894
rect 14924 44830 14926 44882
rect 14978 44830 14980 44882
rect 14924 43540 14980 44830
rect 14924 43474 14980 43484
rect 15484 42084 15540 45164
rect 15596 45154 15652 45164
rect 15820 45220 15876 45230
rect 15820 44882 15876 45164
rect 15932 45106 15988 45388
rect 16156 45778 16212 45790
rect 16156 45726 16158 45778
rect 16210 45726 16212 45778
rect 16156 45332 16212 45726
rect 16380 45332 16436 45342
rect 16156 45276 16380 45332
rect 16380 45238 16436 45276
rect 16604 45218 16660 46508
rect 16604 45166 16606 45218
rect 16658 45166 16660 45218
rect 16604 45108 16660 45166
rect 16716 45780 16772 45790
rect 16716 45218 16772 45724
rect 16716 45166 16718 45218
rect 16770 45166 16772 45218
rect 16716 45154 16772 45166
rect 15932 45054 15934 45106
rect 15986 45054 15988 45106
rect 15932 45042 15988 45054
rect 16044 45052 16660 45108
rect 15820 44830 15822 44882
rect 15874 44830 15876 44882
rect 15820 44322 15876 44830
rect 15820 44270 15822 44322
rect 15874 44270 15876 44322
rect 15820 44258 15876 44270
rect 15484 42018 15540 42028
rect 15596 43650 15652 43662
rect 15596 43598 15598 43650
rect 15650 43598 15652 43650
rect 15596 42868 15652 43598
rect 15708 43538 15764 43550
rect 15708 43486 15710 43538
rect 15762 43486 15764 43538
rect 15708 43428 15764 43486
rect 15708 43362 15764 43372
rect 15708 42868 15764 42878
rect 15596 42866 15764 42868
rect 15596 42814 15710 42866
rect 15762 42814 15764 42866
rect 15596 42812 15764 42814
rect 15372 41972 15428 41982
rect 15372 41878 15428 41916
rect 15484 41858 15540 41870
rect 15484 41806 15486 41858
rect 15538 41806 15540 41858
rect 15484 39730 15540 41806
rect 15596 41746 15652 42812
rect 15708 42802 15764 42812
rect 15596 41694 15598 41746
rect 15650 41694 15652 41746
rect 15596 41682 15652 41694
rect 15932 41186 15988 41198
rect 15932 41134 15934 41186
rect 15986 41134 15988 41186
rect 15484 39678 15486 39730
rect 15538 39678 15540 39730
rect 14924 39394 14980 39406
rect 14924 39342 14926 39394
rect 14978 39342 14980 39394
rect 14924 38948 14980 39342
rect 14924 38882 14980 38892
rect 15372 38836 15428 38874
rect 15372 38770 15428 38780
rect 14812 38612 14868 38622
rect 15036 38612 15092 38622
rect 14868 38610 15092 38612
rect 14868 38558 15038 38610
rect 15090 38558 15092 38610
rect 14868 38556 15092 38558
rect 14812 38546 14868 38556
rect 15036 38164 15092 38556
rect 15372 38610 15428 38622
rect 15372 38558 15374 38610
rect 15426 38558 15428 38610
rect 15036 38108 15316 38164
rect 15260 38050 15316 38108
rect 15260 37998 15262 38050
rect 15314 37998 15316 38050
rect 15260 37986 15316 37998
rect 15036 37940 15092 37950
rect 15092 37884 15204 37940
rect 15036 37874 15092 37884
rect 15148 37266 15204 37884
rect 15372 37604 15428 38558
rect 15372 37538 15428 37548
rect 15148 37214 15150 37266
rect 15202 37214 15204 37266
rect 15148 37202 15204 37214
rect 15484 37154 15540 39678
rect 15596 40404 15652 40414
rect 15932 40404 15988 41134
rect 15596 40402 15988 40404
rect 15596 40350 15598 40402
rect 15650 40350 15988 40402
rect 15596 40348 15988 40350
rect 15596 38162 15652 40348
rect 16044 40292 16100 45052
rect 17500 44996 17556 47292
rect 17612 45778 17668 47516
rect 17724 47506 17780 47516
rect 17948 47458 18004 47470
rect 17948 47406 17950 47458
rect 18002 47406 18004 47458
rect 17948 47348 18004 47406
rect 17948 47282 18004 47292
rect 18060 46898 18116 48972
rect 18508 48962 18564 48972
rect 18844 49026 19348 49028
rect 18844 48974 19294 49026
rect 19346 48974 19348 49026
rect 18844 48972 19348 48974
rect 18844 48914 18900 48972
rect 18844 48862 18846 48914
rect 18898 48862 18900 48914
rect 18844 48850 18900 48862
rect 18732 48804 18788 48814
rect 18732 48466 18788 48748
rect 18732 48414 18734 48466
rect 18786 48414 18788 48466
rect 18732 48402 18788 48414
rect 19292 48468 19348 48972
rect 19404 48914 19460 48926
rect 19404 48862 19406 48914
rect 19458 48862 19460 48914
rect 19404 48804 19460 48862
rect 19516 48916 19572 48926
rect 19516 48822 19572 48860
rect 19404 48738 19460 48748
rect 19628 48468 19684 49646
rect 19964 49250 20020 49756
rect 20524 49718 20580 49756
rect 19964 49198 19966 49250
rect 20018 49198 20020 49250
rect 19964 49186 20020 49198
rect 20188 49026 20244 49038
rect 20188 48974 20190 49026
rect 20242 48974 20244 49026
rect 20188 48916 20244 48974
rect 20188 48850 20244 48860
rect 20748 48914 20804 49980
rect 20860 49970 20916 49980
rect 21196 50708 21252 50718
rect 21196 48916 21252 50652
rect 21532 49924 21588 51326
rect 21756 51380 21812 53454
rect 21980 52276 22036 53678
rect 22316 53730 22372 53742
rect 22316 53678 22318 53730
rect 22370 53678 22372 53730
rect 21980 52210 22036 52220
rect 22092 52836 22148 52846
rect 22316 52836 22372 53678
rect 22540 53506 22596 53518
rect 22540 53454 22542 53506
rect 22594 53454 22596 53506
rect 22092 52834 22372 52836
rect 22092 52782 22094 52834
rect 22146 52782 22372 52834
rect 22092 52780 22372 52782
rect 22428 53058 22484 53070
rect 22428 53006 22430 53058
rect 22482 53006 22484 53058
rect 21868 52162 21924 52174
rect 21868 52110 21870 52162
rect 21922 52110 21924 52162
rect 21868 51828 21924 52110
rect 21980 52052 22036 52062
rect 21980 51958 22036 51996
rect 21868 51762 21924 51772
rect 21868 51604 21924 51614
rect 22092 51604 22148 52780
rect 21868 51602 22148 51604
rect 21868 51550 21870 51602
rect 21922 51550 22148 51602
rect 21868 51548 22148 51550
rect 22316 52612 22372 52622
rect 21868 51538 21924 51548
rect 22204 51380 22260 51390
rect 21756 51378 22260 51380
rect 21756 51326 22206 51378
rect 22258 51326 22260 51378
rect 21756 51324 22260 51326
rect 22204 51314 22260 51324
rect 22316 51266 22372 52556
rect 22316 51214 22318 51266
rect 22370 51214 22372 51266
rect 22316 51202 22372 51214
rect 22428 50820 22484 53006
rect 22540 52164 22596 53454
rect 22652 53060 22708 53790
rect 23884 53620 23940 53630
rect 24108 53620 24164 53630
rect 23660 53508 23716 53518
rect 22652 52994 22708 53004
rect 23548 53506 23716 53508
rect 23548 53454 23662 53506
rect 23714 53454 23716 53506
rect 23548 53452 23716 53454
rect 23436 52836 23492 52846
rect 23548 52836 23604 53452
rect 23660 53442 23716 53452
rect 23660 53060 23716 53070
rect 23660 52946 23716 53004
rect 23660 52894 23662 52946
rect 23714 52894 23716 52946
rect 23660 52882 23716 52894
rect 23492 52780 23604 52836
rect 22876 52164 22932 52174
rect 22540 52162 22932 52164
rect 22540 52110 22878 52162
rect 22930 52110 22932 52162
rect 22540 52108 22932 52110
rect 22876 52098 22932 52108
rect 23100 52162 23156 52174
rect 23100 52110 23102 52162
rect 23154 52110 23156 52162
rect 22540 51940 22596 51950
rect 22540 51490 22596 51884
rect 23100 51940 23156 52110
rect 23100 51874 23156 51884
rect 23324 52162 23380 52174
rect 23324 52110 23326 52162
rect 23378 52110 23380 52162
rect 22540 51438 22542 51490
rect 22594 51438 22596 51490
rect 22540 51426 22596 51438
rect 22540 50820 22596 50830
rect 23324 50820 23380 52110
rect 22428 50818 23380 50820
rect 22428 50766 22542 50818
rect 22594 50766 23380 50818
rect 22428 50764 23380 50766
rect 22540 50754 22596 50764
rect 21868 50652 22372 50708
rect 21868 50482 21924 50652
rect 21868 50430 21870 50482
rect 21922 50430 21924 50482
rect 21532 49858 21588 49868
rect 21644 50370 21700 50382
rect 21644 50318 21646 50370
rect 21698 50318 21700 50370
rect 21644 49922 21700 50318
rect 21644 49870 21646 49922
rect 21698 49870 21700 49922
rect 21644 49858 21700 49870
rect 20748 48862 20750 48914
rect 20802 48862 20804 48914
rect 20748 48850 20804 48862
rect 21084 48860 21252 48916
rect 21420 49698 21476 49710
rect 21420 49646 21422 49698
rect 21474 49646 21476 49698
rect 20524 48804 20580 48814
rect 20524 48710 20580 48748
rect 20860 48802 20916 48814
rect 20860 48750 20862 48802
rect 20914 48750 20916 48802
rect 19836 48636 20100 48646
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 19836 48570 20100 48580
rect 19292 48402 19348 48412
rect 19404 48412 19684 48468
rect 19852 48468 19908 48478
rect 18508 48242 18564 48254
rect 18508 48190 18510 48242
rect 18562 48190 18564 48242
rect 18508 47572 18564 48190
rect 18508 47506 18564 47516
rect 19292 48242 19348 48254
rect 19292 48190 19294 48242
rect 19346 48190 19348 48242
rect 18620 47348 18676 47358
rect 18620 47254 18676 47292
rect 19292 47348 19348 48190
rect 19292 47282 19348 47292
rect 18060 46846 18062 46898
rect 18114 46846 18116 46898
rect 17724 46676 17780 46686
rect 17724 46582 17780 46620
rect 17612 45726 17614 45778
rect 17666 45726 17668 45778
rect 17612 45220 17668 45726
rect 17836 45778 17892 45790
rect 17836 45726 17838 45778
rect 17890 45726 17892 45778
rect 17612 45154 17668 45164
rect 17724 45332 17780 45342
rect 17724 45218 17780 45276
rect 17724 45166 17726 45218
rect 17778 45166 17780 45218
rect 17724 45154 17780 45166
rect 17388 44994 17556 44996
rect 17388 44942 17502 44994
rect 17554 44942 17556 44994
rect 17388 44940 17556 44942
rect 16604 44884 16660 44894
rect 16604 43650 16660 44828
rect 17388 44546 17444 44940
rect 17500 44930 17556 44940
rect 17388 44494 17390 44546
rect 17442 44494 17444 44546
rect 17388 44482 17444 44494
rect 17836 44548 17892 45726
rect 17836 44482 17892 44492
rect 17500 44434 17556 44446
rect 17500 44382 17502 44434
rect 17554 44382 17556 44434
rect 16828 44322 16884 44334
rect 16828 44270 16830 44322
rect 16882 44270 16884 44322
rect 16828 43988 16884 44270
rect 16828 43922 16884 43932
rect 16604 43598 16606 43650
rect 16658 43598 16660 43650
rect 16268 43428 16324 43438
rect 16268 43426 16548 43428
rect 16268 43374 16270 43426
rect 16322 43374 16548 43426
rect 16268 43372 16548 43374
rect 16268 43362 16324 43372
rect 16268 42644 16324 42654
rect 16380 42644 16436 42654
rect 16268 42642 16380 42644
rect 16268 42590 16270 42642
rect 16322 42590 16380 42642
rect 16268 42588 16380 42590
rect 16268 42578 16324 42588
rect 16380 42194 16436 42588
rect 16380 42142 16382 42194
rect 16434 42142 16436 42194
rect 16380 42130 16436 42142
rect 16492 42196 16548 43372
rect 16492 42130 16548 42140
rect 16604 42194 16660 43598
rect 17500 43652 17556 44382
rect 17500 43596 18004 43652
rect 17388 43316 17444 43326
rect 16604 42142 16606 42194
rect 16658 42142 16660 42194
rect 16604 41524 16660 42142
rect 16716 42196 16772 42206
rect 16716 42082 16772 42140
rect 16716 42030 16718 42082
rect 16770 42030 16772 42082
rect 16716 42018 16772 42030
rect 16604 41468 16884 41524
rect 16716 41300 16772 41310
rect 16716 41206 16772 41244
rect 16492 41074 16548 41086
rect 16492 41022 16494 41074
rect 16546 41022 16548 41074
rect 16492 40516 16548 41022
rect 16044 40226 16100 40236
rect 16156 40460 16548 40516
rect 16604 41076 16660 41086
rect 16828 41076 16884 41468
rect 16156 40404 16212 40460
rect 16604 40404 16660 41020
rect 16156 39620 16212 40348
rect 16268 40348 16660 40404
rect 16716 41020 16884 41076
rect 16268 40290 16324 40348
rect 16268 40238 16270 40290
rect 16322 40238 16324 40290
rect 16268 40226 16324 40238
rect 16156 39554 16212 39564
rect 15820 39506 15876 39518
rect 15820 39454 15822 39506
rect 15874 39454 15876 39506
rect 15820 39172 15876 39454
rect 16268 39508 16324 39518
rect 15820 39116 16100 39172
rect 16044 39058 16100 39116
rect 16044 39006 16046 39058
rect 16098 39006 16100 39058
rect 16044 38994 16100 39006
rect 16268 39058 16324 39452
rect 16716 39172 16772 41020
rect 17388 40180 17444 43260
rect 17500 41858 17556 43596
rect 17948 43538 18004 43596
rect 17948 43486 17950 43538
rect 18002 43486 18004 43538
rect 17948 43474 18004 43486
rect 17724 43428 17780 43438
rect 17612 42644 17668 42654
rect 17724 42644 17780 43372
rect 18060 43316 18116 46846
rect 19068 47236 19124 47246
rect 18732 45780 18788 45790
rect 18732 45686 18788 45724
rect 19068 45668 19124 47180
rect 19404 47012 19460 48412
rect 19628 48244 19684 48254
rect 19628 48150 19684 48188
rect 19292 46956 19460 47012
rect 19516 48018 19572 48030
rect 19852 48020 19908 48412
rect 20860 48468 20916 48750
rect 20860 48402 20916 48412
rect 20972 48804 21028 48814
rect 20972 48466 21028 48748
rect 20972 48414 20974 48466
rect 21026 48414 21028 48466
rect 20972 48402 21028 48414
rect 19516 47966 19518 48018
rect 19570 47966 19572 48018
rect 19292 46564 19348 46956
rect 19404 46788 19460 46798
rect 19516 46788 19572 47966
rect 19628 47964 19908 48020
rect 19964 48244 20020 48254
rect 19628 47458 19684 47964
rect 19964 47572 20020 48188
rect 19628 47406 19630 47458
rect 19682 47406 19684 47458
rect 19628 47394 19684 47406
rect 19740 47516 20020 47572
rect 19740 47458 19796 47516
rect 19740 47406 19742 47458
rect 19794 47406 19796 47458
rect 19740 47236 19796 47406
rect 19852 47348 19908 47358
rect 19852 47254 19908 47292
rect 20300 47348 20356 47358
rect 20300 47254 20356 47292
rect 19740 47170 19796 47180
rect 19836 47068 20100 47078
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 19836 47002 20100 47012
rect 20300 46900 20356 46910
rect 19628 46788 19684 46798
rect 19516 46732 19628 46788
rect 19404 46694 19460 46732
rect 19628 46694 19684 46732
rect 20300 46786 20356 46844
rect 20300 46734 20302 46786
rect 20354 46734 20356 46786
rect 20300 46722 20356 46734
rect 20748 46788 20804 46798
rect 20748 46694 20804 46732
rect 20076 46676 20132 46686
rect 20188 46676 20244 46686
rect 20076 46674 20188 46676
rect 20076 46622 20078 46674
rect 20130 46622 20188 46674
rect 20076 46620 20188 46622
rect 20076 46610 20132 46620
rect 19852 46564 19908 46574
rect 19292 46562 19908 46564
rect 19292 46510 19854 46562
rect 19906 46510 19908 46562
rect 19292 46508 19908 46510
rect 19852 46498 19908 46508
rect 19068 45574 19124 45612
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 19516 45330 19572 45342
rect 19516 45278 19518 45330
rect 19570 45278 19572 45330
rect 18956 45220 19012 45230
rect 18956 45106 19012 45164
rect 18956 45054 18958 45106
rect 19010 45054 19012 45106
rect 18956 45042 19012 45054
rect 19404 44548 19460 44558
rect 19404 44322 19460 44492
rect 19404 44270 19406 44322
rect 19458 44270 19460 44322
rect 19404 44258 19460 44270
rect 19292 44100 19348 44110
rect 18620 43428 18676 43438
rect 18620 43334 18676 43372
rect 19180 43426 19236 43438
rect 19180 43374 19182 43426
rect 19234 43374 19236 43426
rect 17948 43260 18116 43316
rect 17612 42642 17780 42644
rect 17612 42590 17614 42642
rect 17666 42590 17780 42642
rect 17612 42588 17780 42590
rect 17836 42642 17892 42654
rect 17836 42590 17838 42642
rect 17890 42590 17892 42642
rect 17612 42532 17668 42588
rect 17612 42466 17668 42476
rect 17500 41806 17502 41858
rect 17554 41806 17556 41858
rect 17500 41300 17556 41806
rect 17500 41234 17556 41244
rect 17612 41186 17668 41198
rect 17612 41134 17614 41186
rect 17666 41134 17668 41186
rect 17612 41076 17668 41134
rect 17612 41010 17668 41020
rect 17836 40964 17892 42590
rect 17948 41188 18004 43260
rect 18060 42644 18116 42654
rect 18060 42082 18116 42588
rect 19180 42644 19236 43374
rect 19292 42866 19348 44044
rect 19516 43652 19572 45278
rect 20076 45332 20132 45342
rect 20188 45332 20244 46620
rect 20524 46676 20580 46686
rect 20524 46582 20580 46620
rect 20860 46676 20916 46686
rect 20860 46582 20916 46620
rect 21084 45556 21140 48860
rect 21420 48804 21476 49646
rect 21868 49364 21924 50430
rect 21980 50484 22036 50494
rect 22316 50484 22372 50652
rect 22652 50596 22708 50606
rect 22652 50502 22708 50540
rect 22540 50484 22596 50494
rect 21980 50482 22260 50484
rect 21980 50430 21982 50482
rect 22034 50430 22260 50482
rect 21980 50428 22260 50430
rect 22316 50482 22596 50484
rect 22316 50430 22542 50482
rect 22594 50430 22596 50482
rect 22316 50428 22596 50430
rect 21980 50418 22036 50428
rect 21868 49308 22148 49364
rect 21868 49138 21924 49150
rect 21868 49086 21870 49138
rect 21922 49086 21924 49138
rect 21868 49028 21924 49086
rect 21868 48962 21924 48972
rect 21980 49140 22036 49150
rect 21980 49026 22036 49084
rect 21980 48974 21982 49026
rect 22034 48974 22036 49026
rect 21980 48962 22036 48974
rect 21420 48738 21476 48748
rect 21532 48802 21588 48814
rect 21532 48750 21534 48802
rect 21586 48750 21588 48802
rect 21196 48468 21252 48478
rect 21532 48468 21588 48750
rect 21252 48412 21588 48468
rect 21756 48802 21812 48814
rect 21756 48750 21758 48802
rect 21810 48750 21812 48802
rect 21756 48468 21812 48750
rect 21756 48412 21924 48468
rect 21196 48374 21252 48412
rect 21868 48356 21924 48412
rect 21980 48356 22036 48366
rect 21868 48354 22036 48356
rect 21868 48302 21982 48354
rect 22034 48302 22036 48354
rect 21868 48300 22036 48302
rect 21308 48244 21364 48254
rect 21756 48244 21812 48254
rect 21308 48242 21812 48244
rect 21308 48190 21310 48242
rect 21362 48190 21758 48242
rect 21810 48190 21812 48242
rect 21308 48188 21812 48190
rect 21308 48178 21364 48188
rect 21756 47570 21812 48188
rect 21756 47518 21758 47570
rect 21810 47518 21812 47570
rect 21756 47506 21812 47518
rect 21196 47460 21252 47470
rect 21196 47366 21252 47404
rect 21644 47458 21700 47470
rect 21644 47406 21646 47458
rect 21698 47406 21700 47458
rect 21532 47348 21588 47358
rect 21644 47348 21700 47406
rect 21588 47292 21700 47348
rect 21532 47282 21588 47292
rect 21868 47234 21924 47246
rect 21868 47182 21870 47234
rect 21922 47182 21924 47234
rect 21868 47124 21924 47182
rect 21980 47236 22036 48300
rect 21980 47170 22036 47180
rect 21532 47068 21924 47124
rect 21420 45778 21476 45790
rect 21420 45726 21422 45778
rect 21474 45726 21476 45778
rect 21084 45500 21252 45556
rect 20076 45330 20244 45332
rect 20076 45278 20078 45330
rect 20130 45278 20244 45330
rect 20076 45276 20244 45278
rect 20524 45444 20580 45454
rect 20076 45266 20132 45276
rect 20412 45218 20468 45230
rect 20412 45166 20414 45218
rect 20466 45166 20468 45218
rect 19964 45106 20020 45118
rect 19964 45054 19966 45106
rect 20018 45054 20020 45106
rect 19964 44548 20020 45054
rect 19740 44492 20020 44548
rect 20188 45106 20244 45118
rect 20188 45054 20190 45106
rect 20242 45054 20244 45106
rect 19516 43586 19572 43596
rect 19628 44324 19684 44334
rect 19740 44324 19796 44492
rect 19628 44322 19796 44324
rect 19628 44270 19630 44322
rect 19682 44270 19796 44322
rect 19628 44268 19796 44270
rect 19852 44322 19908 44334
rect 19852 44270 19854 44322
rect 19906 44270 19908 44322
rect 19404 43428 19460 43438
rect 19404 42978 19460 43372
rect 19628 43204 19684 44268
rect 19852 44100 19908 44270
rect 19964 44324 20020 44334
rect 19964 44230 20020 44268
rect 20188 44100 20244 45054
rect 20412 44548 20468 45166
rect 20412 44482 20468 44492
rect 19908 44044 20244 44100
rect 19852 44034 19908 44044
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 20524 43762 20580 45388
rect 20524 43710 20526 43762
rect 20578 43710 20580 43762
rect 20524 43698 20580 43710
rect 20076 43652 20132 43662
rect 20076 43558 20132 43596
rect 20412 43538 20468 43550
rect 20412 43486 20414 43538
rect 20466 43486 20468 43538
rect 19740 43428 19796 43438
rect 19740 43334 19796 43372
rect 20412 43428 20468 43486
rect 19404 42926 19406 42978
rect 19458 42926 19460 42978
rect 19404 42914 19460 42926
rect 19516 43148 19684 43204
rect 19292 42814 19294 42866
rect 19346 42814 19348 42866
rect 19292 42802 19348 42814
rect 19180 42550 19236 42588
rect 18060 42030 18062 42082
rect 18114 42030 18116 42082
rect 18060 42018 18116 42030
rect 18956 42532 19012 42542
rect 18956 41970 19012 42476
rect 18956 41918 18958 41970
rect 19010 41918 19012 41970
rect 18956 41906 19012 41918
rect 18508 41188 18564 41198
rect 17948 41094 18004 41132
rect 18172 41186 18564 41188
rect 18172 41134 18510 41186
rect 18562 41134 18564 41186
rect 18172 41132 18564 41134
rect 17836 40898 17892 40908
rect 18172 40962 18228 41132
rect 18508 41122 18564 41132
rect 18732 41188 18788 41198
rect 18732 41094 18788 41132
rect 18844 41076 18900 41086
rect 18844 40982 18900 41020
rect 19292 41076 19348 41086
rect 19292 40982 19348 41020
rect 18172 40910 18174 40962
rect 18226 40910 18228 40962
rect 17388 40114 17444 40124
rect 17724 40292 17780 40302
rect 16828 39620 16884 39630
rect 16828 39526 16884 39564
rect 17500 39620 17556 39630
rect 17500 39526 17556 39564
rect 16268 39006 16270 39058
rect 16322 39006 16324 39058
rect 15932 38948 15988 38958
rect 15932 38854 15988 38892
rect 15596 38110 15598 38162
rect 15650 38110 15652 38162
rect 15596 38098 15652 38110
rect 15932 38050 15988 38062
rect 15932 37998 15934 38050
rect 15986 37998 15988 38050
rect 15596 37828 15652 37838
rect 15596 37268 15652 37772
rect 15932 37492 15988 37998
rect 15932 37426 15988 37436
rect 15596 37174 15652 37212
rect 15708 37378 15764 37390
rect 15708 37326 15710 37378
rect 15762 37326 15764 37378
rect 15484 37102 15486 37154
rect 15538 37102 15540 37154
rect 15484 37090 15540 37102
rect 15708 37156 15764 37326
rect 16268 37380 16324 39006
rect 16380 39116 16996 39172
rect 16380 38948 16436 39116
rect 16940 39060 16996 39116
rect 17388 39060 17444 39070
rect 16940 39058 17388 39060
rect 16940 39006 16942 39058
rect 16994 39006 17388 39058
rect 16940 39004 17388 39006
rect 16940 38994 16996 39004
rect 17388 38966 17444 39004
rect 16380 38854 16436 38892
rect 17724 38948 17780 40236
rect 18172 39732 18228 40910
rect 18284 40962 18340 40974
rect 18284 40910 18286 40962
rect 18338 40910 18340 40962
rect 18284 40516 18340 40910
rect 19068 40964 19124 40974
rect 19068 40628 19124 40908
rect 18284 40450 18340 40460
rect 18620 40514 18676 40526
rect 18620 40462 18622 40514
rect 18674 40462 18676 40514
rect 17836 39508 17892 39518
rect 17836 39414 17892 39452
rect 18172 39506 18228 39676
rect 18508 40402 18564 40414
rect 18508 40350 18510 40402
rect 18562 40350 18564 40402
rect 18508 39620 18564 40350
rect 18620 39620 18676 40462
rect 19068 40514 19124 40572
rect 19516 40626 19572 43148
rect 20412 43092 20468 43372
rect 20748 43538 20804 43550
rect 20748 43486 20750 43538
rect 20802 43486 20804 43538
rect 20412 43036 20692 43092
rect 20524 42644 20580 42654
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 20524 42084 20580 42588
rect 20636 42642 20692 43036
rect 20636 42590 20638 42642
rect 20690 42590 20692 42642
rect 20636 42578 20692 42590
rect 20748 42532 20804 43486
rect 21084 43428 21140 43438
rect 20860 43426 21140 43428
rect 20860 43374 21086 43426
rect 21138 43374 21140 43426
rect 20860 43372 21140 43374
rect 20860 42754 20916 43372
rect 21084 43362 21140 43372
rect 20860 42702 20862 42754
rect 20914 42702 20916 42754
rect 20860 42690 20916 42702
rect 20748 42466 20804 42476
rect 20076 42028 20580 42084
rect 19628 41858 19684 41870
rect 19628 41806 19630 41858
rect 19682 41806 19684 41858
rect 19628 41186 19684 41806
rect 20076 41298 20132 42028
rect 20076 41246 20078 41298
rect 20130 41246 20132 41298
rect 20076 41234 20132 41246
rect 19628 41134 19630 41186
rect 19682 41134 19684 41186
rect 19628 41122 19684 41134
rect 19964 41076 20020 41086
rect 19964 40982 20020 41020
rect 20188 40962 20244 40974
rect 20188 40910 20190 40962
rect 20242 40910 20244 40962
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 19516 40574 19518 40626
rect 19570 40574 19572 40626
rect 19516 40562 19572 40574
rect 19852 40628 19908 40638
rect 20188 40628 20244 40910
rect 21196 40740 21252 45500
rect 21308 44324 21364 44334
rect 21308 44230 21364 44268
rect 21420 42756 21476 45726
rect 21532 45444 21588 47068
rect 22092 47012 22148 49308
rect 22204 48692 22260 50428
rect 22540 50418 22596 50428
rect 23436 50148 23492 52780
rect 23884 52612 23940 53564
rect 23996 53618 24164 53620
rect 23996 53566 24110 53618
rect 24162 53566 24164 53618
rect 23996 53564 24164 53566
rect 23996 52836 24052 53564
rect 24108 53554 24164 53564
rect 24444 53618 24500 53630
rect 24444 53566 24446 53618
rect 24498 53566 24500 53618
rect 24332 53508 24388 53518
rect 24332 53414 24388 53452
rect 24444 52946 24500 53566
rect 24556 53284 24612 56142
rect 24668 55522 24724 57372
rect 24892 56754 24948 59200
rect 24892 56702 24894 56754
rect 24946 56702 24948 56754
rect 24892 56306 24948 56702
rect 24892 56254 24894 56306
rect 24946 56254 24948 56306
rect 24892 56242 24948 56254
rect 25116 56642 25172 56654
rect 25116 56590 25118 56642
rect 25170 56590 25172 56642
rect 24668 55470 24670 55522
rect 24722 55470 24724 55522
rect 24668 55458 24724 55470
rect 25004 53732 25060 53742
rect 24780 53730 25060 53732
rect 24780 53678 25006 53730
rect 25058 53678 25060 53730
rect 24780 53676 25060 53678
rect 24556 53228 24724 53284
rect 24444 52894 24446 52946
rect 24498 52894 24500 52946
rect 23996 52770 24052 52780
rect 24108 52836 24164 52846
rect 24108 52834 24388 52836
rect 24108 52782 24110 52834
rect 24162 52782 24388 52834
rect 24108 52780 24388 52782
rect 24108 52770 24164 52780
rect 23884 52546 23940 52556
rect 22204 48356 22260 48636
rect 22428 50092 23492 50148
rect 24220 52162 24276 52174
rect 24220 52110 24222 52162
rect 24274 52110 24276 52162
rect 24220 50594 24276 52110
rect 24332 52164 24388 52780
rect 24444 52612 24500 52894
rect 24556 53058 24612 53070
rect 24556 53006 24558 53058
rect 24610 53006 24612 53058
rect 24556 52836 24612 53006
rect 24556 52770 24612 52780
rect 24668 52612 24724 53228
rect 24780 53170 24836 53676
rect 25004 53666 25060 53676
rect 25116 53508 25172 56590
rect 25564 55970 25620 59200
rect 25564 55918 25566 55970
rect 25618 55918 25620 55970
rect 25564 55906 25620 55918
rect 26236 54740 26292 59200
rect 26908 55468 26964 59200
rect 27580 55972 27636 59200
rect 27804 56084 27860 56094
rect 27804 56082 27972 56084
rect 27804 56030 27806 56082
rect 27858 56030 27972 56082
rect 27804 56028 27972 56030
rect 27804 56018 27860 56028
rect 27580 55906 27636 55916
rect 26908 55412 27412 55468
rect 27468 55412 27524 55422
rect 27356 55356 27468 55412
rect 27020 55300 27076 55310
rect 27020 55298 27188 55300
rect 27020 55246 27022 55298
rect 27074 55246 27188 55298
rect 27020 55244 27188 55246
rect 27020 55234 27076 55244
rect 26460 54740 26516 54750
rect 26236 54738 26516 54740
rect 26236 54686 26238 54738
rect 26290 54686 26462 54738
rect 26514 54686 26516 54738
rect 26236 54684 26516 54686
rect 26236 54674 26292 54684
rect 26460 54674 26516 54684
rect 26908 54404 26964 54414
rect 27132 54404 27188 55244
rect 27468 55298 27524 55356
rect 27468 55246 27470 55298
rect 27522 55246 27524 55298
rect 27468 55234 27524 55246
rect 27692 55074 27748 55086
rect 27692 55022 27694 55074
rect 27746 55022 27748 55074
rect 27468 54404 27524 54414
rect 26908 54402 27076 54404
rect 26908 54350 26910 54402
rect 26962 54350 27076 54402
rect 26908 54348 27076 54350
rect 27132 54402 27524 54404
rect 27132 54350 27470 54402
rect 27522 54350 27524 54402
rect 27132 54348 27524 54350
rect 26908 54338 26964 54348
rect 25228 53842 25284 53854
rect 25228 53790 25230 53842
rect 25282 53790 25284 53842
rect 25228 53620 25284 53790
rect 25228 53554 25284 53564
rect 25900 53620 25956 53630
rect 25900 53618 26292 53620
rect 25900 53566 25902 53618
rect 25954 53566 26292 53618
rect 25900 53564 26292 53566
rect 25900 53554 25956 53564
rect 24780 53118 24782 53170
rect 24834 53118 24836 53170
rect 24780 53106 24836 53118
rect 25004 53452 25172 53508
rect 25676 53508 25732 53518
rect 24444 52556 24612 52612
rect 24668 52556 24836 52612
rect 24444 52164 24500 52174
rect 24332 52162 24500 52164
rect 24332 52110 24446 52162
rect 24498 52110 24500 52162
rect 24332 52108 24500 52110
rect 24332 50706 24388 52108
rect 24444 52098 24500 52108
rect 24556 52164 24612 52556
rect 24668 52388 24724 52398
rect 24668 52294 24724 52332
rect 24556 51940 24612 52108
rect 24444 51884 24612 51940
rect 24444 51490 24500 51884
rect 24780 51716 24836 52556
rect 24668 51660 24836 51716
rect 24444 51438 24446 51490
rect 24498 51438 24500 51490
rect 24444 51426 24500 51438
rect 24556 51490 24612 51502
rect 24556 51438 24558 51490
rect 24610 51438 24612 51490
rect 24332 50654 24334 50706
rect 24386 50654 24388 50706
rect 24332 50642 24388 50654
rect 24220 50542 24222 50594
rect 24274 50542 24276 50594
rect 22428 49026 22484 50092
rect 22428 48974 22430 49026
rect 22482 48974 22484 49026
rect 22316 48356 22372 48366
rect 22204 48354 22372 48356
rect 22204 48302 22318 48354
rect 22370 48302 22372 48354
rect 22204 48300 22372 48302
rect 22316 48290 22372 48300
rect 21644 46956 22148 47012
rect 21644 46674 21700 46956
rect 21644 46622 21646 46674
rect 21698 46622 21700 46674
rect 21644 46610 21700 46622
rect 21756 45778 21812 46956
rect 21756 45726 21758 45778
rect 21810 45726 21812 45778
rect 21756 45714 21812 45726
rect 21868 46786 21924 46798
rect 21868 46734 21870 46786
rect 21922 46734 21924 46786
rect 21868 45780 21924 46734
rect 22092 46002 22148 46956
rect 22316 47236 22372 47246
rect 22428 47236 22484 48974
rect 22652 49924 22708 49934
rect 22652 49026 22708 49868
rect 22988 49810 23044 49822
rect 22988 49758 22990 49810
rect 23042 49758 23044 49810
rect 22988 49140 23044 49758
rect 23548 49700 23604 49710
rect 23548 49698 24164 49700
rect 23548 49646 23550 49698
rect 23602 49646 24164 49698
rect 23548 49644 24164 49646
rect 23548 49634 23604 49644
rect 22988 49074 23044 49084
rect 22652 48974 22654 49026
rect 22706 48974 22708 49026
rect 22652 48962 22708 48974
rect 22876 49028 22932 49038
rect 22876 48934 22932 48972
rect 23324 49028 23380 49038
rect 23548 49028 23604 49038
rect 24108 49028 24164 49644
rect 24220 49138 24276 50542
rect 24556 50484 24612 51438
rect 24556 50418 24612 50428
rect 24220 49086 24222 49138
rect 24274 49086 24276 49138
rect 24220 49074 24276 49086
rect 23324 49026 23604 49028
rect 23324 48974 23326 49026
rect 23378 48974 23550 49026
rect 23602 48974 23604 49026
rect 23324 48972 23604 48974
rect 23324 48962 23380 48972
rect 23548 48962 23604 48972
rect 23996 49026 24164 49028
rect 23996 48974 24110 49026
rect 24162 48974 24164 49026
rect 23996 48972 24164 48974
rect 22540 48914 22596 48926
rect 22540 48862 22542 48914
rect 22594 48862 22596 48914
rect 22540 48468 22596 48862
rect 22652 48468 22708 48478
rect 22540 48412 22652 48468
rect 22652 48374 22708 48412
rect 23996 47570 24052 48972
rect 24108 48962 24164 48972
rect 23996 47518 23998 47570
rect 24050 47518 24052 47570
rect 23996 47506 24052 47518
rect 24220 48914 24276 48926
rect 24220 48862 24222 48914
rect 24274 48862 24276 48914
rect 22764 47460 22820 47470
rect 22316 47234 22484 47236
rect 22316 47182 22318 47234
rect 22370 47182 22484 47234
rect 22316 47180 22484 47182
rect 22540 47458 22820 47460
rect 22540 47406 22766 47458
rect 22818 47406 22820 47458
rect 22540 47404 22820 47406
rect 22204 46676 22260 46686
rect 22204 46582 22260 46620
rect 22316 46452 22372 47180
rect 22428 46898 22484 46910
rect 22428 46846 22430 46898
rect 22482 46846 22484 46898
rect 22428 46564 22484 46846
rect 22540 46900 22596 47404
rect 22764 47394 22820 47404
rect 24220 47458 24276 48862
rect 24220 47406 24222 47458
rect 24274 47406 24276 47458
rect 22540 46834 22596 46844
rect 22652 47236 22708 47246
rect 22652 47124 22708 47180
rect 23100 47234 23156 47246
rect 23324 47236 23380 47246
rect 23100 47182 23102 47234
rect 23154 47182 23156 47234
rect 23100 47124 23156 47182
rect 22652 47068 23156 47124
rect 23212 47234 23380 47236
rect 23212 47182 23326 47234
rect 23378 47182 23380 47234
rect 23212 47180 23380 47182
rect 22428 46498 22484 46508
rect 22540 46676 22596 46686
rect 22652 46676 22708 47068
rect 23212 46900 23268 47180
rect 23324 47170 23380 47180
rect 23436 47234 23492 47246
rect 23436 47182 23438 47234
rect 23490 47182 23492 47234
rect 22540 46674 22708 46676
rect 22540 46622 22542 46674
rect 22594 46622 22708 46674
rect 22540 46620 22708 46622
rect 22764 46844 23268 46900
rect 22764 46786 22820 46844
rect 22764 46734 22766 46786
rect 22818 46734 22820 46786
rect 22092 45950 22094 46002
rect 22146 45950 22148 46002
rect 22092 45938 22148 45950
rect 22204 46396 22372 46452
rect 22204 45780 22260 46396
rect 21868 45724 22260 45780
rect 22316 45890 22372 45902
rect 22316 45838 22318 45890
rect 22370 45838 22372 45890
rect 21532 44546 21588 45388
rect 21868 45332 21924 45724
rect 22316 45668 22372 45838
rect 22316 45602 22372 45612
rect 21868 45266 21924 45276
rect 22540 45108 22596 46620
rect 22652 46116 22708 46126
rect 22764 46116 22820 46734
rect 22652 46114 22820 46116
rect 22652 46062 22654 46114
rect 22706 46062 22820 46114
rect 22652 46060 22820 46062
rect 22652 46050 22708 46060
rect 23100 46002 23156 46844
rect 23100 45950 23102 46002
rect 23154 45950 23156 46002
rect 23100 45938 23156 45950
rect 23324 46676 23380 46686
rect 23100 45108 23156 45118
rect 22540 45106 23156 45108
rect 22540 45054 23102 45106
rect 23154 45054 23156 45106
rect 22540 45052 23156 45054
rect 23100 45042 23156 45052
rect 23324 45106 23380 46620
rect 23436 46674 23492 47182
rect 24220 46786 24276 47406
rect 24220 46734 24222 46786
rect 24274 46734 24276 46786
rect 24220 46722 24276 46734
rect 23436 46622 23438 46674
rect 23490 46622 23492 46674
rect 23436 46610 23492 46622
rect 23772 46674 23828 46686
rect 23772 46622 23774 46674
rect 23826 46622 23828 46674
rect 23660 46564 23716 46574
rect 23660 46470 23716 46508
rect 23324 45054 23326 45106
rect 23378 45054 23380 45106
rect 23324 45042 23380 45054
rect 23436 46452 23492 46462
rect 21532 44494 21534 44546
rect 21586 44494 21588 44546
rect 21532 44482 21588 44494
rect 21756 44322 21812 44334
rect 21756 44270 21758 44322
rect 21810 44270 21812 44322
rect 21644 43652 21700 43662
rect 21756 43652 21812 44270
rect 21868 44324 21924 44334
rect 23100 44324 23156 44334
rect 21868 44322 23156 44324
rect 21868 44270 21870 44322
rect 21922 44270 23102 44322
rect 23154 44270 23156 44322
rect 21868 44268 23156 44270
rect 21868 44258 21924 44268
rect 23100 44258 23156 44268
rect 21644 43650 21812 43652
rect 21644 43598 21646 43650
rect 21698 43598 21812 43650
rect 21644 43596 21812 43598
rect 22540 43652 22596 43662
rect 21644 42756 21700 43596
rect 22540 43538 22596 43596
rect 22540 43486 22542 43538
rect 22594 43486 22596 43538
rect 22540 43474 22596 43486
rect 22988 43092 23044 43102
rect 21868 42756 21924 42766
rect 21644 42754 21924 42756
rect 21644 42702 21870 42754
rect 21922 42702 21924 42754
rect 21644 42700 21924 42702
rect 21308 42644 21364 42654
rect 21308 42550 21364 42588
rect 21308 40740 21364 40750
rect 21196 40684 21308 40740
rect 21308 40674 21364 40684
rect 19068 40462 19070 40514
rect 19122 40462 19124 40514
rect 19068 40450 19124 40462
rect 19292 40516 19348 40526
rect 19292 40422 19348 40460
rect 18844 40404 18900 40414
rect 18844 40310 18900 40348
rect 19740 40404 19796 40414
rect 19740 40310 19796 40348
rect 19852 40402 19908 40572
rect 19852 40350 19854 40402
rect 19906 40350 19908 40402
rect 19852 40338 19908 40350
rect 19964 40572 20244 40628
rect 20524 40628 20580 40638
rect 19964 40180 20020 40572
rect 20524 40534 20580 40572
rect 20412 40516 20468 40526
rect 20412 40422 20468 40460
rect 20188 40404 20244 40414
rect 20188 40310 20244 40348
rect 21308 40404 21364 40414
rect 21420 40404 21476 42700
rect 21868 42690 21924 42700
rect 22092 42756 22148 42766
rect 22092 42642 22148 42700
rect 22092 42590 22094 42642
rect 22146 42590 22148 42642
rect 22092 42578 22148 42590
rect 22204 42642 22260 42654
rect 22204 42590 22206 42642
rect 22258 42590 22260 42642
rect 21644 42532 21700 42542
rect 22204 42532 22260 42590
rect 22652 42532 22708 42542
rect 22204 42530 22708 42532
rect 22204 42478 22654 42530
rect 22706 42478 22708 42530
rect 22204 42476 22708 42478
rect 21644 41972 21700 42476
rect 22652 42420 22708 42476
rect 22652 42354 22708 42364
rect 22876 42196 22932 42206
rect 22092 42194 22932 42196
rect 22092 42142 22878 42194
rect 22930 42142 22932 42194
rect 22092 42140 22932 42142
rect 22092 41972 22148 42140
rect 21532 41300 21588 41310
rect 21644 41300 21700 41916
rect 21868 41970 22148 41972
rect 21868 41918 22094 41970
rect 22146 41918 22148 41970
rect 21868 41916 22148 41918
rect 21532 41298 21700 41300
rect 21532 41246 21534 41298
rect 21586 41246 21700 41298
rect 21532 41244 21700 41246
rect 21756 41524 21812 41534
rect 21532 41234 21588 41244
rect 21756 41186 21812 41468
rect 21756 41134 21758 41186
rect 21810 41134 21812 41186
rect 21756 40628 21812 41134
rect 21756 40562 21812 40572
rect 21868 40626 21924 41916
rect 22092 41906 22148 41916
rect 22204 41972 22260 41982
rect 22204 41878 22260 41916
rect 22540 41970 22596 41982
rect 22540 41918 22542 41970
rect 22594 41918 22596 41970
rect 22428 41858 22484 41870
rect 22428 41806 22430 41858
rect 22482 41806 22484 41858
rect 22428 41300 22484 41806
rect 22540 41524 22596 41918
rect 22540 41458 22596 41468
rect 22428 41244 22596 41300
rect 22540 41186 22596 41244
rect 22540 41134 22542 41186
rect 22594 41134 22596 41186
rect 22540 41122 22596 41134
rect 22764 41186 22820 41198
rect 22764 41134 22766 41186
rect 22818 41134 22820 41186
rect 22092 40964 22148 40974
rect 22092 40870 22148 40908
rect 21868 40574 21870 40626
rect 21922 40574 21924 40626
rect 21868 40562 21924 40574
rect 21308 40402 21476 40404
rect 21308 40350 21310 40402
rect 21362 40350 21476 40402
rect 21308 40348 21476 40350
rect 21308 40338 21364 40348
rect 19516 40124 20020 40180
rect 20524 40180 20580 40190
rect 19516 39842 19572 40124
rect 19516 39790 19518 39842
rect 19570 39790 19572 39842
rect 19516 39778 19572 39790
rect 20412 39956 20468 39966
rect 18956 39620 19012 39630
rect 18620 39618 19012 39620
rect 18620 39566 18958 39618
rect 19010 39566 19012 39618
rect 18620 39564 19012 39566
rect 18508 39554 18564 39564
rect 18172 39454 18174 39506
rect 18226 39454 18228 39506
rect 18172 39442 18228 39454
rect 18956 39396 19012 39564
rect 18956 39330 19012 39340
rect 19180 39620 19236 39630
rect 17724 38854 17780 38892
rect 18060 39060 18116 39070
rect 18060 38946 18116 39004
rect 18060 38894 18062 38946
rect 18114 38894 18116 38946
rect 18060 38882 18116 38894
rect 18172 38948 18228 38958
rect 18172 38946 18340 38948
rect 18172 38894 18174 38946
rect 18226 38894 18340 38946
rect 18172 38892 18340 38894
rect 18172 38882 18228 38892
rect 17052 38724 17108 38734
rect 16268 37314 16324 37324
rect 16940 38388 16996 38398
rect 14700 36594 14756 36652
rect 14700 36542 14702 36594
rect 14754 36542 14756 36594
rect 14700 36530 14756 36542
rect 15148 36596 15204 36606
rect 15148 36482 15204 36540
rect 15596 36484 15652 36494
rect 15148 36430 15150 36482
rect 15202 36430 15204 36482
rect 15148 36418 15204 36430
rect 15484 36482 15652 36484
rect 15484 36430 15598 36482
rect 15650 36430 15652 36482
rect 15484 36428 15652 36430
rect 15260 36372 15316 36382
rect 14476 35812 14532 35822
rect 14252 35534 14254 35586
rect 14306 35534 14308 35586
rect 14252 35522 14308 35534
rect 14364 35698 14420 35710
rect 14364 35646 14366 35698
rect 14418 35646 14420 35698
rect 14364 35364 14420 35646
rect 13468 35308 14420 35364
rect 13580 35028 13636 35038
rect 13580 34130 13636 34972
rect 14140 34916 14196 34926
rect 13916 34804 13972 34814
rect 13916 34244 13972 34748
rect 13916 34178 13972 34188
rect 13580 34078 13582 34130
rect 13634 34078 13636 34130
rect 13468 32564 13524 32574
rect 13468 32470 13524 32508
rect 13580 32450 13636 34078
rect 14140 34130 14196 34860
rect 14252 34244 14308 34254
rect 14364 34244 14420 35308
rect 14476 34356 14532 35756
rect 15036 35698 15092 35710
rect 15036 35646 15038 35698
rect 15090 35646 15092 35698
rect 15036 35028 15092 35646
rect 15036 34962 15092 34972
rect 15148 34916 15204 34926
rect 15148 34822 15204 34860
rect 14476 34290 14532 34300
rect 15260 34354 15316 36316
rect 15484 35812 15540 36428
rect 15596 36418 15652 36428
rect 15372 35700 15428 35710
rect 15372 35606 15428 35644
rect 15260 34302 15262 34354
rect 15314 34302 15316 34354
rect 15260 34290 15316 34302
rect 14252 34242 14420 34244
rect 14252 34190 14254 34242
rect 14306 34190 14420 34242
rect 14252 34188 14420 34190
rect 14252 34178 14308 34188
rect 14140 34078 14142 34130
rect 14194 34078 14196 34130
rect 14140 34066 14196 34078
rect 14924 34130 14980 34142
rect 14924 34078 14926 34130
rect 14978 34078 14980 34130
rect 14476 33460 14532 33470
rect 13580 32398 13582 32450
rect 13634 32398 13636 32450
rect 13580 32386 13636 32398
rect 14364 33346 14420 33358
rect 14364 33294 14366 33346
rect 14418 33294 14420 33346
rect 13916 32004 13972 32014
rect 13692 31892 13748 31902
rect 13692 31798 13748 31836
rect 13244 30790 13300 30828
rect 13916 31778 13972 31948
rect 13916 31726 13918 31778
rect 13970 31726 13972 31778
rect 12460 30324 12516 30334
rect 12460 30230 12516 30268
rect 13916 30324 13972 31726
rect 14252 31780 14308 31790
rect 14252 31686 14308 31724
rect 14364 31556 14420 33294
rect 14476 32562 14532 33404
rect 14924 32676 14980 34078
rect 15260 33348 15316 33358
rect 15484 33348 15540 35756
rect 15708 35586 15764 37100
rect 15820 36596 15876 36606
rect 15820 36370 15876 36540
rect 15820 36318 15822 36370
rect 15874 36318 15876 36370
rect 15820 36306 15876 36318
rect 16156 36372 16212 36382
rect 16156 36278 16212 36316
rect 16380 36258 16436 36270
rect 16380 36206 16382 36258
rect 16434 36206 16436 36258
rect 16380 35698 16436 36206
rect 16380 35646 16382 35698
rect 16434 35646 16436 35698
rect 15708 35534 15710 35586
rect 15762 35534 15764 35586
rect 15708 35522 15764 35534
rect 16044 35586 16100 35598
rect 16044 35534 16046 35586
rect 16098 35534 16100 35586
rect 15708 34916 15764 34926
rect 16044 34916 16100 35534
rect 16156 35028 16212 35038
rect 16156 34934 16212 34972
rect 15708 34914 16044 34916
rect 15708 34862 15710 34914
rect 15762 34862 16044 34914
rect 15708 34860 16044 34862
rect 15708 34850 15764 34860
rect 16044 34822 16100 34860
rect 16380 34914 16436 35646
rect 16380 34862 16382 34914
rect 16434 34862 16436 34914
rect 16380 34804 16436 34862
rect 16380 34738 16436 34748
rect 15596 34356 15652 34366
rect 15596 34262 15652 34300
rect 16940 34356 16996 38332
rect 17052 38050 17108 38668
rect 18172 38612 18228 38622
rect 18060 38610 18228 38612
rect 18060 38558 18174 38610
rect 18226 38558 18228 38610
rect 18060 38556 18228 38558
rect 17388 38164 17444 38174
rect 17388 38070 17444 38108
rect 17052 37998 17054 38050
rect 17106 37998 17108 38050
rect 17052 37986 17108 37998
rect 17948 37828 18004 37838
rect 17388 37716 17444 37726
rect 17164 36708 17220 36718
rect 17164 36594 17220 36652
rect 17164 36542 17166 36594
rect 17218 36542 17220 36594
rect 17164 35700 17220 36542
rect 17388 36036 17444 37660
rect 17500 37156 17556 37166
rect 17500 37062 17556 37100
rect 17948 36482 18004 37772
rect 18060 37378 18116 38556
rect 18172 38546 18228 38556
rect 18284 38052 18340 38892
rect 19180 38722 19236 39564
rect 19404 39508 19460 39518
rect 19852 39508 19908 39518
rect 19404 38834 19460 39452
rect 19628 39506 19908 39508
rect 19628 39454 19854 39506
rect 19906 39454 19908 39506
rect 19628 39452 19908 39454
rect 19404 38782 19406 38834
rect 19458 38782 19460 38834
rect 19404 38770 19460 38782
rect 19516 38948 19572 38958
rect 19180 38670 19182 38722
rect 19234 38670 19236 38722
rect 19180 38658 19236 38670
rect 18284 37986 18340 37996
rect 18732 38050 18788 38062
rect 18732 37998 18734 38050
rect 18786 37998 18788 38050
rect 18060 37326 18062 37378
rect 18114 37326 18116 37378
rect 18060 36708 18116 37326
rect 18060 36642 18116 36652
rect 18172 37604 18228 37614
rect 17948 36430 17950 36482
rect 18002 36430 18004 36482
rect 17948 36418 18004 36430
rect 18172 36482 18228 37548
rect 18620 37604 18676 37614
rect 18508 36708 18564 36718
rect 18508 36614 18564 36652
rect 18620 36706 18676 37548
rect 18732 37156 18788 37998
rect 19068 37938 19124 37950
rect 19068 37886 19070 37938
rect 19122 37886 19124 37938
rect 18956 37828 19012 37838
rect 18956 37734 19012 37772
rect 19068 37268 19124 37886
rect 19516 37380 19572 38892
rect 19628 37604 19684 39452
rect 19852 39442 19908 39452
rect 20188 39508 20244 39518
rect 20188 39414 20244 39452
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 19964 38836 20020 38846
rect 20412 38836 20468 39900
rect 19964 38742 20020 38780
rect 20188 38834 20468 38836
rect 20188 38782 20414 38834
rect 20466 38782 20468 38834
rect 20188 38780 20468 38782
rect 20188 38668 20244 38780
rect 20412 38770 20468 38780
rect 20076 38612 20244 38668
rect 20524 38668 20580 40124
rect 20636 40068 20692 40078
rect 20636 38948 20692 40012
rect 21308 39396 21364 39406
rect 21308 39302 21364 39340
rect 21420 39284 21476 40348
rect 22652 40516 22708 40526
rect 22764 40516 22820 41134
rect 22652 40514 22820 40516
rect 22652 40462 22654 40514
rect 22706 40462 22820 40514
rect 22652 40460 22820 40462
rect 21532 40178 21588 40190
rect 21532 40126 21534 40178
rect 21586 40126 21588 40178
rect 21532 39620 21588 40126
rect 21532 39554 21588 39564
rect 21644 39508 21700 39518
rect 21644 39414 21700 39452
rect 21420 39228 21700 39284
rect 20636 38834 20692 38892
rect 20636 38782 20638 38834
rect 20690 38782 20692 38834
rect 20636 38770 20692 38782
rect 21420 38948 21476 38958
rect 20972 38724 21028 38734
rect 21308 38724 21364 38762
rect 20972 38722 21308 38724
rect 20972 38670 20974 38722
rect 21026 38670 21308 38722
rect 20972 38668 21308 38670
rect 20524 38612 20916 38668
rect 20972 38658 21028 38668
rect 21308 38658 21364 38668
rect 19740 38052 19796 38062
rect 19740 37958 19796 37996
rect 20076 37938 20132 38612
rect 20076 37886 20078 37938
rect 20130 37886 20132 37938
rect 20076 37874 20132 37886
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 19628 37538 19684 37548
rect 19964 37380 20020 37390
rect 19516 37378 20020 37380
rect 19516 37326 19966 37378
rect 20018 37326 20020 37378
rect 19516 37324 20020 37326
rect 19964 37314 20020 37324
rect 20076 37380 20132 37390
rect 20188 37380 20244 37390
rect 20076 37378 20188 37380
rect 20076 37326 20078 37378
rect 20130 37326 20188 37378
rect 20076 37324 20188 37326
rect 20076 37314 20132 37324
rect 19068 37174 19124 37212
rect 18732 37090 18788 37100
rect 19628 37154 19684 37166
rect 19628 37102 19630 37154
rect 19682 37102 19684 37154
rect 18956 37044 19012 37054
rect 18956 36708 19012 36988
rect 18620 36654 18622 36706
rect 18674 36654 18676 36706
rect 18620 36642 18676 36654
rect 18844 36706 19012 36708
rect 18844 36654 18958 36706
rect 19010 36654 19012 36706
rect 18844 36652 19012 36654
rect 19628 36708 19684 37102
rect 20076 37044 20132 37054
rect 20076 36950 20132 36988
rect 19628 36652 20020 36708
rect 18732 36596 18788 36606
rect 18732 36502 18788 36540
rect 18172 36430 18174 36482
rect 18226 36430 18228 36482
rect 18172 36418 18228 36430
rect 17612 36260 17668 36270
rect 17388 35980 17556 36036
rect 17388 35812 17444 35822
rect 17388 35718 17444 35756
rect 17164 35634 17220 35644
rect 17500 35140 17556 35980
rect 17612 35810 17668 36204
rect 17612 35758 17614 35810
rect 17666 35758 17668 35810
rect 17612 35746 17668 35758
rect 18844 35812 18900 36652
rect 18956 36642 19012 36652
rect 19964 36596 20020 36652
rect 19964 36502 20020 36540
rect 19180 36484 19236 36494
rect 19852 36484 19908 36494
rect 17948 35700 18004 35710
rect 17948 35606 18004 35644
rect 17836 35588 17892 35598
rect 17836 35494 17892 35532
rect 17724 35140 17780 35150
rect 17500 35084 17668 35140
rect 17164 35026 17220 35038
rect 17164 34974 17166 35026
rect 17218 34974 17220 35026
rect 17164 34916 17220 34974
rect 17164 34850 17220 34860
rect 17500 34916 17556 34926
rect 17500 34822 17556 34860
rect 16940 34290 16996 34300
rect 17276 34468 17332 34478
rect 15708 34244 15764 34254
rect 15708 34150 15764 34188
rect 15260 33346 15540 33348
rect 15260 33294 15262 33346
rect 15314 33294 15540 33346
rect 15260 33292 15540 33294
rect 15260 33282 15316 33292
rect 14924 32610 14980 32620
rect 14476 32510 14478 32562
rect 14530 32510 14532 32562
rect 14476 32498 14532 32510
rect 15260 32562 15316 32574
rect 15260 32510 15262 32562
rect 15314 32510 15316 32562
rect 15148 32450 15204 32462
rect 15148 32398 15150 32450
rect 15202 32398 15204 32450
rect 15148 31948 15204 32398
rect 14588 31892 14644 31902
rect 14812 31892 15204 31948
rect 15260 32004 15316 32510
rect 14644 31836 14868 31892
rect 14588 31778 14644 31836
rect 14588 31726 14590 31778
rect 14642 31726 14644 31778
rect 14588 31714 14644 31726
rect 14924 31780 14980 31790
rect 15260 31780 15316 31948
rect 16380 31892 16436 31902
rect 16828 31892 16884 31902
rect 16380 31798 16436 31836
rect 16716 31890 16884 31892
rect 16716 31838 16830 31890
rect 16882 31838 16884 31890
rect 16716 31836 16884 31838
rect 14924 31778 15316 31780
rect 14924 31726 14926 31778
rect 14978 31726 15316 31778
rect 14924 31724 15316 31726
rect 16156 31780 16212 31790
rect 14924 31714 14980 31724
rect 16156 31686 16212 31724
rect 16604 31780 16660 31790
rect 16604 31686 16660 31724
rect 14812 31668 14868 31678
rect 14812 31556 14868 31612
rect 14364 31554 14868 31556
rect 14364 31502 14814 31554
rect 14866 31502 14868 31554
rect 14364 31500 14868 31502
rect 14812 31490 14868 31500
rect 16156 30996 16212 31006
rect 16604 30996 16660 31006
rect 16156 30994 16604 30996
rect 16156 30942 16158 30994
rect 16210 30942 16604 30994
rect 16156 30940 16604 30942
rect 16156 30930 16212 30940
rect 16604 30902 16660 30940
rect 15260 30884 15316 30894
rect 15260 30436 15316 30828
rect 13916 30258 13972 30268
rect 14700 30324 14756 30334
rect 11452 30118 11508 30156
rect 14476 30212 14532 30222
rect 14476 30118 14532 30156
rect 10668 30034 10724 30044
rect 14700 30098 14756 30268
rect 14700 30046 14702 30098
rect 14754 30046 14756 30098
rect 14700 30034 14756 30046
rect 15260 30100 15316 30380
rect 15372 30882 15428 30894
rect 15372 30830 15374 30882
rect 15426 30830 15428 30882
rect 15372 30324 15428 30830
rect 16604 30772 16660 30782
rect 16044 30436 16100 30446
rect 16044 30342 16100 30380
rect 15372 30258 15428 30268
rect 15708 30212 15764 30222
rect 15708 30118 15764 30156
rect 15372 30100 15428 30110
rect 15260 30098 15428 30100
rect 15260 30046 15374 30098
rect 15426 30046 15428 30098
rect 15260 30044 15428 30046
rect 15372 30034 15428 30044
rect 16604 30098 16660 30716
rect 16604 30046 16606 30098
rect 16658 30046 16660 30098
rect 16604 30034 16660 30046
rect 9660 29698 9716 29708
rect 13468 29988 13524 29998
rect 8988 29650 9156 29652
rect 8988 29598 8990 29650
rect 9042 29598 9156 29650
rect 8988 29596 9156 29598
rect 8988 29586 9044 29596
rect 8316 29486 8318 29538
rect 8370 29486 8372 29538
rect 8316 29474 8372 29486
rect 7868 29428 7924 29438
rect 7644 29426 7924 29428
rect 7644 29374 7870 29426
rect 7922 29374 7924 29426
rect 7644 29372 7924 29374
rect 7532 29362 7588 29372
rect 6636 29204 6692 29214
rect 6636 29110 6692 29148
rect 7868 29204 7924 29372
rect 8428 29428 8484 29438
rect 8428 29334 8484 29372
rect 8540 29426 8596 29438
rect 8540 29374 8542 29426
rect 8594 29374 8596 29426
rect 7868 29138 7924 29148
rect 8540 29204 8596 29374
rect 13468 29316 13524 29932
rect 14588 29538 14644 29550
rect 14588 29486 14590 29538
rect 14642 29486 14644 29538
rect 14364 29428 14420 29438
rect 14364 29334 14420 29372
rect 8540 29138 8596 29148
rect 9996 29204 10052 29214
rect 5964 28814 5966 28866
rect 6018 28814 6020 28866
rect 5964 28802 6020 28814
rect 5852 28478 5854 28530
rect 5906 28478 5908 28530
rect 5852 28466 5908 28478
rect 6636 28644 6692 28654
rect 3612 28030 3614 28082
rect 3666 28030 3668 28082
rect 3612 27860 3668 28030
rect 3612 27794 3668 27804
rect 6636 27860 6692 28588
rect 6636 27794 6692 27804
rect 3164 27746 3220 27758
rect 3164 27694 3166 27746
rect 3218 27694 3220 27746
rect 3164 27636 3220 27694
rect 3164 27570 3220 27580
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 2716 26962 2996 26964
rect 2716 26910 2718 26962
rect 2770 26910 2996 26962
rect 2716 26908 2996 26910
rect 3164 27074 3220 27086
rect 3164 27022 3166 27074
rect 3218 27022 3220 27074
rect 2716 26898 2772 26908
rect 2044 26516 2100 26526
rect 2044 26422 2100 26460
rect 1820 26404 1876 26414
rect 1820 26290 1876 26348
rect 1820 26238 1822 26290
rect 1874 26238 1876 26290
rect 1820 26226 1876 26238
rect 2380 26290 2436 26302
rect 2380 26238 2382 26290
rect 2434 26238 2436 26290
rect 2380 26068 2436 26238
rect 2492 26292 2548 26796
rect 3164 26852 3220 27022
rect 3612 27076 3668 27086
rect 3612 26982 3668 27020
rect 5068 27076 5124 27086
rect 5068 26908 5124 27020
rect 6860 27074 6916 27086
rect 6860 27022 6862 27074
rect 6914 27022 6916 27074
rect 6524 26962 6580 26974
rect 6524 26910 6526 26962
rect 6578 26910 6580 26962
rect 6524 26908 6580 26910
rect 3164 26786 3220 26796
rect 4956 26852 5124 26908
rect 6300 26852 6580 26908
rect 3388 26740 3444 26750
rect 2716 26628 2772 26638
rect 2716 26514 2772 26572
rect 2716 26462 2718 26514
rect 2770 26462 2772 26514
rect 2716 26450 2772 26462
rect 3388 26514 3444 26684
rect 3388 26462 3390 26514
rect 3442 26462 3444 26514
rect 3388 26450 3444 26462
rect 4732 26404 4788 26414
rect 4732 26310 4788 26348
rect 2492 26226 2548 26236
rect 3052 26290 3108 26302
rect 3052 26238 3054 26290
rect 3106 26238 3108 26290
rect 3052 26180 3108 26238
rect 3052 26114 3108 26124
rect 3836 26180 3892 26190
rect 3836 26086 3892 26124
rect 4284 26180 4340 26190
rect 4284 26086 4340 26124
rect 1932 25618 1988 25630
rect 1932 25566 1934 25618
rect 1986 25566 1988 25618
rect 1932 24948 1988 25566
rect 1932 24882 1988 24892
rect 2044 24722 2100 24734
rect 2044 24670 2046 24722
rect 2098 24670 2100 24722
rect 2044 23940 2100 24670
rect 2380 24276 2436 26012
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 4844 25732 4900 25742
rect 4284 25508 4340 25518
rect 4284 24946 4340 25452
rect 4844 25506 4900 25676
rect 4844 25454 4846 25506
rect 4898 25454 4900 25506
rect 4284 24894 4286 24946
rect 4338 24894 4340 24946
rect 4284 24882 4340 24894
rect 4620 25396 4676 25406
rect 3276 24834 3332 24846
rect 4620 24836 4676 25340
rect 3276 24782 3278 24834
rect 3330 24782 3332 24834
rect 3052 24724 3108 24734
rect 3052 24722 3220 24724
rect 3052 24670 3054 24722
rect 3106 24670 3220 24722
rect 3052 24668 3220 24670
rect 3052 24658 3108 24668
rect 2380 24210 2436 24220
rect 2492 24610 2548 24622
rect 2828 24612 2884 24622
rect 2492 24558 2494 24610
rect 2546 24558 2548 24610
rect 2380 24052 2436 24062
rect 2044 23938 2212 23940
rect 2044 23886 2046 23938
rect 2098 23886 2212 23938
rect 2044 23884 2212 23886
rect 2044 23874 2100 23884
rect 2156 23828 2212 23884
rect 1932 23604 1988 23614
rect 1988 23548 2100 23604
rect 1932 23538 1988 23548
rect 1820 23044 1876 23054
rect 1820 23042 1988 23044
rect 1820 22990 1822 23042
rect 1874 22990 1988 23042
rect 1820 22988 1988 22990
rect 1820 22978 1876 22988
rect 1708 22932 1764 22942
rect 1708 21812 1764 22876
rect 1820 21812 1876 21822
rect 1708 21810 1876 21812
rect 1708 21758 1822 21810
rect 1874 21758 1876 21810
rect 1708 21756 1876 21758
rect 1708 21362 1764 21374
rect 1708 21310 1710 21362
rect 1762 21310 1764 21362
rect 1708 20804 1764 21310
rect 1708 20710 1764 20748
rect 1708 20244 1764 20254
rect 1708 17666 1764 20188
rect 1820 19234 1876 21756
rect 1820 19182 1822 19234
rect 1874 19182 1876 19234
rect 1820 19170 1876 19182
rect 1932 21588 1988 22988
rect 2044 21698 2100 23548
rect 2044 21646 2046 21698
rect 2098 21646 2100 21698
rect 2044 21634 2100 21646
rect 1820 18452 1876 18462
rect 1932 18452 1988 21532
rect 2044 21364 2100 21374
rect 2044 20690 2100 21308
rect 2044 20638 2046 20690
rect 2098 20638 2100 20690
rect 2044 20626 2100 20638
rect 2156 20468 2212 23772
rect 2268 23156 2324 23166
rect 2268 22820 2324 23100
rect 2268 22754 2324 22764
rect 2044 20412 2212 20468
rect 2268 21588 2324 21598
rect 2380 21588 2436 23996
rect 2492 22596 2548 24558
rect 2604 24610 2884 24612
rect 2604 24558 2830 24610
rect 2882 24558 2884 24610
rect 2604 24556 2884 24558
rect 2604 24052 2660 24556
rect 2828 24546 2884 24556
rect 2604 23986 2660 23996
rect 2716 23940 2772 23950
rect 2492 22540 2660 22596
rect 2268 21586 2436 21588
rect 2268 21534 2270 21586
rect 2322 21534 2436 21586
rect 2268 21532 2436 21534
rect 2492 22370 2548 22382
rect 2492 22318 2494 22370
rect 2546 22318 2548 22370
rect 2492 21586 2548 22318
rect 2604 22036 2660 22540
rect 2716 22484 2772 23884
rect 2828 23938 2884 23950
rect 2828 23886 2830 23938
rect 2882 23886 2884 23938
rect 2828 23716 2884 23886
rect 2940 23828 2996 23838
rect 2940 23734 2996 23772
rect 3164 23826 3220 24668
rect 3164 23774 3166 23826
rect 3218 23774 3220 23826
rect 2828 23268 2884 23660
rect 2828 23212 2996 23268
rect 2828 23044 2884 23054
rect 2828 22950 2884 22988
rect 2716 22428 2884 22484
rect 2716 22260 2772 22270
rect 2716 22166 2772 22204
rect 2604 21970 2660 21980
rect 2492 21534 2494 21586
rect 2546 21534 2548 21586
rect 2044 19122 2100 20412
rect 2268 20132 2324 21532
rect 2492 21140 2548 21534
rect 2716 21588 2772 21598
rect 2716 21494 2772 21532
rect 2828 21588 2884 22428
rect 2940 21812 2996 23212
rect 3164 23156 3220 23774
rect 3164 23090 3220 23100
rect 3276 21924 3332 24782
rect 4396 24780 4788 24836
rect 3388 24722 3444 24734
rect 3388 24670 3390 24722
rect 3442 24670 3444 24722
rect 3388 23940 3444 24670
rect 3836 24724 3892 24734
rect 4396 24724 4452 24780
rect 3836 24722 4452 24724
rect 3836 24670 3838 24722
rect 3890 24670 4452 24722
rect 3836 24668 4452 24670
rect 4732 24722 4788 24780
rect 4732 24670 4734 24722
rect 4786 24670 4788 24722
rect 3836 24658 3892 24668
rect 4732 24658 4788 24670
rect 4508 24610 4564 24622
rect 4508 24558 4510 24610
rect 4562 24558 4564 24610
rect 4508 24500 4564 24558
rect 4844 24500 4900 25454
rect 4956 25508 5012 26852
rect 5404 26402 5460 26414
rect 5404 26350 5406 26402
rect 5458 26350 5460 26402
rect 4956 25442 5012 25452
rect 5180 26290 5236 26302
rect 5180 26238 5182 26290
rect 5234 26238 5236 26290
rect 5180 25396 5236 26238
rect 5404 25508 5460 26350
rect 6300 26402 6356 26852
rect 6300 26350 6302 26402
rect 6354 26350 6356 26402
rect 5404 25442 5460 25452
rect 5740 25844 5796 25854
rect 5180 25330 5236 25340
rect 5628 25396 5684 25406
rect 5628 25302 5684 25340
rect 5068 25282 5124 25294
rect 5068 25230 5070 25282
rect 5122 25230 5124 25282
rect 3836 24444 4900 24500
rect 4956 24498 5012 24510
rect 4956 24446 4958 24498
rect 5010 24446 5012 24498
rect 3836 24162 3892 24444
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 3836 24110 3838 24162
rect 3890 24110 3892 24162
rect 3836 24098 3892 24110
rect 3388 23846 3444 23884
rect 4620 23938 4676 23950
rect 4620 23886 4622 23938
rect 4674 23886 4676 23938
rect 4620 23828 4676 23886
rect 4676 23772 4788 23828
rect 4620 23762 4676 23772
rect 4060 23716 4116 23726
rect 4060 23622 4116 23660
rect 3724 23266 3780 23278
rect 3724 23214 3726 23266
rect 3778 23214 3780 23266
rect 3612 23156 3668 23166
rect 3612 22258 3668 23100
rect 3612 22206 3614 22258
rect 3666 22206 3668 22258
rect 3276 21858 3332 21868
rect 3500 22148 3556 22158
rect 2940 21756 3220 21812
rect 2828 21586 3108 21588
rect 2828 21534 2830 21586
rect 2882 21534 3108 21586
rect 2828 21532 3108 21534
rect 2828 21522 2884 21532
rect 2492 21084 2772 21140
rect 2492 20914 2548 20926
rect 2492 20862 2494 20914
rect 2546 20862 2548 20914
rect 2380 20804 2436 20814
rect 2492 20804 2548 20862
rect 2436 20748 2548 20804
rect 2380 20738 2436 20748
rect 2492 20132 2548 20142
rect 2268 20076 2492 20132
rect 2492 20066 2548 20076
rect 2044 19070 2046 19122
rect 2098 19070 2100 19122
rect 2044 19058 2100 19070
rect 2156 20018 2212 20030
rect 2156 19966 2158 20018
rect 2210 19966 2212 20018
rect 1820 18450 1988 18452
rect 1820 18398 1822 18450
rect 1874 18398 1988 18450
rect 1820 18396 1988 18398
rect 2044 18562 2100 18574
rect 2044 18510 2046 18562
rect 2098 18510 2100 18562
rect 1820 18386 1876 18396
rect 1820 18228 1876 18238
rect 2044 18228 2100 18510
rect 1876 18172 2100 18228
rect 1820 18162 1876 18172
rect 1708 17614 1710 17666
rect 1762 17614 1764 17666
rect 1708 17108 1764 17614
rect 1820 17556 1876 17566
rect 2044 17556 2100 17566
rect 1876 17500 1988 17556
rect 1820 17490 1876 17500
rect 1708 17042 1764 17052
rect 1820 17332 1876 17342
rect 1820 16882 1876 17276
rect 1820 16830 1822 16882
rect 1874 16830 1876 16882
rect 1820 16818 1876 16830
rect 1932 16996 1988 17500
rect 2044 17462 2100 17500
rect 2156 17444 2212 19966
rect 2604 20020 2660 20030
rect 2604 19926 2660 19964
rect 2716 19908 2772 21084
rect 2828 20580 2884 20590
rect 2828 20486 2884 20524
rect 2716 19842 2772 19852
rect 2716 19460 2772 19470
rect 2380 19124 2436 19134
rect 2380 19030 2436 19068
rect 2716 19122 2772 19404
rect 3052 19124 3108 21532
rect 2716 19070 2718 19122
rect 2770 19070 2772 19122
rect 2716 19058 2772 19070
rect 2828 19068 3108 19124
rect 2716 18562 2772 18574
rect 2716 18510 2718 18562
rect 2770 18510 2772 18562
rect 2492 18450 2548 18462
rect 2492 18398 2494 18450
rect 2546 18398 2548 18450
rect 2492 18340 2548 18398
rect 2716 18452 2772 18510
rect 2716 18386 2772 18396
rect 2380 17554 2436 17566
rect 2380 17502 2382 17554
rect 2434 17502 2436 17554
rect 2380 17444 2436 17502
rect 2156 17388 2436 17444
rect 2044 17108 2100 17118
rect 2156 17108 2212 17388
rect 2044 17106 2212 17108
rect 2044 17054 2046 17106
rect 2098 17054 2212 17106
rect 2044 17052 2212 17054
rect 2380 17220 2436 17230
rect 2380 17106 2436 17164
rect 2380 17054 2382 17106
rect 2434 17054 2436 17106
rect 2044 17042 2100 17052
rect 2380 17042 2436 17054
rect 1708 15988 1764 15998
rect 1932 15988 1988 16940
rect 1708 15986 1988 15988
rect 1708 15934 1710 15986
rect 1762 15934 1988 15986
rect 1708 15932 1988 15934
rect 2044 16660 2100 16670
rect 2044 15986 2100 16604
rect 2492 16210 2548 18284
rect 2828 18228 2884 19068
rect 2716 18172 2884 18228
rect 2940 18900 2996 18910
rect 2492 16158 2494 16210
rect 2546 16158 2548 16210
rect 2492 16146 2548 16158
rect 2604 18116 2660 18126
rect 2604 16882 2660 18060
rect 2716 17554 2772 18172
rect 2940 17780 2996 18844
rect 3052 18562 3108 19068
rect 3052 18510 3054 18562
rect 3106 18510 3108 18562
rect 3052 18498 3108 18510
rect 2940 17668 2996 17724
rect 3052 17668 3108 17678
rect 2940 17666 3108 17668
rect 2940 17614 3054 17666
rect 3106 17614 3108 17666
rect 2940 17612 3108 17614
rect 3052 17602 3108 17612
rect 2716 17502 2718 17554
rect 2770 17502 2772 17554
rect 2716 17490 2772 17502
rect 3052 17108 3108 17118
rect 3164 17108 3220 21756
rect 3276 21474 3332 21486
rect 3276 21422 3278 21474
rect 3330 21422 3332 21474
rect 3276 21252 3332 21422
rect 3276 21186 3332 21196
rect 3276 20914 3332 20926
rect 3276 20862 3278 20914
rect 3330 20862 3332 20914
rect 3276 20130 3332 20862
rect 3276 20078 3278 20130
rect 3330 20078 3332 20130
rect 3276 19908 3332 20078
rect 3276 18676 3332 19852
rect 3276 18610 3332 18620
rect 3388 20580 3444 20590
rect 3388 18674 3444 20524
rect 3500 19124 3556 22092
rect 3612 22036 3668 22206
rect 3612 21970 3668 21980
rect 3724 22260 3780 23214
rect 4732 23266 4788 23772
rect 4732 23214 4734 23266
rect 4786 23214 4788 23266
rect 4732 23202 4788 23214
rect 3612 21588 3668 21598
rect 3612 20692 3668 21532
rect 3612 19796 3668 20636
rect 3724 20802 3780 22204
rect 3724 20750 3726 20802
rect 3778 20750 3780 20802
rect 3724 20020 3780 20750
rect 4172 23154 4228 23166
rect 4172 23102 4174 23154
rect 4226 23102 4228 23154
rect 4172 23044 4228 23102
rect 4844 23156 4900 23166
rect 4844 23062 4900 23100
rect 4172 21812 4228 22988
rect 4172 20804 4228 21756
rect 4284 23042 4340 23054
rect 4284 22990 4286 23042
rect 4338 22990 4340 23042
rect 4284 21698 4340 22990
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4284 21646 4286 21698
rect 4338 21646 4340 21698
rect 4284 21634 4340 21646
rect 4508 22482 4564 22494
rect 4508 22430 4510 22482
rect 4562 22430 4564 22482
rect 4508 21586 4564 22430
rect 4508 21534 4510 21586
rect 4562 21534 4564 21586
rect 4508 21522 4564 21534
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 4844 20916 4900 20926
rect 4956 20916 5012 24446
rect 5068 23716 5124 25230
rect 5404 25284 5460 25294
rect 5404 24946 5460 25228
rect 5404 24894 5406 24946
rect 5458 24894 5460 24946
rect 5404 24882 5460 24894
rect 5740 24836 5796 25788
rect 5852 25732 5908 25742
rect 5852 25508 5908 25676
rect 5964 25732 6020 25742
rect 6300 25732 6356 26350
rect 6860 26292 6916 27022
rect 7756 27074 7812 27086
rect 7756 27022 7758 27074
rect 7810 27022 7812 27074
rect 6860 26290 7028 26292
rect 6860 26238 6862 26290
rect 6914 26238 7028 26290
rect 6860 26236 7028 26238
rect 6860 26226 6916 26236
rect 5964 25730 6356 25732
rect 5964 25678 5966 25730
rect 6018 25678 6356 25730
rect 5964 25676 6356 25678
rect 6636 25844 6692 25854
rect 5964 25666 6020 25676
rect 5964 25508 6020 25518
rect 5852 25506 6020 25508
rect 5852 25454 5966 25506
rect 6018 25454 6020 25506
rect 5852 25452 6020 25454
rect 5964 25396 6020 25452
rect 5964 25330 6020 25340
rect 6300 25508 6356 25518
rect 5740 24780 5908 24836
rect 5740 24610 5796 24622
rect 5740 24558 5742 24610
rect 5794 24558 5796 24610
rect 5740 24500 5796 24558
rect 5740 24434 5796 24444
rect 5852 23940 5908 24780
rect 6300 24722 6356 25452
rect 6636 25506 6692 25788
rect 6636 25454 6638 25506
rect 6690 25454 6692 25506
rect 6636 25442 6692 25454
rect 6748 25618 6804 25630
rect 6748 25566 6750 25618
rect 6802 25566 6804 25618
rect 6300 24670 6302 24722
rect 6354 24670 6356 24722
rect 6300 24658 6356 24670
rect 5628 23938 5908 23940
rect 5628 23886 5854 23938
rect 5906 23886 5908 23938
rect 5628 23884 5908 23886
rect 5180 23716 5236 23726
rect 5068 23660 5180 23716
rect 5180 23622 5236 23660
rect 5068 22370 5124 22382
rect 5068 22318 5070 22370
rect 5122 22318 5124 22370
rect 5068 21812 5124 22318
rect 5068 21746 5124 21756
rect 5628 21588 5684 23884
rect 5852 23874 5908 23884
rect 6076 24610 6132 24622
rect 6076 24558 6078 24610
rect 6130 24558 6132 24610
rect 6076 24500 6132 24558
rect 6524 24500 6580 24510
rect 6076 23716 6132 24444
rect 6412 24498 6580 24500
rect 6412 24446 6526 24498
rect 6578 24446 6580 24498
rect 6412 24444 6580 24446
rect 5852 23660 6076 23716
rect 5852 22482 5908 23660
rect 6076 23650 6132 23660
rect 6188 23940 6244 23950
rect 6412 23940 6468 24444
rect 6524 24434 6580 24444
rect 6748 24498 6804 25566
rect 6748 24446 6750 24498
rect 6802 24446 6804 24498
rect 6244 23884 6468 23940
rect 6524 23938 6580 23950
rect 6524 23886 6526 23938
rect 6578 23886 6580 23938
rect 6188 23714 6244 23884
rect 6188 23662 6190 23714
rect 6242 23662 6244 23714
rect 5852 22430 5854 22482
rect 5906 22430 5908 22482
rect 5852 22418 5908 22430
rect 6076 22708 6132 22718
rect 5628 21494 5684 21532
rect 5180 21474 5236 21486
rect 5180 21422 5182 21474
rect 5234 21422 5236 21474
rect 5180 21028 5236 21422
rect 5180 20962 5236 20972
rect 4844 20914 5012 20916
rect 4844 20862 4846 20914
rect 4898 20862 5012 20914
rect 4844 20860 5012 20862
rect 4844 20850 4900 20860
rect 4284 20804 4340 20814
rect 4172 20802 4340 20804
rect 4172 20750 4286 20802
rect 4338 20750 4340 20802
rect 4172 20748 4340 20750
rect 4284 20738 4340 20748
rect 3836 20692 3892 20702
rect 3836 20598 3892 20636
rect 4956 20692 5012 20702
rect 4060 20580 4116 20590
rect 3948 20578 4116 20580
rect 3948 20526 4062 20578
rect 4114 20526 4116 20578
rect 3948 20524 4116 20526
rect 3724 19926 3780 19964
rect 3836 20356 3892 20366
rect 3612 19740 3780 19796
rect 3500 19058 3556 19068
rect 3612 19236 3668 19246
rect 3388 18622 3390 18674
rect 3442 18622 3444 18674
rect 3388 17892 3444 18622
rect 3612 18340 3668 19180
rect 3724 18900 3780 19740
rect 3836 19012 3892 20300
rect 3948 19460 4004 20524
rect 4060 20514 4116 20524
rect 4508 20580 4564 20590
rect 4508 20486 4564 20524
rect 4732 20580 4788 20590
rect 4732 20486 4788 20524
rect 4844 20578 4900 20590
rect 4844 20526 4846 20578
rect 4898 20526 4900 20578
rect 4844 20468 4900 20526
rect 4844 20402 4900 20412
rect 4956 20130 5012 20636
rect 5964 20578 6020 20590
rect 5964 20526 5966 20578
rect 6018 20526 6020 20578
rect 5964 20356 6020 20526
rect 5964 20290 6020 20300
rect 5852 20244 5908 20254
rect 4956 20078 4958 20130
rect 5010 20078 5012 20130
rect 4956 20066 5012 20078
rect 5516 20132 5572 20142
rect 5068 20020 5124 20030
rect 5068 19926 5124 19964
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4620 19460 4676 19470
rect 3948 19458 4676 19460
rect 3948 19406 4622 19458
rect 4674 19406 4676 19458
rect 3948 19404 4676 19406
rect 3948 19234 4004 19404
rect 4620 19394 4676 19404
rect 4956 19346 5012 19358
rect 4956 19294 4958 19346
rect 5010 19294 5012 19346
rect 3948 19182 3950 19234
rect 4002 19182 4004 19234
rect 3948 19170 4004 19182
rect 4172 19236 4228 19246
rect 4396 19236 4452 19246
rect 4956 19236 5012 19294
rect 4228 19234 4452 19236
rect 4228 19182 4398 19234
rect 4450 19182 4452 19234
rect 4228 19180 4452 19182
rect 4172 19170 4228 19180
rect 4396 19170 4452 19180
rect 4732 19180 4956 19236
rect 4060 19122 4116 19134
rect 4060 19070 4062 19122
rect 4114 19070 4116 19122
rect 4060 19012 4116 19070
rect 3836 18956 4116 19012
rect 3724 18844 4004 18900
rect 3724 18676 3780 18686
rect 3724 18582 3780 18620
rect 3388 17826 3444 17836
rect 3500 18284 3668 18340
rect 3836 18340 3892 18350
rect 3388 17668 3444 17678
rect 3388 17554 3444 17612
rect 3388 17502 3390 17554
rect 3442 17502 3444 17554
rect 3388 17490 3444 17502
rect 3052 17106 3220 17108
rect 3052 17054 3054 17106
rect 3106 17054 3220 17106
rect 3052 17052 3220 17054
rect 3052 17042 3108 17052
rect 2604 16830 2606 16882
rect 2658 16830 2660 16882
rect 2604 15988 2660 16830
rect 2940 16996 2996 17006
rect 2940 16436 2996 16940
rect 3164 16884 3220 16894
rect 3276 16884 3332 16894
rect 3500 16884 3556 18284
rect 3220 16882 3444 16884
rect 3220 16830 3278 16882
rect 3330 16830 3444 16882
rect 3220 16828 3444 16830
rect 3164 16818 3220 16828
rect 3276 16790 3332 16828
rect 2940 16380 3332 16436
rect 3164 16212 3220 16222
rect 2044 15934 2046 15986
rect 2098 15934 2100 15986
rect 1708 15922 1764 15932
rect 2044 15922 2100 15934
rect 2492 15932 2660 15988
rect 2940 15988 2996 15998
rect 1708 15764 1764 15774
rect 1708 15204 1764 15708
rect 1708 13858 1764 15148
rect 2268 15764 2324 15774
rect 1932 15092 1988 15102
rect 1932 14998 1988 15036
rect 2044 14756 2100 14766
rect 1820 14530 1876 14542
rect 1820 14478 1822 14530
rect 1874 14478 1876 14530
rect 1820 13972 1876 14478
rect 1820 13906 1876 13916
rect 2044 13970 2100 14700
rect 2268 14642 2324 15708
rect 2492 15092 2548 15932
rect 2828 15876 2884 15886
rect 2492 15026 2548 15036
rect 2604 15428 2660 15438
rect 2268 14590 2270 14642
rect 2322 14590 2324 14642
rect 2268 14578 2324 14590
rect 2604 14644 2660 15372
rect 2828 15148 2884 15820
rect 2604 14530 2660 14588
rect 2604 14478 2606 14530
rect 2658 14478 2660 14530
rect 2604 14466 2660 14478
rect 2716 15092 2884 15148
rect 2044 13918 2046 13970
rect 2098 13918 2100 13970
rect 2044 13906 2100 13918
rect 2716 13970 2772 15092
rect 2716 13918 2718 13970
rect 2770 13918 2772 13970
rect 2716 13906 2772 13918
rect 2828 14532 2884 14542
rect 1708 13806 1710 13858
rect 1762 13806 1764 13858
rect 1708 13794 1764 13806
rect 2044 13748 2100 13758
rect 1708 12852 1764 12862
rect 1708 12758 1764 12796
rect 2044 12850 2100 13692
rect 2380 13746 2436 13758
rect 2380 13694 2382 13746
rect 2434 13694 2436 13746
rect 2380 13524 2436 13694
rect 2380 13458 2436 13468
rect 2044 12798 2046 12850
rect 2098 12798 2100 12850
rect 2044 12786 2100 12798
rect 2492 12962 2548 12974
rect 2492 12910 2494 12962
rect 2546 12910 2548 12962
rect 1596 12572 1988 12628
rect 1932 12404 1988 12572
rect 2044 12404 2100 12414
rect 1932 12402 2100 12404
rect 1932 12350 2046 12402
rect 2098 12350 2100 12402
rect 1932 12348 2100 12350
rect 2044 12338 2100 12348
rect 1708 12178 1764 12190
rect 1708 12126 1710 12178
rect 1762 12126 1764 12178
rect 1708 11508 1764 12126
rect 2492 12180 2548 12910
rect 2716 12852 2772 12862
rect 2828 12852 2884 14476
rect 2940 14418 2996 15932
rect 3164 15986 3220 16156
rect 3164 15934 3166 15986
rect 3218 15934 3220 15986
rect 3164 15922 3220 15934
rect 2940 14366 2942 14418
rect 2994 14366 2996 14418
rect 2940 14354 2996 14366
rect 3052 15204 3108 15214
rect 3052 13076 3108 15148
rect 3164 13972 3220 13982
rect 3276 13972 3332 16380
rect 3388 14642 3444 16828
rect 3500 16818 3556 16828
rect 3612 17556 3668 17566
rect 3500 16212 3556 16222
rect 3612 16212 3668 17500
rect 3836 17106 3892 18284
rect 3836 17054 3838 17106
rect 3890 17054 3892 17106
rect 3836 17042 3892 17054
rect 3948 17666 4004 18844
rect 4060 18676 4116 18686
rect 4060 18582 4116 18620
rect 4508 18450 4564 18462
rect 4508 18398 4510 18450
rect 4562 18398 4564 18450
rect 4508 18340 4564 18398
rect 4732 18450 4788 19180
rect 4956 19170 5012 19180
rect 5292 19236 5348 19246
rect 5180 18900 5236 18910
rect 4732 18398 4734 18450
rect 4786 18398 4788 18450
rect 4732 18386 4788 18398
rect 5068 18564 5124 18574
rect 5068 18450 5124 18508
rect 5068 18398 5070 18450
rect 5122 18398 5124 18450
rect 5068 18386 5124 18398
rect 4508 18274 4564 18284
rect 4844 18338 4900 18350
rect 4844 18286 4846 18338
rect 4898 18286 4900 18338
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 3948 17614 3950 17666
rect 4002 17614 4004 17666
rect 3948 17108 4004 17614
rect 4396 17892 4452 17902
rect 4172 17444 4228 17454
rect 4172 17350 4228 17388
rect 4396 17108 4452 17836
rect 4844 17780 4900 18286
rect 4844 17724 5012 17780
rect 4508 17556 4564 17566
rect 4844 17556 4900 17566
rect 4508 17462 4564 17500
rect 4732 17500 4844 17556
rect 4508 17108 4564 17118
rect 3948 17052 4116 17108
rect 3500 16210 3668 16212
rect 3500 16158 3502 16210
rect 3554 16158 3668 16210
rect 3500 16156 3668 16158
rect 3724 16882 3780 16894
rect 3724 16830 3726 16882
rect 3778 16830 3780 16882
rect 3500 16146 3556 16156
rect 3612 15988 3668 15998
rect 3724 15988 3780 16830
rect 3836 16884 3892 16894
rect 3836 16658 3892 16828
rect 3836 16606 3838 16658
rect 3890 16606 3892 16658
rect 3836 16594 3892 16606
rect 3612 15986 3780 15988
rect 3612 15934 3614 15986
rect 3666 15934 3780 15986
rect 3612 15932 3780 15934
rect 3948 15988 4004 15998
rect 3612 15876 3668 15932
rect 3948 15894 4004 15932
rect 3612 15810 3668 15820
rect 4060 15764 4116 17052
rect 4396 17106 4564 17108
rect 4396 17054 4510 17106
rect 4562 17054 4564 17106
rect 4396 17052 4564 17054
rect 4284 16884 4340 16894
rect 4172 16882 4340 16884
rect 4172 16830 4286 16882
rect 4338 16830 4340 16882
rect 4172 16828 4340 16830
rect 4172 16212 4228 16828
rect 4284 16818 4340 16828
rect 4396 16660 4452 17052
rect 4508 16996 4564 17052
rect 4732 17108 4788 17500
rect 4844 17462 4900 17500
rect 4956 17108 5012 17724
rect 5180 17668 5236 18844
rect 5292 18450 5348 19180
rect 5292 18398 5294 18450
rect 5346 18398 5348 18450
rect 5292 18386 5348 18398
rect 5516 18564 5572 20076
rect 5852 20130 5908 20188
rect 5852 20078 5854 20130
rect 5906 20078 5908 20130
rect 5852 20066 5908 20078
rect 6076 19460 6132 22652
rect 6188 20804 6244 23662
rect 6524 23604 6580 23886
rect 6748 23604 6804 24446
rect 6972 24052 7028 26236
rect 7756 26290 7812 27022
rect 9100 26962 9156 26974
rect 9100 26910 9102 26962
rect 9154 26910 9156 26962
rect 7756 26238 7758 26290
rect 7810 26238 7812 26290
rect 7532 25508 7588 25518
rect 7196 25394 7252 25406
rect 7196 25342 7198 25394
rect 7250 25342 7252 25394
rect 7196 24724 7252 25342
rect 7532 24948 7588 25452
rect 7644 25396 7700 25406
rect 7644 25302 7700 25340
rect 7532 24882 7588 24892
rect 7756 24724 7812 26238
rect 8204 26292 8260 26302
rect 8204 26198 8260 26236
rect 9100 25956 9156 26910
rect 9660 26964 9716 26974
rect 9100 25890 9156 25900
rect 9324 26404 9380 26414
rect 7868 25508 7924 25518
rect 7868 25414 7924 25452
rect 8876 25508 8932 25518
rect 8876 25414 8932 25452
rect 8428 25396 8484 25406
rect 8428 25302 8484 25340
rect 8092 25284 8148 25294
rect 7980 25228 8092 25284
rect 7868 24724 7924 24734
rect 7196 24722 7924 24724
rect 7196 24670 7870 24722
rect 7922 24670 7924 24722
rect 7196 24668 7924 24670
rect 7868 24658 7924 24668
rect 7196 24500 7252 24510
rect 7196 24498 7588 24500
rect 7196 24446 7198 24498
rect 7250 24446 7588 24498
rect 7196 24444 7588 24446
rect 7196 24434 7252 24444
rect 6972 23986 7028 23996
rect 6860 23940 6916 23950
rect 6860 23846 6916 23884
rect 7084 23940 7140 23950
rect 7084 23938 7476 23940
rect 7084 23886 7086 23938
rect 7138 23886 7476 23938
rect 7084 23884 7476 23886
rect 7084 23874 7140 23884
rect 6972 23716 7028 23726
rect 6972 23622 7028 23660
rect 7196 23716 7252 23726
rect 7420 23716 7476 23884
rect 7532 23938 7588 24444
rect 7868 23940 7924 23950
rect 7532 23886 7534 23938
rect 7586 23886 7588 23938
rect 7532 23874 7588 23886
rect 7644 23938 7924 23940
rect 7644 23886 7870 23938
rect 7922 23886 7924 23938
rect 7644 23884 7924 23886
rect 7644 23716 7700 23884
rect 7868 23874 7924 23884
rect 7420 23660 7700 23716
rect 7868 23716 7924 23726
rect 7980 23716 8036 25228
rect 8092 25218 8148 25228
rect 9324 25282 9380 26348
rect 9548 26290 9604 26302
rect 9548 26238 9550 26290
rect 9602 26238 9604 26290
rect 9324 25230 9326 25282
rect 9378 25230 9380 25282
rect 9324 25218 9380 25230
rect 9436 25506 9492 25518
rect 9436 25454 9438 25506
rect 9490 25454 9492 25506
rect 9436 25172 9492 25454
rect 9548 25284 9604 26238
rect 9548 25218 9604 25228
rect 7868 23714 8036 23716
rect 7868 23662 7870 23714
rect 7922 23662 8036 23714
rect 7868 23660 8036 23662
rect 8092 24948 8148 24958
rect 8092 24722 8148 24892
rect 8092 24670 8094 24722
rect 8146 24670 8148 24722
rect 8092 23716 8148 24670
rect 8316 24722 8372 24734
rect 8316 24670 8318 24722
rect 8370 24670 8372 24722
rect 8316 24500 8372 24670
rect 9100 24724 9156 24734
rect 9100 24630 9156 24668
rect 8316 24434 8372 24444
rect 9212 24052 9268 24062
rect 9436 24052 9492 25116
rect 9212 24050 9492 24052
rect 9212 23998 9214 24050
rect 9266 23998 9492 24050
rect 9212 23996 9492 23998
rect 9212 23986 9268 23996
rect 8204 23940 8260 23950
rect 8204 23846 8260 23884
rect 8540 23938 8596 23950
rect 8540 23886 8542 23938
rect 8594 23886 8596 23938
rect 7196 23622 7252 23660
rect 7868 23650 7924 23660
rect 8092 23650 8148 23660
rect 6524 23548 6804 23604
rect 6636 22932 6692 22942
rect 6636 22258 6692 22876
rect 6748 22708 6804 23548
rect 7308 23604 7364 23614
rect 7308 23378 7364 23548
rect 7308 23326 7310 23378
rect 7362 23326 7364 23378
rect 7308 23314 7364 23326
rect 7756 23604 7812 23614
rect 6860 23268 6916 23278
rect 6860 23174 6916 23212
rect 7084 23156 7140 23166
rect 6748 22652 6916 22708
rect 6636 22206 6638 22258
rect 6690 22206 6692 22258
rect 6636 22194 6692 22206
rect 6748 22370 6804 22382
rect 6748 22318 6750 22370
rect 6802 22318 6804 22370
rect 6524 21588 6580 21598
rect 6188 20710 6244 20748
rect 6412 21028 6468 21038
rect 6412 20802 6468 20972
rect 6412 20750 6414 20802
rect 6466 20750 6468 20802
rect 6412 20738 6468 20750
rect 6300 20578 6356 20590
rect 6300 20526 6302 20578
rect 6354 20526 6356 20578
rect 6300 20132 6356 20526
rect 6300 20066 6356 20076
rect 6524 20018 6580 21532
rect 6748 20242 6804 22318
rect 6748 20190 6750 20242
rect 6802 20190 6804 20242
rect 6748 20178 6804 20190
rect 6860 21586 6916 22652
rect 7084 22372 7140 23100
rect 7756 23154 7812 23548
rect 8540 23604 8596 23886
rect 8876 23828 8932 23838
rect 8876 23734 8932 23772
rect 8540 23538 8596 23548
rect 8764 23268 8820 23278
rect 8764 23266 8932 23268
rect 8764 23214 8766 23266
rect 8818 23214 8932 23266
rect 8764 23212 8932 23214
rect 8764 23202 8820 23212
rect 7756 23102 7758 23154
rect 7810 23102 7812 23154
rect 7084 22306 7140 22316
rect 7644 22370 7700 22382
rect 7644 22318 7646 22370
rect 7698 22318 7700 22370
rect 6860 21534 6862 21586
rect 6914 21534 6916 21586
rect 6860 20244 6916 21534
rect 7196 21588 7252 21598
rect 7196 21028 7252 21532
rect 7084 20972 7196 21028
rect 6972 20804 7028 20814
rect 6972 20710 7028 20748
rect 6860 20178 6916 20188
rect 6524 19966 6526 20018
rect 6578 19966 6580 20018
rect 6524 19954 6580 19966
rect 6860 20020 6916 20030
rect 7084 20020 7140 20972
rect 7196 20934 7252 20972
rect 7420 20804 7476 20814
rect 7644 20804 7700 22318
rect 7420 20802 7700 20804
rect 7420 20750 7422 20802
rect 7474 20750 7700 20802
rect 7420 20748 7700 20750
rect 7420 20356 7476 20748
rect 7420 20290 7476 20300
rect 7196 20132 7252 20142
rect 7196 20038 7252 20076
rect 7532 20130 7588 20142
rect 7532 20078 7534 20130
rect 7586 20078 7588 20130
rect 6860 20018 7140 20020
rect 6860 19966 6862 20018
rect 6914 19966 7140 20018
rect 6860 19964 7140 19966
rect 6860 19954 6916 19964
rect 6076 19394 6132 19404
rect 6300 19908 6356 19918
rect 5964 19348 6020 19358
rect 5740 19124 5796 19134
rect 5740 19030 5796 19068
rect 5852 18676 5908 18686
rect 5516 18450 5572 18508
rect 5516 18398 5518 18450
rect 5570 18398 5572 18450
rect 5516 18386 5572 18398
rect 5740 18620 5852 18676
rect 5740 18004 5796 18620
rect 5852 18610 5908 18620
rect 5852 18452 5908 18462
rect 5852 18358 5908 18396
rect 5740 17948 5908 18004
rect 5740 17780 5796 17790
rect 5740 17686 5796 17724
rect 5180 17602 5236 17612
rect 4732 17106 4900 17108
rect 4732 17054 4734 17106
rect 4786 17054 4900 17106
rect 4732 17052 4900 17054
rect 4956 17052 5124 17108
rect 4732 17042 4788 17052
rect 4508 16930 4564 16940
rect 4620 16772 4676 16782
rect 4620 16678 4676 16716
rect 4172 16146 4228 16156
rect 4284 16604 4452 16660
rect 4284 16098 4340 16604
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 4284 16046 4286 16098
rect 4338 16046 4340 16098
rect 4284 16034 4340 16046
rect 4508 16100 4564 16110
rect 4508 16006 4564 16044
rect 4732 15988 4788 15998
rect 4732 15894 4788 15932
rect 4060 15698 4116 15708
rect 4284 15876 4340 15886
rect 4284 15314 4340 15820
rect 4284 15262 4286 15314
rect 4338 15262 4340 15314
rect 3388 14590 3390 14642
rect 3442 14590 3444 14642
rect 3388 14578 3444 14590
rect 3836 15092 3892 15102
rect 3836 14642 3892 15036
rect 4284 14756 4340 15262
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 4284 14700 4676 14756
rect 3836 14590 3838 14642
rect 3890 14590 3892 14642
rect 3836 14578 3892 14590
rect 4620 14642 4676 14700
rect 4620 14590 4622 14642
rect 4674 14590 4676 14642
rect 4620 14578 4676 14590
rect 3164 13970 3332 13972
rect 3164 13918 3166 13970
rect 3218 13918 3332 13970
rect 3164 13916 3332 13918
rect 3612 13972 3668 13982
rect 3164 13906 3220 13916
rect 3612 13878 3668 13916
rect 4060 13636 4116 13646
rect 4060 13542 4116 13580
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 3164 13076 3220 13086
rect 3052 13074 3220 13076
rect 3052 13022 3166 13074
rect 3218 13022 3220 13074
rect 3052 13020 3220 13022
rect 3164 13010 3220 13020
rect 4844 12964 4900 17052
rect 4956 16882 5012 16894
rect 4956 16830 4958 16882
rect 5010 16830 5012 16882
rect 4956 15988 5012 16830
rect 5068 16212 5124 17052
rect 5292 16996 5348 17006
rect 5852 16996 5908 17948
rect 5292 16902 5348 16940
rect 5516 16940 5908 16996
rect 5068 16156 5236 16212
rect 5068 15988 5124 15998
rect 4956 15986 5124 15988
rect 4956 15934 5070 15986
rect 5122 15934 5124 15986
rect 4956 15932 5124 15934
rect 4956 15540 5012 15550
rect 4956 15446 5012 15484
rect 4956 14644 5012 14654
rect 4956 14550 5012 14588
rect 2716 12850 2884 12852
rect 2716 12798 2718 12850
rect 2770 12798 2884 12850
rect 2716 12796 2884 12798
rect 3612 12852 3668 12862
rect 2716 12786 2772 12796
rect 3612 12758 3668 12796
rect 4844 12404 4900 12908
rect 4956 12404 5012 12414
rect 4844 12402 5012 12404
rect 4844 12350 4958 12402
rect 5010 12350 5012 12402
rect 4844 12348 5012 12350
rect 4956 12338 5012 12348
rect 2492 12086 2548 12124
rect 4844 12178 4900 12190
rect 4844 12126 4846 12178
rect 4898 12126 4900 12178
rect 1708 11442 1764 11452
rect 2940 12066 2996 12078
rect 2940 12014 2942 12066
rect 2994 12014 2996 12066
rect 2940 11508 2996 12014
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 2940 11442 2996 11452
rect 1260 11218 1316 11228
rect 1708 11282 1764 11294
rect 1708 11230 1710 11282
rect 1762 11230 1764 11282
rect 1708 10836 1764 11230
rect 2044 11284 2100 11294
rect 2044 11190 2100 11228
rect 2492 11170 2548 11182
rect 2492 11118 2494 11170
rect 2546 11118 2548 11170
rect 1708 10770 1764 10780
rect 2044 10948 2100 10958
rect 2044 10834 2100 10892
rect 2044 10782 2046 10834
rect 2098 10782 2100 10834
rect 2044 10770 2100 10782
rect 2492 10836 2548 11118
rect 2492 10770 2548 10780
rect 4844 10724 4900 12126
rect 5068 11284 5124 15932
rect 5180 15540 5236 16156
rect 5516 15876 5572 16940
rect 5852 16882 5908 16940
rect 5852 16830 5854 16882
rect 5906 16830 5908 16882
rect 5852 16818 5908 16830
rect 5628 16772 5684 16782
rect 5684 16716 5796 16772
rect 5628 16706 5684 16716
rect 5740 16324 5796 16716
rect 5852 16324 5908 16334
rect 5740 16322 5908 16324
rect 5740 16270 5854 16322
rect 5906 16270 5908 16322
rect 5740 16268 5908 16270
rect 5852 16258 5908 16268
rect 5628 16100 5684 16110
rect 5628 16006 5684 16044
rect 5964 15876 6020 19292
rect 6076 19236 6132 19246
rect 6076 19142 6132 19180
rect 6300 19234 6356 19852
rect 7532 19908 7588 20078
rect 7532 19842 7588 19852
rect 6300 19182 6302 19234
rect 6354 19182 6356 19234
rect 6300 19170 6356 19182
rect 6860 19236 6916 19246
rect 6860 19142 6916 19180
rect 6412 19122 6468 19134
rect 7756 19124 7812 23102
rect 8204 23156 8260 23166
rect 8204 23062 8260 23100
rect 8652 23156 8708 23166
rect 8652 23062 8708 23100
rect 8764 22932 8820 22942
rect 8764 22838 8820 22876
rect 8204 21698 8260 21710
rect 8204 21646 8206 21698
rect 8258 21646 8260 21698
rect 8092 21474 8148 21486
rect 8092 21422 8094 21474
rect 8146 21422 8148 21474
rect 7868 20804 7924 20814
rect 7868 20710 7924 20748
rect 8092 20468 8148 21422
rect 8092 20402 8148 20412
rect 8204 20580 8260 21646
rect 8428 21586 8484 21598
rect 8652 21588 8708 21598
rect 8428 21534 8430 21586
rect 8482 21534 8484 21586
rect 8428 21028 8484 21534
rect 8316 20972 8484 21028
rect 8540 21586 8708 21588
rect 8540 21534 8654 21586
rect 8706 21534 8708 21586
rect 8540 21532 8708 21534
rect 8316 20580 8372 20972
rect 8428 20804 8484 20814
rect 8540 20804 8596 21532
rect 8652 21522 8708 21532
rect 8428 20802 8540 20804
rect 8428 20750 8430 20802
rect 8482 20750 8540 20802
rect 8428 20748 8540 20750
rect 8428 20738 8484 20748
rect 8540 20738 8596 20748
rect 8540 20580 8596 20590
rect 8316 20578 8596 20580
rect 8316 20526 8542 20578
rect 8594 20526 8596 20578
rect 8316 20524 8596 20526
rect 6412 19070 6414 19122
rect 6466 19070 6468 19122
rect 6300 18340 6356 18350
rect 6412 18340 6468 19070
rect 7532 19068 7812 19124
rect 6356 18284 6468 18340
rect 6300 18246 6356 18284
rect 6412 17780 6468 18284
rect 6972 18562 7028 18574
rect 6972 18510 6974 18562
rect 7026 18510 7028 18562
rect 6972 18004 7028 18510
rect 6524 17780 6580 17790
rect 6188 17778 6580 17780
rect 6188 17726 6526 17778
rect 6578 17726 6580 17778
rect 6188 17724 6580 17726
rect 6188 16322 6244 17724
rect 6524 17714 6580 17724
rect 6972 17554 7028 17948
rect 6972 17502 6974 17554
rect 7026 17502 7028 17554
rect 6972 17490 7028 17502
rect 6748 17332 6804 17342
rect 6300 17108 6356 17118
rect 6300 17014 6356 17052
rect 6748 17106 6804 17276
rect 6748 17054 6750 17106
rect 6802 17054 6804 17106
rect 6748 17042 6804 17054
rect 7532 16884 7588 19068
rect 7756 18452 7812 18462
rect 7812 18396 8036 18452
rect 7756 18358 7812 18396
rect 7644 18004 7700 18014
rect 7644 17106 7700 17948
rect 7980 17666 8036 18396
rect 7980 17614 7982 17666
rect 8034 17614 8036 17666
rect 7980 17602 8036 17614
rect 7644 17054 7646 17106
rect 7698 17054 7700 17106
rect 7644 17042 7700 17054
rect 7756 17444 7812 17454
rect 7756 16994 7812 17388
rect 7756 16942 7758 16994
rect 7810 16942 7812 16994
rect 7756 16930 7812 16942
rect 7532 16882 7700 16884
rect 7532 16830 7534 16882
rect 7586 16830 7700 16882
rect 7532 16828 7700 16830
rect 7532 16818 7588 16828
rect 7644 16772 7700 16828
rect 7644 16716 8036 16772
rect 6972 16324 7028 16334
rect 6188 16270 6190 16322
rect 6242 16270 6244 16322
rect 6188 16258 6244 16270
rect 6748 16268 6972 16324
rect 6636 16100 6692 16110
rect 5516 15820 5684 15876
rect 5180 15474 5236 15484
rect 5516 15204 5572 15242
rect 5516 15138 5572 15148
rect 5180 12180 5236 12190
rect 5180 12086 5236 12124
rect 5180 11396 5236 11406
rect 5628 11396 5684 15820
rect 5964 15810 6020 15820
rect 6412 16044 6636 16100
rect 5964 15540 6020 15550
rect 5964 13970 6020 15484
rect 6076 15202 6132 15214
rect 6076 15150 6078 15202
rect 6130 15150 6132 15202
rect 6076 14868 6132 15150
rect 6076 14802 6132 14812
rect 6412 14644 6468 16044
rect 6636 16006 6692 16044
rect 6524 15876 6580 15886
rect 6524 15426 6580 15820
rect 6524 15374 6526 15426
rect 6578 15374 6580 15426
rect 6524 15362 6580 15374
rect 6636 15204 6692 15214
rect 6748 15148 6804 16268
rect 6972 16230 7028 16268
rect 7420 16212 7476 16222
rect 6860 15874 6916 15886
rect 6860 15822 6862 15874
rect 6914 15822 6916 15874
rect 6860 15540 6916 15822
rect 7196 15876 7252 15886
rect 7196 15782 7252 15820
rect 7420 15874 7476 16156
rect 7980 16100 8036 16716
rect 7980 16006 8036 16044
rect 7532 15988 7588 15998
rect 7532 15986 7924 15988
rect 7532 15934 7534 15986
rect 7586 15934 7924 15986
rect 7532 15932 7924 15934
rect 7532 15922 7588 15932
rect 7420 15822 7422 15874
rect 7474 15822 7476 15874
rect 7420 15764 7476 15822
rect 7868 15876 7924 15932
rect 8204 15876 8260 20524
rect 8540 19908 8596 20524
rect 8764 20580 8820 20590
rect 8764 20486 8820 20524
rect 8876 20468 8932 23212
rect 9548 23156 9604 23166
rect 9100 23154 9604 23156
rect 9100 23102 9550 23154
rect 9602 23102 9604 23154
rect 9100 23100 9604 23102
rect 8988 22596 9044 22606
rect 8988 22502 9044 22540
rect 9100 21810 9156 23100
rect 9548 23090 9604 23100
rect 9100 21758 9102 21810
rect 9154 21758 9156 21810
rect 9100 21746 9156 21758
rect 9436 21588 9492 21598
rect 9100 21586 9492 21588
rect 9100 21534 9438 21586
rect 9490 21534 9492 21586
rect 9100 21532 9492 21534
rect 9100 20914 9156 21532
rect 9436 21522 9492 21532
rect 9660 21140 9716 26908
rect 9996 26740 10052 29148
rect 13468 28754 13524 29260
rect 13468 28702 13470 28754
rect 13522 28702 13524 28754
rect 13468 28690 13524 28702
rect 14588 28756 14644 29486
rect 14588 28690 14644 28700
rect 15148 29540 15204 29550
rect 15148 28980 15204 29484
rect 16716 29538 16772 31836
rect 16828 31826 16884 31836
rect 16940 31780 16996 31790
rect 16828 31668 16884 31678
rect 16940 31668 16996 31724
rect 16828 31666 16996 31668
rect 16828 31614 16830 31666
rect 16882 31614 16996 31666
rect 16828 31612 16996 31614
rect 16828 31602 16884 31612
rect 17052 31554 17108 31566
rect 17052 31502 17054 31554
rect 17106 31502 17108 31554
rect 17052 31332 17108 31502
rect 17052 31266 17108 31276
rect 16716 29486 16718 29538
rect 16770 29486 16772 29538
rect 16716 29474 16772 29486
rect 16828 30210 16884 30222
rect 16828 30158 16830 30210
rect 16882 30158 16884 30210
rect 16828 29540 16884 30158
rect 15596 29428 15652 29438
rect 15596 29334 15652 29372
rect 16604 29426 16660 29438
rect 16604 29374 16606 29426
rect 16658 29374 16660 29426
rect 15932 29316 15988 29326
rect 16604 29316 16660 29374
rect 16828 29316 16884 29484
rect 16604 29260 16884 29316
rect 15932 29222 15988 29260
rect 15148 27186 15204 28924
rect 15596 28756 15652 28766
rect 15596 28662 15652 28700
rect 16268 28644 16324 28654
rect 16268 27970 16324 28588
rect 16380 28642 16436 28654
rect 16380 28590 16382 28642
rect 16434 28590 16436 28642
rect 16380 28084 16436 28590
rect 17052 28644 17108 28654
rect 17052 28550 17108 28588
rect 17276 28308 17332 34412
rect 17612 34020 17668 35084
rect 17724 35046 17780 35084
rect 18844 35026 18900 35756
rect 18956 36482 19236 36484
rect 18956 36430 19182 36482
rect 19234 36430 19236 36482
rect 18956 36428 19236 36430
rect 18956 35810 19012 36428
rect 19180 36418 19236 36428
rect 19292 36482 19908 36484
rect 19292 36430 19854 36482
rect 19906 36430 19908 36482
rect 19292 36428 19908 36430
rect 18956 35758 18958 35810
rect 19010 35758 19012 35810
rect 18956 35308 19012 35758
rect 19180 35812 19236 35822
rect 19180 35718 19236 35756
rect 19292 35586 19348 36428
rect 19852 36418 19908 36428
rect 20188 36372 20244 37324
rect 20748 37268 20804 37278
rect 20748 36482 20804 37212
rect 20748 36430 20750 36482
rect 20802 36430 20804 36482
rect 20748 36418 20804 36430
rect 20188 36306 20244 36316
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 20860 35812 20916 38612
rect 21420 38050 21476 38892
rect 21532 38836 21588 38846
rect 21532 38742 21588 38780
rect 21420 37998 21422 38050
rect 21474 37998 21476 38050
rect 21420 37986 21476 37998
rect 21644 37940 21700 39228
rect 22428 38836 22484 38846
rect 22204 38724 22260 38762
rect 22428 38742 22484 38780
rect 21532 37938 21700 37940
rect 21532 37886 21646 37938
rect 21698 37886 21700 37938
rect 21532 37884 21700 37886
rect 21532 37828 21588 37884
rect 21644 37874 21700 37884
rect 21868 38610 21924 38622
rect 21868 38558 21870 38610
rect 21922 38558 21924 38610
rect 21420 37772 21588 37828
rect 21196 37380 21252 37390
rect 21196 37268 21252 37324
rect 21420 37378 21476 37772
rect 21420 37326 21422 37378
rect 21474 37326 21476 37378
rect 21420 37314 21476 37326
rect 21532 37268 21588 37278
rect 21196 37266 21364 37268
rect 21196 37214 21198 37266
rect 21250 37214 21364 37266
rect 21196 37212 21364 37214
rect 21196 37202 21252 37212
rect 21308 36482 21364 37212
rect 21868 37268 21924 38558
rect 22204 38162 22260 38668
rect 22204 38110 22206 38162
rect 22258 38110 22260 38162
rect 22204 38098 22260 38110
rect 22540 37938 22596 37950
rect 22540 37886 22542 37938
rect 22594 37886 22596 37938
rect 22540 37378 22596 37886
rect 22540 37326 22542 37378
rect 22594 37326 22596 37378
rect 22428 37268 22484 37278
rect 21868 37266 22484 37268
rect 21868 37214 22430 37266
rect 22482 37214 22484 37266
rect 21868 37212 22484 37214
rect 21532 37174 21588 37212
rect 22428 37202 22484 37212
rect 21980 37044 22036 37054
rect 22540 37044 22596 37326
rect 22652 37154 22708 40460
rect 22876 40402 22932 42140
rect 22876 40350 22878 40402
rect 22930 40350 22932 40402
rect 22876 40338 22932 40350
rect 22764 38612 22820 38622
rect 22764 38518 22820 38556
rect 22988 37268 23044 43036
rect 23100 41972 23156 41982
rect 23100 41878 23156 41916
rect 23324 41970 23380 41982
rect 23324 41918 23326 41970
rect 23378 41918 23380 41970
rect 23212 41746 23268 41758
rect 23212 41694 23214 41746
rect 23266 41694 23268 41746
rect 23212 41188 23268 41694
rect 23324 41524 23380 41918
rect 23324 41458 23380 41468
rect 23436 41412 23492 46396
rect 23772 46116 23828 46622
rect 23548 46060 23828 46116
rect 23548 45778 23604 46060
rect 24556 45892 24612 45902
rect 23548 45726 23550 45778
rect 23602 45726 23604 45778
rect 23548 44434 23604 45726
rect 23772 45890 24612 45892
rect 23772 45838 24558 45890
rect 24610 45838 24612 45890
rect 23772 45836 24612 45838
rect 23660 45332 23716 45342
rect 23772 45332 23828 45836
rect 24556 45826 24612 45836
rect 23660 45330 23828 45332
rect 23660 45278 23662 45330
rect 23714 45278 23828 45330
rect 23660 45276 23828 45278
rect 24332 45332 24388 45342
rect 23660 45266 23716 45276
rect 23548 44382 23550 44434
rect 23602 44382 23604 44434
rect 23548 44370 23604 44382
rect 23884 44322 23940 44334
rect 23884 44270 23886 44322
rect 23938 44270 23940 44322
rect 23772 44210 23828 44222
rect 23772 44158 23774 44210
rect 23826 44158 23828 44210
rect 23772 42866 23828 44158
rect 23772 42814 23774 42866
rect 23826 42814 23828 42866
rect 23660 41412 23716 41422
rect 23772 41412 23828 42814
rect 23884 43650 23940 44270
rect 23884 43598 23886 43650
rect 23938 43598 23940 43650
rect 23884 42756 23940 43598
rect 23884 41858 23940 42700
rect 24220 43652 24276 43662
rect 24220 42642 24276 43596
rect 24220 42590 24222 42642
rect 24274 42590 24276 42642
rect 23884 41806 23886 41858
rect 23938 41806 23940 41858
rect 23884 41794 23940 41806
rect 23996 41970 24052 41982
rect 23996 41918 23998 41970
rect 24050 41918 24052 41970
rect 23996 41412 24052 41918
rect 23436 41356 23604 41412
rect 23436 41188 23492 41198
rect 23212 41186 23492 41188
rect 23212 41134 23438 41186
rect 23490 41134 23492 41186
rect 23212 41132 23492 41134
rect 23436 41122 23492 41132
rect 23548 40964 23604 41356
rect 23660 41410 24052 41412
rect 23660 41358 23662 41410
rect 23714 41358 24052 41410
rect 23660 41356 24052 41358
rect 23660 41346 23716 41356
rect 23436 40908 23604 40964
rect 23772 40964 23828 40974
rect 23324 38612 23380 38622
rect 22988 37212 23156 37268
rect 22652 37102 22654 37154
rect 22706 37102 22708 37154
rect 22652 37090 22708 37102
rect 23100 37156 23156 37212
rect 23324 37266 23380 38556
rect 23324 37214 23326 37266
rect 23378 37214 23380 37266
rect 23324 37202 23380 37214
rect 23100 37100 23268 37156
rect 21980 37042 22596 37044
rect 21980 36990 21982 37042
rect 22034 36990 22596 37042
rect 21980 36988 22596 36990
rect 21980 36978 22036 36988
rect 22540 36708 22596 36988
rect 22876 37044 22932 37054
rect 22764 36708 22820 36718
rect 22540 36706 22820 36708
rect 22540 36654 22766 36706
rect 22818 36654 22820 36706
rect 22540 36652 22820 36654
rect 22764 36642 22820 36652
rect 21308 36430 21310 36482
rect 21362 36430 21364 36482
rect 21308 36418 21364 36430
rect 21644 36260 21700 36270
rect 21644 36166 21700 36204
rect 20860 35756 21252 35812
rect 19292 35534 19294 35586
rect 19346 35534 19348 35586
rect 18956 35252 19124 35308
rect 19068 35140 19124 35252
rect 19068 35046 19124 35084
rect 18844 34974 18846 35026
rect 18898 34974 18900 35026
rect 18844 34962 18900 34974
rect 19292 35028 19348 35534
rect 21084 35586 21140 35598
rect 21084 35534 21086 35586
rect 21138 35534 21140 35586
rect 19292 34962 19348 34972
rect 20188 35028 20244 35038
rect 20188 34934 20244 34972
rect 20412 35028 20468 35038
rect 19404 34916 19460 34926
rect 19740 34916 19796 34926
rect 19404 34914 19796 34916
rect 19404 34862 19406 34914
rect 19458 34862 19742 34914
rect 19794 34862 19796 34914
rect 19404 34860 19796 34862
rect 19404 34850 19460 34860
rect 19740 34850 19796 34860
rect 19964 34916 20020 34926
rect 19964 34914 20132 34916
rect 19964 34862 19966 34914
rect 20018 34862 20132 34914
rect 19964 34860 20132 34862
rect 19964 34850 20020 34860
rect 20076 34692 20132 34860
rect 20412 34914 20468 34972
rect 20412 34862 20414 34914
rect 20466 34862 20468 34914
rect 20412 34850 20468 34862
rect 20076 34636 20244 34692
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 20188 34356 20244 34636
rect 20076 34300 20244 34356
rect 20524 34690 20580 34702
rect 20524 34638 20526 34690
rect 20578 34638 20580 34690
rect 19740 34244 19796 34254
rect 19740 34150 19796 34188
rect 17612 33926 17668 33964
rect 19180 34020 19236 34030
rect 17724 33460 17780 33470
rect 17388 33012 17444 33022
rect 17388 32562 17444 32956
rect 17724 32564 17780 33404
rect 19180 33458 19236 33964
rect 19852 34020 19908 34030
rect 19516 33684 19572 33694
rect 19516 33570 19572 33628
rect 19516 33518 19518 33570
rect 19570 33518 19572 33570
rect 19516 33506 19572 33518
rect 19852 33570 19908 33964
rect 19852 33518 19854 33570
rect 19906 33518 19908 33570
rect 19852 33506 19908 33518
rect 19180 33406 19182 33458
rect 19234 33406 19236 33458
rect 19180 33394 19236 33406
rect 20076 33460 20132 34300
rect 20412 34132 20468 34142
rect 20076 33394 20132 33404
rect 20300 34076 20412 34132
rect 17836 33124 17892 33134
rect 17836 32786 17892 33068
rect 17836 32734 17838 32786
rect 17890 32734 17892 32786
rect 17836 32722 17892 32734
rect 18732 33124 18788 33134
rect 18732 32786 18788 33068
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 18732 32734 18734 32786
rect 18786 32734 18788 32786
rect 18732 32722 18788 32734
rect 19180 32788 19236 32798
rect 17388 32510 17390 32562
rect 17442 32510 17444 32562
rect 17388 32498 17444 32510
rect 17500 32562 17780 32564
rect 17500 32510 17726 32562
rect 17778 32510 17780 32562
rect 17500 32508 17780 32510
rect 17500 32002 17556 32508
rect 17724 32498 17780 32508
rect 18060 32562 18116 32574
rect 18060 32510 18062 32562
rect 18114 32510 18116 32562
rect 17948 32452 18004 32462
rect 17500 31950 17502 32002
rect 17554 31950 17556 32002
rect 17500 31892 17556 31950
rect 17500 31826 17556 31836
rect 17836 32450 18004 32452
rect 17836 32398 17950 32450
rect 18002 32398 18004 32450
rect 17836 32396 18004 32398
rect 17724 31778 17780 31790
rect 17724 31726 17726 31778
rect 17778 31726 17780 31778
rect 17388 31444 17444 31454
rect 17388 30882 17444 31388
rect 17724 31108 17780 31726
rect 17724 31042 17780 31052
rect 17388 30830 17390 30882
rect 17442 30830 17444 30882
rect 17388 30436 17444 30830
rect 17836 30772 17892 32396
rect 17948 32386 18004 32396
rect 18060 31780 18116 32510
rect 17948 31724 18116 31780
rect 19180 31890 19236 32732
rect 19180 31838 19182 31890
rect 19234 31838 19236 31890
rect 19180 31780 19236 31838
rect 17948 31554 18004 31724
rect 19180 31714 19236 31724
rect 18172 31668 18228 31678
rect 18172 31574 18228 31612
rect 18732 31668 18788 31678
rect 18732 31574 18788 31612
rect 17948 31502 17950 31554
rect 18002 31502 18004 31554
rect 17948 31332 18004 31502
rect 17948 31108 18004 31276
rect 17948 31042 18004 31052
rect 18060 31554 18116 31566
rect 18060 31502 18062 31554
rect 18114 31502 18116 31554
rect 17836 30706 17892 30716
rect 17388 30370 17444 30380
rect 17948 29540 18004 29550
rect 17388 28980 17444 28990
rect 17388 28866 17444 28924
rect 17388 28814 17390 28866
rect 17442 28814 17444 28866
rect 17388 28802 17444 28814
rect 17948 28642 18004 29484
rect 17948 28590 17950 28642
rect 18002 28590 18004 28642
rect 17948 28578 18004 28590
rect 18060 28530 18116 31502
rect 20300 31554 20356 34076
rect 20412 34038 20468 34076
rect 20524 33234 20580 34638
rect 20636 34692 20692 34702
rect 21084 34692 21140 35534
rect 20636 34690 21140 34692
rect 20636 34638 20638 34690
rect 20690 34638 21140 34690
rect 20636 34636 21140 34638
rect 20636 34626 20692 34636
rect 20524 33182 20526 33234
rect 20578 33182 20580 33234
rect 20524 33170 20580 33182
rect 20636 33346 20692 33358
rect 20636 33294 20638 33346
rect 20690 33294 20692 33346
rect 20636 33236 20692 33294
rect 20524 32788 20580 32798
rect 20636 32788 20692 33180
rect 20524 32786 20692 32788
rect 20524 32734 20526 32786
rect 20578 32734 20692 32786
rect 20524 32732 20692 32734
rect 20524 32722 20580 32732
rect 20300 31502 20302 31554
rect 20354 31502 20356 31554
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 20188 30996 20244 31006
rect 20300 30996 20356 31502
rect 20748 31554 20804 34636
rect 20860 34244 20916 34254
rect 20860 34150 20916 34188
rect 21084 34130 21140 34142
rect 21084 34078 21086 34130
rect 21138 34078 21140 34130
rect 21084 33684 21140 34078
rect 21084 33618 21140 33628
rect 20860 33236 20916 33246
rect 20860 32674 20916 33180
rect 20860 32622 20862 32674
rect 20914 32622 20916 32674
rect 20860 32610 20916 32622
rect 21196 31892 21252 35756
rect 21868 35028 21924 35038
rect 21868 34934 21924 34972
rect 21420 34690 21476 34702
rect 21420 34638 21422 34690
rect 21474 34638 21476 34690
rect 21420 34132 21476 34638
rect 21420 34066 21476 34076
rect 21756 34356 21812 34366
rect 21756 34020 21812 34300
rect 21756 34018 22260 34020
rect 21756 33966 21758 34018
rect 21810 33966 22260 34018
rect 21756 33964 22260 33966
rect 21756 33954 21812 33964
rect 21532 33572 21588 33582
rect 21588 33516 21700 33572
rect 21532 33506 21588 33516
rect 21420 33460 21476 33470
rect 21420 33234 21476 33404
rect 21420 33182 21422 33234
rect 21474 33182 21476 33234
rect 21420 33170 21476 33182
rect 20748 31502 20750 31554
rect 20802 31502 20804 31554
rect 20748 31444 20804 31502
rect 20244 30940 20356 30996
rect 20636 31220 20692 31230
rect 20636 30994 20692 31164
rect 20636 30942 20638 30994
rect 20690 30942 20692 30994
rect 20188 30902 20244 30940
rect 20636 30930 20692 30942
rect 19516 30884 19572 30894
rect 18508 30882 19572 30884
rect 18508 30830 19518 30882
rect 19570 30830 19572 30882
rect 18508 30828 19572 30830
rect 18284 30210 18340 30222
rect 18284 30158 18286 30210
rect 18338 30158 18340 30210
rect 18284 30100 18340 30158
rect 18284 30034 18340 30044
rect 18508 30098 18564 30828
rect 19516 30818 19572 30828
rect 20076 30884 20132 30894
rect 19404 30436 19460 30446
rect 19404 30342 19460 30380
rect 18508 30046 18510 30098
rect 18562 30046 18564 30098
rect 18508 30034 18564 30046
rect 19068 30100 19124 30110
rect 19068 30006 19124 30044
rect 20076 30098 20132 30828
rect 20748 30772 20804 31388
rect 20748 30706 20804 30716
rect 20860 31836 21252 31892
rect 21308 32562 21364 32574
rect 21308 32510 21310 32562
rect 21362 32510 21364 32562
rect 20188 30212 20244 30222
rect 20860 30212 20916 31836
rect 21308 31780 21364 32510
rect 21644 32452 21700 33516
rect 21756 33348 21812 33358
rect 21756 33254 21812 33292
rect 21756 32452 21812 32462
rect 21644 32396 21756 32452
rect 21756 32358 21812 32396
rect 22204 31892 22260 33964
rect 22876 33236 22932 36988
rect 23100 36932 23156 36942
rect 23100 36706 23156 36876
rect 23100 36654 23102 36706
rect 23154 36654 23156 36706
rect 23100 36642 23156 36654
rect 22988 36482 23044 36494
rect 22988 36430 22990 36482
rect 23042 36430 23044 36482
rect 22988 35812 23044 36430
rect 23100 36260 23156 36270
rect 23100 36166 23156 36204
rect 22988 33348 23044 35756
rect 22988 33282 23044 33292
rect 23100 33796 23156 33806
rect 22876 33170 22932 33180
rect 22204 31798 22260 31836
rect 22764 32452 22820 32462
rect 22764 31890 22820 32396
rect 22764 31838 22766 31890
rect 22818 31838 22820 31890
rect 22764 31826 22820 31838
rect 20188 30210 20356 30212
rect 20188 30158 20190 30210
rect 20242 30158 20356 30210
rect 20188 30156 20356 30158
rect 20188 30146 20244 30156
rect 20076 30046 20078 30098
rect 20130 30046 20132 30098
rect 20076 30034 20132 30046
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 20076 29652 20132 29662
rect 20076 29558 20132 29596
rect 20300 29540 20356 30156
rect 20860 30146 20916 30156
rect 20972 31724 21364 31780
rect 22988 31780 23044 31790
rect 23100 31780 23156 33740
rect 23212 33684 23268 37100
rect 23436 35812 23492 40908
rect 23772 40402 23828 40908
rect 23772 40350 23774 40402
rect 23826 40350 23828 40402
rect 23772 40338 23828 40350
rect 24108 39844 24164 39854
rect 24220 39844 24276 42590
rect 24332 40180 24388 45276
rect 24668 43708 24724 51660
rect 24780 51492 24836 51502
rect 24780 51398 24836 51436
rect 24892 50482 24948 50494
rect 24892 50430 24894 50482
rect 24946 50430 24948 50482
rect 24892 48804 24948 50430
rect 24892 48738 24948 48748
rect 24780 47346 24836 47358
rect 24780 47294 24782 47346
rect 24834 47294 24836 47346
rect 24780 45108 24836 47294
rect 24780 45042 24836 45052
rect 24556 43652 24724 43708
rect 24444 40404 24500 40414
rect 24444 40310 24500 40348
rect 24332 40124 24500 40180
rect 24108 39842 24276 39844
rect 24108 39790 24110 39842
rect 24162 39790 24276 39842
rect 24108 39788 24276 39790
rect 24108 39778 24164 39788
rect 23996 39620 24052 39630
rect 23996 39526 24052 39564
rect 23772 39394 23828 39406
rect 23772 39342 23774 39394
rect 23826 39342 23828 39394
rect 23772 39284 23828 39342
rect 24108 39394 24164 39406
rect 24108 39342 24110 39394
rect 24162 39342 24164 39394
rect 24108 39284 24164 39342
rect 23772 39228 24164 39284
rect 23884 39060 23940 39070
rect 23548 38836 23604 38846
rect 23548 38050 23604 38780
rect 23884 38668 23940 39004
rect 23996 38948 24052 38958
rect 24108 38948 24164 39228
rect 24220 38948 24276 38958
rect 23996 38946 24220 38948
rect 23996 38894 23998 38946
rect 24050 38894 24220 38946
rect 23996 38892 24220 38894
rect 23996 38882 24052 38892
rect 24220 38854 24276 38892
rect 24332 38946 24388 38958
rect 24332 38894 24334 38946
rect 24386 38894 24388 38946
rect 24332 38668 24388 38894
rect 23548 37998 23550 38050
rect 23602 37998 23604 38050
rect 23548 37986 23604 37998
rect 23660 38612 23940 38668
rect 24108 38612 24388 38668
rect 23660 36036 23716 38612
rect 23884 37268 23940 37278
rect 23884 37174 23940 37212
rect 24108 37266 24164 38612
rect 24444 38276 24500 40124
rect 24556 39060 24612 43652
rect 24668 43540 24724 43550
rect 24668 41970 24724 43484
rect 24668 41918 24670 41970
rect 24722 41918 24724 41970
rect 24668 41906 24724 41918
rect 24556 38994 24612 39004
rect 25004 39618 25060 53452
rect 25676 52946 25732 53452
rect 25676 52894 25678 52946
rect 25730 52894 25732 52946
rect 25676 52882 25732 52894
rect 26236 52946 26292 53564
rect 26236 52894 26238 52946
rect 26290 52894 26292 52946
rect 25340 52836 25396 52846
rect 25340 52742 25396 52780
rect 26012 52388 26068 52398
rect 26012 52162 26068 52332
rect 26236 52274 26292 52894
rect 26460 53058 26516 53070
rect 26460 53006 26462 53058
rect 26514 53006 26516 53058
rect 26236 52222 26238 52274
rect 26290 52222 26292 52274
rect 26236 52210 26292 52222
rect 26348 52834 26404 52846
rect 26348 52782 26350 52834
rect 26402 52782 26404 52834
rect 26012 52110 26014 52162
rect 26066 52110 26068 52162
rect 26012 52098 26068 52110
rect 26348 52164 26404 52782
rect 26460 52388 26516 53006
rect 27020 52500 27076 54348
rect 27020 52444 27300 52500
rect 26460 52322 26516 52332
rect 27132 52276 27188 52286
rect 25564 51492 25620 51502
rect 25564 51398 25620 51436
rect 25676 51492 25732 51502
rect 26348 51492 26404 52108
rect 26796 52274 27188 52276
rect 26796 52222 27134 52274
rect 27186 52222 27188 52274
rect 26796 52220 27188 52222
rect 26684 52052 26740 52062
rect 25676 51490 26404 51492
rect 25676 51438 25678 51490
rect 25730 51438 26350 51490
rect 26402 51438 26404 51490
rect 25676 51436 26404 51438
rect 25676 51426 25732 51436
rect 26348 51426 26404 51436
rect 26460 52050 26740 52052
rect 26460 51998 26686 52050
rect 26738 51998 26740 52050
rect 26460 51996 26740 51998
rect 26012 51266 26068 51278
rect 26012 51214 26014 51266
rect 26066 51214 26068 51266
rect 25564 51156 25620 51166
rect 25564 51062 25620 51100
rect 26012 50708 26068 51214
rect 26012 50642 26068 50652
rect 25676 50596 25732 50606
rect 25676 50502 25732 50540
rect 25788 50484 25844 50494
rect 25676 50372 25844 50428
rect 25676 49476 25732 50372
rect 26012 50370 26068 50382
rect 26012 50318 26014 50370
rect 26066 50318 26068 50370
rect 25788 49924 25844 49934
rect 26012 49924 26068 50318
rect 25788 49922 26068 49924
rect 25788 49870 25790 49922
rect 25842 49870 26068 49922
rect 25788 49868 26068 49870
rect 26460 50148 26516 51996
rect 26684 51986 26740 51996
rect 26684 50596 26740 50606
rect 26796 50596 26852 52220
rect 27132 52210 27188 52220
rect 27020 52052 27076 52062
rect 27020 51958 27076 51996
rect 26684 50594 26852 50596
rect 26684 50542 26686 50594
rect 26738 50542 26852 50594
rect 26684 50540 26852 50542
rect 27020 51156 27076 51166
rect 27020 50594 27076 51100
rect 27020 50542 27022 50594
rect 27074 50542 27076 50594
rect 26684 50530 26740 50540
rect 27020 50530 27076 50542
rect 27244 50428 27300 52444
rect 27356 52162 27412 52174
rect 27356 52110 27358 52162
rect 27410 52110 27412 52162
rect 27356 51492 27412 52110
rect 27468 51716 27524 54348
rect 27692 53172 27748 55022
rect 27916 54404 27972 56028
rect 28252 55468 28308 59200
rect 28588 55972 28644 55982
rect 28588 55878 28644 55916
rect 28924 55524 28980 59200
rect 29596 55468 29652 59200
rect 28140 55412 28196 55422
rect 28252 55412 28644 55468
rect 28924 55458 28980 55468
rect 29372 55412 29876 55468
rect 28140 55318 28196 55356
rect 28588 55410 28868 55412
rect 28588 55358 28590 55410
rect 28642 55358 28868 55410
rect 28588 55356 28868 55358
rect 28588 55346 28644 55356
rect 28476 55300 28532 55310
rect 28812 55300 28868 55356
rect 29148 55300 29204 55310
rect 28812 55298 29204 55300
rect 28812 55246 29150 55298
rect 29202 55246 29204 55298
rect 28812 55244 29204 55246
rect 28476 54628 28532 55244
rect 29148 55234 29204 55244
rect 29372 55076 29428 55412
rect 28924 55020 29428 55076
rect 29708 55298 29764 55310
rect 29708 55246 29710 55298
rect 29762 55246 29764 55298
rect 28924 54738 28980 55020
rect 29148 54852 29204 54862
rect 28924 54686 28926 54738
rect 28978 54686 28980 54738
rect 28924 54674 28980 54686
rect 29036 54796 29148 54852
rect 28476 54534 28532 54572
rect 27692 53106 27748 53116
rect 27804 54402 27972 54404
rect 27804 54350 27918 54402
rect 27970 54350 27972 54402
rect 27804 54348 27972 54350
rect 27468 51660 27748 51716
rect 27356 51378 27412 51436
rect 27356 51326 27358 51378
rect 27410 51326 27412 51378
rect 27356 51314 27412 51326
rect 27580 51490 27636 51502
rect 27580 51438 27582 51490
rect 27634 51438 27636 51490
rect 25788 49812 25844 49868
rect 25788 49746 25844 49756
rect 25900 49700 25956 49710
rect 25900 49606 25956 49644
rect 26012 49700 26068 49710
rect 26460 49700 26516 50092
rect 27132 50372 27300 50428
rect 27468 50706 27524 50718
rect 27468 50654 27470 50706
rect 27522 50654 27524 50706
rect 26908 49922 26964 49934
rect 26908 49870 26910 49922
rect 26962 49870 26964 49922
rect 26012 49698 26516 49700
rect 26012 49646 26014 49698
rect 26066 49646 26516 49698
rect 26012 49644 26516 49646
rect 26796 49700 26852 49710
rect 26012 49634 26068 49644
rect 25676 49420 25844 49476
rect 25676 48468 25732 48478
rect 25676 48354 25732 48412
rect 25676 48302 25678 48354
rect 25730 48302 25732 48354
rect 25676 48244 25732 48302
rect 25788 48356 25844 49420
rect 26796 49026 26852 49644
rect 26908 49140 26964 49870
rect 26908 49084 27076 49140
rect 26796 48974 26798 49026
rect 26850 48974 26852 49026
rect 26796 48962 26852 48974
rect 27020 49026 27076 49084
rect 27020 48974 27022 49026
rect 27074 48974 27076 49026
rect 26012 48804 26068 48814
rect 27020 48804 27076 48974
rect 25788 48354 25956 48356
rect 25788 48302 25790 48354
rect 25842 48302 25956 48354
rect 25788 48300 25956 48302
rect 25788 48290 25844 48300
rect 25676 47572 25732 48188
rect 25788 48020 25844 48030
rect 25788 47926 25844 47964
rect 25900 47684 25956 48300
rect 25900 47618 25956 47628
rect 25676 47516 25844 47572
rect 25564 47348 25620 47358
rect 25452 47346 25620 47348
rect 25452 47294 25566 47346
rect 25618 47294 25620 47346
rect 25452 47292 25620 47294
rect 25116 45666 25172 45678
rect 25116 45614 25118 45666
rect 25170 45614 25172 45666
rect 25116 43764 25172 45614
rect 25116 43698 25172 43708
rect 25340 43652 25396 43662
rect 25340 43558 25396 43596
rect 25228 43540 25284 43550
rect 25228 43446 25284 43484
rect 25452 42980 25508 47292
rect 25564 47282 25620 47292
rect 25788 46898 25844 47516
rect 26012 47460 26068 48748
rect 26684 48748 27076 48804
rect 25788 46846 25790 46898
rect 25842 46846 25844 46898
rect 25788 46834 25844 46846
rect 25900 47458 26068 47460
rect 25900 47406 26014 47458
rect 26066 47406 26068 47458
rect 25900 47404 26068 47406
rect 25564 46676 25620 46686
rect 25900 46676 25956 47404
rect 26012 47394 26068 47404
rect 26124 48412 26516 48468
rect 25564 46674 25956 46676
rect 25564 46622 25566 46674
rect 25618 46622 25956 46674
rect 25564 46620 25956 46622
rect 26012 46900 26068 46910
rect 26124 46900 26180 48412
rect 26236 48244 26292 48254
rect 26236 48150 26292 48188
rect 26460 48242 26516 48412
rect 26460 48190 26462 48242
rect 26514 48190 26516 48242
rect 26460 48178 26516 48190
rect 26348 48130 26404 48142
rect 26348 48078 26350 48130
rect 26402 48078 26404 48130
rect 26012 46898 26180 46900
rect 26012 46846 26014 46898
rect 26066 46846 26180 46898
rect 26012 46844 26180 46846
rect 26236 47684 26292 47694
rect 25564 46610 25620 46620
rect 26012 45892 26068 46844
rect 26124 46676 26180 46686
rect 26124 46582 26180 46620
rect 26236 46452 26292 47628
rect 26348 46674 26404 48078
rect 26572 46900 26628 46910
rect 26684 46900 26740 48748
rect 26796 48580 26852 48590
rect 26796 48354 26852 48524
rect 26796 48302 26798 48354
rect 26850 48302 26852 48354
rect 26796 48290 26852 48302
rect 27020 48020 27076 48030
rect 27020 47458 27076 47964
rect 27020 47406 27022 47458
rect 27074 47406 27076 47458
rect 27020 47394 27076 47406
rect 27132 46900 27188 50372
rect 27244 49812 27300 49822
rect 27244 48916 27300 49756
rect 27244 48850 27300 48860
rect 26572 46898 26740 46900
rect 26572 46846 26574 46898
rect 26626 46846 26740 46898
rect 26572 46844 26740 46846
rect 27020 46844 27188 46900
rect 27356 47458 27412 47470
rect 27356 47406 27358 47458
rect 27410 47406 27412 47458
rect 26572 46834 26628 46844
rect 26348 46622 26350 46674
rect 26402 46622 26404 46674
rect 26348 46610 26404 46622
rect 26908 46676 26964 46686
rect 26908 46582 26964 46620
rect 27020 46452 27076 46844
rect 27356 46788 27412 47406
rect 26236 46396 26404 46452
rect 26012 45890 26292 45892
rect 26012 45838 26014 45890
rect 26066 45838 26292 45890
rect 26012 45836 26292 45838
rect 25788 44322 25844 44334
rect 25788 44270 25790 44322
rect 25842 44270 25844 44322
rect 25564 43538 25620 43550
rect 25564 43486 25566 43538
rect 25618 43486 25620 43538
rect 25564 43204 25620 43486
rect 25564 43138 25620 43148
rect 25228 42924 25508 42980
rect 25788 42980 25844 44270
rect 26012 44210 26068 45836
rect 26124 45668 26180 45678
rect 26124 45108 26180 45612
rect 26236 45332 26292 45836
rect 26348 45666 26404 46396
rect 27020 46386 27076 46396
rect 27132 46786 27412 46788
rect 27132 46734 27358 46786
rect 27410 46734 27412 46786
rect 27132 46732 27412 46734
rect 27132 46002 27188 46732
rect 27356 46722 27412 46732
rect 27132 45950 27134 46002
rect 27186 45950 27188 46002
rect 27132 45938 27188 45950
rect 27020 45668 27076 45678
rect 26348 45614 26350 45666
rect 26402 45614 26404 45666
rect 26348 45556 26404 45614
rect 26908 45666 27076 45668
rect 26908 45614 27022 45666
rect 27074 45614 27076 45666
rect 26908 45612 27076 45614
rect 26348 45500 26740 45556
rect 26348 45332 26404 45342
rect 26236 45330 26404 45332
rect 26236 45278 26350 45330
rect 26402 45278 26404 45330
rect 26236 45276 26404 45278
rect 26348 45266 26404 45276
rect 26572 45220 26628 45230
rect 26572 45126 26628 45164
rect 26236 45108 26292 45118
rect 26124 45106 26292 45108
rect 26124 45054 26238 45106
rect 26290 45054 26292 45106
rect 26124 45052 26292 45054
rect 26236 45042 26292 45052
rect 26012 44158 26014 44210
rect 26066 44158 26068 44210
rect 26012 44146 26068 44158
rect 26572 44100 26628 44110
rect 26572 44006 26628 44044
rect 26684 43708 26740 45500
rect 26908 45330 26964 45612
rect 27020 45602 27076 45612
rect 27244 45668 27300 45678
rect 27244 45574 27300 45612
rect 27468 45332 27524 50654
rect 27580 50482 27636 51438
rect 27580 50430 27582 50482
rect 27634 50430 27636 50482
rect 27580 49250 27636 50430
rect 27580 49198 27582 49250
rect 27634 49198 27636 49250
rect 27580 49186 27636 49198
rect 27692 46116 27748 51660
rect 27804 46340 27860 54348
rect 27916 54338 27972 54348
rect 28812 53732 28868 53742
rect 28812 50428 28868 53676
rect 28700 50372 28868 50428
rect 27916 50148 27972 50158
rect 27916 49810 27972 50092
rect 27916 49758 27918 49810
rect 27970 49758 27972 49810
rect 27916 49028 27972 49758
rect 28588 49700 28644 49710
rect 28588 49606 28644 49644
rect 27916 48962 27972 48972
rect 28028 49028 28084 49038
rect 28252 49028 28308 49038
rect 28028 49026 28308 49028
rect 28028 48974 28030 49026
rect 28082 48974 28254 49026
rect 28306 48974 28308 49026
rect 28028 48972 28308 48974
rect 28028 48962 28084 48972
rect 28252 48962 28308 48972
rect 28588 49028 28644 49038
rect 28588 48934 28644 48972
rect 28476 48916 28532 48926
rect 28476 48822 28532 48860
rect 27804 46274 27860 46284
rect 27692 46060 27972 46116
rect 26908 45278 26910 45330
rect 26962 45278 26964 45330
rect 26908 45266 26964 45278
rect 27356 45276 27524 45332
rect 27692 45890 27748 45902
rect 27692 45838 27694 45890
rect 27746 45838 27748 45890
rect 27692 45332 27748 45838
rect 27804 45332 27860 45342
rect 27692 45330 27860 45332
rect 27692 45278 27806 45330
rect 27858 45278 27860 45330
rect 27692 45276 27860 45278
rect 27132 45220 27188 45230
rect 26796 45108 26852 45118
rect 26796 44322 26852 45052
rect 27132 45106 27188 45164
rect 27132 45054 27134 45106
rect 27186 45054 27188 45106
rect 27132 45042 27188 45054
rect 26796 44270 26798 44322
rect 26850 44270 26852 44322
rect 26796 44258 26852 44270
rect 26684 43652 27076 43708
rect 26796 43540 26852 43550
rect 26236 43428 26292 43438
rect 25116 41074 25172 41086
rect 25116 41022 25118 41074
rect 25170 41022 25172 41074
rect 25116 40404 25172 41022
rect 25116 40338 25172 40348
rect 25004 39566 25006 39618
rect 25058 39566 25060 39618
rect 25004 38948 25060 39566
rect 25228 39620 25284 42924
rect 25788 42914 25844 42924
rect 26012 43426 26292 43428
rect 26012 43374 26238 43426
rect 26290 43374 26292 43426
rect 26012 43372 26292 43374
rect 25340 42756 25396 42766
rect 25340 42662 25396 42700
rect 25788 42532 25844 42542
rect 26012 42532 26068 43372
rect 26236 43362 26292 43372
rect 26348 43316 26404 43326
rect 26348 43222 26404 43260
rect 26124 43204 26180 43214
rect 26180 43148 26292 43204
rect 26124 43138 26180 43148
rect 25788 42530 26068 42532
rect 25788 42478 25790 42530
rect 25842 42478 26068 42530
rect 25788 42476 26068 42478
rect 26124 42980 26180 42990
rect 25788 41970 25844 42476
rect 26124 42196 26180 42924
rect 26236 42754 26292 43148
rect 26796 42866 26852 43484
rect 26796 42814 26798 42866
rect 26850 42814 26852 42866
rect 26796 42802 26852 42814
rect 26908 43316 26964 43326
rect 26236 42702 26238 42754
rect 26290 42702 26292 42754
rect 26236 42690 26292 42702
rect 26908 42754 26964 43260
rect 26908 42702 26910 42754
rect 26962 42702 26964 42754
rect 26908 42690 26964 42702
rect 26684 42532 26740 42542
rect 25788 41918 25790 41970
rect 25842 41918 25844 41970
rect 25788 41906 25844 41918
rect 25900 42140 26180 42196
rect 26348 42530 26740 42532
rect 26348 42478 26686 42530
rect 26738 42478 26740 42530
rect 26348 42476 26740 42478
rect 25676 41860 25732 41870
rect 25676 41766 25732 41804
rect 25900 41636 25956 42140
rect 26348 41972 26404 42476
rect 26684 42466 26740 42476
rect 26796 42532 26852 42542
rect 25564 41580 25956 41636
rect 26012 41970 26404 41972
rect 26012 41918 26350 41970
rect 26402 41918 26404 41970
rect 26012 41916 26404 41918
rect 25564 41074 25620 41580
rect 26012 41298 26068 41916
rect 26348 41906 26404 41916
rect 26796 41300 26852 42476
rect 26012 41246 26014 41298
rect 26066 41246 26068 41298
rect 26012 41234 26068 41246
rect 26572 41244 26852 41300
rect 25564 41022 25566 41074
rect 25618 41022 25620 41074
rect 25340 40964 25396 40974
rect 25340 40870 25396 40908
rect 25564 40852 25620 41022
rect 25676 41076 25732 41086
rect 25900 41076 25956 41086
rect 25676 41074 25956 41076
rect 25676 41022 25678 41074
rect 25730 41022 25902 41074
rect 25954 41022 25956 41074
rect 25676 41020 25956 41022
rect 25676 41010 25732 41020
rect 25900 41010 25956 41020
rect 26236 41076 26292 41086
rect 26236 41074 26404 41076
rect 26236 41022 26238 41074
rect 26290 41022 26404 41074
rect 26236 41020 26404 41022
rect 26236 41010 26292 41020
rect 26012 40964 26068 40974
rect 25900 40852 25956 40862
rect 25564 40796 25732 40852
rect 25676 40516 25732 40796
rect 25900 40626 25956 40796
rect 25900 40574 25902 40626
rect 25954 40574 25956 40626
rect 25900 40562 25956 40574
rect 25676 40514 25844 40516
rect 25676 40462 25678 40514
rect 25730 40462 25844 40514
rect 25676 40460 25844 40462
rect 25676 40450 25732 40460
rect 25564 40404 25620 40414
rect 25564 40180 25620 40348
rect 25564 40124 25732 40180
rect 25228 39564 25396 39620
rect 25228 39396 25284 39406
rect 25228 39302 25284 39340
rect 25340 39172 25396 39564
rect 25004 38882 25060 38892
rect 25228 39116 25396 39172
rect 25564 39506 25620 39518
rect 25564 39454 25566 39506
rect 25618 39454 25620 39506
rect 24556 38834 24612 38846
rect 24556 38782 24558 38834
rect 24610 38782 24612 38834
rect 24556 38668 24612 38782
rect 24556 38612 24836 38668
rect 24444 38220 24724 38276
rect 24556 38050 24612 38062
rect 24556 37998 24558 38050
rect 24610 37998 24612 38050
rect 24220 37940 24276 37950
rect 24556 37940 24612 37998
rect 24220 37938 24612 37940
rect 24220 37886 24222 37938
rect 24274 37886 24612 37938
rect 24220 37884 24612 37886
rect 24220 37874 24276 37884
rect 24556 37604 24612 37884
rect 24556 37538 24612 37548
rect 24444 37380 24500 37390
rect 24668 37380 24724 38220
rect 24108 37214 24110 37266
rect 24162 37214 24164 37266
rect 24108 36372 24164 37214
rect 24108 36306 24164 36316
rect 24220 37378 24724 37380
rect 24220 37326 24446 37378
rect 24498 37326 24724 37378
rect 24220 37324 24724 37326
rect 24780 38050 24836 38612
rect 25116 38276 25172 38286
rect 25116 38182 25172 38220
rect 24780 37998 24782 38050
rect 24834 37998 24836 38050
rect 23772 36258 23828 36270
rect 23772 36206 23774 36258
rect 23826 36206 23828 36258
rect 23772 36148 23828 36206
rect 24220 36148 24276 37324
rect 24444 37314 24500 37324
rect 24332 37154 24388 37166
rect 24332 37102 24334 37154
rect 24386 37102 24388 37154
rect 24332 37044 24388 37102
rect 24332 36978 24388 36988
rect 24780 36706 24836 37998
rect 25116 38052 25172 38062
rect 24780 36654 24782 36706
rect 24834 36654 24836 36706
rect 24780 36642 24836 36654
rect 25004 37604 25060 37614
rect 25004 36370 25060 37548
rect 25116 36706 25172 37996
rect 25116 36654 25118 36706
rect 25170 36654 25172 36706
rect 25116 36642 25172 36654
rect 25004 36318 25006 36370
rect 25058 36318 25060 36370
rect 25004 36306 25060 36318
rect 23772 36092 24276 36148
rect 23212 33618 23268 33628
rect 23324 35756 23492 35812
rect 23548 35980 23716 36036
rect 23324 32788 23380 35756
rect 23436 35588 23492 35598
rect 23436 35494 23492 35532
rect 23548 34356 23604 35980
rect 23660 35812 23716 35822
rect 23660 35718 23716 35756
rect 25228 35698 25284 39116
rect 25340 38948 25396 38958
rect 25340 38854 25396 38892
rect 25564 38500 25620 39454
rect 25676 39508 25732 40124
rect 25788 39732 25844 40460
rect 26012 40404 26068 40908
rect 26348 40628 26404 41020
rect 26460 41074 26516 41086
rect 26460 41022 26462 41074
rect 26514 41022 26516 41074
rect 26460 40852 26516 41022
rect 26460 40786 26516 40796
rect 26348 40572 26516 40628
rect 26348 40404 26404 40414
rect 25900 40402 26068 40404
rect 25900 40350 26014 40402
rect 26066 40350 26068 40402
rect 25900 40348 26068 40350
rect 25900 39956 25956 40348
rect 26012 40338 26068 40348
rect 26124 40402 26404 40404
rect 26124 40350 26350 40402
rect 26402 40350 26404 40402
rect 26124 40348 26404 40350
rect 25900 39890 25956 39900
rect 25788 39676 25956 39732
rect 25788 39508 25844 39518
rect 25676 39506 25844 39508
rect 25676 39454 25790 39506
rect 25842 39454 25844 39506
rect 25676 39452 25844 39454
rect 25788 39442 25844 39452
rect 25900 39396 25956 39676
rect 25900 39330 25956 39340
rect 26012 39060 26068 39070
rect 26124 39060 26180 40348
rect 26348 40338 26404 40348
rect 26460 39508 26516 40572
rect 26460 39442 26516 39452
rect 26012 39058 26180 39060
rect 26012 39006 26014 39058
rect 26066 39006 26180 39058
rect 26012 39004 26180 39006
rect 26012 38668 26068 39004
rect 25564 38434 25620 38444
rect 25788 38612 26068 38668
rect 25340 38388 25396 38398
rect 25340 37380 25396 38332
rect 25452 38052 25508 38090
rect 25452 37986 25508 37996
rect 25676 38052 25732 38090
rect 25676 37986 25732 37996
rect 25676 37716 25732 37726
rect 25564 37660 25676 37716
rect 25340 37324 25508 37380
rect 25228 35646 25230 35698
rect 25282 35646 25284 35698
rect 25228 35634 25284 35646
rect 25340 37154 25396 37166
rect 25340 37102 25342 37154
rect 25394 37102 25396 37154
rect 24668 35586 24724 35598
rect 24668 35534 24670 35586
rect 24722 35534 24724 35586
rect 23772 35476 23828 35486
rect 23772 35474 24276 35476
rect 23772 35422 23774 35474
rect 23826 35422 24276 35474
rect 23772 35420 24276 35422
rect 23772 35410 23828 35420
rect 23996 34916 24052 34926
rect 23996 34822 24052 34860
rect 24220 34914 24276 35420
rect 24220 34862 24222 34914
rect 24274 34862 24276 34914
rect 24220 34850 24276 34862
rect 24556 35252 24612 35262
rect 24556 34914 24612 35196
rect 24556 34862 24558 34914
rect 24610 34862 24612 34914
rect 24556 34850 24612 34862
rect 24668 34916 24724 35534
rect 25340 35588 25396 37102
rect 25340 35364 25396 35532
rect 25116 35308 25396 35364
rect 25004 34916 25060 34926
rect 25116 34916 25172 35308
rect 24668 34914 25172 34916
rect 24668 34862 25006 34914
rect 25058 34862 25172 34914
rect 24668 34860 25172 34862
rect 24332 34690 24388 34702
rect 24332 34638 24334 34690
rect 24386 34638 24388 34690
rect 24332 34356 24388 34638
rect 24444 34692 24500 34702
rect 24444 34598 24500 34636
rect 23548 34300 23716 34356
rect 23548 34132 23604 34142
rect 23548 33458 23604 34076
rect 23548 33406 23550 33458
rect 23602 33406 23604 33458
rect 23548 33394 23604 33406
rect 23436 32788 23492 32798
rect 23324 32732 23436 32788
rect 23436 32722 23492 32732
rect 23660 31890 23716 34300
rect 24332 34290 24388 34300
rect 24556 34132 24612 34142
rect 23884 34020 23940 34030
rect 23884 33926 23940 33964
rect 23996 33012 24052 33022
rect 23884 32450 23940 32462
rect 23884 32398 23886 32450
rect 23938 32398 23940 32450
rect 23884 32002 23940 32398
rect 23884 31950 23886 32002
rect 23938 31950 23940 32002
rect 23884 31938 23940 31950
rect 23660 31838 23662 31890
rect 23714 31838 23716 31890
rect 23100 31724 23268 31780
rect 20300 29446 20356 29484
rect 20412 29988 20468 29998
rect 18060 28478 18062 28530
rect 18114 28478 18116 28530
rect 18060 28466 18116 28478
rect 18172 29314 18228 29326
rect 18172 29262 18174 29314
rect 18226 29262 18228 29314
rect 17276 28242 17332 28252
rect 18060 28308 18116 28318
rect 16380 28018 16436 28028
rect 17948 28084 18004 28094
rect 16268 27918 16270 27970
rect 16322 27918 16324 27970
rect 16268 27906 16324 27918
rect 16604 27970 16660 27982
rect 16604 27918 16606 27970
rect 16658 27918 16660 27970
rect 15148 27134 15150 27186
rect 15202 27134 15204 27186
rect 15148 27122 15204 27134
rect 16604 27188 16660 27918
rect 17612 27972 17668 27982
rect 16604 27122 16660 27132
rect 17276 27188 17332 27198
rect 17276 27094 17332 27132
rect 17612 26908 17668 27916
rect 17948 27074 18004 28028
rect 18060 28082 18116 28252
rect 18172 28196 18228 29262
rect 19628 29314 19684 29326
rect 19628 29262 19630 29314
rect 19682 29262 19684 29314
rect 19628 29204 19684 29262
rect 19628 29138 19684 29148
rect 19068 28868 19124 28878
rect 19068 28756 19124 28812
rect 19068 28754 19572 28756
rect 19068 28702 19070 28754
rect 19122 28702 19572 28754
rect 19068 28700 19572 28702
rect 19068 28690 19124 28700
rect 19292 28532 19348 28542
rect 19180 28530 19348 28532
rect 19180 28478 19294 28530
rect 19346 28478 19348 28530
rect 19180 28476 19348 28478
rect 18172 28130 18228 28140
rect 18508 28196 18564 28206
rect 19180 28196 19236 28476
rect 19292 28466 19348 28476
rect 19516 28530 19572 28700
rect 19516 28478 19518 28530
rect 19570 28478 19572 28530
rect 19516 28466 19572 28478
rect 19628 28754 19684 28766
rect 19628 28702 19630 28754
rect 19682 28702 19684 28754
rect 18060 28030 18062 28082
rect 18114 28030 18116 28082
rect 18060 27748 18116 28030
rect 18508 28082 18564 28140
rect 18508 28030 18510 28082
rect 18562 28030 18564 28082
rect 18508 28018 18564 28030
rect 18732 28140 19236 28196
rect 18732 28082 18788 28140
rect 18732 28030 18734 28082
rect 18786 28030 18788 28082
rect 18732 28018 18788 28030
rect 19068 27972 19124 27982
rect 19068 27878 19124 27916
rect 18060 27682 18116 27692
rect 18396 27858 18452 27870
rect 18396 27806 18398 27858
rect 18450 27806 18452 27858
rect 17948 27022 17950 27074
rect 18002 27022 18004 27074
rect 17948 27010 18004 27022
rect 18396 26908 18452 27806
rect 19292 27858 19348 27870
rect 19292 27806 19294 27858
rect 19346 27806 19348 27858
rect 18956 27748 19012 27758
rect 18844 27746 19012 27748
rect 18844 27694 18958 27746
rect 19010 27694 19012 27746
rect 18844 27692 19012 27694
rect 9996 26674 10052 26684
rect 15148 26852 15204 26862
rect 12684 26516 12740 26526
rect 12684 26422 12740 26460
rect 14364 26516 14420 26526
rect 9884 26404 9940 26414
rect 9884 26290 9940 26348
rect 11116 26404 11172 26414
rect 9884 26238 9886 26290
rect 9938 26238 9940 26290
rect 9884 26226 9940 26238
rect 10108 26292 10164 26302
rect 10108 26198 10164 26236
rect 11116 26290 11172 26348
rect 12460 26402 12516 26414
rect 12460 26350 12462 26402
rect 12514 26350 12516 26402
rect 11116 26238 11118 26290
rect 11170 26238 11172 26290
rect 11116 26226 11172 26238
rect 11452 26290 11508 26302
rect 11452 26238 11454 26290
rect 11506 26238 11508 26290
rect 9996 26178 10052 26190
rect 9996 26126 9998 26178
rect 10050 26126 10052 26178
rect 9996 25732 10052 26126
rect 11452 25956 11508 26238
rect 11564 26292 11620 26302
rect 11564 26198 11620 26236
rect 12348 26292 12404 26302
rect 12348 26198 12404 26236
rect 12460 26180 12516 26350
rect 13804 26404 13860 26414
rect 13804 26310 13860 26348
rect 14028 26404 14084 26414
rect 14028 26310 14084 26348
rect 13132 26292 13188 26302
rect 13132 26198 13188 26236
rect 14364 26290 14420 26460
rect 14924 26516 14980 26526
rect 15148 26516 15204 26796
rect 17500 26852 17668 26908
rect 18172 26852 18452 26908
rect 18620 26964 18676 27002
rect 18844 26964 18900 27692
rect 18956 27682 19012 27692
rect 18956 27300 19012 27310
rect 19292 27300 19348 27806
rect 19628 27858 19684 28702
rect 20188 28420 20244 28430
rect 20188 28418 20356 28420
rect 20188 28366 20190 28418
rect 20242 28366 20356 28418
rect 20188 28364 20356 28366
rect 20188 28354 20244 28364
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 20300 27970 20356 28364
rect 20300 27918 20302 27970
rect 20354 27918 20356 27970
rect 20188 27860 20244 27870
rect 19628 27806 19630 27858
rect 19682 27806 19684 27858
rect 19628 27794 19684 27806
rect 20076 27804 20188 27860
rect 19964 27636 20020 27646
rect 19964 27542 20020 27580
rect 18956 27298 19348 27300
rect 18956 27246 18958 27298
rect 19010 27246 19348 27298
rect 18956 27244 19348 27246
rect 18956 27234 19012 27244
rect 20076 27186 20132 27804
rect 20188 27766 20244 27804
rect 20188 27412 20244 27422
rect 20300 27412 20356 27918
rect 20244 27356 20356 27412
rect 20188 27346 20244 27356
rect 20076 27134 20078 27186
rect 20130 27134 20132 27186
rect 20076 27122 20132 27134
rect 18676 26908 18900 26964
rect 19068 27074 19124 27086
rect 19068 27022 19070 27074
rect 19122 27022 19124 27074
rect 18620 26898 18676 26908
rect 15484 26516 15540 26526
rect 14924 26514 15540 26516
rect 14924 26462 14926 26514
rect 14978 26462 15486 26514
rect 15538 26462 15540 26514
rect 14924 26460 15540 26462
rect 14924 26450 14980 26460
rect 15484 26450 15540 26460
rect 14700 26292 14756 26302
rect 16492 26292 16548 26302
rect 14364 26238 14366 26290
rect 14418 26238 14420 26290
rect 14364 26226 14420 26238
rect 14588 26290 14756 26292
rect 14588 26238 14702 26290
rect 14754 26238 14756 26290
rect 14588 26236 14756 26238
rect 12908 26180 12964 26190
rect 12460 26178 12964 26180
rect 12460 26126 12910 26178
rect 12962 26126 12964 26178
rect 12460 26124 12964 26126
rect 11452 25890 11508 25900
rect 12684 25956 12740 25966
rect 9996 25676 10164 25732
rect 9772 25506 9828 25518
rect 9772 25454 9774 25506
rect 9826 25454 9828 25506
rect 9772 25396 9828 25454
rect 9996 25508 10052 25518
rect 9996 25414 10052 25452
rect 9772 25330 9828 25340
rect 9772 24724 9828 24734
rect 9772 24630 9828 24668
rect 10108 23828 10164 25676
rect 11452 25508 11508 25518
rect 11452 25506 11620 25508
rect 11452 25454 11454 25506
rect 11506 25454 11620 25506
rect 11452 25452 11620 25454
rect 11452 25442 11508 25452
rect 10668 25396 10724 25406
rect 10668 25302 10724 25340
rect 10332 25282 10388 25294
rect 10332 25230 10334 25282
rect 10386 25230 10388 25282
rect 10332 25172 10388 25230
rect 10780 25282 10836 25294
rect 10780 25230 10782 25282
rect 10834 25230 10836 25282
rect 10780 25172 10836 25230
rect 11004 25284 11060 25294
rect 11004 25190 11060 25228
rect 10332 25116 10836 25172
rect 10556 24610 10612 24622
rect 10556 24558 10558 24610
rect 10610 24558 10612 24610
rect 10108 23772 10388 23828
rect 10108 23492 10164 23502
rect 10108 23154 10164 23436
rect 10108 23102 10110 23154
rect 10162 23102 10164 23154
rect 10108 22596 10164 23102
rect 10108 22530 10164 22540
rect 10332 21586 10388 23772
rect 10444 23716 10500 23726
rect 10444 23622 10500 23660
rect 10556 23268 10612 24558
rect 10780 24612 10836 25116
rect 10780 24546 10836 24556
rect 11564 25172 11620 25452
rect 11564 24610 11620 25116
rect 11564 24558 11566 24610
rect 11618 24558 11620 24610
rect 10780 24052 10836 24062
rect 10332 21534 10334 21586
rect 10386 21534 10388 21586
rect 10332 21522 10388 21534
rect 10444 23212 10612 23268
rect 10668 23996 10780 24052
rect 10668 23266 10724 23996
rect 10780 23958 10836 23996
rect 11564 24052 11620 24558
rect 11564 23986 11620 23996
rect 11676 25506 11732 25518
rect 11676 25454 11678 25506
rect 11730 25454 11732 25506
rect 10668 23214 10670 23266
rect 10722 23214 10724 23266
rect 10444 21588 10500 23212
rect 10668 23202 10724 23214
rect 11228 23826 11284 23838
rect 11228 23774 11230 23826
rect 11282 23774 11284 23826
rect 11228 23156 11284 23774
rect 11228 23090 11284 23100
rect 11340 23716 11396 23726
rect 11340 23154 11396 23660
rect 11676 23604 11732 25454
rect 12348 25396 12404 25406
rect 12236 25394 12404 25396
rect 12236 25342 12350 25394
rect 12402 25342 12404 25394
rect 12236 25340 12404 25342
rect 12012 25282 12068 25294
rect 12012 25230 12014 25282
rect 12066 25230 12068 25282
rect 11788 24722 11844 24734
rect 11788 24670 11790 24722
rect 11842 24670 11844 24722
rect 11788 23940 11844 24670
rect 11788 23874 11844 23884
rect 11676 23538 11732 23548
rect 11676 23380 11732 23390
rect 11676 23286 11732 23324
rect 11340 23102 11342 23154
rect 11394 23102 11396 23154
rect 10556 23044 10612 23054
rect 10556 23042 10724 23044
rect 10556 22990 10558 23042
rect 10610 22990 10724 23042
rect 10556 22988 10724 22990
rect 10556 22978 10612 22988
rect 10668 22372 10724 22988
rect 10668 22278 10724 22316
rect 10444 21522 10500 21532
rect 10556 22258 10612 22270
rect 10556 22206 10558 22258
rect 10610 22206 10612 22258
rect 9100 20862 9102 20914
rect 9154 20862 9156 20914
rect 9100 20850 9156 20862
rect 9436 21084 9716 21140
rect 10108 21474 10164 21486
rect 10108 21422 10110 21474
rect 10162 21422 10164 21474
rect 9324 20804 9380 20814
rect 9324 20710 9380 20748
rect 8988 20692 9044 20702
rect 8988 20598 9044 20636
rect 8876 20402 8932 20412
rect 9436 20356 9492 21084
rect 10108 21028 10164 21422
rect 9884 20972 10164 21028
rect 10444 21362 10500 21374
rect 10444 21310 10446 21362
rect 10498 21310 10500 21362
rect 9884 20914 9940 20972
rect 9884 20862 9886 20914
rect 9938 20862 9940 20914
rect 9884 20850 9940 20862
rect 9772 20692 9828 20702
rect 9772 20598 9828 20636
rect 10332 20690 10388 20702
rect 10332 20638 10334 20690
rect 10386 20638 10388 20690
rect 9548 20578 9604 20590
rect 9548 20526 9550 20578
rect 9602 20526 9604 20578
rect 9548 20468 9604 20526
rect 9884 20580 9940 20590
rect 9884 20486 9940 20524
rect 10332 20468 10388 20638
rect 9548 20412 9828 20468
rect 9436 20300 9716 20356
rect 8540 19842 8596 19852
rect 9100 20020 9156 20030
rect 8316 19236 8372 19246
rect 8316 19142 8372 19180
rect 8876 19234 8932 19246
rect 8876 19182 8878 19234
rect 8930 19182 8932 19234
rect 8764 19124 8820 19134
rect 8652 17780 8708 17790
rect 8764 17780 8820 19068
rect 8652 17778 8820 17780
rect 8652 17726 8654 17778
rect 8706 17726 8820 17778
rect 8652 17724 8820 17726
rect 8652 17714 8708 17724
rect 8876 17444 8932 19182
rect 8988 19236 9044 19246
rect 8988 17666 9044 19180
rect 9100 18450 9156 19964
rect 9100 18398 9102 18450
rect 9154 18398 9156 18450
rect 9100 18386 9156 18398
rect 9548 20018 9604 20030
rect 9548 19966 9550 20018
rect 9602 19966 9604 20018
rect 9436 18004 9492 18014
rect 9436 17890 9492 17948
rect 9436 17838 9438 17890
rect 9490 17838 9492 17890
rect 9436 17826 9492 17838
rect 9548 17890 9604 19966
rect 9548 17838 9550 17890
rect 9602 17838 9604 17890
rect 9548 17826 9604 17838
rect 8988 17614 8990 17666
rect 9042 17614 9044 17666
rect 8988 17602 9044 17614
rect 9212 17666 9268 17678
rect 9212 17614 9214 17666
rect 9266 17614 9268 17666
rect 9212 17444 9268 17614
rect 8876 17388 9268 17444
rect 8876 16324 8932 17388
rect 8876 16258 8932 16268
rect 8652 16100 8708 16110
rect 8652 16006 8708 16044
rect 8316 15876 8372 15886
rect 8988 15876 9044 15886
rect 7868 15874 8372 15876
rect 7868 15822 8318 15874
rect 8370 15822 8372 15874
rect 7868 15820 8372 15822
rect 8316 15810 8372 15820
rect 8764 15874 9044 15876
rect 8764 15822 8990 15874
rect 9042 15822 9044 15874
rect 8764 15820 9044 15822
rect 7644 15764 7700 15774
rect 7420 15708 7588 15764
rect 6860 15474 6916 15484
rect 7532 15316 7588 15708
rect 7532 15250 7588 15260
rect 6636 15092 6804 15148
rect 5964 13918 5966 13970
rect 6018 13918 6020 13970
rect 5964 13906 6020 13918
rect 6188 14642 6468 14644
rect 6188 14590 6414 14642
rect 6466 14590 6468 14642
rect 6188 14588 6468 14590
rect 6188 13970 6244 14588
rect 6412 14578 6468 14588
rect 6524 14868 6580 14878
rect 6188 13918 6190 13970
rect 6242 13918 6244 13970
rect 6188 13906 6244 13918
rect 6524 13748 6580 14812
rect 6636 14754 6692 15092
rect 6636 14702 6638 14754
rect 6690 14702 6692 14754
rect 6636 14690 6692 14702
rect 6860 14868 6916 14878
rect 6860 14754 6916 14812
rect 6860 14702 6862 14754
rect 6914 14702 6916 14754
rect 6860 14690 6916 14702
rect 7644 14756 7700 15708
rect 7756 15540 7812 15550
rect 8764 15540 8820 15820
rect 8988 15810 9044 15820
rect 7756 15314 7812 15484
rect 7756 15262 7758 15314
rect 7810 15262 7812 15314
rect 7756 15250 7812 15262
rect 8428 15484 8820 15540
rect 7644 14690 7700 14700
rect 8092 14530 8148 14542
rect 8092 14478 8094 14530
rect 8146 14478 8148 14530
rect 7308 14308 7364 14318
rect 7308 14214 7364 14252
rect 8092 14308 8148 14478
rect 8428 14530 8484 15484
rect 9212 15428 9268 15438
rect 8428 14478 8430 14530
rect 8482 14478 8484 14530
rect 8092 13860 8148 14252
rect 8204 14306 8260 14318
rect 8204 14254 8206 14306
rect 8258 14254 8260 14306
rect 8204 14084 8260 14254
rect 8204 14018 8260 14028
rect 8316 13860 8372 13870
rect 8092 13804 8316 13860
rect 8316 13766 8372 13804
rect 6412 13746 6580 13748
rect 6412 13694 6526 13746
rect 6578 13694 6580 13746
rect 6412 13692 6580 13694
rect 6076 13634 6132 13646
rect 6076 13582 6078 13634
rect 6130 13582 6132 13634
rect 5740 12964 5796 12974
rect 5740 12870 5796 12908
rect 6076 12964 6132 13582
rect 6300 13076 6356 13086
rect 6300 12982 6356 13020
rect 6076 12898 6132 12908
rect 6412 12290 6468 13692
rect 6524 13682 6580 13692
rect 7420 13748 7476 13758
rect 6860 13076 6916 13086
rect 6748 12964 6804 12974
rect 6412 12238 6414 12290
rect 6466 12238 6468 12290
rect 6412 12226 6468 12238
rect 6524 12908 6748 12964
rect 5964 12178 6020 12190
rect 5964 12126 5966 12178
rect 6018 12126 6020 12178
rect 5964 12068 6020 12126
rect 6188 12180 6244 12190
rect 6188 12086 6244 12124
rect 5180 11394 5684 11396
rect 5180 11342 5182 11394
rect 5234 11342 5630 11394
rect 5682 11342 5684 11394
rect 5180 11340 5684 11342
rect 5180 11330 5236 11340
rect 5068 11218 5124 11228
rect 5628 10836 5684 11340
rect 5740 11732 5796 11742
rect 5740 11284 5796 11676
rect 5964 11394 6020 12012
rect 6524 11618 6580 12908
rect 6748 12870 6804 12908
rect 6748 12068 6804 12078
rect 6748 11974 6804 12012
rect 6860 11788 6916 13020
rect 7084 12738 7140 12750
rect 7084 12686 7086 12738
rect 7138 12686 7140 12738
rect 7084 12628 7140 12686
rect 7420 12628 7476 13692
rect 8428 13412 8484 14478
rect 8540 15316 8596 15326
rect 8540 13972 8596 15260
rect 8764 15204 8820 15242
rect 8764 15138 8820 15148
rect 9212 15148 9268 15372
rect 9212 15092 9380 15148
rect 8764 14532 8820 14542
rect 8988 14532 9044 14542
rect 8764 14530 9044 14532
rect 8764 14478 8766 14530
rect 8818 14478 8990 14530
rect 9042 14478 9044 14530
rect 8764 14476 9044 14478
rect 8764 14466 8820 14476
rect 8988 14466 9044 14476
rect 8652 14418 8708 14430
rect 8652 14366 8654 14418
rect 8706 14366 8708 14418
rect 8652 14308 8708 14366
rect 9324 14308 9380 15092
rect 9548 14644 9604 14654
rect 8652 14252 9380 14308
rect 8764 13972 8820 13982
rect 8540 13970 9044 13972
rect 8540 13918 8766 13970
rect 8818 13918 9044 13970
rect 8540 13916 9044 13918
rect 8764 13906 8820 13916
rect 8540 13748 8596 13758
rect 8540 13654 8596 13692
rect 8764 13748 8820 13758
rect 8764 13634 8820 13692
rect 8764 13582 8766 13634
rect 8818 13582 8820 13634
rect 8764 13570 8820 13582
rect 8876 13746 8932 13758
rect 8876 13694 8878 13746
rect 8930 13694 8932 13746
rect 8876 13412 8932 13694
rect 8428 13356 8932 13412
rect 7084 12572 7476 12628
rect 6972 12180 7028 12190
rect 6972 12086 7028 12124
rect 6524 11566 6526 11618
rect 6578 11566 6580 11618
rect 5964 11342 5966 11394
rect 6018 11342 6020 11394
rect 5964 11330 6020 11342
rect 6300 11396 6356 11406
rect 6300 11302 6356 11340
rect 5740 11190 5796 11228
rect 5740 10836 5796 10846
rect 6076 10836 6132 10846
rect 5628 10834 6076 10836
rect 5628 10782 5742 10834
rect 5794 10782 6076 10834
rect 5628 10780 6076 10782
rect 5740 10770 5796 10780
rect 4844 10658 4900 10668
rect 6076 10722 6132 10780
rect 6076 10670 6078 10722
rect 6130 10670 6132 10722
rect 6076 10658 6132 10670
rect 6188 10724 6244 10734
rect 1708 10610 1764 10622
rect 1708 10558 1710 10610
rect 1762 10558 1764 10610
rect 1708 10164 1764 10558
rect 1708 10098 1764 10108
rect 2492 10498 2548 10510
rect 2492 10446 2494 10498
rect 2546 10446 2548 10498
rect 2492 10164 2548 10446
rect 6188 10388 6244 10668
rect 5964 10332 6244 10388
rect 6412 10610 6468 10622
rect 6412 10558 6414 10610
rect 6466 10558 6468 10610
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 2492 10098 2548 10108
rect 5628 9268 5684 9278
rect 5628 9174 5684 9212
rect 2044 9156 2100 9166
rect 2044 9062 2100 9100
rect 1708 9042 1764 9054
rect 1708 8990 1710 9042
rect 1762 8990 1764 9042
rect 1708 8820 1764 8990
rect 5964 9042 6020 10332
rect 6412 9826 6468 10558
rect 6524 10610 6580 11566
rect 6524 10558 6526 10610
rect 6578 10558 6580 10610
rect 6524 10546 6580 10558
rect 6636 11732 6916 11788
rect 7308 11954 7364 11966
rect 7308 11902 7310 11954
rect 7362 11902 7364 11954
rect 6636 10164 6692 11732
rect 6860 11508 6916 11518
rect 6860 11414 6916 11452
rect 6972 11396 7028 11406
rect 6860 10834 6916 10846
rect 6860 10782 6862 10834
rect 6914 10782 6916 10834
rect 6636 10108 6804 10164
rect 6412 9774 6414 9826
rect 6466 9774 6468 9826
rect 6300 9268 6356 9278
rect 5964 8990 5966 9042
rect 6018 8990 6020 9042
rect 5964 8978 6020 8990
rect 6188 9154 6244 9166
rect 6188 9102 6190 9154
rect 6242 9102 6244 9154
rect 1708 8754 1764 8764
rect 2492 8930 2548 8942
rect 2492 8878 2494 8930
rect 2546 8878 2548 8930
rect 2492 8820 2548 8878
rect 2492 8754 2548 8764
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 6188 8484 6244 9102
rect 6300 8932 6356 9212
rect 6412 9156 6468 9774
rect 6636 9938 6692 9950
rect 6636 9886 6638 9938
rect 6690 9886 6692 9938
rect 6524 9156 6580 9166
rect 6412 9154 6580 9156
rect 6412 9102 6526 9154
rect 6578 9102 6580 9154
rect 6412 9100 6580 9102
rect 6524 9090 6580 9100
rect 6300 8876 6580 8932
rect 6188 8418 6244 8428
rect 6524 8370 6580 8876
rect 6524 8318 6526 8370
rect 6578 8318 6580 8370
rect 6524 8036 6580 8318
rect 6636 8260 6692 9886
rect 6748 9268 6804 10108
rect 6860 9380 6916 10782
rect 6972 10722 7028 11340
rect 7308 11396 7364 11902
rect 7308 11302 7364 11340
rect 7420 11394 7476 12572
rect 8764 12516 8820 13356
rect 8988 12962 9044 13916
rect 8988 12910 8990 12962
rect 9042 12910 9044 12962
rect 8988 12898 9044 12910
rect 9324 12852 9380 14252
rect 9436 14642 9604 14644
rect 9436 14590 9550 14642
rect 9602 14590 9604 14642
rect 9436 14588 9604 14590
rect 9436 13748 9492 14588
rect 9548 14578 9604 14588
rect 9660 14532 9716 20300
rect 9772 19908 9828 20412
rect 10332 20402 10388 20412
rect 10444 20132 10500 21310
rect 10556 21364 10612 22206
rect 11228 21812 11284 21822
rect 11228 21718 11284 21756
rect 11228 21588 11284 21598
rect 11340 21588 11396 23102
rect 11900 23156 11956 23166
rect 11284 21532 11396 21588
rect 11452 22372 11508 22382
rect 10556 21308 10948 21364
rect 10892 20802 10948 21308
rect 10892 20750 10894 20802
rect 10946 20750 10948 20802
rect 10892 20738 10948 20750
rect 10668 20692 10724 20702
rect 10668 20598 10724 20636
rect 11116 20692 11172 20702
rect 11116 20598 11172 20636
rect 11228 20690 11284 21532
rect 11228 20638 11230 20690
rect 11282 20638 11284 20690
rect 11228 20468 11284 20638
rect 10444 20038 10500 20076
rect 11116 20412 11284 20468
rect 10332 20020 10388 20030
rect 10332 19926 10388 19964
rect 9772 19842 9828 19852
rect 9996 19906 10052 19918
rect 9996 19854 9998 19906
rect 10050 19854 10052 19906
rect 9660 14466 9716 14476
rect 9996 17780 10052 19854
rect 10556 19346 10612 19358
rect 10556 19294 10558 19346
rect 10610 19294 10612 19346
rect 10108 19234 10164 19246
rect 10108 19182 10110 19234
rect 10162 19182 10164 19234
rect 10108 18004 10164 19182
rect 10108 17938 10164 17948
rect 10332 18338 10388 18350
rect 10332 18286 10334 18338
rect 10386 18286 10388 18338
rect 10332 17780 10388 18286
rect 9996 17724 10388 17780
rect 10556 17780 10612 19294
rect 10892 18564 10948 18574
rect 10556 17778 10836 17780
rect 10556 17726 10558 17778
rect 10610 17726 10836 17778
rect 10556 17724 10836 17726
rect 9996 14530 10052 17724
rect 10556 17714 10612 17724
rect 10780 17108 10836 17724
rect 10892 17554 10948 18508
rect 10892 17502 10894 17554
rect 10946 17502 10948 17554
rect 10892 17490 10948 17502
rect 10780 17052 11060 17108
rect 10780 16100 10836 16110
rect 10220 15314 10276 15326
rect 10220 15262 10222 15314
rect 10274 15262 10276 15314
rect 10220 15148 10276 15262
rect 10556 15316 10612 15326
rect 10780 15316 10836 16044
rect 11004 16098 11060 17052
rect 11004 16046 11006 16098
rect 11058 16046 11060 16098
rect 11004 15426 11060 16046
rect 11116 15764 11172 20412
rect 11340 20132 11396 20142
rect 11340 20018 11396 20076
rect 11340 19966 11342 20018
rect 11394 19966 11396 20018
rect 11340 19954 11396 19966
rect 11452 19796 11508 22316
rect 11676 22370 11732 22382
rect 11676 22318 11678 22370
rect 11730 22318 11732 22370
rect 11564 21812 11620 21822
rect 11564 21718 11620 21756
rect 11676 20916 11732 22318
rect 11788 21812 11844 21822
rect 11900 21812 11956 23100
rect 12012 22820 12068 25230
rect 12236 23938 12292 25340
rect 12348 25330 12404 25340
rect 12460 25282 12516 25294
rect 12460 25230 12462 25282
rect 12514 25230 12516 25282
rect 12460 24164 12516 25230
rect 12572 25282 12628 25294
rect 12572 25230 12574 25282
rect 12626 25230 12628 25282
rect 12572 25172 12628 25230
rect 12572 25106 12628 25116
rect 12684 24722 12740 25900
rect 12908 25172 12964 26124
rect 13468 26066 13524 26078
rect 13468 26014 13470 26066
rect 13522 26014 13524 26066
rect 13468 25844 13524 26014
rect 14140 26068 14196 26078
rect 14140 25974 14196 26012
rect 14588 25844 14644 26236
rect 14700 26226 14756 26236
rect 15596 26290 16548 26292
rect 15596 26238 16494 26290
rect 16546 26238 16548 26290
rect 15596 26236 16548 26238
rect 14812 26068 14868 26078
rect 14868 26012 14980 26068
rect 14812 26002 14868 26012
rect 13468 25788 14644 25844
rect 12908 25106 12964 25116
rect 13916 25618 13972 25630
rect 13916 25566 13918 25618
rect 13970 25566 13972 25618
rect 12684 24670 12686 24722
rect 12738 24670 12740 24722
rect 12684 24658 12740 24670
rect 13580 25060 13636 25070
rect 13580 24722 13636 25004
rect 13580 24670 13582 24722
rect 13634 24670 13636 24722
rect 13580 24658 13636 24670
rect 13468 24612 13524 24622
rect 13468 24518 13524 24556
rect 12236 23886 12238 23938
rect 12290 23886 12292 23938
rect 12124 23604 12180 23614
rect 12236 23604 12292 23886
rect 12180 23548 12292 23604
rect 12348 24108 12516 24164
rect 12124 23538 12180 23548
rect 12348 23042 12404 24108
rect 12908 24052 12964 24062
rect 13916 24052 13972 25566
rect 12908 23958 12964 23996
rect 13804 23996 13916 24052
rect 13468 23940 13524 23950
rect 12572 23380 12628 23390
rect 12348 22990 12350 23042
rect 12402 22990 12404 23042
rect 12348 22978 12404 22990
rect 12460 23154 12516 23166
rect 12460 23102 12462 23154
rect 12514 23102 12516 23154
rect 12460 22820 12516 23102
rect 12012 22764 12516 22820
rect 12236 22484 12292 22494
rect 11788 21810 11956 21812
rect 11788 21758 11790 21810
rect 11842 21758 11956 21810
rect 11788 21756 11956 21758
rect 12012 21812 12068 21822
rect 11788 21746 11844 21756
rect 12012 21718 12068 21756
rect 12124 21588 12180 21598
rect 12124 21494 12180 21532
rect 12236 21364 12292 22428
rect 12572 21700 12628 23324
rect 13468 23268 13524 23884
rect 13692 23938 13748 23950
rect 13692 23886 13694 23938
rect 13746 23886 13748 23938
rect 13692 23828 13748 23886
rect 13692 23762 13748 23772
rect 13468 23266 13748 23268
rect 13468 23214 13470 23266
rect 13522 23214 13748 23266
rect 13468 23212 13748 23214
rect 13468 23202 13524 23212
rect 12684 23156 12740 23166
rect 12684 23062 12740 23100
rect 13692 22820 13748 23212
rect 13804 23154 13860 23996
rect 13916 23986 13972 23996
rect 14028 25506 14084 25788
rect 14028 25454 14030 25506
rect 14082 25454 14084 25506
rect 13916 23716 13972 23726
rect 13916 23622 13972 23660
rect 13804 23102 13806 23154
rect 13858 23102 13860 23154
rect 13804 23090 13860 23102
rect 14028 23042 14084 25454
rect 14700 25508 14756 25518
rect 14924 25508 14980 26012
rect 15036 26066 15092 26078
rect 15036 26014 15038 26066
rect 15090 26014 15092 26066
rect 15036 25956 15092 26014
rect 15036 25900 15316 25956
rect 15036 25508 15092 25518
rect 14924 25506 15092 25508
rect 14924 25454 15038 25506
rect 15090 25454 15092 25506
rect 14924 25452 15092 25454
rect 14700 25414 14756 25452
rect 15036 25442 15092 25452
rect 15148 25284 15204 25294
rect 15148 25190 15204 25228
rect 14140 25172 14196 25182
rect 14140 23938 14196 25116
rect 15260 24836 15316 25900
rect 15372 25284 15428 25294
rect 15372 25190 15428 25228
rect 15596 24948 15652 26236
rect 16492 26226 16548 26236
rect 16604 26066 16660 26078
rect 16604 26014 16606 26066
rect 16658 26014 16660 26066
rect 16604 25508 16660 26014
rect 16604 25506 16772 25508
rect 16604 25454 16606 25506
rect 16658 25454 16772 25506
rect 16604 25452 16772 25454
rect 16604 25442 16660 25452
rect 16268 25394 16324 25406
rect 16268 25342 16270 25394
rect 16322 25342 16324 25394
rect 15484 24892 15652 24948
rect 15708 25284 15764 25294
rect 15372 24836 15428 24846
rect 15260 24780 15372 24836
rect 15372 24770 15428 24780
rect 15372 24610 15428 24622
rect 15372 24558 15374 24610
rect 15426 24558 15428 24610
rect 14140 23886 14142 23938
rect 14194 23886 14196 23938
rect 14140 23874 14196 23886
rect 14924 23940 14980 23950
rect 14364 23828 14420 23838
rect 14364 23734 14420 23772
rect 14476 23826 14532 23838
rect 14476 23774 14478 23826
rect 14530 23774 14532 23826
rect 14476 23380 14532 23774
rect 14476 23314 14532 23324
rect 14924 23266 14980 23884
rect 14924 23214 14926 23266
rect 14978 23214 14980 23266
rect 14924 23202 14980 23214
rect 15372 23492 15428 24558
rect 14028 22990 14030 23042
rect 14082 22990 14084 23042
rect 14028 22978 14084 22990
rect 14812 23156 14868 23166
rect 13692 22764 14084 22820
rect 12908 22596 12964 22606
rect 12908 22502 12964 22540
rect 13804 22596 13860 22606
rect 13804 22502 13860 22540
rect 14028 22482 14084 22764
rect 14812 22596 14868 23100
rect 15036 23156 15092 23166
rect 15372 23156 15428 23436
rect 15484 23826 15540 24892
rect 15596 24722 15652 24734
rect 15596 24670 15598 24722
rect 15650 24670 15652 24722
rect 15596 23940 15652 24670
rect 15596 23846 15652 23884
rect 15484 23774 15486 23826
rect 15538 23774 15540 23826
rect 15484 23378 15540 23774
rect 15708 23716 15764 25228
rect 16268 24836 16324 25342
rect 16716 24946 16772 25452
rect 16716 24894 16718 24946
rect 16770 24894 16772 24946
rect 16716 24882 16772 24894
rect 16604 24836 16660 24846
rect 16268 24834 16660 24836
rect 16268 24782 16270 24834
rect 16322 24782 16606 24834
rect 16658 24782 16660 24834
rect 16268 24780 16660 24782
rect 16268 24770 16324 24780
rect 16604 24770 16660 24780
rect 16940 24724 16996 24734
rect 17276 24724 17332 24734
rect 16940 24722 17332 24724
rect 16940 24670 16942 24722
rect 16994 24670 17278 24722
rect 17330 24670 17332 24722
rect 16940 24668 17332 24670
rect 16940 24658 16996 24668
rect 17276 24658 17332 24668
rect 17164 24052 17220 24062
rect 17164 23958 17220 23996
rect 15484 23326 15486 23378
rect 15538 23326 15540 23378
rect 15484 23314 15540 23326
rect 15596 23660 15764 23716
rect 16492 23938 16548 23950
rect 16492 23886 16494 23938
rect 16546 23886 16548 23938
rect 15092 23100 15428 23156
rect 15036 23090 15092 23100
rect 14812 22530 14868 22540
rect 14924 22930 14980 22942
rect 14924 22878 14926 22930
rect 14978 22878 14980 22930
rect 14028 22430 14030 22482
rect 14082 22430 14084 22482
rect 14028 22418 14084 22430
rect 13468 22148 13524 22158
rect 12236 21298 12292 21308
rect 12460 21644 12628 21700
rect 13356 22146 13524 22148
rect 13356 22094 13470 22146
rect 13522 22094 13524 22146
rect 13356 22092 13524 22094
rect 11564 20860 11732 20916
rect 11564 20020 11620 20860
rect 12460 20804 12516 21644
rect 12572 21476 12628 21486
rect 12572 21382 12628 21420
rect 11788 20748 12516 20804
rect 11676 20692 11732 20702
rect 11676 20598 11732 20636
rect 11564 19906 11620 19964
rect 11564 19854 11566 19906
rect 11618 19854 11620 19906
rect 11564 19842 11620 19854
rect 11340 19740 11508 19796
rect 11340 19346 11396 19740
rect 11340 19294 11342 19346
rect 11394 19294 11396 19346
rect 11340 19282 11396 19294
rect 11228 19234 11284 19246
rect 11228 19182 11230 19234
rect 11282 19182 11284 19234
rect 11228 19124 11284 19182
rect 11228 19058 11284 19068
rect 11788 17106 11844 20748
rect 11900 20580 11956 20590
rect 11900 18676 11956 20524
rect 12012 20580 12068 20590
rect 12012 20578 12180 20580
rect 12012 20526 12014 20578
rect 12066 20526 12180 20578
rect 12012 20524 12180 20526
rect 12012 20514 12068 20524
rect 11900 18610 11956 18620
rect 12012 19906 12068 19918
rect 12012 19854 12014 19906
rect 12066 19854 12068 19906
rect 11788 17054 11790 17106
rect 11842 17054 11844 17106
rect 11676 15988 11732 15998
rect 11676 15894 11732 15932
rect 11116 15698 11172 15708
rect 11004 15374 11006 15426
rect 11058 15374 11060 15426
rect 11004 15362 11060 15374
rect 11676 15428 11732 15438
rect 11676 15334 11732 15372
rect 11788 15426 11844 17054
rect 11900 18450 11956 18462
rect 11900 18398 11902 18450
rect 11954 18398 11956 18450
rect 11900 17666 11956 18398
rect 12012 18452 12068 19854
rect 12124 18788 12180 20524
rect 12460 20356 12516 20748
rect 12796 20692 12852 20702
rect 12796 20598 12852 20636
rect 12908 20692 12964 20702
rect 13356 20692 13412 22092
rect 13468 22082 13524 22092
rect 14476 21698 14532 21710
rect 14476 21646 14478 21698
rect 14530 21646 14532 21698
rect 13580 21476 13636 21486
rect 13580 20914 13636 21420
rect 13580 20862 13582 20914
rect 13634 20862 13636 20914
rect 13580 20850 13636 20862
rect 14028 21474 14084 21486
rect 14028 21422 14030 21474
rect 14082 21422 14084 21474
rect 12908 20690 13412 20692
rect 12908 20638 12910 20690
rect 12962 20638 13412 20690
rect 12908 20636 13412 20638
rect 14028 20692 14084 21422
rect 12684 20578 12740 20590
rect 12684 20526 12686 20578
rect 12738 20526 12740 20578
rect 12460 20300 12628 20356
rect 12460 20130 12516 20142
rect 12460 20078 12462 20130
rect 12514 20078 12516 20130
rect 12124 18722 12180 18732
rect 12236 20018 12292 20030
rect 12236 19966 12238 20018
rect 12290 19966 12292 20018
rect 12236 18564 12292 19966
rect 12236 18498 12292 18508
rect 12012 18386 12068 18396
rect 11900 17614 11902 17666
rect 11954 17614 11956 17666
rect 11900 16100 11956 17614
rect 11900 16034 11956 16044
rect 12124 17892 12180 17902
rect 12124 16994 12180 17836
rect 12460 17444 12516 20078
rect 12572 20130 12628 20300
rect 12572 20078 12574 20130
rect 12626 20078 12628 20130
rect 12572 20066 12628 20078
rect 12684 20132 12740 20526
rect 12684 20066 12740 20076
rect 12908 20018 12964 20636
rect 13132 20132 13188 20142
rect 13132 20038 13188 20076
rect 12908 19966 12910 20018
rect 12962 19966 12964 20018
rect 12908 19236 12964 19966
rect 13468 20018 13524 20030
rect 13468 19966 13470 20018
rect 13522 19966 13524 20018
rect 12908 19170 12964 19180
rect 13020 19906 13076 19918
rect 13020 19854 13022 19906
rect 13074 19854 13076 19906
rect 12572 18228 12628 18238
rect 12572 17778 12628 18172
rect 12572 17726 12574 17778
rect 12626 17726 12628 17778
rect 12572 17714 12628 17726
rect 12460 17106 12516 17388
rect 12460 17054 12462 17106
rect 12514 17054 12516 17106
rect 12460 17042 12516 17054
rect 12124 16942 12126 16994
rect 12178 16942 12180 16994
rect 11788 15374 11790 15426
rect 11842 15374 11844 15426
rect 11788 15362 11844 15374
rect 10556 15314 10836 15316
rect 10556 15262 10558 15314
rect 10610 15262 10836 15314
rect 10556 15260 10836 15262
rect 11452 15314 11508 15326
rect 11452 15262 11454 15314
rect 11506 15262 11508 15314
rect 10556 15204 10612 15260
rect 10220 15092 10500 15148
rect 10556 15138 10612 15148
rect 11004 15202 11060 15214
rect 11004 15150 11006 15202
rect 11058 15150 11060 15202
rect 9996 14478 9998 14530
rect 10050 14478 10052 14530
rect 9996 14466 10052 14478
rect 10332 14420 10388 14430
rect 10332 14326 10388 14364
rect 10444 13972 10500 15092
rect 10780 14642 10836 14654
rect 10780 14590 10782 14642
rect 10834 14590 10836 14642
rect 10780 14420 10836 14590
rect 10836 14364 10948 14420
rect 10780 14354 10836 14364
rect 10556 13972 10612 13982
rect 10444 13970 10612 13972
rect 10444 13918 10558 13970
rect 10610 13918 10612 13970
rect 10444 13916 10612 13918
rect 10556 13906 10612 13916
rect 10108 13860 10164 13870
rect 9436 13682 9492 13692
rect 9772 13746 9828 13758
rect 9772 13694 9774 13746
rect 9826 13694 9828 13746
rect 9548 13634 9604 13646
rect 9548 13582 9550 13634
rect 9602 13582 9604 13634
rect 9548 12852 9604 13582
rect 9380 12796 9604 12852
rect 9772 12964 9828 13694
rect 9884 13746 9940 13758
rect 9884 13694 9886 13746
rect 9938 13694 9940 13746
rect 9884 13636 9940 13694
rect 10108 13746 10164 13804
rect 10108 13694 10110 13746
rect 10162 13694 10164 13746
rect 10108 13682 10164 13694
rect 9884 13570 9940 13580
rect 9772 12908 10052 12964
rect 9324 12758 9380 12796
rect 9660 12738 9716 12750
rect 9660 12686 9662 12738
rect 9714 12686 9716 12738
rect 9660 12516 9716 12686
rect 8764 12460 9716 12516
rect 8428 12290 8484 12302
rect 8428 12238 8430 12290
rect 8482 12238 8484 12290
rect 8428 11732 8484 12238
rect 8764 12178 8820 12460
rect 9772 12404 9828 12908
rect 9996 12850 10052 12908
rect 9996 12798 9998 12850
rect 10050 12798 10052 12850
rect 9996 12786 10052 12798
rect 9324 12348 9828 12404
rect 8764 12126 8766 12178
rect 8818 12126 8820 12178
rect 8764 12114 8820 12126
rect 8988 12180 9044 12190
rect 8428 11666 8484 11676
rect 8988 12066 9044 12124
rect 8988 12014 8990 12066
rect 9042 12014 9044 12066
rect 8652 11508 8708 11518
rect 8428 11452 8652 11508
rect 7420 11342 7422 11394
rect 7474 11342 7476 11394
rect 7420 11330 7476 11342
rect 7532 11396 7588 11406
rect 7532 10836 7588 11340
rect 7980 11284 8036 11294
rect 7980 11190 8036 11228
rect 7196 10780 7588 10836
rect 7644 10836 7700 10846
rect 7700 10780 7812 10836
rect 7196 10724 7252 10780
rect 7644 10742 7700 10780
rect 6972 10670 6974 10722
rect 7026 10670 7028 10722
rect 6972 10658 7028 10670
rect 7084 10722 7252 10724
rect 7084 10670 7198 10722
rect 7250 10670 7252 10722
rect 7084 10668 7252 10670
rect 7084 9938 7140 10668
rect 7196 10658 7252 10668
rect 7084 9886 7086 9938
rect 7138 9886 7140 9938
rect 7084 9874 7140 9886
rect 7644 9714 7700 9726
rect 7644 9662 7646 9714
rect 7698 9662 7700 9714
rect 6860 9324 7476 9380
rect 6748 9154 6804 9212
rect 7420 9266 7476 9324
rect 7420 9214 7422 9266
rect 7474 9214 7476 9266
rect 6748 9102 6750 9154
rect 6802 9102 6804 9154
rect 6748 9090 6804 9102
rect 7084 9156 7140 9166
rect 6972 8930 7028 8942
rect 6972 8878 6974 8930
rect 7026 8878 7028 8930
rect 6748 8260 6804 8270
rect 6636 8258 6804 8260
rect 6636 8206 6750 8258
rect 6802 8206 6804 8258
rect 6636 8204 6804 8206
rect 6748 8194 6804 8204
rect 6972 8260 7028 8878
rect 6972 8194 7028 8204
rect 7084 8258 7140 9100
rect 7420 8482 7476 9214
rect 7644 9156 7700 9662
rect 7756 9714 7812 10780
rect 8428 9938 8484 11452
rect 8652 11414 8708 11452
rect 8428 9886 8430 9938
rect 8482 9886 8484 9938
rect 8428 9874 8484 9886
rect 8988 11282 9044 12014
rect 8988 11230 8990 11282
rect 9042 11230 9044 11282
rect 7756 9662 7758 9714
rect 7810 9662 7812 9714
rect 7756 9650 7812 9662
rect 8876 9716 8932 9726
rect 8988 9716 9044 11230
rect 8876 9714 9044 9716
rect 8876 9662 8878 9714
rect 8930 9662 9044 9714
rect 8876 9660 9044 9662
rect 8876 9650 8932 9660
rect 7980 9604 8036 9614
rect 7980 9602 8372 9604
rect 7980 9550 7982 9602
rect 8034 9550 8372 9602
rect 7980 9548 8372 9550
rect 7980 9538 8036 9548
rect 7644 9090 7700 9100
rect 7980 9268 8036 9278
rect 7980 9042 8036 9212
rect 7980 8990 7982 9042
rect 8034 8990 8036 9042
rect 7980 8978 8036 8990
rect 7420 8430 7422 8482
rect 7474 8430 7476 8482
rect 7420 8418 7476 8430
rect 7756 8372 7812 8382
rect 8204 8372 8260 8382
rect 7756 8370 8260 8372
rect 7756 8318 7758 8370
rect 7810 8318 8206 8370
rect 8258 8318 8260 8370
rect 7756 8316 8260 8318
rect 7756 8306 7812 8316
rect 8204 8306 8260 8316
rect 7084 8206 7086 8258
rect 7138 8206 7140 8258
rect 7084 8194 7140 8206
rect 7644 8260 7700 8270
rect 7644 8146 7700 8204
rect 7644 8094 7646 8146
rect 7698 8094 7700 8146
rect 7644 8082 7700 8094
rect 8316 8148 8372 9548
rect 9100 9268 9156 9278
rect 8652 9156 8708 9166
rect 8652 9062 8708 9100
rect 8988 9154 9044 9166
rect 8988 9102 8990 9154
rect 9042 9102 9044 9154
rect 8876 9044 8932 9054
rect 6972 8036 7028 8046
rect 6524 8034 7028 8036
rect 6524 7982 6974 8034
rect 7026 7982 7028 8034
rect 6524 7980 7028 7982
rect 6972 7970 7028 7980
rect 8316 7476 8372 8092
rect 8652 8372 8708 8382
rect 8652 8146 8708 8316
rect 8652 8094 8654 8146
rect 8706 8094 8708 8146
rect 8652 8082 8708 8094
rect 8764 8260 8820 8270
rect 8764 7700 8820 8204
rect 8764 7606 8820 7644
rect 8876 7698 8932 8988
rect 8988 7924 9044 9102
rect 8988 7858 9044 7868
rect 8876 7646 8878 7698
rect 8930 7646 8932 7698
rect 8876 7634 8932 7646
rect 8988 7700 9044 7710
rect 9100 7700 9156 9212
rect 8988 7698 9156 7700
rect 8988 7646 8990 7698
rect 9042 7646 9156 7698
rect 8988 7644 9156 7646
rect 8988 7634 9044 7644
rect 8428 7476 8484 7486
rect 8316 7474 8484 7476
rect 8316 7422 8430 7474
rect 8482 7422 8484 7474
rect 8316 7420 8484 7422
rect 8428 7410 8484 7420
rect 9100 7252 9156 7644
rect 9100 7186 9156 7196
rect 9212 8484 9268 8494
rect 9212 8036 9268 8428
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 9212 6692 9268 7980
rect 9324 7588 9380 12348
rect 9772 12178 9828 12190
rect 9772 12126 9774 12178
rect 9826 12126 9828 12178
rect 9660 12068 9716 12078
rect 9548 12012 9660 12068
rect 9548 10388 9604 12012
rect 9660 12002 9716 12012
rect 9772 11284 9828 12126
rect 9660 10612 9716 10622
rect 9772 10612 9828 11228
rect 9660 10610 9828 10612
rect 9660 10558 9662 10610
rect 9714 10558 9828 10610
rect 9660 10556 9828 10558
rect 9996 12180 10052 12190
rect 9660 10546 9716 10556
rect 9772 10388 9828 10398
rect 9548 10386 9828 10388
rect 9548 10334 9774 10386
rect 9826 10334 9828 10386
rect 9548 10332 9828 10334
rect 9548 9268 9604 10332
rect 9772 10322 9828 10332
rect 9996 10386 10052 12124
rect 10220 12068 10276 12078
rect 10220 11974 10276 12012
rect 10892 11956 10948 14364
rect 11004 13636 11060 15150
rect 11452 15148 11508 15262
rect 11228 15092 11508 15148
rect 12124 15148 12180 16942
rect 12796 16994 12852 17006
rect 12796 16942 12798 16994
rect 12850 16942 12852 16994
rect 12796 16100 12852 16942
rect 13020 16882 13076 19854
rect 13468 19124 13524 19966
rect 14028 19906 14084 20636
rect 14028 19854 14030 19906
rect 14082 19854 14084 19906
rect 14028 19842 14084 19854
rect 14252 20132 14308 20142
rect 13244 19068 13468 19124
rect 13132 18564 13188 18574
rect 13244 18564 13300 19068
rect 13468 19030 13524 19068
rect 14252 19346 14308 20076
rect 14476 20130 14532 21646
rect 14924 20188 14980 22878
rect 15484 21586 15540 21598
rect 15484 21534 15486 21586
rect 15538 21534 15540 21586
rect 15372 21026 15428 21038
rect 15372 20974 15374 21026
rect 15426 20974 15428 21026
rect 15372 20914 15428 20974
rect 15372 20862 15374 20914
rect 15426 20862 15428 20914
rect 15372 20850 15428 20862
rect 14924 20132 15204 20188
rect 14476 20078 14478 20130
rect 14530 20078 14532 20130
rect 14476 19460 14532 20078
rect 14476 19394 14532 19404
rect 14252 19294 14254 19346
rect 14306 19294 14308 19346
rect 13132 18562 13300 18564
rect 13132 18510 13134 18562
rect 13186 18510 13300 18562
rect 13132 18508 13300 18510
rect 13468 18788 13524 18798
rect 13132 18498 13188 18508
rect 13356 18452 13412 18462
rect 13356 17668 13412 18396
rect 13468 18452 13524 18732
rect 14252 18674 14308 19294
rect 14476 19236 14532 19246
rect 14476 19142 14532 19180
rect 15036 19124 15092 19134
rect 15036 19030 15092 19068
rect 14252 18622 14254 18674
rect 14306 18622 14308 18674
rect 14252 18610 14308 18622
rect 15148 18562 15204 20132
rect 15372 20018 15428 20030
rect 15372 19966 15374 20018
rect 15426 19966 15428 20018
rect 15260 19572 15316 19582
rect 15260 19348 15316 19516
rect 15260 19282 15316 19292
rect 15148 18510 15150 18562
rect 15202 18510 15204 18562
rect 15148 18498 15204 18510
rect 13468 18450 13636 18452
rect 13468 18398 13470 18450
rect 13522 18398 13636 18450
rect 13468 18396 13636 18398
rect 13468 18386 13524 18396
rect 13468 17668 13524 17678
rect 13356 17666 13524 17668
rect 13356 17614 13470 17666
rect 13522 17614 13524 17666
rect 13356 17612 13524 17614
rect 13468 17602 13524 17612
rect 13020 16830 13022 16882
rect 13074 16830 13076 16882
rect 13020 16818 13076 16830
rect 13132 17444 13188 17454
rect 13580 17444 13636 18396
rect 13692 18450 13748 18462
rect 13692 18398 13694 18450
rect 13746 18398 13748 18450
rect 13692 17892 13748 18398
rect 13804 18452 13860 18462
rect 13804 18358 13860 18396
rect 14588 18450 14644 18462
rect 14812 18452 14868 18462
rect 14588 18398 14590 18450
rect 14642 18398 14644 18450
rect 14588 18228 14644 18398
rect 14588 18162 14644 18172
rect 14700 18450 14868 18452
rect 14700 18398 14814 18450
rect 14866 18398 14868 18450
rect 14700 18396 14868 18398
rect 14700 18004 14756 18396
rect 14812 18386 14868 18396
rect 15372 18452 15428 19966
rect 15484 19124 15540 21534
rect 15484 19058 15540 19068
rect 15372 18386 15428 18396
rect 15036 18340 15092 18350
rect 15036 18246 15092 18284
rect 15484 18340 15540 18350
rect 13692 17826 13748 17836
rect 14028 17948 14756 18004
rect 15148 18228 15204 18238
rect 14028 17890 14084 17948
rect 14028 17838 14030 17890
rect 14082 17838 14084 17890
rect 14028 17826 14084 17838
rect 14476 17780 14532 17790
rect 13692 17668 13748 17678
rect 13692 17666 14084 17668
rect 13692 17614 13694 17666
rect 13746 17614 14084 17666
rect 13692 17612 14084 17614
rect 13692 17602 13748 17612
rect 14028 17556 14084 17612
rect 14476 17666 14532 17724
rect 14476 17614 14478 17666
rect 14530 17614 14532 17666
rect 14476 17602 14532 17614
rect 15148 17778 15204 18172
rect 15148 17726 15150 17778
rect 15202 17726 15204 17778
rect 14252 17556 14308 17566
rect 14028 17554 14308 17556
rect 14028 17502 14254 17554
rect 14306 17502 14308 17554
rect 14028 17500 14308 17502
rect 13916 17444 13972 17454
rect 13580 17442 13972 17444
rect 13580 17390 13918 17442
rect 13970 17390 13972 17442
rect 13580 17388 13972 17390
rect 12796 16034 12852 16044
rect 12908 15316 12964 15326
rect 13132 15316 13188 17388
rect 13916 17378 13972 17388
rect 13356 16882 13412 16894
rect 13580 16884 13636 16894
rect 13356 16830 13358 16882
rect 13410 16830 13412 16882
rect 13244 16772 13300 16782
rect 13244 16678 13300 16716
rect 13356 16100 13412 16830
rect 13244 16044 13412 16100
rect 13468 16882 13636 16884
rect 13468 16830 13582 16882
rect 13634 16830 13636 16882
rect 13468 16828 13636 16830
rect 13244 15538 13300 16044
rect 13244 15486 13246 15538
rect 13298 15486 13300 15538
rect 13244 15474 13300 15486
rect 13356 15426 13412 15438
rect 13356 15374 13358 15426
rect 13410 15374 13412 15426
rect 13356 15316 13412 15374
rect 13132 15260 13412 15316
rect 13468 15316 13524 16828
rect 13580 16818 13636 16828
rect 14028 16212 14084 17500
rect 14252 17490 14308 17500
rect 14364 17444 14420 17454
rect 14364 17106 14420 17388
rect 14364 17054 14366 17106
rect 14418 17054 14420 17106
rect 13916 16156 14084 16212
rect 14140 16994 14196 17006
rect 14140 16942 14142 16994
rect 14194 16942 14196 16994
rect 14140 16884 14196 16942
rect 13692 16100 13748 16110
rect 13692 16006 13748 16044
rect 13916 16098 13972 16156
rect 13916 16046 13918 16098
rect 13970 16046 13972 16098
rect 13916 15652 13972 16046
rect 13692 15596 13972 15652
rect 14028 15988 14084 15998
rect 13580 15540 13636 15550
rect 13692 15540 13748 15596
rect 13580 15538 13748 15540
rect 13580 15486 13582 15538
rect 13634 15486 13748 15538
rect 13580 15484 13748 15486
rect 13580 15474 13636 15484
rect 13580 15316 13636 15326
rect 13468 15260 13580 15316
rect 12124 15092 12516 15148
rect 11228 14418 11284 15092
rect 11228 14366 11230 14418
rect 11282 14366 11284 14418
rect 11228 13860 11284 14366
rect 11340 13860 11396 13870
rect 11228 13858 11396 13860
rect 11228 13806 11342 13858
rect 11394 13806 11396 13858
rect 11228 13804 11396 13806
rect 11340 13794 11396 13804
rect 11676 13746 11732 13758
rect 11676 13694 11678 13746
rect 11730 13694 11732 13746
rect 11676 13636 11732 13694
rect 11004 13580 11732 13636
rect 11340 12180 11396 12190
rect 11676 12180 11732 13580
rect 12348 12180 12404 12190
rect 11676 12178 12404 12180
rect 11676 12126 12350 12178
rect 12402 12126 12404 12178
rect 11676 12124 12404 12126
rect 12460 12180 12516 15092
rect 12908 14642 12964 15260
rect 13580 15250 13636 15260
rect 12908 14590 12910 14642
rect 12962 14590 12964 14642
rect 12908 14578 12964 14590
rect 12572 14418 12628 14430
rect 12572 14366 12574 14418
rect 12626 14366 12628 14418
rect 12572 13748 12628 14366
rect 12572 13746 12740 13748
rect 12572 13694 12574 13746
rect 12626 13694 12740 13746
rect 12572 13692 12740 13694
rect 12572 13682 12628 13692
rect 12572 12852 12628 12862
rect 12572 12758 12628 12796
rect 12460 12124 12628 12180
rect 11340 12086 11396 12124
rect 12348 12114 12404 12124
rect 10892 11900 11396 11956
rect 10444 11732 10500 11742
rect 10220 11396 10276 11406
rect 10108 10612 10164 10622
rect 10108 10518 10164 10556
rect 9996 10334 9998 10386
rect 10050 10334 10052 10386
rect 9996 10322 10052 10334
rect 10220 10164 10276 11340
rect 10444 10834 10500 11676
rect 10444 10782 10446 10834
rect 10498 10782 10500 10834
rect 10444 10770 10500 10782
rect 11340 11396 11396 11900
rect 11452 11620 11508 11630
rect 11452 11526 11508 11564
rect 11788 11620 11844 11630
rect 10780 10722 10836 10734
rect 10780 10670 10782 10722
rect 10834 10670 10836 10722
rect 9996 10108 10276 10164
rect 10444 10164 10500 10174
rect 9996 9826 10052 10108
rect 10444 9938 10500 10108
rect 10444 9886 10446 9938
rect 10498 9886 10500 9938
rect 10444 9874 10500 9886
rect 9996 9774 9998 9826
rect 10050 9774 10052 9826
rect 9996 9762 10052 9774
rect 10780 9828 10836 10670
rect 11340 10722 11396 11340
rect 11340 10670 11342 10722
rect 11394 10670 11396 10722
rect 11340 10658 11396 10670
rect 10892 10612 10948 10622
rect 11116 10612 11172 10622
rect 10948 10610 11172 10612
rect 10948 10558 11118 10610
rect 11170 10558 11172 10610
rect 10948 10556 11172 10558
rect 10892 10546 10948 10556
rect 11116 10546 11172 10556
rect 11788 10610 11844 11564
rect 12236 11396 12292 11406
rect 12236 11302 12292 11340
rect 11788 10558 11790 10610
rect 11842 10558 11844 10610
rect 11788 10546 11844 10558
rect 12460 10722 12516 10734
rect 12460 10670 12462 10722
rect 12514 10670 12516 10722
rect 11564 10500 11620 10510
rect 11564 10406 11620 10444
rect 12124 10500 12180 10510
rect 12124 10406 12180 10444
rect 10780 9762 10836 9772
rect 12460 9604 12516 10670
rect 12572 9716 12628 12124
rect 12684 11620 12740 13692
rect 13692 12962 13748 15484
rect 13916 15316 13972 15326
rect 14028 15316 14084 15932
rect 13916 15314 14084 15316
rect 13916 15262 13918 15314
rect 13970 15262 14084 15314
rect 13916 15260 14084 15262
rect 13916 15250 13972 15260
rect 14140 15148 14196 16828
rect 14364 16324 14420 17054
rect 14588 17108 14644 17118
rect 15148 17108 15204 17726
rect 15484 17780 15540 18284
rect 15484 17666 15540 17724
rect 15484 17614 15486 17666
rect 15538 17614 15540 17666
rect 15484 17602 15540 17614
rect 15484 17444 15540 17454
rect 14588 17106 15428 17108
rect 14588 17054 14590 17106
rect 14642 17054 15428 17106
rect 14588 17052 15428 17054
rect 14588 17042 14644 17052
rect 15036 16884 15092 16894
rect 15036 16790 15092 16828
rect 15372 16882 15428 17052
rect 15372 16830 15374 16882
rect 15426 16830 15428 16882
rect 15372 16818 15428 16830
rect 15484 16882 15540 17388
rect 15484 16830 15486 16882
rect 15538 16830 15540 16882
rect 15484 16818 15540 16830
rect 14476 16772 14532 16782
rect 15260 16772 15316 16782
rect 14476 16770 14644 16772
rect 14476 16718 14478 16770
rect 14530 16718 14644 16770
rect 14476 16716 14644 16718
rect 14476 16706 14532 16716
rect 14476 16324 14532 16334
rect 14364 16322 14532 16324
rect 14364 16270 14478 16322
rect 14530 16270 14532 16322
rect 14364 16268 14532 16270
rect 14476 16258 14532 16268
rect 13916 15092 14196 15148
rect 13916 13858 13972 15092
rect 13916 13806 13918 13858
rect 13970 13806 13972 13858
rect 13916 13794 13972 13806
rect 13692 12910 13694 12962
rect 13746 12910 13748 12962
rect 13692 12898 13748 12910
rect 14588 12962 14644 16716
rect 14924 15538 14980 15550
rect 14924 15486 14926 15538
rect 14978 15486 14980 15538
rect 14924 14532 14980 15486
rect 15148 15316 15204 15354
rect 15148 15250 15204 15260
rect 14924 14466 14980 14476
rect 15260 14530 15316 16716
rect 15596 16660 15652 23660
rect 16492 23492 16548 23886
rect 16492 23426 16548 23436
rect 16716 23828 16772 23838
rect 15708 23266 15764 23278
rect 15708 23214 15710 23266
rect 15762 23214 15764 23266
rect 15708 21812 15764 23214
rect 15820 23156 15876 23166
rect 16156 23156 16212 23166
rect 16716 23156 16772 23772
rect 15820 23154 16212 23156
rect 15820 23102 15822 23154
rect 15874 23102 16158 23154
rect 16210 23102 16212 23154
rect 15820 23100 16212 23102
rect 15820 22484 15876 23100
rect 16156 23090 16212 23100
rect 16604 23154 16772 23156
rect 16604 23102 16718 23154
rect 16770 23102 16772 23154
rect 16604 23100 16772 23102
rect 15820 22418 15876 22428
rect 15820 21812 15876 21822
rect 15708 21756 15820 21812
rect 15820 20244 15876 21756
rect 16156 21812 16212 21822
rect 16156 21698 16212 21756
rect 16156 21646 16158 21698
rect 16210 21646 16212 21698
rect 16156 21634 16212 21646
rect 15932 21026 15988 21038
rect 15932 20974 15934 21026
rect 15986 20974 15988 21026
rect 15932 20580 15988 20974
rect 16492 20804 16548 20814
rect 15932 20578 16100 20580
rect 15932 20526 15934 20578
rect 15986 20526 16100 20578
rect 15932 20524 16100 20526
rect 15932 20514 15988 20524
rect 15820 20178 15876 20188
rect 15932 20132 15988 20142
rect 15820 19348 15876 19358
rect 15708 18900 15764 18910
rect 15708 18562 15764 18844
rect 15820 18674 15876 19292
rect 15932 19012 15988 20076
rect 16044 20020 16100 20524
rect 16492 20130 16548 20748
rect 16492 20078 16494 20130
rect 16546 20078 16548 20130
rect 16492 20066 16548 20078
rect 16156 20020 16212 20030
rect 16044 19964 16156 20020
rect 16044 19236 16100 19964
rect 16156 19954 16212 19964
rect 16604 19796 16660 23100
rect 16716 23090 16772 23100
rect 17500 22708 17556 26852
rect 18172 26292 18228 26852
rect 19068 26628 19124 27022
rect 19068 26562 19124 26572
rect 19292 27074 19348 27086
rect 19292 27022 19294 27074
rect 19346 27022 19348 27074
rect 18396 26402 18452 26414
rect 18396 26350 18398 26402
rect 18450 26350 18452 26402
rect 18172 26226 18228 26236
rect 18284 26290 18340 26302
rect 18284 26238 18286 26290
rect 18338 26238 18340 26290
rect 18172 25506 18228 25518
rect 18172 25454 18174 25506
rect 18226 25454 18228 25506
rect 17500 22642 17556 22652
rect 17612 25282 17668 25294
rect 17612 25230 17614 25282
rect 17666 25230 17668 25282
rect 17612 21588 17668 25230
rect 18060 24724 18116 24734
rect 17836 24612 17892 24622
rect 17836 24162 17892 24556
rect 17836 24110 17838 24162
rect 17890 24110 17892 24162
rect 17836 24052 17892 24110
rect 17836 23986 17892 23996
rect 18060 23826 18116 24668
rect 18172 24162 18228 25454
rect 18284 25508 18340 26238
rect 18284 25442 18340 25452
rect 18396 25396 18452 26350
rect 18620 26292 18676 26302
rect 18620 26290 18788 26292
rect 18620 26238 18622 26290
rect 18674 26238 18788 26290
rect 18620 26236 18788 26238
rect 18620 26226 18676 26236
rect 18732 26066 18788 26236
rect 18732 26014 18734 26066
rect 18786 26014 18788 26066
rect 18732 26002 18788 26014
rect 18956 26180 19012 26190
rect 19292 26180 19348 27022
rect 18956 26178 19348 26180
rect 18956 26126 18958 26178
rect 19010 26126 19348 26178
rect 18956 26124 19348 26126
rect 19404 27074 19460 27086
rect 19404 27022 19406 27074
rect 19458 27022 19460 27074
rect 19404 26178 19460 27022
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 20412 26404 20468 29932
rect 20748 29986 20804 29998
rect 20748 29934 20750 29986
rect 20802 29934 20804 29986
rect 20748 29092 20804 29934
rect 20860 29540 20916 29550
rect 20972 29540 21028 31724
rect 21084 31556 21140 31566
rect 21084 31106 21140 31500
rect 21308 31554 21364 31566
rect 21308 31502 21310 31554
rect 21362 31502 21364 31554
rect 21308 31444 21364 31502
rect 21308 31378 21364 31388
rect 21644 31554 21700 31566
rect 21644 31502 21646 31554
rect 21698 31502 21700 31554
rect 21196 31332 21252 31342
rect 21196 31218 21252 31276
rect 21196 31166 21198 31218
rect 21250 31166 21252 31218
rect 21196 31154 21252 31166
rect 21308 31220 21364 31230
rect 21644 31220 21700 31502
rect 22988 31556 23044 31724
rect 23100 31556 23156 31566
rect 22988 31554 23156 31556
rect 22988 31502 23102 31554
rect 23154 31502 23156 31554
rect 22988 31500 23156 31502
rect 23100 31490 23156 31500
rect 22092 31220 22148 31230
rect 21308 31218 21588 31220
rect 21308 31166 21310 31218
rect 21362 31166 21588 31218
rect 21308 31164 21588 31166
rect 21644 31218 22148 31220
rect 21644 31166 22094 31218
rect 22146 31166 22148 31218
rect 21644 31164 22148 31166
rect 21308 31154 21364 31164
rect 21084 31054 21086 31106
rect 21138 31054 21140 31106
rect 21084 31042 21140 31054
rect 20916 29484 21028 29540
rect 21420 30994 21476 31006
rect 21420 30942 21422 30994
rect 21474 30942 21476 30994
rect 20860 29446 20916 29484
rect 21308 29426 21364 29438
rect 21308 29374 21310 29426
rect 21362 29374 21364 29426
rect 21308 29204 21364 29374
rect 21308 29138 21364 29148
rect 20748 29026 20804 29036
rect 21420 29092 21476 30942
rect 21532 30996 21588 31164
rect 21756 31108 21812 31164
rect 22092 31154 22148 31164
rect 22316 31220 22372 31230
rect 22316 31126 22372 31164
rect 21756 31042 21812 31052
rect 21644 30996 21700 31006
rect 21532 30994 21700 30996
rect 21532 30942 21646 30994
rect 21698 30942 21700 30994
rect 21532 30940 21700 30942
rect 21644 30930 21700 30940
rect 22988 30996 23044 31006
rect 22988 30902 23044 30940
rect 22204 30884 22260 30894
rect 22204 30790 22260 30828
rect 21644 30212 21700 30222
rect 21644 29986 21700 30156
rect 21644 29934 21646 29986
rect 21698 29934 21700 29986
rect 21644 29922 21700 29934
rect 21532 29652 21588 29662
rect 21532 29426 21588 29596
rect 23212 29650 23268 31724
rect 23660 31556 23716 31838
rect 23996 31890 24052 32956
rect 24556 32562 24612 34076
rect 25004 34132 25060 34860
rect 25452 34468 25508 37324
rect 25228 34412 25508 34468
rect 25004 34066 25060 34076
rect 25116 34130 25172 34142
rect 25116 34078 25118 34130
rect 25170 34078 25172 34130
rect 25116 34020 25172 34078
rect 25116 33954 25172 33964
rect 24556 32510 24558 32562
rect 24610 32510 24612 32562
rect 24556 32498 24612 32510
rect 24668 33684 24724 33694
rect 23996 31838 23998 31890
rect 24050 31838 24052 31890
rect 23996 31826 24052 31838
rect 24220 32004 24276 32014
rect 23660 31490 23716 31500
rect 23212 29598 23214 29650
rect 23266 29598 23268 29650
rect 22204 29540 22260 29550
rect 22204 29446 22260 29484
rect 21532 29374 21534 29426
rect 21586 29374 21588 29426
rect 21532 29362 21588 29374
rect 22540 29428 22596 29438
rect 22876 29428 22932 29438
rect 22540 29426 22932 29428
rect 22540 29374 22542 29426
rect 22594 29374 22878 29426
rect 22930 29374 22932 29426
rect 22540 29372 22932 29374
rect 21756 29204 21812 29214
rect 21420 29026 21476 29036
rect 21644 29202 21812 29204
rect 21644 29150 21758 29202
rect 21810 29150 21812 29202
rect 21644 29148 21812 29150
rect 21644 28868 21700 29148
rect 21756 29138 21812 29148
rect 21868 29204 21924 29214
rect 21868 29202 22484 29204
rect 21868 29150 21870 29202
rect 21922 29150 22484 29202
rect 21868 29148 22484 29150
rect 20748 28812 21700 28868
rect 20748 28754 20804 28812
rect 20748 28702 20750 28754
rect 20802 28702 20804 28754
rect 20524 28420 20580 28430
rect 20524 27860 20580 28364
rect 20524 27186 20580 27804
rect 20524 27134 20526 27186
rect 20578 27134 20580 27186
rect 20524 27122 20580 27134
rect 20748 26908 20804 28702
rect 21868 28308 21924 29148
rect 21532 28252 21924 28308
rect 22092 28530 22148 28542
rect 22092 28478 22094 28530
rect 22146 28478 22148 28530
rect 21196 27858 21252 27870
rect 21196 27806 21198 27858
rect 21250 27806 21252 27858
rect 21196 27748 21252 27806
rect 21196 27682 21252 27692
rect 21308 27636 21364 27646
rect 21308 27074 21364 27580
rect 21308 27022 21310 27074
rect 21362 27022 21364 27074
rect 21308 27010 21364 27022
rect 21532 27074 21588 28252
rect 21532 27022 21534 27074
rect 21586 27022 21588 27074
rect 21532 27010 21588 27022
rect 21644 28082 21700 28094
rect 21644 28030 21646 28082
rect 21698 28030 21700 28082
rect 21644 27972 21700 28030
rect 22092 28084 22148 28478
rect 22092 28018 22148 28028
rect 22428 28082 22484 29148
rect 22428 28030 22430 28082
rect 22482 28030 22484 28082
rect 22428 28018 22484 28030
rect 21644 27074 21700 27916
rect 21756 27970 21812 27982
rect 21756 27918 21758 27970
rect 21810 27918 21812 27970
rect 21756 27860 21812 27918
rect 22204 27972 22260 27982
rect 22204 27878 22260 27916
rect 21756 27794 21812 27804
rect 22092 27860 22148 27870
rect 22092 27298 22148 27804
rect 22540 27746 22596 29372
rect 22876 29362 22932 29372
rect 23212 28084 23268 29598
rect 23324 31444 23380 31454
rect 23324 30994 23380 31388
rect 23660 31108 23716 31118
rect 23996 31108 24052 31118
rect 24220 31108 24276 31948
rect 24444 31666 24500 31678
rect 24444 31614 24446 31666
rect 24498 31614 24500 31666
rect 24444 31444 24500 31614
rect 24444 31378 24500 31388
rect 23660 31106 24276 31108
rect 23660 31054 23662 31106
rect 23714 31054 23998 31106
rect 24050 31054 24276 31106
rect 23660 31052 24276 31054
rect 23660 31042 23716 31052
rect 23996 31042 24052 31052
rect 23324 30942 23326 30994
rect 23378 30942 23380 30994
rect 23324 29540 23380 30942
rect 24108 30882 24164 30894
rect 24108 30830 24110 30882
rect 24162 30830 24164 30882
rect 24108 30324 24164 30830
rect 24220 30772 24276 31052
rect 24556 31108 24612 31118
rect 24556 31014 24612 31052
rect 24332 30996 24388 31006
rect 24668 30996 24724 33628
rect 25228 33236 25284 34412
rect 25228 33170 25284 33180
rect 25340 34242 25396 34254
rect 25340 34190 25342 34242
rect 25394 34190 25396 34242
rect 25340 32900 25396 34190
rect 25452 34130 25508 34142
rect 25452 34078 25454 34130
rect 25506 34078 25508 34130
rect 25452 33684 25508 34078
rect 25452 33618 25508 33628
rect 25228 32844 25396 32900
rect 25452 33012 25508 33022
rect 25116 32562 25172 32574
rect 25116 32510 25118 32562
rect 25170 32510 25172 32562
rect 25116 32004 25172 32510
rect 25228 32228 25284 32844
rect 25452 32786 25508 32956
rect 25452 32734 25454 32786
rect 25506 32734 25508 32786
rect 25452 32722 25508 32734
rect 25340 32676 25396 32686
rect 25340 32564 25396 32620
rect 25452 32564 25508 32574
rect 25340 32562 25508 32564
rect 25340 32510 25454 32562
rect 25506 32510 25508 32562
rect 25340 32508 25508 32510
rect 25452 32498 25508 32508
rect 25228 32172 25508 32228
rect 25116 31778 25172 31948
rect 25116 31726 25118 31778
rect 25170 31726 25172 31778
rect 25116 31714 25172 31726
rect 25228 31892 25284 31902
rect 25228 31666 25284 31836
rect 25452 31778 25508 32172
rect 25452 31726 25454 31778
rect 25506 31726 25508 31778
rect 25452 31714 25508 31726
rect 25564 31780 25620 37660
rect 25676 37650 25732 37660
rect 25676 36484 25732 36494
rect 25788 36484 25844 38612
rect 25900 38276 25956 38286
rect 25900 38182 25956 38220
rect 26572 38162 26628 41244
rect 26796 41076 26852 41086
rect 26684 41074 26852 41076
rect 26684 41022 26798 41074
rect 26850 41022 26852 41074
rect 26684 41020 26852 41022
rect 26684 40964 26740 41020
rect 26796 41010 26852 41020
rect 26908 41076 26964 41086
rect 27020 41076 27076 43652
rect 27244 43652 27300 43662
rect 27244 43558 27300 43596
rect 27132 43540 27188 43550
rect 27132 43316 27188 43484
rect 27132 43250 27188 43260
rect 27356 43092 27412 45276
rect 27804 45266 27860 45276
rect 27580 45220 27636 45230
rect 27468 45108 27524 45118
rect 27468 45014 27524 45052
rect 27580 44324 27636 45164
rect 27916 45108 27972 46060
rect 27804 45052 27972 45108
rect 28252 45668 28308 45678
rect 27692 44324 27748 44334
rect 27580 44322 27748 44324
rect 27580 44270 27694 44322
rect 27746 44270 27748 44322
rect 27580 44268 27748 44270
rect 27692 44258 27748 44268
rect 27468 43650 27524 43662
rect 27468 43598 27470 43650
rect 27522 43598 27524 43650
rect 27468 43540 27524 43598
rect 27580 43540 27636 43550
rect 27468 43538 27636 43540
rect 27468 43486 27582 43538
rect 27634 43486 27636 43538
rect 27468 43484 27636 43486
rect 27804 43540 27860 45052
rect 28252 44212 28308 45612
rect 27916 44210 28308 44212
rect 27916 44158 28254 44210
rect 28306 44158 28308 44210
rect 27916 44156 28308 44158
rect 27916 43762 27972 44156
rect 28252 44146 28308 44156
rect 27916 43710 27918 43762
rect 27970 43710 27972 43762
rect 27916 43698 27972 43710
rect 28028 43540 28084 43550
rect 27804 43484 27972 43540
rect 27580 43474 27636 43484
rect 27132 43036 27412 43092
rect 27132 42532 27188 43036
rect 27244 42868 27300 42878
rect 27244 42774 27300 42812
rect 27468 42756 27524 42766
rect 27132 42466 27188 42476
rect 27356 42754 27524 42756
rect 27356 42702 27470 42754
rect 27522 42702 27524 42754
rect 27356 42700 27524 42702
rect 27356 42308 27412 42700
rect 27468 42690 27524 42700
rect 27804 42644 27860 42654
rect 27804 42550 27860 42588
rect 27132 42252 27412 42308
rect 27132 42196 27188 42252
rect 27132 42102 27188 42140
rect 26908 41074 27076 41076
rect 26908 41022 26910 41074
rect 26962 41022 27076 41074
rect 26908 41020 27076 41022
rect 27580 41746 27636 41758
rect 27580 41694 27582 41746
rect 27634 41694 27636 41746
rect 26908 41010 26964 41020
rect 27132 40964 27188 40974
rect 26684 40898 26740 40908
rect 27020 40962 27188 40964
rect 27020 40910 27134 40962
rect 27186 40910 27188 40962
rect 27020 40908 27188 40910
rect 27020 39618 27076 40908
rect 27132 40898 27188 40908
rect 27244 40740 27300 40750
rect 27132 40516 27188 40526
rect 27132 40422 27188 40460
rect 27020 39566 27022 39618
rect 27074 39566 27076 39618
rect 27020 39554 27076 39566
rect 27132 39508 27188 39518
rect 27132 39172 27188 39452
rect 26796 39116 27188 39172
rect 26796 38276 26852 39116
rect 26796 38210 26852 38220
rect 26572 38110 26574 38162
rect 26626 38110 26628 38162
rect 26124 38052 26180 38062
rect 26012 37940 26068 37950
rect 25900 37938 26068 37940
rect 25900 37886 26014 37938
rect 26066 37886 26068 37938
rect 25900 37884 26068 37886
rect 25900 37266 25956 37884
rect 26012 37874 26068 37884
rect 25900 37214 25902 37266
rect 25954 37214 25956 37266
rect 25900 37202 25956 37214
rect 26012 37266 26068 37278
rect 26012 37214 26014 37266
rect 26066 37214 26068 37266
rect 25676 36482 25844 36484
rect 25676 36430 25678 36482
rect 25730 36430 25844 36482
rect 25676 36428 25844 36430
rect 25676 35588 25732 36428
rect 25676 35522 25732 35532
rect 25788 35586 25844 35598
rect 25788 35534 25790 35586
rect 25842 35534 25844 35586
rect 25788 35474 25844 35534
rect 25788 35422 25790 35474
rect 25842 35422 25844 35474
rect 25788 35252 25844 35422
rect 25788 35186 25844 35196
rect 25564 31714 25620 31724
rect 25676 35140 25732 35150
rect 25676 34692 25732 35084
rect 26012 35140 26068 37214
rect 26124 35812 26180 37996
rect 26572 37716 26628 38110
rect 26572 37650 26628 37660
rect 26348 37378 26404 37390
rect 26348 37326 26350 37378
rect 26402 37326 26404 37378
rect 26348 37268 26404 37326
rect 26796 37380 26852 37418
rect 26796 37314 26852 37324
rect 26572 37268 26628 37278
rect 26236 37154 26292 37166
rect 26236 37102 26238 37154
rect 26290 37102 26292 37154
rect 26236 37044 26292 37102
rect 26236 36978 26292 36988
rect 26124 35746 26180 35756
rect 26012 35074 26068 35084
rect 25676 33124 25732 34636
rect 25788 34802 25844 34814
rect 25788 34750 25790 34802
rect 25842 34750 25844 34802
rect 25788 34580 25844 34750
rect 26236 34804 26292 34814
rect 25788 34524 26180 34580
rect 26012 34356 26068 34366
rect 26012 34262 26068 34300
rect 26124 34354 26180 34524
rect 26124 34302 26126 34354
rect 26178 34302 26180 34354
rect 26124 34290 26180 34302
rect 26236 34354 26292 34748
rect 26236 34302 26238 34354
rect 26290 34302 26292 34354
rect 26236 34290 26292 34302
rect 26348 34132 26404 37212
rect 26460 37212 26572 37268
rect 26460 36594 26516 37212
rect 26572 37202 26628 37212
rect 26684 37266 26740 37278
rect 26684 37214 26686 37266
rect 26738 37214 26740 37266
rect 26684 37044 26740 37214
rect 26684 36978 26740 36988
rect 26908 37266 26964 37278
rect 26908 37214 26910 37266
rect 26962 37214 26964 37266
rect 26460 36542 26462 36594
rect 26514 36542 26516 36594
rect 26460 36530 26516 36542
rect 26572 36820 26628 36830
rect 26572 35308 26628 36764
rect 26908 35476 26964 37214
rect 27244 35588 27300 40684
rect 27580 37492 27636 41694
rect 27916 38668 27972 43484
rect 28028 42980 28084 43484
rect 28252 43540 28308 43550
rect 28252 43446 28308 43484
rect 28700 43428 28756 50372
rect 28812 43652 28868 43662
rect 28812 43558 28868 43596
rect 28924 43540 28980 43550
rect 28700 43372 28868 43428
rect 28028 42914 28084 42924
rect 28476 43316 28532 43326
rect 28588 43316 28644 43326
rect 28532 43314 28644 43316
rect 28532 43262 28590 43314
rect 28642 43262 28644 43314
rect 28532 43260 28644 43262
rect 28252 41972 28308 41982
rect 28476 41972 28532 43260
rect 28588 43250 28644 43260
rect 28252 41970 28532 41972
rect 28252 41918 28254 41970
rect 28306 41918 28532 41970
rect 28252 41916 28532 41918
rect 28252 41906 28308 41916
rect 28700 39844 28756 39854
rect 28700 39730 28756 39788
rect 28700 39678 28702 39730
rect 28754 39678 28756 39730
rect 28700 39666 28756 39678
rect 27916 38612 28532 38668
rect 28140 38164 28196 38174
rect 27804 38108 28140 38164
rect 27580 37436 27748 37492
rect 27356 37268 27412 37278
rect 27580 37268 27636 37278
rect 27356 37266 27636 37268
rect 27356 37214 27358 37266
rect 27410 37214 27582 37266
rect 27634 37214 27636 37266
rect 27356 37212 27636 37214
rect 27356 37202 27412 37212
rect 27580 37202 27636 37212
rect 27356 36484 27412 36494
rect 27692 36484 27748 37436
rect 27804 37490 27860 38108
rect 28140 38070 28196 38108
rect 27804 37438 27806 37490
rect 27858 37438 27860 37490
rect 27804 37426 27860 37438
rect 27916 37940 27972 37950
rect 27916 37378 27972 37884
rect 27916 37326 27918 37378
rect 27970 37326 27972 37378
rect 27916 37314 27972 37326
rect 28364 37492 28420 37502
rect 28364 37266 28420 37436
rect 28364 37214 28366 37266
rect 28418 37214 28420 37266
rect 28364 37202 28420 37214
rect 27356 35922 27412 36428
rect 27356 35870 27358 35922
rect 27410 35870 27412 35922
rect 27356 35858 27412 35870
rect 27580 36428 27748 36484
rect 27916 36484 27972 36494
rect 27244 35522 27300 35532
rect 26908 35410 26964 35420
rect 27244 35364 27300 35374
rect 26572 35252 26852 35308
rect 25228 31614 25230 31666
rect 25282 31614 25284 31666
rect 25228 31602 25284 31614
rect 25676 31668 25732 33068
rect 26236 34076 26404 34132
rect 26684 34692 26740 34702
rect 26684 34130 26740 34636
rect 26684 34078 26686 34130
rect 26738 34078 26740 34130
rect 25788 32562 25844 32574
rect 25788 32510 25790 32562
rect 25842 32510 25844 32562
rect 25788 32004 25844 32510
rect 25788 31948 26180 32004
rect 26124 31890 26180 31948
rect 26124 31838 26126 31890
rect 26178 31838 26180 31890
rect 26124 31826 26180 31838
rect 26012 31780 26068 31790
rect 26012 31686 26068 31724
rect 25676 31612 25956 31668
rect 24780 31554 24836 31566
rect 24780 31502 24782 31554
rect 24834 31502 24836 31554
rect 24780 31444 24836 31502
rect 24780 31378 24836 31388
rect 25452 31332 25508 31342
rect 25228 31220 25284 31230
rect 25228 31106 25284 31164
rect 25228 31054 25230 31106
rect 25282 31054 25284 31106
rect 25228 31042 25284 31054
rect 25340 31108 25396 31118
rect 25340 31014 25396 31052
rect 25452 31108 25508 31276
rect 25452 31106 25732 31108
rect 25452 31054 25454 31106
rect 25506 31054 25732 31106
rect 25452 31052 25732 31054
rect 25452 31042 25508 31052
rect 24332 30994 24500 30996
rect 24332 30942 24334 30994
rect 24386 30942 24500 30994
rect 24332 30940 24500 30942
rect 24332 30930 24388 30940
rect 24220 30716 24388 30772
rect 23324 29474 23380 29484
rect 23548 30268 24164 30324
rect 23548 29538 23604 30268
rect 24220 30212 24276 30222
rect 23884 30100 23940 30110
rect 23660 30098 23940 30100
rect 23660 30046 23886 30098
rect 23938 30046 23940 30098
rect 23660 30044 23940 30046
rect 23660 29650 23716 30044
rect 23884 30034 23940 30044
rect 23660 29598 23662 29650
rect 23714 29598 23716 29650
rect 23660 29586 23716 29598
rect 24220 29650 24276 30156
rect 24220 29598 24222 29650
rect 24274 29598 24276 29650
rect 24220 29586 24276 29598
rect 23548 29486 23550 29538
rect 23602 29486 23604 29538
rect 23548 29474 23604 29486
rect 23324 28084 23380 28094
rect 23212 28082 23380 28084
rect 23212 28030 23326 28082
rect 23378 28030 23380 28082
rect 23212 28028 23380 28030
rect 22540 27694 22542 27746
rect 22594 27694 22596 27746
rect 22540 27682 22596 27694
rect 22652 27970 22708 27982
rect 22652 27918 22654 27970
rect 22706 27918 22708 27970
rect 22652 27636 22708 27918
rect 22988 27636 23044 27646
rect 22652 27570 22708 27580
rect 22764 27580 22988 27636
rect 22092 27246 22094 27298
rect 22146 27246 22148 27298
rect 22092 27234 22148 27246
rect 22652 27188 22708 27198
rect 22764 27188 22820 27580
rect 22988 27570 23044 27580
rect 22652 27186 22820 27188
rect 22652 27134 22654 27186
rect 22706 27134 22820 27186
rect 22652 27132 22820 27134
rect 22876 27300 22932 27310
rect 22876 27186 22932 27244
rect 22876 27134 22878 27186
rect 22930 27134 22932 27186
rect 22652 27122 22708 27132
rect 22876 27122 22932 27134
rect 21644 27022 21646 27074
rect 21698 27022 21700 27074
rect 21644 27010 21700 27022
rect 20636 26852 20804 26908
rect 20412 26338 20468 26348
rect 20524 26740 20580 26750
rect 19404 26126 19406 26178
rect 19458 26126 19460 26178
rect 18732 25508 18788 25518
rect 18732 25414 18788 25452
rect 18508 25396 18564 25406
rect 18396 25394 18676 25396
rect 18396 25342 18510 25394
rect 18562 25342 18676 25394
rect 18396 25340 18676 25342
rect 18508 25330 18564 25340
rect 18508 24612 18564 24622
rect 18508 24518 18564 24556
rect 18172 24110 18174 24162
rect 18226 24110 18228 24162
rect 18172 24098 18228 24110
rect 18284 24498 18340 24510
rect 18284 24446 18286 24498
rect 18338 24446 18340 24498
rect 18060 23774 18062 23826
rect 18114 23774 18116 23826
rect 18060 23762 18116 23774
rect 18172 23156 18228 23166
rect 18284 23156 18340 24446
rect 18620 24162 18676 25340
rect 18956 25284 19012 26124
rect 19404 25844 19460 26126
rect 19404 25778 19460 25788
rect 19516 26066 19572 26078
rect 19516 26014 19518 26066
rect 19570 26014 19572 26066
rect 19516 25506 19572 26014
rect 20524 25620 20580 26684
rect 19516 25454 19518 25506
rect 19570 25454 19572 25506
rect 19516 25442 19572 25454
rect 20076 25618 20580 25620
rect 20076 25566 20526 25618
rect 20578 25566 20580 25618
rect 20076 25564 20580 25566
rect 20076 25394 20132 25564
rect 20524 25554 20580 25564
rect 20076 25342 20078 25394
rect 20130 25342 20132 25394
rect 20076 25330 20132 25342
rect 18956 25218 19012 25228
rect 19068 25282 19124 25294
rect 19852 25284 19908 25294
rect 19068 25230 19070 25282
rect 19122 25230 19124 25282
rect 19068 24724 19124 25230
rect 19628 25282 19908 25284
rect 19628 25230 19854 25282
rect 19906 25230 19908 25282
rect 19628 25228 19908 25230
rect 19292 24724 19348 24734
rect 19628 24724 19684 25228
rect 19852 25218 19908 25228
rect 20188 25284 20244 25294
rect 20188 25190 20244 25228
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 19068 24668 19292 24724
rect 19348 24668 19684 24724
rect 20188 24724 20244 24734
rect 20524 24724 20580 24734
rect 20188 24722 20580 24724
rect 20188 24670 20190 24722
rect 20242 24670 20526 24722
rect 20578 24670 20580 24722
rect 20188 24668 20580 24670
rect 19292 24630 19348 24668
rect 19740 24612 19796 24622
rect 19740 24518 19796 24556
rect 18620 24110 18622 24162
rect 18674 24110 18676 24162
rect 18620 24098 18676 24110
rect 20188 24162 20244 24668
rect 20524 24658 20580 24668
rect 20188 24110 20190 24162
rect 20242 24110 20244 24162
rect 20188 24098 20244 24110
rect 20636 24052 20692 26852
rect 23212 26516 23268 26526
rect 20412 23996 20692 24052
rect 20748 26180 20804 26190
rect 22988 26180 23044 26190
rect 19740 23940 19796 23950
rect 19964 23940 20020 23950
rect 19740 23938 19964 23940
rect 19740 23886 19742 23938
rect 19794 23886 19964 23938
rect 19740 23884 19964 23886
rect 19740 23874 19796 23884
rect 19964 23846 20020 23884
rect 18508 23828 18564 23838
rect 19404 23828 19460 23838
rect 18508 23734 18564 23772
rect 19292 23826 19460 23828
rect 19292 23774 19406 23826
rect 19458 23774 19460 23826
rect 19292 23772 19460 23774
rect 18620 23716 18676 23726
rect 18620 23622 18676 23660
rect 18060 23154 18340 23156
rect 18060 23102 18174 23154
rect 18226 23102 18340 23154
rect 18060 23100 18340 23102
rect 17836 22930 17892 22942
rect 17836 22878 17838 22930
rect 17890 22878 17892 22930
rect 17836 22372 17892 22878
rect 17836 22306 17892 22316
rect 18060 22372 18116 23100
rect 18172 23090 18228 23100
rect 18732 23044 18788 23054
rect 18732 23042 19012 23044
rect 18732 22990 18734 23042
rect 18786 22990 19012 23042
rect 18732 22988 19012 22990
rect 18732 22978 18788 22988
rect 18172 22930 18228 22942
rect 18172 22878 18174 22930
rect 18226 22878 18228 22930
rect 18172 22596 18228 22878
rect 18172 22540 18564 22596
rect 18172 22372 18228 22382
rect 18060 22370 18228 22372
rect 18060 22318 18174 22370
rect 18226 22318 18228 22370
rect 18060 22316 18228 22318
rect 17948 22258 18004 22270
rect 17948 22206 17950 22258
rect 18002 22206 18004 22258
rect 17948 21700 18004 22206
rect 17948 21634 18004 21644
rect 17612 21494 17668 21532
rect 17724 21474 17780 21486
rect 17724 21422 17726 21474
rect 17778 21422 17780 21474
rect 17276 20916 17332 20926
rect 17276 20914 17556 20916
rect 17276 20862 17278 20914
rect 17330 20862 17556 20914
rect 17276 20860 17556 20862
rect 17276 20850 17332 20860
rect 16828 20802 16884 20814
rect 16828 20750 16830 20802
rect 16882 20750 16884 20802
rect 16716 20132 16772 20142
rect 16828 20132 16884 20750
rect 16772 20076 16884 20132
rect 16716 20066 16772 20076
rect 17388 20020 17444 20030
rect 16492 19740 16660 19796
rect 16828 20018 17444 20020
rect 16828 19966 17390 20018
rect 17442 19966 17444 20018
rect 16828 19964 17444 19966
rect 16492 19236 16548 19740
rect 16044 19170 16100 19180
rect 16380 19234 16548 19236
rect 16380 19182 16494 19234
rect 16546 19182 16548 19234
rect 16380 19180 16548 19182
rect 15932 19010 16324 19012
rect 15932 18958 15934 19010
rect 15986 18958 16324 19010
rect 15932 18956 16324 18958
rect 15932 18946 15988 18956
rect 15820 18622 15822 18674
rect 15874 18622 15876 18674
rect 15820 18610 15876 18622
rect 15708 18510 15710 18562
rect 15762 18510 15764 18562
rect 15708 18498 15764 18510
rect 16044 18564 16100 18574
rect 16044 18450 16100 18508
rect 16044 18398 16046 18450
rect 16098 18398 16100 18450
rect 16044 18386 16100 18398
rect 16268 18450 16324 18956
rect 16268 18398 16270 18450
rect 16322 18398 16324 18450
rect 16268 18386 16324 18398
rect 15932 17780 15988 17790
rect 15932 17686 15988 17724
rect 16380 17668 16436 19180
rect 16492 19170 16548 19180
rect 16716 19460 16772 19470
rect 16604 19122 16660 19134
rect 16604 19070 16606 19122
rect 16658 19070 16660 19122
rect 16604 18788 16660 19070
rect 16604 18722 16660 18732
rect 16492 18452 16548 18462
rect 16492 18358 16548 18396
rect 16716 18450 16772 19404
rect 16828 18562 16884 19964
rect 17388 19954 17444 19964
rect 17052 19460 17108 19470
rect 17052 19346 17108 19404
rect 17052 19294 17054 19346
rect 17106 19294 17108 19346
rect 17052 19282 17108 19294
rect 17500 19236 17556 20860
rect 17724 20804 17780 21422
rect 18060 21252 18116 22316
rect 18172 22306 18228 22316
rect 18396 22372 18452 22382
rect 18396 21812 18452 22316
rect 18172 21476 18228 21486
rect 18172 21382 18228 21420
rect 18060 21196 18228 21252
rect 17724 20738 17780 20748
rect 18060 20802 18116 20814
rect 18060 20750 18062 20802
rect 18114 20750 18116 20802
rect 16828 18510 16830 18562
rect 16882 18510 16884 18562
rect 16828 18498 16884 18510
rect 17388 19180 17556 19236
rect 17836 19906 17892 19918
rect 17836 19854 17838 19906
rect 17890 19854 17892 19906
rect 16716 18398 16718 18450
rect 16770 18398 16772 18450
rect 16716 18386 16772 18398
rect 17388 18452 17444 19180
rect 17500 19010 17556 19022
rect 17500 18958 17502 19010
rect 17554 18958 17556 19010
rect 17500 18788 17556 18958
rect 17500 18722 17556 18732
rect 17388 18386 17444 18396
rect 17836 18338 17892 19854
rect 18060 19460 18116 20750
rect 18172 20130 18228 21196
rect 18172 20078 18174 20130
rect 18226 20078 18228 20130
rect 18172 20066 18228 20078
rect 18396 20018 18452 21756
rect 18508 21588 18564 22540
rect 18732 21588 18788 21598
rect 18508 21586 18788 21588
rect 18508 21534 18734 21586
rect 18786 21534 18788 21586
rect 18508 21532 18788 21534
rect 18732 21522 18788 21532
rect 18620 20914 18676 20926
rect 18620 20862 18622 20914
rect 18674 20862 18676 20914
rect 18396 19966 18398 20018
rect 18450 19966 18452 20018
rect 18396 19954 18452 19966
rect 18508 20020 18564 20030
rect 18060 19394 18116 19404
rect 17948 19348 18004 19358
rect 17948 19254 18004 19292
rect 18508 19234 18564 19964
rect 18508 19182 18510 19234
rect 18562 19182 18564 19234
rect 18508 19170 18564 19182
rect 18060 18564 18116 18574
rect 18060 18470 18116 18508
rect 17836 18286 17838 18338
rect 17890 18286 17892 18338
rect 16380 17602 16436 17612
rect 17164 17668 17220 17678
rect 15596 16594 15652 16604
rect 16044 17442 16100 17454
rect 16044 17390 16046 17442
rect 16098 17390 16100 17442
rect 16044 16098 16100 17390
rect 16156 17444 16212 17454
rect 16156 17350 16212 17388
rect 17052 17442 17108 17454
rect 17052 17390 17054 17442
rect 17106 17390 17108 17442
rect 16044 16046 16046 16098
rect 16098 16046 16100 16098
rect 15932 15988 15988 15998
rect 15932 15894 15988 15932
rect 16044 15314 16100 16046
rect 16044 15262 16046 15314
rect 16098 15262 16100 15314
rect 16044 15250 16100 15262
rect 16268 16882 16324 16894
rect 16268 16830 16270 16882
rect 16322 16830 16324 16882
rect 16268 16212 16324 16830
rect 15708 15204 15764 15214
rect 15596 15092 15764 15148
rect 15596 14642 15652 15092
rect 15596 14590 15598 14642
rect 15650 14590 15652 14642
rect 15596 14578 15652 14590
rect 16268 14642 16324 16156
rect 16940 16884 16996 16894
rect 16268 14590 16270 14642
rect 16322 14590 16324 14642
rect 16268 14578 16324 14590
rect 16380 16100 16436 16110
rect 16380 15204 16436 16044
rect 16940 16098 16996 16828
rect 16940 16046 16942 16098
rect 16994 16046 16996 16098
rect 16940 16034 16996 16046
rect 15260 14478 15262 14530
rect 15314 14478 15316 14530
rect 15260 13858 15316 14478
rect 16380 14530 16436 15148
rect 16492 15988 16548 15998
rect 16492 15426 16548 15932
rect 17052 15988 17108 17390
rect 17052 15922 17108 15932
rect 16492 15374 16494 15426
rect 16546 15374 16548 15426
rect 16492 15148 16548 15374
rect 17164 15148 17220 17612
rect 17276 17554 17332 17566
rect 17276 17502 17278 17554
rect 17330 17502 17332 17554
rect 17276 15876 17332 17502
rect 17276 15810 17332 15820
rect 16492 15092 16660 15148
rect 17164 15092 17668 15148
rect 16380 14478 16382 14530
rect 16434 14478 16436 14530
rect 15260 13806 15262 13858
rect 15314 13806 15316 13858
rect 15260 13794 15316 13806
rect 15484 13858 15540 13870
rect 15484 13806 15486 13858
rect 15538 13806 15540 13858
rect 14588 12910 14590 12962
rect 14642 12910 14644 12962
rect 14588 12898 14644 12910
rect 15036 13074 15092 13086
rect 15036 13022 15038 13074
rect 15090 13022 15092 13074
rect 14364 12850 14420 12862
rect 14364 12798 14366 12850
rect 14418 12798 14420 12850
rect 12908 12740 12964 12750
rect 14028 12740 14084 12750
rect 12908 12738 13412 12740
rect 12908 12686 12910 12738
rect 12962 12686 13412 12738
rect 12908 12684 13412 12686
rect 12908 12674 12964 12684
rect 12684 11394 12740 11564
rect 12684 11342 12686 11394
rect 12738 11342 12740 11394
rect 12684 11330 12740 11342
rect 12796 12178 12852 12190
rect 12796 12126 12798 12178
rect 12850 12126 12852 12178
rect 12796 10164 12852 12126
rect 13020 11954 13076 11966
rect 13020 11902 13022 11954
rect 13074 11902 13076 11954
rect 12908 11284 12964 11294
rect 12908 11190 12964 11228
rect 12796 10098 12852 10108
rect 12796 9828 12852 9838
rect 12796 9734 12852 9772
rect 12684 9716 12740 9726
rect 12572 9714 12740 9716
rect 12572 9662 12686 9714
rect 12738 9662 12740 9714
rect 12572 9660 12740 9662
rect 12684 9604 12740 9660
rect 12460 9602 12628 9604
rect 12460 9550 12462 9602
rect 12514 9550 12628 9602
rect 12460 9548 12628 9550
rect 12684 9548 12852 9604
rect 12460 9538 12516 9548
rect 9548 9202 9604 9212
rect 12572 9154 12628 9548
rect 12572 9102 12574 9154
rect 12626 9102 12628 9154
rect 12572 9090 12628 9102
rect 9548 9042 9604 9054
rect 9548 8990 9550 9042
rect 9602 8990 9604 9042
rect 9548 8372 9604 8990
rect 9548 7924 9604 8316
rect 9884 9042 9940 9054
rect 9884 8990 9886 9042
rect 9938 8990 9940 9042
rect 9660 8258 9716 8270
rect 9660 8206 9662 8258
rect 9714 8206 9716 8258
rect 9660 8148 9716 8206
rect 9716 8092 9828 8148
rect 9660 8082 9716 8092
rect 9548 7868 9716 7924
rect 9324 7028 9380 7532
rect 9548 7700 9604 7710
rect 9548 7474 9604 7644
rect 9548 7422 9550 7474
rect 9602 7422 9604 7474
rect 9548 7410 9604 7422
rect 9324 6972 9604 7028
rect 9324 6692 9380 6702
rect 9212 6690 9380 6692
rect 9212 6638 9326 6690
rect 9378 6638 9380 6690
rect 9212 6636 9380 6638
rect 9324 6626 9380 6636
rect 9436 6580 9492 6590
rect 9548 6580 9604 6972
rect 9660 6690 9716 7868
rect 9772 7700 9828 8092
rect 9884 7812 9940 8990
rect 10108 9044 10164 9054
rect 10108 8950 10164 8988
rect 9996 8930 10052 8942
rect 9996 8878 9998 8930
rect 10050 8878 10052 8930
rect 9996 8372 10052 8878
rect 9996 8306 10052 8316
rect 11228 8372 11284 8382
rect 11004 8260 11060 8270
rect 11004 8166 11060 8204
rect 11228 8258 11284 8316
rect 11228 8206 11230 8258
rect 11282 8206 11284 8258
rect 11228 8194 11284 8206
rect 11676 8370 11732 8382
rect 11676 8318 11678 8370
rect 11730 8318 11732 8370
rect 9884 7756 10500 7812
rect 10444 7700 10500 7756
rect 9772 7644 10052 7700
rect 9996 7474 10052 7644
rect 10444 7698 10836 7700
rect 10444 7646 10446 7698
rect 10498 7646 10836 7698
rect 10444 7644 10836 7646
rect 10444 7634 10500 7644
rect 9996 7422 9998 7474
rect 10050 7422 10052 7474
rect 9996 7410 10052 7422
rect 9772 7252 9828 7262
rect 9772 7158 9828 7196
rect 10668 6914 10724 7644
rect 10780 7474 10836 7644
rect 10780 7422 10782 7474
rect 10834 7422 10836 7474
rect 10780 7410 10836 7422
rect 11004 7476 11060 7486
rect 11564 7476 11620 7486
rect 11004 7474 11620 7476
rect 11004 7422 11006 7474
rect 11058 7422 11566 7474
rect 11618 7422 11620 7474
rect 11004 7420 11620 7422
rect 11004 7410 11060 7420
rect 11564 7410 11620 7420
rect 11004 7252 11060 7262
rect 10668 6862 10670 6914
rect 10722 6862 10724 6914
rect 10668 6850 10724 6862
rect 10892 7196 11004 7252
rect 9660 6638 9662 6690
rect 9714 6638 9716 6690
rect 9660 6626 9716 6638
rect 9436 6578 9604 6580
rect 9436 6526 9438 6578
rect 9490 6526 9604 6578
rect 9436 6524 9604 6526
rect 10892 6578 10948 7196
rect 11004 7186 11060 7196
rect 11340 7252 11396 7262
rect 11340 7250 11620 7252
rect 11340 7198 11342 7250
rect 11394 7198 11620 7250
rect 11340 7196 11620 7198
rect 11340 7186 11396 7196
rect 11004 6804 11060 6814
rect 11340 6804 11396 6814
rect 11004 6802 11396 6804
rect 11004 6750 11006 6802
rect 11058 6750 11342 6802
rect 11394 6750 11396 6802
rect 11004 6748 11396 6750
rect 11004 6738 11060 6748
rect 10892 6526 10894 6578
rect 10946 6526 10948 6578
rect 9436 6514 9492 6524
rect 10892 6514 10948 6526
rect 11340 6580 11396 6748
rect 11340 6514 11396 6524
rect 11564 6578 11620 7196
rect 11676 7028 11732 8318
rect 12348 8372 12404 8382
rect 11788 8260 11844 8270
rect 11788 8166 11844 8204
rect 12348 8146 12404 8316
rect 12348 8094 12350 8146
rect 12402 8094 12404 8146
rect 12348 8082 12404 8094
rect 12684 8146 12740 8158
rect 12684 8094 12686 8146
rect 12738 8094 12740 8146
rect 12684 8036 12740 8094
rect 12796 8146 12852 9548
rect 13020 9042 13076 11902
rect 13356 11396 13412 12684
rect 13692 12738 14084 12740
rect 13692 12686 14030 12738
rect 14082 12686 14084 12738
rect 13692 12684 14084 12686
rect 13468 11396 13524 11406
rect 13356 11340 13468 11396
rect 13468 11302 13524 11340
rect 13692 11282 13748 12684
rect 14028 12674 14084 12684
rect 14252 11508 14308 11518
rect 14252 11414 14308 11452
rect 13692 11230 13694 11282
rect 13746 11230 13748 11282
rect 13020 8990 13022 9042
rect 13074 8990 13076 9042
rect 13020 8372 13076 8990
rect 13580 10610 13636 10622
rect 13580 10558 13582 10610
rect 13634 10558 13636 10610
rect 13580 9044 13636 10558
rect 13692 9716 13748 11230
rect 13804 11284 13860 11294
rect 13804 9828 13860 11228
rect 14252 10836 14308 10846
rect 14140 9828 14196 9838
rect 13804 9826 14196 9828
rect 13804 9774 14142 9826
rect 14194 9774 14196 9826
rect 13804 9772 14196 9774
rect 14140 9762 14196 9772
rect 13692 9650 13748 9660
rect 14252 9266 14308 10780
rect 14364 10050 14420 12798
rect 14588 12068 14644 12078
rect 14588 11974 14644 12012
rect 15036 11956 15092 13022
rect 15036 11890 15092 11900
rect 15260 12962 15316 12974
rect 15260 12910 15262 12962
rect 15314 12910 15316 12962
rect 15260 12178 15316 12910
rect 15260 12126 15262 12178
rect 15314 12126 15316 12178
rect 14364 9998 14366 10050
rect 14418 9998 14420 10050
rect 14364 9986 14420 9998
rect 14700 11396 14756 11406
rect 14476 9716 14532 9726
rect 14476 9622 14532 9660
rect 14700 9714 14756 11340
rect 15036 10836 15092 10846
rect 15260 10836 15316 12126
rect 15372 11508 15428 11518
rect 15484 11508 15540 13806
rect 15596 13524 15652 13534
rect 15596 13522 15988 13524
rect 15596 13470 15598 13522
rect 15650 13470 15988 13522
rect 15596 13468 15988 13470
rect 15596 13458 15652 13468
rect 15932 13074 15988 13468
rect 16380 13076 16436 14478
rect 16604 14530 16660 15092
rect 16604 14478 16606 14530
rect 16658 14478 16660 14530
rect 16604 14466 16660 14478
rect 17612 13970 17668 15092
rect 17836 14642 17892 18286
rect 18620 17668 18676 20862
rect 18956 20020 19012 22988
rect 19068 22372 19124 22382
rect 19068 22278 19124 22316
rect 19068 21588 19124 21598
rect 19068 20802 19124 21532
rect 19180 21476 19236 21486
rect 19180 21382 19236 21420
rect 19068 20750 19070 20802
rect 19122 20750 19124 20802
rect 19068 20738 19124 20750
rect 19292 20356 19348 23772
rect 19404 23762 19460 23772
rect 19516 23716 19572 23726
rect 19516 23622 19572 23660
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 20412 23044 20468 23996
rect 20524 23714 20580 23726
rect 20524 23662 20526 23714
rect 20578 23662 20580 23714
rect 20524 23268 20580 23662
rect 20748 23716 20804 26124
rect 22876 26178 23044 26180
rect 22876 26126 22990 26178
rect 23042 26126 23044 26178
rect 22876 26124 23044 26126
rect 22876 25282 22932 26124
rect 22988 26114 23044 26124
rect 22988 25732 23044 25742
rect 22988 25638 23044 25676
rect 23212 25730 23268 26460
rect 23324 26292 23380 28028
rect 23548 28084 23604 28094
rect 23436 27300 23492 27310
rect 23436 26852 23492 27244
rect 23548 27076 23604 28028
rect 23660 27970 23716 27982
rect 23660 27918 23662 27970
rect 23714 27918 23716 27970
rect 23660 27636 23716 27918
rect 24108 27970 24164 27982
rect 24108 27918 24110 27970
rect 24162 27918 24164 27970
rect 23660 27570 23716 27580
rect 23884 27858 23940 27870
rect 23884 27806 23886 27858
rect 23938 27806 23940 27858
rect 23548 26908 23604 27020
rect 23548 26852 23716 26908
rect 23436 26786 23492 26796
rect 23324 26226 23380 26236
rect 23660 26404 23716 26852
rect 23884 26628 23940 27806
rect 24108 26908 24164 27918
rect 24220 27858 24276 27870
rect 24220 27806 24222 27858
rect 24274 27806 24276 27858
rect 24220 27636 24276 27806
rect 24220 27570 24276 27580
rect 24108 26852 24276 26908
rect 23884 26562 23940 26572
rect 23660 26348 24164 26404
rect 23660 26290 23716 26348
rect 23660 26238 23662 26290
rect 23714 26238 23716 26290
rect 23660 26226 23716 26238
rect 23212 25678 23214 25730
rect 23266 25678 23268 25730
rect 23212 25666 23268 25678
rect 23660 26068 23716 26078
rect 23660 25506 23716 26012
rect 23884 25956 23940 25966
rect 23772 25900 23884 25956
rect 23772 25730 23828 25900
rect 23884 25890 23940 25900
rect 23772 25678 23774 25730
rect 23826 25678 23828 25730
rect 23772 25666 23828 25678
rect 23660 25454 23662 25506
rect 23714 25454 23716 25506
rect 23660 25442 23716 25454
rect 24108 25508 24164 26348
rect 24220 26180 24276 26852
rect 24220 26086 24276 26124
rect 24332 26068 24388 30716
rect 24444 30212 24500 30940
rect 24444 30146 24500 30156
rect 24556 30210 24612 30222
rect 24556 30158 24558 30210
rect 24610 30158 24612 30210
rect 24556 27076 24612 30158
rect 24668 29652 24724 30940
rect 25228 29988 25284 29998
rect 25228 29894 25284 29932
rect 25564 29986 25620 29998
rect 25564 29934 25566 29986
rect 25618 29934 25620 29986
rect 24780 29652 24836 29662
rect 24668 29650 24836 29652
rect 24668 29598 24782 29650
rect 24834 29598 24836 29650
rect 24668 29596 24836 29598
rect 24780 29586 24836 29596
rect 25452 29652 25508 29662
rect 25452 29558 25508 29596
rect 25564 29428 25620 29934
rect 25340 29372 25620 29428
rect 25116 29092 25172 29102
rect 24668 28084 24724 28094
rect 24668 27746 24724 28028
rect 24668 27694 24670 27746
rect 24722 27694 24724 27746
rect 24668 27412 24724 27694
rect 24668 27346 24724 27356
rect 25004 27188 25060 27198
rect 25004 27094 25060 27132
rect 24556 27010 24612 27020
rect 25116 26964 25172 29036
rect 25116 26290 25172 26908
rect 25116 26238 25118 26290
rect 25170 26238 25172 26290
rect 24332 26002 24388 26012
rect 24892 26180 24948 26190
rect 24444 25956 24500 25966
rect 24220 25508 24276 25518
rect 24108 25506 24388 25508
rect 24108 25454 24222 25506
rect 24274 25454 24388 25506
rect 24108 25452 24388 25454
rect 24220 25442 24276 25452
rect 23548 25396 23604 25406
rect 22876 25230 22878 25282
rect 22930 25230 22932 25282
rect 22876 25218 22932 25230
rect 23212 25284 23268 25294
rect 20860 24948 20916 24958
rect 21644 24948 21700 24958
rect 20860 24946 21140 24948
rect 20860 24894 20862 24946
rect 20914 24894 21140 24946
rect 20860 24892 21140 24894
rect 20860 24882 20916 24892
rect 20860 24722 20916 24734
rect 20860 24670 20862 24722
rect 20914 24670 20916 24722
rect 20860 23940 20916 24670
rect 20860 23874 20916 23884
rect 20748 23660 21028 23716
rect 20524 23212 20916 23268
rect 20860 23154 20916 23212
rect 20860 23102 20862 23154
rect 20914 23102 20916 23154
rect 20412 22978 20468 22988
rect 20524 23042 20580 23054
rect 20524 22990 20526 23042
rect 20578 22990 20580 23042
rect 20412 22260 20468 22270
rect 20524 22260 20580 22990
rect 20412 22258 20580 22260
rect 20412 22206 20414 22258
rect 20466 22206 20580 22258
rect 20412 22204 20580 22206
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 20300 21700 20356 21710
rect 20300 21586 20356 21644
rect 20300 21534 20302 21586
rect 20354 21534 20356 21586
rect 19404 20804 19460 20814
rect 19404 20710 19460 20748
rect 18956 19926 19012 19964
rect 19068 20300 19348 20356
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 19068 19236 19124 20300
rect 19628 20244 19684 20254
rect 19292 20132 19348 20142
rect 19292 20038 19348 20076
rect 19628 20130 19684 20188
rect 20300 20244 20356 21534
rect 20412 21588 20468 22204
rect 20860 21812 20916 23102
rect 20860 21746 20916 21756
rect 20412 21522 20468 21532
rect 20300 20178 20356 20188
rect 19628 20078 19630 20130
rect 19682 20078 19684 20130
rect 19628 20066 19684 20078
rect 20076 20132 20132 20142
rect 20076 20038 20132 20076
rect 20412 20130 20468 20142
rect 20412 20078 20414 20130
rect 20466 20078 20468 20130
rect 20412 19908 20468 20078
rect 20412 19842 20468 19852
rect 20972 19572 21028 23660
rect 21084 20244 21140 24892
rect 21644 24854 21700 24892
rect 22204 24948 22260 24958
rect 22204 24854 22260 24892
rect 21196 24724 21252 24734
rect 21420 24724 21476 24734
rect 21196 24722 21476 24724
rect 21196 24670 21198 24722
rect 21250 24670 21422 24722
rect 21474 24670 21476 24722
rect 21196 24668 21476 24670
rect 21196 24658 21252 24668
rect 21420 24658 21476 24668
rect 21756 24722 21812 24734
rect 21756 24670 21758 24722
rect 21810 24670 21812 24722
rect 21756 23268 21812 24670
rect 23212 23828 23268 25228
rect 23212 23762 23268 23772
rect 23324 24948 23380 24958
rect 23324 23826 23380 24892
rect 23548 24164 23604 25340
rect 24108 24948 24164 24958
rect 24108 24854 24164 24892
rect 23660 24610 23716 24622
rect 23660 24558 23662 24610
rect 23714 24558 23716 24610
rect 23660 24500 23716 24558
rect 23660 24434 23716 24444
rect 24220 24500 24276 24510
rect 23548 24098 23604 24108
rect 24108 24388 24164 24398
rect 23996 23938 24052 23950
rect 23996 23886 23998 23938
rect 24050 23886 24052 23938
rect 23324 23774 23326 23826
rect 23378 23774 23380 23826
rect 23324 23762 23380 23774
rect 23436 23826 23492 23838
rect 23436 23774 23438 23826
rect 23490 23774 23492 23826
rect 22540 23716 22596 23726
rect 22428 23660 22540 23716
rect 22316 23380 22372 23390
rect 22316 23286 22372 23324
rect 21420 23212 21812 23268
rect 21308 23156 21364 23166
rect 21308 23062 21364 23100
rect 21308 21812 21364 21822
rect 21420 21812 21476 23212
rect 21980 23156 22036 23166
rect 21980 23062 22036 23100
rect 21756 23044 21812 23054
rect 21756 22950 21812 22988
rect 21868 22372 21924 22382
rect 21868 22278 21924 22316
rect 22092 22370 22148 22382
rect 22092 22318 22094 22370
rect 22146 22318 22148 22370
rect 21532 22148 21588 22158
rect 22092 22148 22148 22318
rect 22428 22260 22484 23660
rect 22540 23622 22596 23660
rect 22876 23716 22932 23726
rect 22876 23714 23044 23716
rect 22876 23662 22878 23714
rect 22930 23662 23044 23714
rect 22876 23660 23044 23662
rect 22876 23650 22932 23660
rect 22652 23212 22932 23268
rect 22540 23156 22596 23166
rect 22540 23062 22596 23100
rect 22652 23044 22708 23212
rect 22876 23154 22932 23212
rect 22876 23102 22878 23154
rect 22930 23102 22932 23154
rect 22876 23090 22932 23102
rect 22540 22596 22596 22606
rect 22652 22596 22708 22988
rect 22540 22594 22708 22596
rect 22540 22542 22542 22594
rect 22594 22542 22708 22594
rect 22540 22540 22708 22542
rect 22764 23042 22820 23054
rect 22764 22990 22766 23042
rect 22818 22990 22820 23042
rect 22540 22530 22596 22540
rect 22652 22372 22708 22382
rect 22652 22278 22708 22316
rect 22540 22260 22596 22270
rect 22428 22258 22596 22260
rect 22428 22206 22542 22258
rect 22594 22206 22596 22258
rect 22428 22204 22596 22206
rect 22540 22194 22596 22204
rect 21532 22146 21700 22148
rect 21532 22094 21534 22146
rect 21586 22094 21700 22146
rect 21532 22092 21700 22094
rect 21532 22082 21588 22092
rect 21364 21756 21476 21812
rect 21308 21586 21364 21756
rect 21308 21534 21310 21586
rect 21362 21534 21364 21586
rect 21308 21522 21364 21534
rect 21084 20178 21140 20188
rect 21308 20690 21364 20702
rect 21308 20638 21310 20690
rect 21362 20638 21364 20690
rect 21196 20132 21252 20142
rect 21308 20132 21364 20638
rect 21196 20130 21364 20132
rect 21196 20078 21198 20130
rect 21250 20078 21364 20130
rect 21196 20076 21364 20078
rect 21196 20066 21252 20076
rect 20972 19506 21028 19516
rect 21644 20018 21700 22092
rect 22092 22082 22148 22092
rect 21756 21588 21812 21598
rect 21756 21494 21812 21532
rect 21644 19966 21646 20018
rect 21698 19966 21700 20018
rect 19628 19346 19684 19358
rect 19628 19294 19630 19346
rect 19682 19294 19684 19346
rect 18732 19180 19124 19236
rect 18732 19122 18788 19180
rect 18732 19070 18734 19122
rect 18786 19070 18788 19122
rect 18732 19058 18788 19070
rect 19068 18340 19124 19180
rect 19516 19236 19572 19246
rect 19516 19142 19572 19180
rect 19292 18452 19348 18462
rect 19068 18274 19124 18284
rect 19180 18450 19348 18452
rect 19180 18398 19294 18450
rect 19346 18398 19348 18450
rect 19180 18396 19348 18398
rect 19180 17668 19236 18396
rect 19292 18386 19348 18396
rect 19628 18452 19684 19294
rect 20524 19348 20580 19358
rect 20524 19234 20580 19292
rect 21420 19346 21476 19358
rect 21420 19294 21422 19346
rect 21474 19294 21476 19346
rect 20524 19182 20526 19234
rect 20578 19182 20580 19234
rect 19740 19124 19796 19134
rect 19740 19030 19796 19068
rect 20412 19122 20468 19134
rect 20412 19070 20414 19122
rect 20466 19070 20468 19122
rect 20412 19012 20468 19070
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19628 18386 19684 18396
rect 20300 18340 20356 18350
rect 18172 17666 18676 17668
rect 18172 17614 18622 17666
rect 18674 17614 18676 17666
rect 18172 17612 18676 17614
rect 18172 16882 18228 17612
rect 18620 17602 18676 17612
rect 18844 17666 19236 17668
rect 18844 17614 19182 17666
rect 19234 17614 19236 17666
rect 18844 17612 19236 17614
rect 18844 16884 18900 17612
rect 19180 17602 19236 17612
rect 19292 17668 19348 17678
rect 19628 17668 19684 17678
rect 19292 17666 19684 17668
rect 19292 17614 19294 17666
rect 19346 17614 19630 17666
rect 19682 17614 19684 17666
rect 19292 17612 19684 17614
rect 19292 17602 19348 17612
rect 19628 17602 19684 17612
rect 19740 17554 19796 17566
rect 19740 17502 19742 17554
rect 19794 17502 19796 17554
rect 19740 17444 19796 17502
rect 19628 17388 19796 17444
rect 19516 16994 19572 17006
rect 19516 16942 19518 16994
rect 19570 16942 19572 16994
rect 18172 16830 18174 16882
rect 18226 16830 18228 16882
rect 18172 16818 18228 16830
rect 18284 16882 18900 16884
rect 18284 16830 18846 16882
rect 18898 16830 18900 16882
rect 18284 16828 18900 16830
rect 18284 16322 18340 16828
rect 18844 16818 18900 16828
rect 19180 16882 19236 16894
rect 19180 16830 19182 16882
rect 19234 16830 19236 16882
rect 18284 16270 18286 16322
rect 18338 16270 18340 16322
rect 18284 16258 18340 16270
rect 19180 16322 19236 16830
rect 19180 16270 19182 16322
rect 19234 16270 19236 16322
rect 19180 16258 19236 16270
rect 18956 16212 19012 16222
rect 18956 16118 19012 16156
rect 18844 16100 18900 16110
rect 18844 16006 18900 16044
rect 19180 16098 19236 16110
rect 19180 16046 19182 16098
rect 19234 16046 19236 16098
rect 19180 15988 19236 16046
rect 19180 15922 19236 15932
rect 19404 16100 19460 16110
rect 19404 15426 19460 16044
rect 19404 15374 19406 15426
rect 19458 15374 19460 15426
rect 19404 15362 19460 15374
rect 19292 15316 19348 15326
rect 18844 15202 18900 15214
rect 18844 15150 18846 15202
rect 18898 15150 18900 15202
rect 17948 14756 18004 14766
rect 17948 14662 18004 14700
rect 18844 14756 18900 15150
rect 18900 14700 19012 14756
rect 18844 14690 18900 14700
rect 17836 14590 17838 14642
rect 17890 14590 17892 14642
rect 17836 14578 17892 14590
rect 17724 14532 17780 14542
rect 17724 14438 17780 14476
rect 17612 13918 17614 13970
rect 17666 13918 17668 13970
rect 17612 13906 17668 13918
rect 18060 13636 18116 13646
rect 15932 13022 15934 13074
rect 15986 13022 15988 13074
rect 15932 12178 15988 13022
rect 15932 12126 15934 12178
rect 15986 12126 15988 12178
rect 15932 12114 15988 12126
rect 16044 13020 16436 13076
rect 17948 13634 18116 13636
rect 17948 13582 18062 13634
rect 18114 13582 18116 13634
rect 17948 13580 18116 13582
rect 15428 11452 15540 11508
rect 15372 11414 15428 11452
rect 15484 11172 15540 11452
rect 15708 11396 15764 11406
rect 16044 11396 16100 13020
rect 17388 12962 17444 12974
rect 17388 12910 17390 12962
rect 17442 12910 17444 12962
rect 16492 12850 16548 12862
rect 16492 12798 16494 12850
rect 16546 12798 16548 12850
rect 16492 12292 16548 12798
rect 16492 12198 16548 12236
rect 15708 11394 16100 11396
rect 15708 11342 15710 11394
rect 15762 11342 16100 11394
rect 15708 11340 16100 11342
rect 16604 11396 16660 11406
rect 15484 11116 15652 11172
rect 15092 10780 15316 10836
rect 15036 10770 15092 10780
rect 14924 10724 14980 10734
rect 14924 10630 14980 10668
rect 15372 10722 15428 10734
rect 15372 10670 15374 10722
rect 15426 10670 15428 10722
rect 14700 9662 14702 9714
rect 14754 9662 14756 9714
rect 14700 9650 14756 9662
rect 15148 9828 15204 9838
rect 14252 9214 14254 9266
rect 14306 9214 14308 9266
rect 14252 9202 14308 9214
rect 15148 9156 15204 9772
rect 15372 9828 15428 10670
rect 15596 10610 15652 11116
rect 15596 10558 15598 10610
rect 15650 10558 15652 10610
rect 15596 10546 15652 10558
rect 15708 10498 15764 11340
rect 16604 11282 16660 11340
rect 17388 11396 17444 12910
rect 17388 11330 17444 11340
rect 17724 11954 17780 11966
rect 17724 11902 17726 11954
rect 17778 11902 17780 11954
rect 16604 11230 16606 11282
rect 16658 11230 16660 11282
rect 16604 10724 16660 11230
rect 16604 10610 16660 10668
rect 16604 10558 16606 10610
rect 16658 10558 16660 10610
rect 16604 10546 16660 10558
rect 17052 11170 17108 11182
rect 17052 11118 17054 11170
rect 17106 11118 17108 11170
rect 17052 10612 17108 11118
rect 17724 10612 17780 11902
rect 17836 11956 17892 11966
rect 17836 11862 17892 11900
rect 17948 11620 18004 13580
rect 18060 13570 18116 13580
rect 18956 12962 19012 14700
rect 18956 12910 18958 12962
rect 19010 12910 19012 12962
rect 18956 12898 19012 12910
rect 19292 14642 19348 15260
rect 19292 14590 19294 14642
rect 19346 14590 19348 14642
rect 18060 12852 18116 12862
rect 18732 12852 18788 12862
rect 18060 12758 18116 12796
rect 18172 12850 18788 12852
rect 18172 12798 18734 12850
rect 18786 12798 18788 12850
rect 18172 12796 18788 12798
rect 17836 11564 18004 11620
rect 18060 12292 18116 12302
rect 18060 11954 18116 12236
rect 18172 12290 18228 12796
rect 18732 12786 18788 12796
rect 19292 12852 19348 14590
rect 19292 12758 19348 12796
rect 19516 14530 19572 16942
rect 19516 14478 19518 14530
rect 19570 14478 19572 14530
rect 19180 12738 19236 12750
rect 19180 12686 19182 12738
rect 19234 12686 19236 12738
rect 18172 12238 18174 12290
rect 18226 12238 18228 12290
rect 18172 12226 18228 12238
rect 18956 12292 19012 12302
rect 18956 12198 19012 12236
rect 19180 12178 19236 12686
rect 19180 12126 19182 12178
rect 19234 12126 19236 12178
rect 19180 12114 19236 12126
rect 19404 12740 19460 12750
rect 18060 11902 18062 11954
rect 18114 11902 18116 11954
rect 17836 11060 17892 11564
rect 18060 11508 18116 11902
rect 18508 11956 18564 11966
rect 18284 11508 18340 11518
rect 18060 11506 18340 11508
rect 18060 11454 18286 11506
rect 18338 11454 18340 11506
rect 18060 11452 18340 11454
rect 17948 11394 18004 11406
rect 17948 11342 17950 11394
rect 18002 11342 18004 11394
rect 17948 11284 18004 11342
rect 17948 11218 18004 11228
rect 18060 11282 18116 11294
rect 18060 11230 18062 11282
rect 18114 11230 18116 11282
rect 18060 11060 18116 11230
rect 17836 11004 18116 11060
rect 17836 10612 17892 10622
rect 17724 10556 17836 10612
rect 17052 10546 17108 10556
rect 17836 10518 17892 10556
rect 15708 10446 15710 10498
rect 15762 10446 15764 10498
rect 15708 10434 15764 10446
rect 15148 9062 15204 9100
rect 15260 9268 15316 9278
rect 13804 9044 13860 9054
rect 14812 9044 14868 9054
rect 13580 9042 13860 9044
rect 13580 8990 13806 9042
rect 13858 8990 13860 9042
rect 13580 8988 13860 8990
rect 13020 8306 13076 8316
rect 13580 8260 13636 8270
rect 13692 8260 13748 8988
rect 13804 8978 13860 8988
rect 14588 9042 14868 9044
rect 14588 8990 14814 9042
rect 14866 8990 14868 9042
rect 14588 8988 14868 8990
rect 13636 8204 13748 8260
rect 13804 8372 13860 8382
rect 13804 8258 13860 8316
rect 14476 8372 14532 8382
rect 14588 8372 14644 8988
rect 14812 8978 14868 8988
rect 14476 8370 14644 8372
rect 14476 8318 14478 8370
rect 14530 8318 14644 8370
rect 14476 8316 14644 8318
rect 14476 8306 14532 8316
rect 13804 8206 13806 8258
rect 13858 8206 13860 8258
rect 13580 8166 13636 8204
rect 13804 8194 13860 8206
rect 15260 8258 15316 9212
rect 15260 8206 15262 8258
rect 15314 8206 15316 8258
rect 15260 8194 15316 8206
rect 15372 8258 15428 9772
rect 16268 9826 16324 9838
rect 16268 9774 16270 9826
rect 16322 9774 16324 9826
rect 15484 9716 15540 9726
rect 15484 9156 15540 9660
rect 15820 9716 15876 9726
rect 15820 9268 15876 9660
rect 15820 9174 15876 9212
rect 15484 9154 15652 9156
rect 15484 9102 15486 9154
rect 15538 9102 15652 9154
rect 15484 9100 15652 9102
rect 15484 9090 15540 9100
rect 15372 8206 15374 8258
rect 15426 8206 15428 8258
rect 15372 8194 15428 8206
rect 12796 8094 12798 8146
rect 12850 8094 12852 8146
rect 12796 8082 12852 8094
rect 15484 8148 15540 8158
rect 11900 7924 11956 7934
rect 11788 7588 11844 7598
rect 11788 7494 11844 7532
rect 11900 7586 11956 7868
rect 11900 7534 11902 7586
rect 11954 7534 11956 7586
rect 11900 7522 11956 7534
rect 12348 7588 12404 7598
rect 12348 7494 12404 7532
rect 12684 7588 12740 7980
rect 13020 8036 13076 8046
rect 13020 7942 13076 7980
rect 14140 8036 14196 8046
rect 12796 7924 12852 7934
rect 12796 7698 12852 7868
rect 14140 7700 14196 7980
rect 12796 7646 12798 7698
rect 12850 7646 12852 7698
rect 12796 7634 12852 7646
rect 14028 7698 14196 7700
rect 14028 7646 14142 7698
rect 14194 7646 14196 7698
rect 14028 7644 14196 7646
rect 12684 7522 12740 7532
rect 12236 7252 12292 7262
rect 12236 7158 12292 7196
rect 13916 7250 13972 7262
rect 13916 7198 13918 7250
rect 13970 7198 13972 7250
rect 11676 6972 11844 7028
rect 11676 6804 11732 6814
rect 11676 6710 11732 6748
rect 11564 6526 11566 6578
rect 11618 6526 11620 6578
rect 11564 6020 11620 6526
rect 11788 6468 11844 6972
rect 13132 6804 13188 6814
rect 12460 6692 12516 6702
rect 12460 6598 12516 6636
rect 12348 6580 12404 6590
rect 12348 6486 12404 6524
rect 11788 6402 11844 6412
rect 12124 6466 12180 6478
rect 12124 6414 12126 6466
rect 12178 6414 12180 6466
rect 12124 6132 12180 6414
rect 12572 6468 12628 6478
rect 12628 6412 12964 6468
rect 12572 6374 12628 6412
rect 12236 6132 12292 6142
rect 12124 6130 12292 6132
rect 12124 6078 12238 6130
rect 12290 6078 12292 6130
rect 12124 6076 12292 6078
rect 12236 6066 12292 6076
rect 11564 5954 11620 5964
rect 12348 6020 12404 6030
rect 12348 5926 12404 5964
rect 12908 5906 12964 6412
rect 12908 5854 12910 5906
rect 12962 5854 12964 5906
rect 12908 5842 12964 5854
rect 13132 5906 13188 6748
rect 13580 6804 13636 6814
rect 13580 6710 13636 6748
rect 13804 6020 13860 6030
rect 13916 6020 13972 7198
rect 14028 6690 14084 7644
rect 14140 7634 14196 7644
rect 14924 7924 14980 7934
rect 14924 7698 14980 7868
rect 14924 7646 14926 7698
rect 14978 7646 14980 7698
rect 14924 7476 14980 7646
rect 15372 7700 15428 7710
rect 15372 7606 15428 7644
rect 15260 7476 15316 7486
rect 14924 7474 15316 7476
rect 14924 7422 15262 7474
rect 15314 7422 15316 7474
rect 14924 7420 15316 7422
rect 14252 7364 14308 7374
rect 14252 7270 14308 7308
rect 14028 6638 14030 6690
rect 14082 6638 14084 6690
rect 14028 6626 14084 6638
rect 15148 6690 15204 6702
rect 15148 6638 15150 6690
rect 15202 6638 15204 6690
rect 15148 6468 15204 6638
rect 15148 6402 15204 6412
rect 15260 6356 15316 7420
rect 15484 6914 15540 8092
rect 15596 7812 15652 9100
rect 15932 8932 15988 8942
rect 15932 8370 15988 8876
rect 15932 8318 15934 8370
rect 15986 8318 15988 8370
rect 15932 8306 15988 8318
rect 16268 8148 16324 9774
rect 17052 9828 17108 9838
rect 17052 9734 17108 9772
rect 17948 9828 18004 11004
rect 18284 10612 18340 11452
rect 18284 10546 18340 10556
rect 18508 10610 18564 11900
rect 19292 11508 19348 11518
rect 19404 11508 19460 12684
rect 19516 11956 19572 14478
rect 19628 12964 19684 17388
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 20076 16100 20132 16110
rect 20076 16006 20132 16044
rect 20300 15986 20356 18284
rect 20412 17556 20468 18956
rect 20412 17490 20468 17500
rect 20524 18564 20580 19182
rect 20524 17554 20580 18508
rect 20636 19236 20692 19246
rect 20636 18338 20692 19180
rect 20636 18286 20638 18338
rect 20690 18286 20692 18338
rect 20636 18274 20692 18286
rect 20748 19122 20804 19134
rect 20748 19070 20750 19122
rect 20802 19070 20804 19122
rect 20524 17502 20526 17554
rect 20578 17502 20580 17554
rect 20524 17490 20580 17502
rect 20636 17108 20692 17118
rect 20300 15934 20302 15986
rect 20354 15934 20356 15986
rect 20300 15764 20356 15934
rect 20412 15986 20468 15998
rect 20412 15934 20414 15986
rect 20466 15934 20468 15986
rect 20412 15876 20468 15934
rect 20524 15876 20580 15886
rect 20412 15820 20524 15876
rect 20524 15810 20580 15820
rect 19836 15708 20100 15718
rect 20300 15708 20468 15764
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 20300 15316 20356 15326
rect 20300 15222 20356 15260
rect 20076 14644 20132 14654
rect 20076 14550 20132 14588
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 20412 13076 20468 15708
rect 20636 15538 20692 17052
rect 20748 16996 20804 19070
rect 21420 19124 21476 19294
rect 21644 19234 21700 19966
rect 21644 19182 21646 19234
rect 21698 19182 21700 19234
rect 21644 19170 21700 19182
rect 21756 21362 21812 21374
rect 21756 21310 21758 21362
rect 21810 21310 21812 21362
rect 21756 20802 21812 21310
rect 21756 20750 21758 20802
rect 21810 20750 21812 20802
rect 21420 19058 21476 19068
rect 21756 19124 21812 20750
rect 22204 20802 22260 20814
rect 22204 20750 22206 20802
rect 22258 20750 22260 20802
rect 22204 19236 22260 20750
rect 22764 19684 22820 22990
rect 22876 22372 22932 22382
rect 22988 22372 23044 23660
rect 23100 23714 23156 23726
rect 23100 23662 23102 23714
rect 23154 23662 23156 23714
rect 23100 23154 23156 23662
rect 23436 23380 23492 23774
rect 23436 23314 23492 23324
rect 23100 23102 23102 23154
rect 23154 23102 23156 23154
rect 23100 23090 23156 23102
rect 23548 23044 23604 23054
rect 23436 23042 23604 23044
rect 23436 22990 23550 23042
rect 23602 22990 23604 23042
rect 23436 22988 23604 22990
rect 23212 22372 23268 22382
rect 23436 22372 23492 22988
rect 23548 22978 23604 22988
rect 23772 23044 23828 23054
rect 23996 23044 24052 23886
rect 24108 23378 24164 24332
rect 24220 24162 24276 24444
rect 24220 24110 24222 24162
rect 24274 24110 24276 24162
rect 24220 24098 24276 24110
rect 24332 23940 24388 25452
rect 24444 24948 24500 25900
rect 24892 25618 24948 26124
rect 24892 25566 24894 25618
rect 24946 25566 24948 25618
rect 24892 25554 24948 25566
rect 24444 24882 24500 24892
rect 25116 24948 25172 26238
rect 25116 24882 25172 24892
rect 25340 28196 25396 29372
rect 25676 28756 25732 31052
rect 25788 30770 25844 30782
rect 25788 30718 25790 30770
rect 25842 30718 25844 30770
rect 25788 30324 25844 30718
rect 25788 30258 25844 30268
rect 24444 24052 24500 24062
rect 24444 23958 24500 23996
rect 25116 24052 25172 24062
rect 25340 24052 25396 28140
rect 25452 28700 25676 28756
rect 25452 26908 25508 28700
rect 25676 28690 25732 28700
rect 25788 29426 25844 29438
rect 25788 29374 25790 29426
rect 25842 29374 25844 29426
rect 25788 28980 25844 29374
rect 25900 29316 25956 31612
rect 26012 31444 26068 31454
rect 26012 31108 26068 31388
rect 26012 30994 26068 31052
rect 26012 30942 26014 30994
rect 26066 30942 26068 30994
rect 26012 30930 26068 30942
rect 26012 29540 26068 29550
rect 26012 29446 26068 29484
rect 26236 29428 26292 34076
rect 26684 34066 26740 34078
rect 26796 33572 26852 35252
rect 27132 35252 27188 35262
rect 27020 34130 27076 34142
rect 27020 34078 27022 34130
rect 27074 34078 27076 34130
rect 26684 33516 26852 33572
rect 26908 33908 26964 33918
rect 26572 33012 26628 33022
rect 26572 32786 26628 32956
rect 26684 32900 26740 33516
rect 26684 32834 26740 32844
rect 26796 33346 26852 33358
rect 26796 33294 26798 33346
rect 26850 33294 26852 33346
rect 26572 32734 26574 32786
rect 26626 32734 26628 32786
rect 26572 32722 26628 32734
rect 26348 32564 26404 32574
rect 26348 32562 26516 32564
rect 26348 32510 26350 32562
rect 26402 32510 26516 32562
rect 26348 32508 26516 32510
rect 26348 32498 26404 32508
rect 26348 31778 26404 31790
rect 26348 31726 26350 31778
rect 26402 31726 26404 31778
rect 26348 30322 26404 31726
rect 26460 31780 26516 32508
rect 26572 32116 26628 32126
rect 26572 32002 26628 32060
rect 26572 31950 26574 32002
rect 26626 31950 26628 32002
rect 26572 31938 26628 31950
rect 26572 31780 26628 31790
rect 26460 31778 26628 31780
rect 26460 31726 26574 31778
rect 26626 31726 26628 31778
rect 26460 31724 26628 31726
rect 26572 31218 26628 31724
rect 26572 31166 26574 31218
rect 26626 31166 26628 31218
rect 26572 31108 26628 31166
rect 26572 31042 26628 31052
rect 26796 30884 26852 33294
rect 26908 31218 26964 33852
rect 27020 33796 27076 34078
rect 27020 33730 27076 33740
rect 26908 31166 26910 31218
rect 26962 31166 26964 31218
rect 26908 31154 26964 31166
rect 27020 32450 27076 32462
rect 27020 32398 27022 32450
rect 27074 32398 27076 32450
rect 27020 31556 27076 32398
rect 26348 30270 26350 30322
rect 26402 30270 26404 30322
rect 26348 30212 26404 30270
rect 26348 30146 26404 30156
rect 26684 30828 26796 30884
rect 26348 29428 26404 29438
rect 26236 29426 26404 29428
rect 26236 29374 26350 29426
rect 26402 29374 26404 29426
rect 26236 29372 26404 29374
rect 25900 29260 26292 29316
rect 25564 28084 25620 28094
rect 25564 27990 25620 28028
rect 25788 27972 25844 28924
rect 25788 27906 25844 27916
rect 25676 27860 25732 27870
rect 25676 27766 25732 27804
rect 26124 27858 26180 27870
rect 26124 27806 26126 27858
rect 26178 27806 26180 27858
rect 25564 27636 25620 27646
rect 25564 27634 25956 27636
rect 25564 27582 25566 27634
rect 25618 27582 25956 27634
rect 25564 27580 25956 27582
rect 25564 27570 25620 27580
rect 25676 27412 25732 27422
rect 25676 27076 25732 27356
rect 25900 27076 25956 27580
rect 26012 27524 26068 27534
rect 26124 27524 26180 27806
rect 26068 27468 26180 27524
rect 26012 27458 26068 27468
rect 26012 27076 26068 27086
rect 25900 27074 26068 27076
rect 25900 27022 26014 27074
rect 26066 27022 26068 27074
rect 25900 27020 26068 27022
rect 25676 27010 25732 27020
rect 26012 27010 26068 27020
rect 26236 26908 26292 29260
rect 26348 28644 26404 29372
rect 26572 29428 26628 29438
rect 26572 29334 26628 29372
rect 26460 29316 26516 29326
rect 26460 29222 26516 29260
rect 26348 28578 26404 28588
rect 26684 28642 26740 30828
rect 26796 30818 26852 30828
rect 27020 30324 27076 31500
rect 26796 30268 27076 30324
rect 26796 30210 26852 30268
rect 26796 30158 26798 30210
rect 26850 30158 26852 30210
rect 26796 30146 26852 30158
rect 27020 29986 27076 29998
rect 27020 29934 27022 29986
rect 27074 29934 27076 29986
rect 26796 29540 26852 29550
rect 26796 29446 26852 29484
rect 27020 29316 27076 29934
rect 27132 29988 27188 35196
rect 27244 34804 27300 35308
rect 27244 33012 27300 34748
rect 27356 35140 27412 35150
rect 27356 34354 27412 35084
rect 27356 34302 27358 34354
rect 27410 34302 27412 34354
rect 27356 34290 27412 34302
rect 27244 31444 27300 32956
rect 27468 32788 27524 32798
rect 27468 32450 27524 32732
rect 27468 32398 27470 32450
rect 27522 32398 27524 32450
rect 27468 32338 27524 32398
rect 27468 32286 27470 32338
rect 27522 32286 27524 32338
rect 27468 32274 27524 32286
rect 27580 31780 27636 36428
rect 27692 36260 27748 36270
rect 27692 35810 27748 36204
rect 27692 35758 27694 35810
rect 27746 35758 27748 35810
rect 27692 35746 27748 35758
rect 27916 35364 27972 36428
rect 28140 36260 28196 36270
rect 28140 35922 28196 36204
rect 28476 36036 28532 38612
rect 28812 38164 28868 43372
rect 28924 43426 28980 43484
rect 28924 43374 28926 43426
rect 28978 43374 28980 43426
rect 28924 43362 28980 43374
rect 29036 38668 29092 54796
rect 29148 54786 29204 54796
rect 29708 54852 29764 55246
rect 29708 54786 29764 54796
rect 29820 54738 29876 55412
rect 30268 55412 30324 59200
rect 30940 56980 30996 59200
rect 30940 56924 31444 56980
rect 31276 56196 31332 56206
rect 30716 56194 31332 56196
rect 30716 56142 31278 56194
rect 31330 56142 31332 56194
rect 30716 56140 31332 56142
rect 30604 56082 30660 56094
rect 30604 56030 30606 56082
rect 30658 56030 30660 56082
rect 30268 55410 30548 55412
rect 30268 55358 30270 55410
rect 30322 55358 30548 55410
rect 30268 55356 30548 55358
rect 30268 55346 30324 55356
rect 30492 55298 30548 55356
rect 30492 55246 30494 55298
rect 30546 55246 30548 55298
rect 30492 55234 30548 55246
rect 29820 54686 29822 54738
rect 29874 54686 29876 54738
rect 29820 54674 29876 54686
rect 29148 54628 29204 54638
rect 29148 54534 29204 54572
rect 29484 54628 29540 54638
rect 29484 54626 29764 54628
rect 29484 54574 29486 54626
rect 29538 54574 29764 54626
rect 29484 54572 29764 54574
rect 29484 54562 29540 54572
rect 29708 53284 29764 54572
rect 30156 54626 30212 54638
rect 30156 54574 30158 54626
rect 30210 54574 30212 54626
rect 29932 53508 29988 53518
rect 29932 53414 29988 53452
rect 29708 53228 30100 53284
rect 29148 53172 29204 53182
rect 29148 53078 29204 53116
rect 29708 52836 29764 52846
rect 29708 52742 29764 52780
rect 29708 52276 29764 52286
rect 29708 51380 29764 52220
rect 29820 52162 29876 53228
rect 30044 53170 30100 53228
rect 30044 53118 30046 53170
rect 30098 53118 30100 53170
rect 30044 53106 30100 53118
rect 29820 52110 29822 52162
rect 29874 52110 29876 52162
rect 29820 52098 29876 52110
rect 29932 53060 29988 53070
rect 29932 52164 29988 53004
rect 29932 52070 29988 52108
rect 30044 52164 30100 52174
rect 30156 52164 30212 54574
rect 30604 53956 30660 56030
rect 30604 53890 30660 53900
rect 30268 53732 30324 53742
rect 30716 53732 30772 56140
rect 31276 56130 31332 56140
rect 31388 56084 31444 56924
rect 31612 56308 31668 59200
rect 31612 56242 31668 56252
rect 31500 56084 31556 56094
rect 31388 56082 31556 56084
rect 31388 56030 31502 56082
rect 31554 56030 31556 56082
rect 31388 56028 31556 56030
rect 31388 55468 31444 56028
rect 31500 56018 31556 56028
rect 32172 56082 32228 56094
rect 32172 56030 32174 56082
rect 32226 56030 32228 56082
rect 32172 55468 32228 56030
rect 31276 55412 31444 55468
rect 32060 55412 32228 55468
rect 32284 55412 32340 59200
rect 31276 55410 31332 55412
rect 31276 55358 31278 55410
rect 31330 55358 31332 55410
rect 31276 55346 31332 55358
rect 30828 55076 30884 55086
rect 31724 55076 31780 55086
rect 30828 55074 30996 55076
rect 30828 55022 30830 55074
rect 30882 55022 30996 55074
rect 30828 55020 30996 55022
rect 30828 55010 30884 55020
rect 30268 53730 30772 53732
rect 30268 53678 30270 53730
rect 30322 53678 30718 53730
rect 30770 53678 30772 53730
rect 30268 53676 30772 53678
rect 30268 53666 30324 53676
rect 30716 53666 30772 53676
rect 30044 52162 30212 52164
rect 30044 52110 30046 52162
rect 30098 52110 30212 52162
rect 30044 52108 30212 52110
rect 30044 52098 30100 52108
rect 30156 52052 30212 52108
rect 30268 53508 30324 53518
rect 30268 52276 30324 53452
rect 30940 53060 30996 55020
rect 31612 55074 31780 55076
rect 31612 55022 31726 55074
rect 31778 55022 31780 55074
rect 31612 55020 31780 55022
rect 31276 54404 31332 54414
rect 31164 53620 31220 53630
rect 31164 53526 31220 53564
rect 30268 52162 30324 52220
rect 30268 52110 30270 52162
rect 30322 52110 30324 52162
rect 30268 52098 30324 52110
rect 30380 53004 30996 53060
rect 30156 51986 30212 51996
rect 30380 51490 30436 53004
rect 30492 52836 30548 52846
rect 30492 52276 30548 52780
rect 30604 52834 30660 52846
rect 30604 52782 30606 52834
rect 30658 52782 30660 52834
rect 30604 52500 30660 52782
rect 30604 52434 30660 52444
rect 30492 52220 30660 52276
rect 30380 51438 30382 51490
rect 30434 51438 30436 51490
rect 30380 51426 30436 51438
rect 30492 52052 30548 52062
rect 30492 51490 30548 51996
rect 30604 51716 30660 52220
rect 30940 52162 30996 53004
rect 31164 52500 31220 52510
rect 30940 52110 30942 52162
rect 30994 52110 30996 52162
rect 30940 52098 30996 52110
rect 31052 52164 31108 52174
rect 30716 51940 30772 51950
rect 30716 51938 30884 51940
rect 30716 51886 30718 51938
rect 30770 51886 30884 51938
rect 30716 51884 30884 51886
rect 30716 51874 30772 51884
rect 30604 51660 30772 51716
rect 30492 51438 30494 51490
rect 30546 51438 30548 51490
rect 29932 51380 29988 51390
rect 29708 51378 29988 51380
rect 29708 51326 29934 51378
rect 29986 51326 29988 51378
rect 29708 51324 29988 51326
rect 29932 51314 29988 51324
rect 29708 51154 29764 51166
rect 29708 51102 29710 51154
rect 29762 51102 29764 51154
rect 29708 49812 29764 51102
rect 30492 50594 30548 51438
rect 30716 51378 30772 51660
rect 30716 51326 30718 51378
rect 30770 51326 30772 51378
rect 30716 51314 30772 51326
rect 30492 50542 30494 50594
rect 30546 50542 30548 50594
rect 30380 50036 30436 50046
rect 30156 49980 30380 50036
rect 29372 49698 29428 49710
rect 29372 49646 29374 49698
rect 29426 49646 29428 49698
rect 29372 49364 29428 49646
rect 29372 49298 29428 49308
rect 29708 49028 29764 49756
rect 29820 49810 29876 49822
rect 30156 49812 30212 49980
rect 30380 49970 30436 49980
rect 29820 49758 29822 49810
rect 29874 49758 29876 49810
rect 29820 49252 29876 49758
rect 30044 49810 30212 49812
rect 30044 49758 30158 49810
rect 30210 49758 30212 49810
rect 30044 49756 30212 49758
rect 29820 49186 29876 49196
rect 29932 49700 29988 49710
rect 29820 49028 29876 49038
rect 29708 49026 29876 49028
rect 29708 48974 29822 49026
rect 29874 48974 29876 49026
rect 29708 48972 29876 48974
rect 29596 48916 29652 48926
rect 29596 46676 29652 48860
rect 29708 48354 29764 48972
rect 29820 48962 29876 48972
rect 29708 48302 29710 48354
rect 29762 48302 29764 48354
rect 29708 48290 29764 48302
rect 29820 48130 29876 48142
rect 29820 48078 29822 48130
rect 29874 48078 29876 48130
rect 29260 46674 29652 46676
rect 29260 46622 29598 46674
rect 29650 46622 29652 46674
rect 29260 46620 29652 46622
rect 29260 46002 29316 46620
rect 29596 46610 29652 46620
rect 29708 46788 29764 46798
rect 29820 46788 29876 48078
rect 29708 46786 29876 46788
rect 29708 46734 29710 46786
rect 29762 46734 29876 46786
rect 29708 46732 29876 46734
rect 29260 45950 29262 46002
rect 29314 45950 29316 46002
rect 29260 45938 29316 45950
rect 29372 46340 29428 46350
rect 29148 43652 29204 43662
rect 29148 42644 29204 43596
rect 29148 41858 29204 42588
rect 29260 42980 29316 42990
rect 29260 41970 29316 42924
rect 29260 41918 29262 41970
rect 29314 41918 29316 41970
rect 29260 41906 29316 41918
rect 29148 41806 29150 41858
rect 29202 41806 29204 41858
rect 29148 41794 29204 41806
rect 29148 40962 29204 40974
rect 29148 40910 29150 40962
rect 29202 40910 29204 40962
rect 29148 40516 29204 40910
rect 29148 40450 29204 40460
rect 29260 40290 29316 40302
rect 29260 40238 29262 40290
rect 29314 40238 29316 40290
rect 29260 39844 29316 40238
rect 29260 39778 29316 39788
rect 28588 38108 28812 38164
rect 28588 36594 28644 38108
rect 28812 38098 28868 38108
rect 28924 38612 29092 38668
rect 28588 36542 28590 36594
rect 28642 36542 28644 36594
rect 28588 36530 28644 36542
rect 28924 36148 28980 38612
rect 29036 37156 29092 37166
rect 29036 37154 29316 37156
rect 29036 37102 29038 37154
rect 29090 37102 29316 37154
rect 29036 37100 29316 37102
rect 29036 37090 29092 37100
rect 29260 36594 29316 37100
rect 29260 36542 29262 36594
rect 29314 36542 29316 36594
rect 29260 36530 29316 36542
rect 29372 36484 29428 46284
rect 29708 45778 29764 46732
rect 29708 45726 29710 45778
rect 29762 45726 29764 45778
rect 29708 45714 29764 45726
rect 29932 43708 29988 49644
rect 30044 48242 30100 49756
rect 30156 49746 30212 49756
rect 30380 49812 30436 49822
rect 30380 49718 30436 49756
rect 30492 49588 30548 50542
rect 30604 51268 30660 51278
rect 30604 49810 30660 51212
rect 30604 49758 30606 49810
rect 30658 49758 30660 49810
rect 30604 49746 30660 49758
rect 30828 50036 30884 51884
rect 31052 51602 31108 52108
rect 31052 51550 31054 51602
rect 31106 51550 31108 51602
rect 31052 51538 31108 51550
rect 31052 50596 31108 50606
rect 31052 50502 31108 50540
rect 31164 50484 31220 52444
rect 31164 50418 31220 50428
rect 30492 49532 30660 49588
rect 30604 48914 30660 49532
rect 30604 48862 30606 48914
rect 30658 48862 30660 48914
rect 30604 48850 30660 48862
rect 30044 48190 30046 48242
rect 30098 48190 30100 48242
rect 30044 48178 30100 48190
rect 30156 48802 30212 48814
rect 30156 48750 30158 48802
rect 30210 48750 30212 48802
rect 30156 48020 30212 48750
rect 30828 48468 30884 49980
rect 31276 49812 31332 54348
rect 31612 53732 31668 55020
rect 31724 55010 31780 55020
rect 31612 53666 31668 53676
rect 31724 54628 31780 54638
rect 31612 53060 31668 53070
rect 31500 53004 31612 53060
rect 31724 53060 31780 54572
rect 31836 54404 31892 54414
rect 32060 54404 32116 55412
rect 32284 55346 32340 55356
rect 32508 55298 32564 55310
rect 32508 55246 32510 55298
rect 32562 55246 32564 55298
rect 31892 54348 32116 54404
rect 32172 55076 32228 55086
rect 32508 55076 32564 55246
rect 32172 55074 32564 55076
rect 32172 55022 32174 55074
rect 32226 55022 32564 55074
rect 32172 55020 32564 55022
rect 31836 54310 31892 54348
rect 31836 53060 31892 53070
rect 31724 53058 31892 53060
rect 31724 53006 31838 53058
rect 31890 53006 31892 53058
rect 31724 53004 31892 53006
rect 31388 52946 31444 52958
rect 31388 52894 31390 52946
rect 31442 52894 31444 52946
rect 31388 52836 31444 52894
rect 31388 52770 31444 52780
rect 31500 52274 31556 53004
rect 31612 52966 31668 53004
rect 31836 52994 31892 53004
rect 31500 52222 31502 52274
rect 31554 52222 31556 52274
rect 31500 52210 31556 52222
rect 32060 52946 32116 52958
rect 32060 52894 32062 52946
rect 32114 52894 32116 52946
rect 32060 52276 32116 52894
rect 32060 52210 32116 52220
rect 31724 51940 31780 51950
rect 31612 51492 31668 51502
rect 31612 51398 31668 51436
rect 31724 50708 31780 51884
rect 32172 51940 32228 55020
rect 32956 54740 33012 59200
rect 33628 56980 33684 59200
rect 33628 56924 33796 56980
rect 33180 56308 33236 56318
rect 33180 56214 33236 56252
rect 33516 55412 33572 55422
rect 33516 55318 33572 55356
rect 33740 55412 33796 56924
rect 34300 55972 34356 59200
rect 34300 55906 34356 55916
rect 33740 55346 33796 55356
rect 34972 55300 35028 59200
rect 35644 57428 35700 59200
rect 35644 57372 36148 57428
rect 34972 55234 35028 55244
rect 35084 56194 35140 56206
rect 35084 56142 35086 56194
rect 35138 56142 35140 56194
rect 32956 54674 33012 54684
rect 34188 54740 34244 54750
rect 34188 54646 34244 54684
rect 32396 54628 32452 54638
rect 32284 54514 32340 54526
rect 32284 54462 32286 54514
rect 32338 54462 32340 54514
rect 32284 53620 32340 54462
rect 32396 53956 32452 54572
rect 32620 54514 32676 54526
rect 32620 54462 32622 54514
rect 32674 54462 32676 54514
rect 32620 54404 32676 54462
rect 33180 54516 33236 54526
rect 33180 54422 33236 54460
rect 32620 54338 32676 54348
rect 32396 53890 32452 53900
rect 33516 53842 33572 53854
rect 35084 53844 35140 56142
rect 35420 56084 35476 56094
rect 35420 56082 35588 56084
rect 35420 56030 35422 56082
rect 35474 56030 35588 56082
rect 35420 56028 35588 56030
rect 35420 56018 35476 56028
rect 35196 55692 35460 55702
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35196 55626 35460 55636
rect 35532 55468 35588 56028
rect 35532 55412 35812 55468
rect 35532 55346 35588 55356
rect 35644 55298 35700 55310
rect 35644 55246 35646 55298
rect 35698 55246 35700 55298
rect 35420 55188 35476 55198
rect 35420 55186 35588 55188
rect 35420 55134 35422 55186
rect 35474 55134 35588 55186
rect 35420 55132 35588 55134
rect 35420 55122 35476 55132
rect 35196 54124 35460 54134
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35196 54058 35460 54068
rect 33516 53790 33518 53842
rect 33570 53790 33572 53842
rect 32844 53730 32900 53742
rect 32844 53678 32846 53730
rect 32898 53678 32900 53730
rect 32396 53620 32452 53630
rect 32284 53564 32396 53620
rect 32396 52948 32452 53564
rect 32844 53060 32900 53678
rect 32844 52994 32900 53004
rect 33292 53618 33348 53630
rect 33292 53566 33294 53618
rect 33346 53566 33348 53618
rect 32396 52882 32452 52892
rect 32396 52722 32452 52734
rect 32396 52670 32398 52722
rect 32450 52670 32452 52722
rect 32396 52164 32452 52670
rect 32172 51874 32228 51884
rect 32284 52108 32396 52164
rect 30156 47572 30212 47964
rect 30492 48466 30884 48468
rect 30492 48414 30830 48466
rect 30882 48414 30884 48466
rect 30492 48412 30884 48414
rect 30156 47516 30436 47572
rect 30380 47458 30436 47516
rect 30380 47406 30382 47458
rect 30434 47406 30436 47458
rect 30380 47394 30436 47406
rect 30492 47346 30548 48412
rect 30828 48402 30884 48412
rect 30940 49756 31332 49812
rect 31612 50652 31780 50708
rect 32284 51378 32340 52108
rect 32396 52098 32452 52108
rect 32620 52050 32676 52062
rect 32620 51998 32622 52050
rect 32674 51998 32676 52050
rect 32508 51492 32564 51502
rect 32508 51398 32564 51436
rect 32284 51326 32286 51378
rect 32338 51326 32340 51378
rect 30940 47684 30996 49756
rect 31500 49700 31556 49710
rect 31052 49588 31108 49598
rect 31052 49586 31332 49588
rect 31052 49534 31054 49586
rect 31106 49534 31332 49586
rect 31052 49532 31332 49534
rect 31052 49522 31108 49532
rect 31052 49028 31108 49066
rect 31052 48962 31108 48972
rect 31164 48916 31220 48926
rect 31164 48822 31220 48860
rect 31164 48354 31220 48366
rect 31164 48302 31166 48354
rect 31218 48302 31220 48354
rect 31164 48132 31220 48302
rect 31164 48066 31220 48076
rect 30940 47628 31220 47684
rect 30492 47294 30494 47346
rect 30546 47294 30548 47346
rect 30492 47282 30548 47294
rect 30604 47572 30660 47582
rect 29932 43652 30324 43708
rect 29484 41076 29540 41086
rect 29484 41074 29876 41076
rect 29484 41022 29486 41074
rect 29538 41022 29876 41074
rect 29484 41020 29876 41022
rect 29484 41010 29540 41020
rect 29596 40402 29652 40414
rect 29596 40350 29598 40402
rect 29650 40350 29652 40402
rect 29484 39394 29540 39406
rect 29484 39342 29486 39394
rect 29538 39342 29540 39394
rect 29484 39060 29540 39342
rect 29484 37156 29540 39004
rect 29596 37492 29652 40350
rect 29820 39842 29876 41020
rect 29820 39790 29822 39842
rect 29874 39790 29876 39842
rect 29820 39778 29876 39790
rect 30156 39844 30212 39854
rect 30156 39750 30212 39788
rect 30268 38668 30324 43652
rect 30604 43204 30660 47516
rect 31052 47458 31108 47470
rect 31052 47406 31054 47458
rect 31106 47406 31108 47458
rect 30716 47236 30772 47246
rect 31052 47236 31108 47406
rect 30716 47234 31108 47236
rect 30716 47182 30718 47234
rect 30770 47182 31108 47234
rect 30716 47180 31108 47182
rect 30716 47170 30772 47180
rect 30940 46788 30996 46798
rect 30940 45890 30996 46732
rect 31052 46116 31108 47180
rect 31052 46050 31108 46060
rect 30940 45838 30942 45890
rect 30994 45838 30996 45890
rect 30940 45826 30996 45838
rect 31164 44660 31220 47628
rect 31276 47346 31332 49532
rect 31500 49364 31556 49644
rect 31500 49026 31556 49308
rect 31500 48974 31502 49026
rect 31554 48974 31556 49026
rect 31500 48962 31556 48974
rect 31388 47572 31444 47582
rect 31388 47478 31444 47516
rect 31612 47460 31668 50652
rect 31724 50484 31780 50494
rect 31724 48914 31780 50428
rect 32172 50036 32228 50046
rect 31836 49586 31892 49598
rect 31836 49534 31838 49586
rect 31890 49534 31892 49586
rect 31836 49476 31892 49534
rect 31836 49420 32004 49476
rect 31724 48862 31726 48914
rect 31778 48862 31780 48914
rect 31724 47684 31780 48862
rect 31724 47618 31780 47628
rect 31276 47294 31278 47346
rect 31330 47294 31332 47346
rect 31276 47236 31332 47294
rect 31276 47170 31332 47180
rect 31500 47404 31668 47460
rect 31388 47124 31444 47134
rect 31388 46002 31444 47068
rect 31388 45950 31390 46002
rect 31442 45950 31444 46002
rect 31388 45938 31444 45950
rect 30940 44604 31220 44660
rect 30604 43138 30660 43148
rect 30716 43426 30772 43438
rect 30716 43374 30718 43426
rect 30770 43374 30772 43426
rect 30492 42642 30548 42654
rect 30492 42590 30494 42642
rect 30546 42590 30548 42642
rect 30492 41972 30548 42590
rect 30604 42644 30660 42654
rect 30604 42550 30660 42588
rect 30716 41972 30772 43374
rect 30492 41916 30716 41972
rect 30716 41906 30772 41916
rect 30828 42530 30884 42542
rect 30828 42478 30830 42530
rect 30882 42478 30884 42530
rect 30828 41188 30884 42478
rect 30828 41122 30884 41132
rect 30828 40964 30884 40974
rect 30380 40962 30884 40964
rect 30380 40910 30830 40962
rect 30882 40910 30884 40962
rect 30380 40908 30884 40910
rect 30380 40514 30436 40908
rect 30828 40898 30884 40908
rect 30940 40740 30996 44604
rect 31388 43538 31444 43550
rect 31388 43486 31390 43538
rect 31442 43486 31444 43538
rect 31388 43204 31444 43486
rect 31388 43138 31444 43148
rect 31500 41412 31556 47404
rect 31612 47236 31668 47246
rect 31668 47180 31780 47236
rect 31612 47170 31668 47180
rect 31724 46002 31780 47180
rect 31948 46788 32004 49420
rect 32172 49028 32228 49980
rect 32284 49810 32340 51326
rect 32620 50706 32676 51998
rect 32732 51940 32788 51950
rect 32732 51938 32900 51940
rect 32732 51886 32734 51938
rect 32786 51886 32900 51938
rect 32732 51884 32900 51886
rect 32732 51874 32788 51884
rect 32620 50654 32622 50706
rect 32674 50654 32676 50706
rect 32620 50642 32676 50654
rect 32844 50708 32900 51884
rect 33180 51604 33236 51614
rect 33292 51604 33348 53566
rect 33236 51548 33348 51604
rect 33404 53060 33460 53070
rect 33068 51490 33124 51502
rect 33068 51438 33070 51490
rect 33122 51438 33124 51490
rect 33068 51380 33124 51438
rect 33068 51314 33124 51324
rect 32844 50642 32900 50652
rect 33180 50594 33236 51548
rect 33404 51490 33460 53004
rect 33516 52162 33572 53790
rect 34748 53788 35140 53844
rect 35420 53956 35476 53966
rect 34636 53732 34692 53742
rect 34524 53730 34692 53732
rect 34524 53678 34638 53730
rect 34690 53678 34692 53730
rect 34524 53676 34692 53678
rect 33852 52948 33908 52958
rect 33516 52110 33518 52162
rect 33570 52110 33572 52162
rect 33516 52098 33572 52110
rect 33740 52388 33796 52398
rect 33404 51438 33406 51490
rect 33458 51438 33460 51490
rect 33404 51426 33460 51438
rect 33180 50542 33182 50594
rect 33234 50542 33236 50594
rect 33180 50530 33236 50542
rect 32956 50484 33012 50494
rect 33740 50428 33796 52332
rect 32956 50390 33012 50428
rect 33180 50372 33796 50428
rect 33852 50482 33908 52892
rect 33964 52164 34020 52174
rect 33964 52070 34020 52108
rect 34524 51716 34580 53676
rect 34636 53666 34692 53676
rect 34188 51660 34580 51716
rect 34636 51828 34692 51838
rect 33852 50430 33854 50482
rect 33906 50430 33908 50482
rect 33852 50418 33908 50430
rect 34076 51492 34132 51502
rect 34076 50428 34132 51436
rect 34188 51378 34244 51660
rect 34636 51602 34692 51772
rect 34636 51550 34638 51602
rect 34690 51550 34692 51602
rect 34636 51538 34692 51550
rect 34188 51326 34190 51378
rect 34242 51326 34244 51378
rect 34188 50596 34244 51326
rect 34412 51378 34468 51390
rect 34412 51326 34414 51378
rect 34466 51326 34468 51378
rect 34412 50820 34468 51326
rect 34524 51268 34580 51278
rect 34524 51174 34580 51212
rect 34412 50754 34468 50764
rect 34412 50596 34468 50606
rect 34244 50594 34468 50596
rect 34244 50542 34414 50594
rect 34466 50542 34468 50594
rect 34244 50540 34468 50542
rect 34188 50502 34244 50540
rect 34076 50372 34356 50428
rect 33180 50036 33236 50372
rect 32284 49758 32286 49810
rect 32338 49758 32340 49810
rect 32284 49028 32340 49758
rect 32508 49980 33236 50036
rect 32508 49810 32564 49980
rect 33404 49924 33460 49934
rect 32508 49758 32510 49810
rect 32562 49758 32564 49810
rect 32508 49746 32564 49758
rect 32620 49922 33460 49924
rect 32620 49870 33406 49922
rect 33458 49870 33460 49922
rect 32620 49868 33460 49870
rect 32508 49028 32564 49038
rect 32284 49026 32564 49028
rect 32284 48974 32510 49026
rect 32562 48974 32564 49026
rect 32284 48972 32564 48974
rect 31948 46722 32004 46732
rect 32060 48802 32116 48814
rect 32060 48750 32062 48802
rect 32114 48750 32116 48802
rect 32060 47458 32116 48750
rect 32172 48356 32228 48972
rect 32508 48962 32564 48972
rect 32620 48466 32676 49868
rect 33404 49858 33460 49868
rect 33180 49700 33236 49710
rect 32732 49698 33236 49700
rect 32732 49646 33182 49698
rect 33234 49646 33236 49698
rect 32732 49644 33236 49646
rect 32732 49138 32788 49644
rect 33180 49634 33236 49644
rect 32732 49086 32734 49138
rect 32786 49086 32788 49138
rect 32732 49074 32788 49086
rect 32844 49140 32900 49150
rect 32844 49046 32900 49084
rect 33516 49028 33572 50372
rect 34300 49138 34356 50372
rect 34300 49086 34302 49138
rect 34354 49086 34356 49138
rect 33516 48972 33796 49028
rect 33180 48916 33236 48926
rect 33180 48822 33236 48860
rect 33404 48914 33460 48926
rect 33404 48862 33406 48914
rect 33458 48862 33460 48914
rect 33292 48804 33348 48814
rect 33292 48692 33348 48748
rect 32620 48414 32622 48466
rect 32674 48414 32676 48466
rect 32620 48402 32676 48414
rect 33180 48636 33348 48692
rect 32284 48356 32340 48366
rect 32172 48354 32340 48356
rect 32172 48302 32286 48354
rect 32338 48302 32340 48354
rect 32172 48300 32340 48302
rect 32284 48290 32340 48300
rect 32396 48356 32452 48366
rect 32396 48262 32452 48300
rect 32844 48244 32900 48254
rect 32284 47684 32340 47694
rect 32340 47628 32452 47684
rect 32284 47618 32340 47628
rect 32060 47406 32062 47458
rect 32114 47406 32116 47458
rect 32060 47012 32116 47406
rect 31724 45950 31726 46002
rect 31778 45950 31780 46002
rect 31724 45938 31780 45950
rect 31836 46564 31892 46574
rect 31836 45556 31892 46508
rect 31948 46116 32004 46126
rect 31948 46022 32004 46060
rect 31612 45500 31892 45556
rect 31612 43538 31668 45500
rect 32060 45218 32116 46956
rect 32284 46676 32340 46686
rect 32284 46116 32340 46620
rect 32172 46114 32340 46116
rect 32172 46062 32286 46114
rect 32338 46062 32340 46114
rect 32172 46060 32340 46062
rect 32172 45330 32228 46060
rect 32284 46050 32340 46060
rect 32172 45278 32174 45330
rect 32226 45278 32228 45330
rect 32172 45266 32228 45278
rect 32060 45166 32062 45218
rect 32114 45166 32116 45218
rect 32060 45154 32116 45166
rect 32172 44884 32228 44894
rect 32060 44882 32228 44884
rect 32060 44830 32174 44882
rect 32226 44830 32228 44882
rect 32060 44828 32228 44830
rect 32060 43764 32116 44828
rect 32172 44818 32228 44828
rect 32396 44660 32452 47628
rect 32844 47682 32900 48188
rect 32844 47630 32846 47682
rect 32898 47630 32900 47682
rect 32844 47618 32900 47630
rect 33068 48132 33124 48142
rect 33068 47236 33124 48076
rect 33180 47458 33236 48636
rect 33292 48020 33348 48030
rect 33292 47926 33348 47964
rect 33404 47570 33460 48862
rect 33516 48804 33572 48814
rect 33516 48242 33572 48748
rect 33516 48190 33518 48242
rect 33570 48190 33572 48242
rect 33516 48178 33572 48190
rect 33628 48802 33684 48814
rect 33628 48750 33630 48802
rect 33682 48750 33684 48802
rect 33404 47518 33406 47570
rect 33458 47518 33460 47570
rect 33404 47506 33460 47518
rect 33516 48020 33572 48030
rect 33628 48020 33684 48750
rect 33740 48244 33796 48972
rect 33852 49026 33908 49038
rect 33852 48974 33854 49026
rect 33906 48974 33908 49026
rect 33852 48692 33908 48974
rect 34300 48804 34356 49086
rect 34300 48738 34356 48748
rect 34412 48692 34468 50540
rect 34636 50596 34692 50606
rect 34636 50428 34692 50540
rect 34524 50372 34692 50428
rect 34524 49140 34580 50372
rect 34748 50036 34804 53788
rect 35084 53618 35140 53630
rect 35084 53566 35086 53618
rect 35138 53566 35140 53618
rect 34860 51380 34916 51390
rect 35084 51380 35140 53566
rect 35420 53058 35476 53900
rect 35532 53732 35588 55132
rect 35644 54404 35700 55246
rect 35756 55188 35812 55412
rect 36092 55412 36148 57372
rect 36316 56308 36372 59200
rect 36316 56242 36372 56252
rect 36988 56196 37044 59200
rect 36988 56130 37044 56140
rect 36204 55972 36260 55982
rect 36204 55878 36260 55916
rect 36092 55346 36148 55356
rect 37212 55412 37268 55422
rect 37212 55318 37268 55356
rect 35756 55122 35812 55132
rect 36428 55188 36484 55198
rect 36428 55094 36484 55132
rect 35980 55076 36036 55086
rect 35980 54982 36036 55020
rect 36764 55076 36820 55086
rect 36092 54626 36148 54638
rect 36092 54574 36094 54626
rect 36146 54574 36148 54626
rect 35700 54348 35924 54404
rect 35644 54310 35700 54348
rect 35868 53842 35924 54348
rect 35868 53790 35870 53842
rect 35922 53790 35924 53842
rect 35868 53778 35924 53790
rect 35756 53732 35812 53742
rect 35532 53730 35812 53732
rect 35532 53678 35758 53730
rect 35810 53678 35812 53730
rect 35532 53676 35812 53678
rect 35420 53006 35422 53058
rect 35474 53006 35476 53058
rect 35420 52994 35476 53006
rect 35308 52946 35364 52958
rect 35308 52894 35310 52946
rect 35362 52894 35364 52946
rect 35308 52836 35364 52894
rect 35308 52770 35364 52780
rect 35196 52556 35460 52566
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35196 52490 35460 52500
rect 35532 52388 35588 52398
rect 34860 50484 34916 51324
rect 34860 50418 34916 50428
rect 34972 51378 35140 51380
rect 34972 51326 35086 51378
rect 35138 51326 35140 51378
rect 34972 51324 35140 51326
rect 34748 49970 34804 49980
rect 34972 49812 35028 51324
rect 35084 51314 35140 51324
rect 35196 52276 35252 52286
rect 35196 51156 35252 52220
rect 35532 52162 35588 52332
rect 35532 52110 35534 52162
rect 35586 52110 35588 52162
rect 35532 52098 35588 52110
rect 35756 52164 35812 53676
rect 36092 53060 36148 54574
rect 36316 54516 36372 54526
rect 36092 52994 36148 53004
rect 36204 54514 36372 54516
rect 36204 54462 36318 54514
rect 36370 54462 36372 54514
rect 36204 54460 36372 54462
rect 36204 53956 36260 54460
rect 36316 54450 36372 54460
rect 35980 52834 36036 52846
rect 35980 52782 35982 52834
rect 36034 52782 36036 52834
rect 35980 52388 36036 52782
rect 35980 52322 36036 52332
rect 36092 52164 36148 52174
rect 35756 52162 36148 52164
rect 35756 52110 36094 52162
rect 36146 52110 36148 52162
rect 35756 52108 36148 52110
rect 36092 52098 36148 52108
rect 36204 51940 36260 53900
rect 36764 53844 36820 55020
rect 37548 54626 37604 54638
rect 37548 54574 37550 54626
rect 37602 54574 37604 54626
rect 37212 54402 37268 54414
rect 37212 54350 37214 54402
rect 37266 54350 37268 54402
rect 36764 52946 36820 53788
rect 36764 52894 36766 52946
rect 36818 52894 36820 52946
rect 36764 52882 36820 52894
rect 36876 54180 36932 54190
rect 36316 52836 36372 52846
rect 36316 52050 36372 52780
rect 36876 52724 36932 54124
rect 37212 53844 37268 54350
rect 37436 54068 37492 54078
rect 37100 53842 37268 53844
rect 37100 53790 37214 53842
rect 37266 53790 37268 53842
rect 37100 53788 37268 53790
rect 37100 53620 37156 53788
rect 37212 53778 37268 53788
rect 37324 54012 37436 54068
rect 36764 52668 36932 52724
rect 36988 53060 37044 53070
rect 36316 51998 36318 52050
rect 36370 51998 36372 52050
rect 36316 51986 36372 51998
rect 36428 52050 36484 52062
rect 36428 51998 36430 52050
rect 36482 51998 36484 52050
rect 35980 51884 36260 51940
rect 36428 51940 36484 51998
rect 35644 51604 35700 51614
rect 35980 51604 36036 51884
rect 36428 51874 36484 51884
rect 36540 52052 36596 52062
rect 36316 51828 36372 51838
rect 35644 51602 36036 51604
rect 35644 51550 35646 51602
rect 35698 51550 36036 51602
rect 35644 51548 36036 51550
rect 36092 51772 36316 51828
rect 36092 51602 36148 51772
rect 36316 51762 36372 51772
rect 36092 51550 36094 51602
rect 36146 51550 36148 51602
rect 35644 51538 35700 51548
rect 36092 51538 36148 51550
rect 36316 51604 36372 51614
rect 35532 51492 35588 51502
rect 35532 51398 35588 51436
rect 35084 51100 35252 51156
rect 35756 51378 35812 51390
rect 35756 51326 35758 51378
rect 35810 51326 35812 51378
rect 35084 50594 35140 51100
rect 35196 50988 35460 50998
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35196 50922 35460 50932
rect 35084 50542 35086 50594
rect 35138 50542 35140 50594
rect 35084 50530 35140 50542
rect 35420 50820 35476 50830
rect 35420 50482 35476 50764
rect 35756 50596 35812 51326
rect 36316 51378 36372 51548
rect 36316 51326 36318 51378
rect 36370 51326 36372 51378
rect 36316 51314 36372 51326
rect 36428 51492 36484 51502
rect 35756 50530 35812 50540
rect 35420 50430 35422 50482
rect 35474 50430 35476 50482
rect 35420 50418 35476 50430
rect 35532 50484 35588 50494
rect 34748 49810 35028 49812
rect 34748 49758 34974 49810
rect 35026 49758 35028 49810
rect 34748 49756 35028 49758
rect 34748 49250 34804 49756
rect 34972 49746 35028 49756
rect 35196 49420 35460 49430
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35196 49354 35460 49364
rect 34748 49198 34750 49250
rect 34802 49198 34804 49250
rect 34748 49186 34804 49198
rect 34524 49046 34580 49084
rect 35196 49028 35252 49038
rect 35196 48934 35252 48972
rect 35532 49026 35588 50428
rect 36204 50482 36260 50494
rect 36204 50430 36206 50482
rect 36258 50430 36260 50482
rect 35532 48974 35534 49026
rect 35586 48974 35588 49026
rect 35420 48692 35476 48702
rect 33852 48636 34244 48692
rect 34412 48636 34580 48692
rect 34188 48354 34244 48636
rect 34188 48302 34190 48354
rect 34242 48302 34244 48354
rect 34188 48290 34244 48302
rect 33740 48150 33796 48188
rect 34412 48242 34468 48254
rect 34412 48190 34414 48242
rect 34466 48190 34468 48242
rect 34412 48020 34468 48190
rect 33628 47964 34468 48020
rect 33180 47406 33182 47458
rect 33234 47406 33236 47458
rect 33180 47394 33236 47406
rect 33516 47458 33572 47964
rect 33516 47406 33518 47458
rect 33570 47406 33572 47458
rect 33516 47348 33572 47406
rect 33404 47292 33572 47348
rect 33292 47236 33348 47246
rect 33068 47234 33348 47236
rect 33068 47182 33294 47234
rect 33346 47182 33348 47234
rect 33068 47180 33348 47182
rect 32732 46788 32788 46798
rect 32732 46002 32788 46732
rect 33068 46676 33124 46686
rect 33068 46582 33124 46620
rect 32732 45950 32734 46002
rect 32786 45950 32788 46002
rect 32732 45938 32788 45950
rect 33180 45892 33236 47180
rect 33292 47170 33348 47180
rect 33292 47012 33348 47022
rect 33292 46674 33348 46956
rect 33292 46622 33294 46674
rect 33346 46622 33348 46674
rect 33292 46610 33348 46622
rect 33068 45890 33236 45892
rect 33068 45838 33182 45890
rect 33234 45838 33236 45890
rect 33068 45836 33236 45838
rect 33404 45892 33460 47292
rect 33516 46676 33572 46686
rect 33516 46114 33572 46620
rect 33516 46062 33518 46114
rect 33570 46062 33572 46114
rect 33516 46050 33572 46062
rect 33516 45892 33572 45902
rect 33404 45890 33572 45892
rect 33404 45838 33518 45890
rect 33570 45838 33572 45890
rect 33404 45836 33572 45838
rect 33068 44772 33124 45836
rect 33180 45826 33236 45836
rect 33516 45826 33572 45836
rect 34412 45892 34468 45902
rect 34524 45892 34580 48636
rect 34636 48242 34692 48254
rect 34636 48190 34638 48242
rect 34690 48190 34692 48242
rect 34636 47572 34692 48190
rect 34860 48244 34916 48254
rect 34860 48150 34916 48188
rect 35084 48242 35140 48254
rect 35084 48190 35086 48242
rect 35138 48190 35140 48242
rect 34636 47506 34692 47516
rect 34972 47458 35028 47470
rect 34972 47406 34974 47458
rect 35026 47406 35028 47458
rect 34860 46674 34916 46686
rect 34860 46622 34862 46674
rect 34914 46622 34916 46674
rect 34860 46564 34916 46622
rect 34860 46498 34916 46508
rect 34972 46562 35028 47406
rect 35084 47124 35140 48190
rect 35420 48020 35476 48636
rect 35532 48356 35588 48974
rect 35644 49924 35700 49934
rect 35644 48914 35700 49868
rect 36204 49924 36260 50430
rect 36316 50484 36372 50494
rect 36428 50484 36484 51436
rect 36540 50594 36596 51996
rect 36764 51602 36820 52668
rect 36988 52388 37044 53004
rect 37100 53058 37156 53564
rect 37100 53006 37102 53058
rect 37154 53006 37156 53058
rect 37100 52994 37156 53006
rect 36988 52332 37156 52388
rect 36988 52162 37044 52174
rect 36988 52110 36990 52162
rect 37042 52110 37044 52162
rect 36988 51828 37044 52110
rect 36764 51550 36766 51602
rect 36818 51550 36820 51602
rect 36764 51538 36820 51550
rect 36876 51772 37044 51828
rect 36876 51604 36932 51772
rect 37100 51716 37156 52332
rect 37212 52164 37268 52174
rect 37324 52164 37380 54012
rect 37436 54002 37492 54012
rect 37548 53620 37604 54574
rect 37660 54628 37716 59200
rect 38332 56754 38388 59200
rect 40348 59108 40404 59200
rect 40572 59108 40628 59276
rect 40348 59052 40628 59108
rect 38332 56702 38334 56754
rect 38386 56702 38388 56754
rect 38332 56690 38388 56702
rect 40236 56754 40292 56766
rect 40236 56702 40238 56754
rect 40290 56702 40292 56754
rect 38892 56194 38948 56206
rect 38892 56142 38894 56194
rect 38946 56142 38948 56194
rect 38556 56082 38612 56094
rect 38556 56030 38558 56082
rect 38610 56030 38612 56082
rect 38556 55972 38612 56030
rect 38556 55468 38612 55916
rect 37660 54562 37716 54572
rect 38108 55412 38612 55468
rect 37660 53620 37716 53630
rect 37548 53618 37828 53620
rect 37548 53566 37662 53618
rect 37714 53566 37828 53618
rect 37548 53564 37828 53566
rect 37660 53554 37716 53564
rect 37548 52724 37604 52734
rect 37548 52722 37716 52724
rect 37548 52670 37550 52722
rect 37602 52670 37716 52722
rect 37548 52668 37716 52670
rect 37548 52658 37604 52668
rect 37212 52162 37380 52164
rect 37212 52110 37214 52162
rect 37266 52110 37380 52162
rect 37212 52108 37380 52110
rect 37212 52098 37268 52108
rect 36876 51538 36932 51548
rect 36988 51660 37156 51716
rect 37324 51940 37380 52108
rect 37436 52164 37492 52174
rect 37436 52050 37492 52108
rect 37436 51998 37438 52050
rect 37490 51998 37492 52050
rect 37436 51986 37492 51998
rect 37548 52162 37604 52174
rect 37548 52110 37550 52162
rect 37602 52110 37604 52162
rect 36540 50542 36542 50594
rect 36594 50542 36596 50594
rect 36540 50530 36596 50542
rect 36988 50484 37044 51660
rect 37100 51492 37156 51502
rect 37100 51490 37268 51492
rect 37100 51438 37102 51490
rect 37154 51438 37268 51490
rect 37100 51436 37268 51438
rect 37100 51426 37156 51436
rect 37212 50820 37268 51436
rect 37324 51380 37380 51884
rect 37548 51940 37604 52110
rect 37436 51492 37492 51502
rect 37436 51398 37492 51436
rect 37324 51314 37380 51324
rect 37548 50820 37604 51884
rect 37660 51156 37716 52668
rect 37772 51716 37828 53564
rect 37996 53060 38052 53070
rect 37884 52946 37940 52958
rect 37884 52894 37886 52946
rect 37938 52894 37940 52946
rect 37884 51940 37940 52894
rect 37996 52386 38052 53004
rect 37996 52334 37998 52386
rect 38050 52334 38052 52386
rect 37996 52322 38052 52334
rect 37884 51874 37940 51884
rect 37772 51660 37940 51716
rect 37772 51380 37828 51418
rect 37772 51314 37828 51324
rect 37772 51156 37828 51166
rect 37660 51100 37772 51156
rect 37772 51090 37828 51100
rect 36316 50482 36484 50484
rect 36316 50430 36318 50482
rect 36370 50430 36484 50482
rect 36316 50428 36484 50430
rect 36652 50428 37044 50484
rect 37100 50764 37492 50820
rect 36316 50418 36372 50428
rect 36652 50372 36820 50428
rect 36204 49858 36260 49868
rect 36316 49810 36372 49822
rect 36316 49758 36318 49810
rect 36370 49758 36372 49810
rect 35644 48862 35646 48914
rect 35698 48862 35700 48914
rect 35644 48850 35700 48862
rect 35756 49698 35812 49710
rect 35756 49646 35758 49698
rect 35810 49646 35812 49698
rect 35756 48692 35812 49646
rect 35980 49476 36036 49486
rect 35756 48626 35812 48636
rect 35868 49252 35924 49262
rect 35756 48466 35812 48478
rect 35756 48414 35758 48466
rect 35810 48414 35812 48466
rect 35644 48356 35700 48366
rect 35756 48356 35812 48414
rect 35532 48300 35644 48356
rect 35700 48300 35812 48356
rect 35644 48290 35700 48300
rect 35420 47964 35588 48020
rect 35196 47852 35460 47862
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35196 47786 35460 47796
rect 35420 47460 35476 47470
rect 35532 47460 35588 47964
rect 35420 47458 35700 47460
rect 35420 47406 35422 47458
rect 35474 47406 35700 47458
rect 35420 47404 35700 47406
rect 35420 47394 35476 47404
rect 35084 47058 35140 47068
rect 35532 47124 35588 47134
rect 34972 46510 34974 46562
rect 35026 46510 35028 46562
rect 34412 45890 34580 45892
rect 34412 45838 34414 45890
rect 34466 45838 34580 45890
rect 34412 45836 34580 45838
rect 34412 45826 34468 45836
rect 34636 45666 34692 45678
rect 34636 45614 34638 45666
rect 34690 45614 34692 45666
rect 34636 45220 34692 45614
rect 34748 45220 34804 45230
rect 34636 45218 34804 45220
rect 34636 45166 34750 45218
rect 34802 45166 34804 45218
rect 34636 45164 34804 45166
rect 33740 45108 33796 45118
rect 33740 45014 33796 45052
rect 33180 44996 33236 45006
rect 33516 44996 33572 45006
rect 33180 44994 33348 44996
rect 33180 44942 33182 44994
rect 33234 44942 33348 44994
rect 33180 44940 33348 44942
rect 33180 44930 33236 44940
rect 33068 44716 33236 44772
rect 32060 43698 32116 43708
rect 32172 44604 33124 44660
rect 32172 43650 32228 44604
rect 32172 43598 32174 43650
rect 32226 43598 32228 43650
rect 32172 43586 32228 43598
rect 32284 44436 32340 44446
rect 32284 43650 32340 44380
rect 32284 43598 32286 43650
rect 32338 43598 32340 43650
rect 32284 43586 32340 43598
rect 32396 44210 32452 44222
rect 32396 44158 32398 44210
rect 32450 44158 32452 44210
rect 31948 43540 32004 43550
rect 31612 43486 31614 43538
rect 31666 43486 31668 43538
rect 31612 43474 31668 43486
rect 31724 43538 32004 43540
rect 31724 43486 31950 43538
rect 32002 43486 32004 43538
rect 31724 43484 32004 43486
rect 31724 42644 31780 43484
rect 31948 43474 32004 43484
rect 31612 42084 31668 42094
rect 31724 42084 31780 42588
rect 32172 42866 32228 42878
rect 32172 42814 32174 42866
rect 32226 42814 32228 42866
rect 32172 42196 32228 42814
rect 32396 42754 32452 44158
rect 33068 43650 33124 44604
rect 33068 43598 33070 43650
rect 33122 43598 33124 43650
rect 33068 43586 33124 43598
rect 33180 43428 33236 44716
rect 32396 42702 32398 42754
rect 32450 42702 32452 42754
rect 32172 42194 32340 42196
rect 32172 42142 32174 42194
rect 32226 42142 32340 42194
rect 32172 42140 32340 42142
rect 32172 42130 32228 42140
rect 31612 42082 31780 42084
rect 31612 42030 31614 42082
rect 31666 42030 31780 42082
rect 31612 42028 31780 42030
rect 31612 42018 31668 42028
rect 31836 41972 31892 41982
rect 31836 41878 31892 41916
rect 30380 40462 30382 40514
rect 30434 40462 30436 40514
rect 30380 40450 30436 40462
rect 30492 40684 30996 40740
rect 31052 41356 31556 41412
rect 30268 38612 30436 38668
rect 29820 37940 29876 37950
rect 29596 37426 29652 37436
rect 29708 37884 29820 37940
rect 29484 37090 29540 37100
rect 29372 36418 29428 36428
rect 29148 36260 29204 36270
rect 29148 36166 29204 36204
rect 29372 36260 29428 36270
rect 29372 36258 29540 36260
rect 29372 36206 29374 36258
rect 29426 36206 29540 36258
rect 29372 36204 29540 36206
rect 29372 36194 29428 36204
rect 28924 36092 29092 36148
rect 28476 35980 28980 36036
rect 28140 35870 28142 35922
rect 28194 35870 28196 35922
rect 28140 35858 28196 35870
rect 28924 35922 28980 35980
rect 28924 35870 28926 35922
rect 28978 35870 28980 35922
rect 27916 35026 27972 35308
rect 27916 34974 27918 35026
rect 27970 34974 27972 35026
rect 27916 34962 27972 34974
rect 28028 35698 28084 35710
rect 28028 35646 28030 35698
rect 28082 35646 28084 35698
rect 27916 34804 27972 34814
rect 27916 34018 27972 34748
rect 27916 33966 27918 34018
rect 27970 33966 27972 34018
rect 27916 33954 27972 33966
rect 27804 33460 27860 33470
rect 27692 32004 27748 32014
rect 27692 31910 27748 31948
rect 27804 31892 27860 33404
rect 28028 33236 28084 35646
rect 28252 35698 28308 35710
rect 28252 35646 28254 35698
rect 28306 35646 28308 35698
rect 28252 35588 28308 35646
rect 28140 34692 28196 34702
rect 28140 34598 28196 34636
rect 28140 33236 28196 33246
rect 28028 33234 28196 33236
rect 28028 33182 28142 33234
rect 28194 33182 28196 33234
rect 28028 33180 28196 33182
rect 28028 33124 28084 33180
rect 28140 33170 28196 33180
rect 28028 33058 28084 33068
rect 28252 33012 28308 35532
rect 28924 35474 28980 35870
rect 28924 35422 28926 35474
rect 28978 35422 28980 35474
rect 28924 35410 28980 35422
rect 28364 35364 28420 35374
rect 28364 34802 28420 35308
rect 28476 35140 28532 35150
rect 28476 34914 28532 35084
rect 28476 34862 28478 34914
rect 28530 34862 28532 34914
rect 28476 34850 28532 34862
rect 28364 34750 28366 34802
rect 28418 34750 28420 34802
rect 28364 34738 28420 34750
rect 29036 33572 29092 36092
rect 29372 35588 29428 35598
rect 29372 35494 29428 35532
rect 29260 35474 29316 35486
rect 29260 35422 29262 35474
rect 29314 35422 29316 35474
rect 29260 35364 29316 35422
rect 29484 35476 29540 36204
rect 29484 35410 29540 35420
rect 29596 35700 29652 35710
rect 29260 35308 29428 35364
rect 29260 35140 29316 35150
rect 29260 34914 29316 35084
rect 29260 34862 29262 34914
rect 29314 34862 29316 34914
rect 29260 34850 29316 34862
rect 29372 34804 29428 35308
rect 29596 35252 29652 35644
rect 29372 34710 29428 34748
rect 29484 35196 29652 35252
rect 29036 33516 29316 33572
rect 29036 33460 29092 33516
rect 29036 33394 29092 33404
rect 29260 33458 29316 33516
rect 29260 33406 29262 33458
rect 29314 33406 29316 33458
rect 29260 33394 29316 33406
rect 29484 33236 29540 35196
rect 29708 35140 29764 37884
rect 29820 37846 29876 37884
rect 29932 37828 29988 37838
rect 30156 37828 30212 37838
rect 29932 37734 29988 37772
rect 30044 37826 30212 37828
rect 30044 37774 30158 37826
rect 30210 37774 30212 37826
rect 30044 37772 30212 37774
rect 29820 36484 29876 36494
rect 30044 36484 30100 37772
rect 30156 37762 30212 37772
rect 29820 36482 30100 36484
rect 29820 36430 29822 36482
rect 29874 36430 30100 36482
rect 29820 36428 30100 36430
rect 29820 36418 29876 36428
rect 29708 35074 29764 35084
rect 30268 35812 30324 35822
rect 29596 34916 29652 34926
rect 29596 34914 29988 34916
rect 29596 34862 29598 34914
rect 29650 34862 29988 34914
rect 29596 34860 29988 34862
rect 29596 34850 29652 34860
rect 29932 34802 29988 34860
rect 29932 34750 29934 34802
rect 29986 34750 29988 34802
rect 29932 34738 29988 34750
rect 30044 34804 30100 34814
rect 30044 34802 30212 34804
rect 30044 34750 30046 34802
rect 30098 34750 30212 34802
rect 30044 34748 30212 34750
rect 30044 34738 30100 34748
rect 29708 34692 29764 34702
rect 29708 34690 29876 34692
rect 29708 34638 29710 34690
rect 29762 34638 29876 34690
rect 29708 34636 29876 34638
rect 29708 34626 29764 34636
rect 29820 34356 29876 34636
rect 29820 34300 30100 34356
rect 30044 34242 30100 34300
rect 30044 34190 30046 34242
rect 30098 34190 30100 34242
rect 30044 34178 30100 34190
rect 30156 33460 30212 34748
rect 30156 33394 30212 33404
rect 29260 33180 29540 33236
rect 30156 33236 30212 33246
rect 28140 32956 28308 33012
rect 28476 33122 28532 33134
rect 28476 33070 28478 33122
rect 28530 33070 28532 33122
rect 27916 32450 27972 32462
rect 27916 32398 27918 32450
rect 27970 32398 27972 32450
rect 27916 32338 27972 32398
rect 27916 32286 27918 32338
rect 27970 32286 27972 32338
rect 27916 32228 27972 32286
rect 27916 32162 27972 32172
rect 28028 31892 28084 31902
rect 27804 31836 28028 31892
rect 27468 31724 27636 31780
rect 27692 31780 27748 31790
rect 27804 31780 27860 31836
rect 28028 31798 28084 31836
rect 27692 31778 27860 31780
rect 27692 31726 27694 31778
rect 27746 31726 27860 31778
rect 27692 31724 27860 31726
rect 27356 31668 27412 31678
rect 27356 31574 27412 31612
rect 27244 31388 27412 31444
rect 27244 30996 27300 31006
rect 27356 30996 27412 31388
rect 27468 31220 27524 31724
rect 27692 31714 27748 31724
rect 27468 31154 27524 31164
rect 27356 30940 27524 30996
rect 27244 30902 27300 30940
rect 27356 30436 27412 30446
rect 27356 30210 27412 30380
rect 27356 30158 27358 30210
rect 27410 30158 27412 30210
rect 27356 30146 27412 30158
rect 27468 29988 27524 30940
rect 27692 30212 27748 30222
rect 27580 30100 27636 30110
rect 27580 30006 27636 30044
rect 27132 29932 27412 29988
rect 27132 29540 27188 29550
rect 27132 29426 27188 29484
rect 27132 29374 27134 29426
rect 27186 29374 27188 29426
rect 27132 29362 27188 29374
rect 27020 29250 27076 29260
rect 26684 28590 26686 28642
rect 26738 28590 26740 28642
rect 26684 28578 26740 28590
rect 27132 28532 27188 28542
rect 27356 28532 27412 29932
rect 27468 29922 27524 29932
rect 27692 29540 27748 30156
rect 28028 30210 28084 30222
rect 28028 30158 28030 30210
rect 28082 30158 28084 30210
rect 28028 30100 28084 30158
rect 28028 30034 28084 30044
rect 27692 29474 27748 29484
rect 27804 29876 27860 29886
rect 28140 29876 28196 32956
rect 28476 32788 28532 33070
rect 28476 32722 28532 32732
rect 28700 32562 28756 32574
rect 28700 32510 28702 32562
rect 28754 32510 28756 32562
rect 28252 32450 28308 32462
rect 28252 32398 28254 32450
rect 28306 32398 28308 32450
rect 28252 31778 28308 32398
rect 28252 31726 28254 31778
rect 28306 31726 28308 31778
rect 28252 31668 28308 31726
rect 28252 31602 28308 31612
rect 28364 32338 28420 32350
rect 28364 32286 28366 32338
rect 28418 32286 28420 32338
rect 28364 31780 28420 32286
rect 28252 30436 28308 30446
rect 28364 30436 28420 31724
rect 28252 30434 28420 30436
rect 28252 30382 28254 30434
rect 28306 30382 28420 30434
rect 28252 30380 28420 30382
rect 28476 31892 28532 31902
rect 28252 30370 28308 30380
rect 28476 30322 28532 31836
rect 28476 30270 28478 30322
rect 28530 30270 28532 30322
rect 28476 30258 28532 30270
rect 28588 31556 28644 31566
rect 28700 31556 28756 32510
rect 28588 31554 28756 31556
rect 28588 31502 28590 31554
rect 28642 31502 28756 31554
rect 28588 31500 28756 31502
rect 29036 32562 29092 32574
rect 29036 32510 29038 32562
rect 29090 32510 29092 32562
rect 29036 32228 29092 32510
rect 28588 30212 28644 31500
rect 28588 30146 28644 30156
rect 27860 29820 28196 29876
rect 27580 29426 27636 29438
rect 27580 29374 27582 29426
rect 27634 29374 27636 29426
rect 27580 29316 27636 29374
rect 27804 29426 27860 29820
rect 28588 29652 28644 29662
rect 28140 29650 28644 29652
rect 28140 29598 28590 29650
rect 28642 29598 28644 29650
rect 28140 29596 28644 29598
rect 27804 29374 27806 29426
rect 27858 29374 27860 29426
rect 27804 29362 27860 29374
rect 28028 29428 28084 29438
rect 27580 28644 27636 29260
rect 27692 29314 27748 29326
rect 27692 29262 27694 29314
rect 27746 29262 27748 29314
rect 27692 28868 27748 29262
rect 27692 28802 27748 28812
rect 27692 28644 27748 28654
rect 27580 28642 27748 28644
rect 27580 28590 27694 28642
rect 27746 28590 27748 28642
rect 27580 28588 27748 28590
rect 27692 28578 27748 28588
rect 28028 28642 28084 29372
rect 28028 28590 28030 28642
rect 28082 28590 28084 28642
rect 28028 28578 28084 28590
rect 27468 28532 27524 28542
rect 27356 28530 27524 28532
rect 27356 28478 27470 28530
rect 27522 28478 27524 28530
rect 27356 28476 27524 28478
rect 26348 28420 26404 28430
rect 26348 27076 26404 28364
rect 26796 27748 26852 27758
rect 26796 27654 26852 27692
rect 26796 27524 26852 27534
rect 26572 27188 26628 27198
rect 26572 27094 26628 27132
rect 26348 27020 26516 27076
rect 25452 26852 25732 26908
rect 25564 26516 25620 26526
rect 25564 26422 25620 26460
rect 25452 26290 25508 26302
rect 25452 26238 25454 26290
rect 25506 26238 25508 26290
rect 25452 24388 25508 26238
rect 25676 26290 25732 26852
rect 26124 26852 26292 26908
rect 26460 26962 26516 27020
rect 26460 26910 26462 26962
rect 26514 26910 26516 26962
rect 26460 26898 26516 26910
rect 26684 26852 26740 26862
rect 26796 26852 26852 27468
rect 27132 27186 27188 28476
rect 27132 27134 27134 27186
rect 27186 27134 27188 27186
rect 27132 27122 27188 27134
rect 27356 28084 27412 28094
rect 26124 26402 26180 26852
rect 26684 26850 26852 26852
rect 26684 26798 26686 26850
rect 26738 26798 26852 26850
rect 26684 26796 26852 26798
rect 26684 26786 26740 26796
rect 26460 26516 26516 26526
rect 26460 26422 26516 26460
rect 26684 26516 26740 26526
rect 26684 26422 26740 26460
rect 26124 26350 26126 26402
rect 26178 26350 26180 26402
rect 26124 26338 26180 26350
rect 25676 26238 25678 26290
rect 25730 26238 25732 26290
rect 25676 26226 25732 26238
rect 27132 26290 27188 26302
rect 27132 26238 27134 26290
rect 27186 26238 27188 26290
rect 25900 26180 25956 26190
rect 25452 24322 25508 24332
rect 25788 26178 25956 26180
rect 25788 26126 25902 26178
rect 25954 26126 25956 26178
rect 25788 26124 25956 26126
rect 25172 23996 25396 24052
rect 25116 23958 25172 23996
rect 24332 23874 24388 23884
rect 25452 23940 25508 23950
rect 25452 23846 25508 23884
rect 24556 23826 24612 23838
rect 24556 23774 24558 23826
rect 24610 23774 24612 23826
rect 24108 23326 24110 23378
rect 24162 23326 24164 23378
rect 24108 23314 24164 23326
rect 24444 23380 24500 23390
rect 23996 22988 24276 23044
rect 23772 22950 23828 22988
rect 23660 22484 23716 22494
rect 23660 22390 23716 22428
rect 24220 22484 24276 22988
rect 24220 22418 24276 22428
rect 22988 22370 23492 22372
rect 22988 22318 23214 22370
rect 23266 22318 23492 22370
rect 22988 22316 23492 22318
rect 24444 22372 24500 23324
rect 24556 22596 24612 23774
rect 24668 23044 24724 23054
rect 24724 22988 25172 23044
rect 24668 22950 24724 22988
rect 24556 22530 24612 22540
rect 25116 22482 25172 22988
rect 25116 22430 25118 22482
rect 25170 22430 25172 22482
rect 25116 22418 25172 22430
rect 25564 22372 25620 22382
rect 24444 22316 24612 22372
rect 22876 21026 22932 22316
rect 23212 22260 23268 22316
rect 23548 22260 23604 22270
rect 24332 22260 24388 22270
rect 23212 22194 23268 22204
rect 23436 22258 23604 22260
rect 23436 22206 23550 22258
rect 23602 22206 23604 22258
rect 23436 22204 23604 22206
rect 23324 22146 23380 22158
rect 23324 22094 23326 22146
rect 23378 22094 23380 22146
rect 22876 20974 22878 21026
rect 22930 20974 22932 21026
rect 22876 20914 22932 20974
rect 22876 20862 22878 20914
rect 22930 20862 22932 20914
rect 22876 20850 22932 20862
rect 23100 21028 23156 21038
rect 22876 20132 22932 20142
rect 22876 20038 22932 20076
rect 23100 20018 23156 20972
rect 23324 20580 23380 22094
rect 23436 21364 23492 22204
rect 23548 22036 23604 22204
rect 24220 22258 24388 22260
rect 24220 22206 24334 22258
rect 24386 22206 24388 22258
rect 24220 22204 24388 22206
rect 23660 22148 23716 22186
rect 23660 22082 23716 22092
rect 23548 21970 23604 21980
rect 24220 21812 24276 22204
rect 24332 22194 24388 22204
rect 24556 22258 24612 22316
rect 25564 22278 25620 22316
rect 24556 22206 24558 22258
rect 24610 22206 24612 22258
rect 23660 21756 24276 21812
rect 24444 22146 24500 22158
rect 24444 22094 24446 22146
rect 24498 22094 24500 22146
rect 23548 21588 23604 21598
rect 23548 21494 23604 21532
rect 23660 21474 23716 21756
rect 23660 21422 23662 21474
rect 23714 21422 23716 21474
rect 23436 21308 23604 21364
rect 23324 20486 23380 20524
rect 23436 21026 23492 21038
rect 23436 20974 23438 21026
rect 23490 20974 23492 21026
rect 23436 20132 23492 20974
rect 23548 20916 23604 21308
rect 23548 20850 23604 20860
rect 23548 20132 23604 20142
rect 23436 20130 23604 20132
rect 23436 20078 23550 20130
rect 23602 20078 23604 20130
rect 23436 20076 23604 20078
rect 23100 19966 23102 20018
rect 23154 19966 23156 20018
rect 23100 19954 23156 19966
rect 22764 19618 22820 19628
rect 22204 19170 22260 19180
rect 22876 19236 22932 19246
rect 22876 19142 22932 19180
rect 21756 19058 21812 19068
rect 23548 19124 23604 20076
rect 23660 19346 23716 21422
rect 24332 21700 24388 21710
rect 24332 21474 24388 21644
rect 24332 21422 24334 21474
rect 24386 21422 24388 21474
rect 24332 21410 24388 21422
rect 24444 21028 24500 22094
rect 24556 21588 24612 22206
rect 24556 21522 24612 21532
rect 24780 22148 24836 22158
rect 24444 20962 24500 20972
rect 24220 20802 24276 20814
rect 24220 20750 24222 20802
rect 24274 20750 24276 20802
rect 24220 20242 24276 20750
rect 24556 20804 24612 20814
rect 24556 20802 24724 20804
rect 24556 20750 24558 20802
rect 24610 20750 24724 20802
rect 24556 20748 24724 20750
rect 24556 20738 24612 20748
rect 24220 20190 24222 20242
rect 24274 20190 24276 20242
rect 24220 20178 24276 20190
rect 24444 20130 24500 20142
rect 24444 20078 24446 20130
rect 24498 20078 24500 20130
rect 24444 20020 24500 20078
rect 24668 20132 24724 20748
rect 24444 19460 24500 19964
rect 24556 20018 24612 20030
rect 24556 19966 24558 20018
rect 24610 19966 24612 20018
rect 24556 19908 24612 19966
rect 24556 19842 24612 19852
rect 23660 19294 23662 19346
rect 23714 19294 23716 19346
rect 23660 19282 23716 19294
rect 24220 19404 24500 19460
rect 23548 19068 23940 19124
rect 23436 19012 23492 19022
rect 23548 19012 23604 19068
rect 23492 18956 23604 19012
rect 23436 18946 23492 18956
rect 21084 18562 21140 18574
rect 21084 18510 21086 18562
rect 21138 18510 21140 18562
rect 20972 18452 21028 18462
rect 20860 18450 21028 18452
rect 20860 18398 20974 18450
rect 21026 18398 21028 18450
rect 20860 18396 21028 18398
rect 20860 17780 20916 18396
rect 20972 18386 21028 18396
rect 21084 18452 21140 18510
rect 23212 18562 23268 18574
rect 23212 18510 23214 18562
rect 23266 18510 23268 18562
rect 21084 17892 21140 18396
rect 22764 18450 22820 18462
rect 22764 18398 22766 18450
rect 22818 18398 22820 18450
rect 21084 17836 21364 17892
rect 20860 17778 21252 17780
rect 20860 17726 20862 17778
rect 20914 17726 21252 17778
rect 20860 17724 21252 17726
rect 20860 17714 20916 17724
rect 20748 16930 20804 16940
rect 20972 17556 21028 17566
rect 20972 17106 21028 17500
rect 21196 17332 21252 17724
rect 21308 17554 21364 17836
rect 21644 17668 21700 17678
rect 21980 17668 22036 17678
rect 22204 17668 22260 17678
rect 21644 17666 22148 17668
rect 21644 17614 21646 17666
rect 21698 17614 21982 17666
rect 22034 17614 22148 17666
rect 21644 17612 22148 17614
rect 21644 17602 21700 17612
rect 21980 17602 22036 17612
rect 21308 17502 21310 17554
rect 21362 17502 21364 17554
rect 21308 17490 21364 17502
rect 21420 17442 21476 17454
rect 21420 17390 21422 17442
rect 21474 17390 21476 17442
rect 21420 17332 21476 17390
rect 21196 17276 21476 17332
rect 20972 17054 20974 17106
rect 21026 17054 21028 17106
rect 20972 16884 21028 17054
rect 21756 16996 21812 17006
rect 21756 16902 21812 16940
rect 20972 16818 21028 16828
rect 22092 16882 22148 17612
rect 22204 17574 22260 17612
rect 22316 17554 22372 17566
rect 22316 17502 22318 17554
rect 22370 17502 22372 17554
rect 22092 16830 22094 16882
rect 22146 16830 22148 16882
rect 22092 16818 22148 16830
rect 22204 16884 22260 16894
rect 20636 15486 20638 15538
rect 20690 15486 20692 15538
rect 20636 15474 20692 15486
rect 21420 16098 21476 16110
rect 21420 16046 21422 16098
rect 21474 16046 21476 16098
rect 21308 14756 21364 14766
rect 21420 14756 21476 16046
rect 21308 14754 21476 14756
rect 21308 14702 21310 14754
rect 21362 14702 21476 14754
rect 21308 14700 21476 14702
rect 21644 16100 21700 16110
rect 21308 14644 21364 14700
rect 21308 14578 21364 14588
rect 21644 14530 21700 16044
rect 21644 14478 21646 14530
rect 21698 14478 21700 14530
rect 21644 14466 21700 14478
rect 21420 14308 21476 14318
rect 21420 14214 21476 14252
rect 19628 12898 19684 12908
rect 19964 13020 20468 13076
rect 19964 12850 20020 13020
rect 20412 12962 20468 13020
rect 20412 12910 20414 12962
rect 20466 12910 20468 12962
rect 20412 12898 20468 12910
rect 20636 13636 20692 13646
rect 19964 12798 19966 12850
rect 20018 12798 20020 12850
rect 19964 12786 20020 12798
rect 20076 12852 20132 12862
rect 20076 12758 20132 12796
rect 19740 12740 19796 12750
rect 19628 12738 19796 12740
rect 19628 12686 19742 12738
rect 19794 12686 19796 12738
rect 19628 12684 19796 12686
rect 19628 12292 19684 12684
rect 19740 12674 19796 12684
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 20636 12402 20692 13580
rect 21756 13188 21812 13198
rect 21644 13132 21756 13188
rect 20748 12964 20804 12974
rect 20748 12850 20804 12908
rect 20748 12798 20750 12850
rect 20802 12798 20804 12850
rect 20748 12786 20804 12798
rect 21420 12964 21476 12974
rect 20636 12350 20638 12402
rect 20690 12350 20692 12402
rect 20636 12338 20692 12350
rect 19628 12226 19684 12236
rect 20188 12180 20244 12190
rect 20076 12178 20244 12180
rect 20076 12126 20190 12178
rect 20242 12126 20244 12178
rect 20076 12124 20244 12126
rect 19628 11956 19684 11966
rect 19516 11900 19628 11956
rect 19628 11890 19684 11900
rect 19292 11506 19460 11508
rect 19292 11454 19294 11506
rect 19346 11454 19460 11506
rect 19292 11452 19460 11454
rect 19292 11442 19348 11452
rect 19852 11396 19908 11406
rect 20076 11396 20132 12124
rect 20188 12114 20244 12124
rect 20972 12068 21028 12078
rect 20412 11956 20468 11966
rect 19852 11394 20132 11396
rect 19852 11342 19854 11394
rect 19906 11342 20132 11394
rect 19852 11340 20132 11342
rect 20300 11394 20356 11406
rect 20300 11342 20302 11394
rect 20354 11342 20356 11394
rect 18732 11284 18788 11294
rect 18732 11190 18788 11228
rect 19852 11172 19908 11340
rect 19628 11116 19908 11172
rect 18508 10558 18510 10610
rect 18562 10558 18564 10610
rect 18508 10546 18564 10558
rect 19404 10612 19460 10622
rect 19404 10518 19460 10556
rect 17948 9772 18340 9828
rect 16940 9716 16996 9726
rect 16940 9622 16996 9660
rect 17836 9714 17892 9726
rect 17836 9662 17838 9714
rect 17890 9662 17892 9714
rect 16268 8082 16324 8092
rect 16380 9604 16436 9614
rect 15596 7746 15652 7756
rect 15596 7476 15652 7486
rect 16044 7476 16100 7486
rect 15596 7474 15764 7476
rect 15596 7422 15598 7474
rect 15650 7422 15764 7474
rect 15596 7420 15764 7422
rect 15596 7410 15652 7420
rect 15484 6862 15486 6914
rect 15538 6862 15540 6914
rect 15484 6850 15540 6862
rect 15708 6804 15764 7420
rect 16044 7382 16100 7420
rect 16380 7474 16436 9548
rect 16716 9604 16772 9614
rect 17724 9604 17780 9614
rect 16716 9602 16884 9604
rect 16716 9550 16718 9602
rect 16770 9550 16884 9602
rect 16716 9548 16884 9550
rect 16716 9538 16772 9548
rect 16716 8820 16772 8830
rect 16716 8146 16772 8764
rect 16828 8260 16884 9548
rect 17724 9042 17780 9548
rect 17836 9268 17892 9662
rect 17948 9714 18004 9772
rect 17948 9662 17950 9714
rect 18002 9662 18004 9714
rect 17948 9650 18004 9662
rect 17836 9202 17892 9212
rect 18172 9602 18228 9614
rect 18172 9550 18174 9602
rect 18226 9550 18228 9602
rect 17724 8990 17726 9042
rect 17778 8990 17780 9042
rect 17724 8978 17780 8990
rect 17948 9044 18004 9054
rect 18172 9044 18228 9550
rect 17948 9042 18228 9044
rect 17948 8990 17950 9042
rect 18002 8990 18228 9042
rect 17948 8988 18228 8990
rect 17500 8932 17556 8942
rect 17500 8838 17556 8876
rect 17948 8820 18004 8988
rect 17948 8754 18004 8764
rect 16940 8260 16996 8270
rect 16828 8258 16996 8260
rect 16828 8206 16942 8258
rect 16994 8206 16996 8258
rect 16828 8204 16996 8206
rect 16940 8194 16996 8204
rect 17836 8258 17892 8270
rect 17836 8206 17838 8258
rect 17890 8206 17892 8258
rect 16716 8094 16718 8146
rect 16770 8094 16772 8146
rect 16716 8082 16772 8094
rect 17836 8148 17892 8206
rect 17836 8082 17892 8092
rect 18284 8036 18340 9772
rect 18732 9826 18788 9838
rect 18732 9774 18734 9826
rect 18786 9774 18788 9826
rect 18732 9266 18788 9774
rect 19292 9828 19348 9838
rect 19628 9828 19684 11116
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 20300 10388 20356 11342
rect 20412 10610 20468 11900
rect 20748 11396 20804 11406
rect 20748 11302 20804 11340
rect 20412 10558 20414 10610
rect 20466 10558 20468 10610
rect 20412 10546 20468 10558
rect 20972 10610 21028 12012
rect 20972 10558 20974 10610
rect 21026 10558 21028 10610
rect 20972 10546 21028 10558
rect 20524 10388 20580 10398
rect 20300 10386 20580 10388
rect 20300 10334 20526 10386
rect 20578 10334 20580 10386
rect 20300 10332 20580 10334
rect 19292 9826 19684 9828
rect 19292 9774 19294 9826
rect 19346 9774 19684 9826
rect 19292 9772 19684 9774
rect 20188 9938 20244 9950
rect 20188 9886 20190 9938
rect 20242 9886 20244 9938
rect 18732 9214 18734 9266
rect 18786 9214 18788 9266
rect 18732 9202 18788 9214
rect 19180 9268 19236 9278
rect 19180 9174 19236 9212
rect 19180 8484 19236 8494
rect 19292 8484 19348 9772
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 19516 9268 19572 9278
rect 19516 9174 19572 9212
rect 19180 8482 19348 8484
rect 19180 8430 19182 8482
rect 19234 8430 19348 8482
rect 19180 8428 19348 8430
rect 20076 8932 20132 8942
rect 20188 8932 20244 9886
rect 20524 9826 20580 10332
rect 20524 9774 20526 9826
rect 20578 9774 20580 9826
rect 20524 9762 20580 9774
rect 21420 9940 21476 12908
rect 21644 12850 21700 13132
rect 21756 13122 21812 13132
rect 21644 12798 21646 12850
rect 21698 12798 21700 12850
rect 21644 12786 21700 12798
rect 21756 12962 21812 12974
rect 21756 12910 21758 12962
rect 21810 12910 21812 12962
rect 21756 12852 21812 12910
rect 21756 11732 21812 12796
rect 22092 12850 22148 12862
rect 22092 12798 22094 12850
rect 22146 12798 22148 12850
rect 22092 12740 22148 12798
rect 22092 12674 22148 12684
rect 22204 12404 22260 16828
rect 22316 16884 22372 17502
rect 22764 17108 22820 18398
rect 23212 17780 23268 18510
rect 23660 18562 23716 18574
rect 23660 18510 23662 18562
rect 23714 18510 23716 18562
rect 23324 17780 23380 17790
rect 23100 17778 23380 17780
rect 23100 17726 23326 17778
rect 23378 17726 23380 17778
rect 23100 17724 23380 17726
rect 22876 17668 22932 17678
rect 22876 17574 22932 17612
rect 22764 17042 22820 17052
rect 22988 16884 23044 16894
rect 22316 16882 23044 16884
rect 22316 16830 22990 16882
rect 23042 16830 23044 16882
rect 22316 16828 23044 16830
rect 22316 16210 22372 16828
rect 22988 16818 23044 16828
rect 22988 16324 23044 16334
rect 23100 16324 23156 17724
rect 23324 17714 23380 17724
rect 23660 16548 23716 18510
rect 23884 18450 23940 19068
rect 23884 18398 23886 18450
rect 23938 18398 23940 18450
rect 23884 18386 23940 18398
rect 23660 16492 24164 16548
rect 22988 16322 23156 16324
rect 22988 16270 22990 16322
rect 23042 16270 23156 16322
rect 22988 16268 23156 16270
rect 22652 16212 22708 16222
rect 22316 16158 22318 16210
rect 22370 16158 22372 16210
rect 22316 16146 22372 16158
rect 22540 16210 22708 16212
rect 22540 16158 22654 16210
rect 22706 16158 22708 16210
rect 22540 16156 22708 16158
rect 22428 15876 22484 15886
rect 22428 15426 22484 15820
rect 22428 15374 22430 15426
rect 22482 15374 22484 15426
rect 22428 15362 22484 15374
rect 22540 15314 22596 16156
rect 22652 16146 22708 16156
rect 22540 15262 22542 15314
rect 22594 15262 22596 15314
rect 22540 15250 22596 15262
rect 22764 15874 22820 15886
rect 22764 15822 22766 15874
rect 22818 15822 22820 15874
rect 22764 14980 22820 15822
rect 22540 14924 22764 14980
rect 22540 14308 22596 14924
rect 22764 14914 22820 14924
rect 22988 14756 23044 16268
rect 23660 16100 23716 16110
rect 23324 15988 23380 15998
rect 23324 15894 23380 15932
rect 23660 15986 23716 16044
rect 23660 15934 23662 15986
rect 23714 15934 23716 15986
rect 23436 15314 23492 15326
rect 23436 15262 23438 15314
rect 23490 15262 23492 15314
rect 22428 13748 22484 13758
rect 22540 13748 22596 14252
rect 22428 13746 22596 13748
rect 22428 13694 22430 13746
rect 22482 13694 22596 13746
rect 22428 13692 22596 13694
rect 22652 14700 23044 14756
rect 23100 14980 23156 14990
rect 22652 14642 22708 14700
rect 22652 14590 22654 14642
rect 22706 14590 22708 14642
rect 22652 13746 22708 14590
rect 23100 14530 23156 14924
rect 23100 14478 23102 14530
rect 23154 14478 23156 14530
rect 23100 14466 23156 14478
rect 23436 14530 23492 15262
rect 23548 14644 23604 14654
rect 23548 14550 23604 14588
rect 23436 14478 23438 14530
rect 23490 14478 23492 14530
rect 22652 13694 22654 13746
rect 22706 13694 22708 13746
rect 22428 13682 22484 13692
rect 22652 13682 22708 13694
rect 23324 13748 23380 13758
rect 23324 13654 23380 13692
rect 22876 13636 22932 13646
rect 22876 13542 22932 13580
rect 23436 13636 23492 14478
rect 23660 13858 23716 15934
rect 24108 15986 24164 16492
rect 24220 16436 24276 19404
rect 24668 19236 24724 20076
rect 24780 19908 24836 22092
rect 25676 21700 25732 21710
rect 25788 21700 25844 26124
rect 25900 26114 25956 26124
rect 26572 26180 26628 26190
rect 26572 26086 26628 26124
rect 27020 25620 27076 25630
rect 26460 24948 26516 24958
rect 26460 24854 26516 24892
rect 26908 24948 26964 24958
rect 26908 24890 26964 24892
rect 26908 24838 26910 24890
rect 26962 24838 26964 24890
rect 26908 24826 26964 24838
rect 27020 24834 27076 25564
rect 27132 24948 27188 26238
rect 27244 24948 27300 24958
rect 27132 24946 27300 24948
rect 27132 24894 27246 24946
rect 27298 24894 27300 24946
rect 27132 24892 27300 24894
rect 27244 24882 27300 24892
rect 27020 24782 27022 24834
rect 27074 24782 27076 24834
rect 27020 24612 27076 24782
rect 26908 24556 27076 24612
rect 26236 23826 26292 23838
rect 26236 23774 26238 23826
rect 26290 23774 26292 23826
rect 26236 23380 26292 23774
rect 26236 23314 26292 23324
rect 26908 22708 26964 24556
rect 27356 23378 27412 28028
rect 27468 26908 27524 28476
rect 27580 28418 27636 28430
rect 27580 28366 27582 28418
rect 27634 28366 27636 28418
rect 27580 27524 27636 28366
rect 28140 28084 28196 29596
rect 28588 29586 28644 29596
rect 28700 29652 28756 29662
rect 28476 29426 28532 29438
rect 28476 29374 28478 29426
rect 28530 29374 28532 29426
rect 28476 29316 28532 29374
rect 28476 29250 28532 29260
rect 28700 29204 28756 29596
rect 29036 29316 29092 32172
rect 29148 30100 29204 30110
rect 29148 29876 29204 30044
rect 29148 29650 29204 29820
rect 29260 29764 29316 33180
rect 30156 33142 30212 33180
rect 29708 33122 29764 33134
rect 29708 33070 29710 33122
rect 29762 33070 29764 33122
rect 29708 32900 29764 33070
rect 29708 32834 29764 32844
rect 29820 32788 29876 32798
rect 29820 32694 29876 32732
rect 29484 32450 29540 32462
rect 29484 32398 29486 32450
rect 29538 32398 29540 32450
rect 29372 31780 29428 31790
rect 29372 31686 29428 31724
rect 29484 30210 29540 32398
rect 29820 32452 29876 32462
rect 29596 32228 29652 32238
rect 29596 31890 29652 32172
rect 29596 31838 29598 31890
rect 29650 31838 29652 31890
rect 29596 31826 29652 31838
rect 29820 31892 29876 32396
rect 30156 32338 30212 32350
rect 30156 32286 30158 32338
rect 30210 32286 30212 32338
rect 30156 32004 30212 32286
rect 30156 31938 30212 31948
rect 29820 31780 29876 31836
rect 29708 31778 29876 31780
rect 29708 31726 29822 31778
rect 29874 31726 29876 31778
rect 29708 31724 29876 31726
rect 29484 30158 29486 30210
rect 29538 30158 29540 30210
rect 29484 29988 29540 30158
rect 29484 29922 29540 29932
rect 29596 31554 29652 31566
rect 29596 31502 29598 31554
rect 29650 31502 29652 31554
rect 29596 30322 29652 31502
rect 29596 30270 29598 30322
rect 29650 30270 29652 30322
rect 29260 29708 29540 29764
rect 29148 29598 29150 29650
rect 29202 29598 29204 29650
rect 29148 29586 29204 29598
rect 29372 29426 29428 29438
rect 29372 29374 29374 29426
rect 29426 29374 29428 29426
rect 29372 29316 29428 29374
rect 29036 29260 29428 29316
rect 28588 29148 28756 29204
rect 28476 28868 28532 28878
rect 28140 28018 28196 28028
rect 28252 28866 28532 28868
rect 28252 28814 28478 28866
rect 28530 28814 28532 28866
rect 28252 28812 28532 28814
rect 27580 27458 27636 27468
rect 27692 27748 27748 27758
rect 27692 27186 27748 27692
rect 27692 27134 27694 27186
rect 27746 27134 27748 27186
rect 27692 27122 27748 27134
rect 27580 27076 27636 27114
rect 27580 27010 27636 27020
rect 28252 27074 28308 28812
rect 28476 28802 28532 28812
rect 28252 27022 28254 27074
rect 28306 27022 28308 27074
rect 28252 27010 28308 27022
rect 28364 28530 28420 28542
rect 28364 28478 28366 28530
rect 28418 28478 28420 28530
rect 28364 27860 28420 28478
rect 28476 28420 28532 28430
rect 28476 28326 28532 28364
rect 28364 26908 28420 27804
rect 28588 27186 28644 29148
rect 28924 28420 28980 28430
rect 28588 27134 28590 27186
rect 28642 27134 28644 27186
rect 28588 27122 28644 27134
rect 28700 27972 28756 27982
rect 27468 26852 27748 26908
rect 27692 26628 27748 26852
rect 27804 26852 27860 26862
rect 27804 26758 27860 26796
rect 28252 26852 28420 26908
rect 27692 26572 28196 26628
rect 28140 26514 28196 26572
rect 28140 26462 28142 26514
rect 28194 26462 28196 26514
rect 28140 26450 28196 26462
rect 27692 26402 27748 26414
rect 27692 26350 27694 26402
rect 27746 26350 27748 26402
rect 27468 26292 27524 26302
rect 27692 26292 27748 26350
rect 28252 26292 28308 26852
rect 27524 26236 27636 26292
rect 27692 26236 28308 26292
rect 27468 26198 27524 26236
rect 27468 25620 27524 25630
rect 27468 25526 27524 25564
rect 27580 25508 27636 26236
rect 27804 25508 27860 25518
rect 27580 25506 27860 25508
rect 27580 25454 27806 25506
rect 27858 25454 27860 25506
rect 27580 25452 27860 25454
rect 27804 25442 27860 25452
rect 27916 25284 27972 26236
rect 28140 25508 28196 25518
rect 28140 25394 28196 25452
rect 28140 25342 28142 25394
rect 28194 25342 28196 25394
rect 28140 25330 28196 25342
rect 27692 25228 27972 25284
rect 27692 24948 27748 25228
rect 27692 24834 27748 24892
rect 27692 24782 27694 24834
rect 27746 24782 27748 24834
rect 27692 24770 27748 24782
rect 27804 24836 27860 24846
rect 27804 24834 27972 24836
rect 27804 24782 27806 24834
rect 27858 24782 27972 24834
rect 27804 24780 27972 24782
rect 27804 24770 27860 24780
rect 27916 24612 27972 24780
rect 28364 24612 28420 24622
rect 27916 24610 28420 24612
rect 27916 24558 28366 24610
rect 28418 24558 28420 24610
rect 27916 24556 28420 24558
rect 27804 24498 27860 24510
rect 27804 24446 27806 24498
rect 27858 24446 27860 24498
rect 27356 23326 27358 23378
rect 27410 23326 27412 23378
rect 27356 23314 27412 23326
rect 27468 23380 27524 23390
rect 27468 23286 27524 23324
rect 27804 23378 27860 24446
rect 28364 24052 28420 24556
rect 28364 24050 28532 24052
rect 28364 23998 28366 24050
rect 28418 23998 28532 24050
rect 28364 23996 28532 23998
rect 28364 23986 28420 23996
rect 27804 23326 27806 23378
rect 27858 23326 27860 23378
rect 27804 23314 27860 23326
rect 27580 23154 27636 23166
rect 27580 23102 27582 23154
rect 27634 23102 27636 23154
rect 26908 22652 27300 22708
rect 26460 22484 26516 22494
rect 26460 22482 26852 22484
rect 26460 22430 26462 22482
rect 26514 22430 26852 22482
rect 26460 22428 26852 22430
rect 26460 22418 26516 22428
rect 26348 22370 26404 22382
rect 26348 22318 26350 22370
rect 26402 22318 26404 22370
rect 25676 21698 25844 21700
rect 25676 21646 25678 21698
rect 25730 21646 25844 21698
rect 25676 21644 25844 21646
rect 26012 22258 26068 22270
rect 26012 22206 26014 22258
rect 26066 22206 26068 22258
rect 26012 21700 26068 22206
rect 26348 22260 26404 22318
rect 26348 22194 26404 22204
rect 26572 22258 26628 22270
rect 26572 22206 26574 22258
rect 26626 22206 26628 22258
rect 25676 21634 25732 21644
rect 26012 21634 26068 21644
rect 26348 21588 26404 21598
rect 26348 21494 26404 21532
rect 26012 21474 26068 21486
rect 26012 21422 26014 21474
rect 26066 21422 26068 21474
rect 26012 20916 26068 21422
rect 26012 20822 26068 20860
rect 25228 20804 25284 20814
rect 24780 19842 24836 19852
rect 25116 20802 25284 20804
rect 25116 20750 25230 20802
rect 25282 20750 25284 20802
rect 25116 20748 25284 20750
rect 24780 19236 24836 19246
rect 24668 19234 24836 19236
rect 24668 19182 24782 19234
rect 24834 19182 24836 19234
rect 24668 19180 24836 19182
rect 24780 18900 24836 19180
rect 24780 18834 24836 18844
rect 25004 19236 25060 19246
rect 25116 19236 25172 20748
rect 25228 20738 25284 20748
rect 25564 20132 25620 20142
rect 25564 20038 25620 20076
rect 26572 20132 26628 22206
rect 26796 21812 26852 22428
rect 26796 21756 27076 21812
rect 26684 21700 26740 21710
rect 26684 21476 26740 21644
rect 27020 21698 27076 21756
rect 27020 21646 27022 21698
rect 27074 21646 27076 21698
rect 27020 21634 27076 21646
rect 27132 21588 27188 21598
rect 27132 21494 27188 21532
rect 26684 21420 26964 21476
rect 26908 20802 26964 21420
rect 27244 21364 27300 22652
rect 26908 20750 26910 20802
rect 26962 20750 26964 20802
rect 26908 20738 26964 20750
rect 27020 21308 27300 21364
rect 27356 22260 27412 22270
rect 27020 20356 27076 21308
rect 27356 20690 27412 22204
rect 27580 22148 27636 23102
rect 28028 22596 28084 22606
rect 28028 22502 28084 22540
rect 27916 22484 27972 22494
rect 27916 22370 27972 22428
rect 27916 22318 27918 22370
rect 27970 22318 27972 22370
rect 27916 22306 27972 22318
rect 28252 22370 28308 22382
rect 28252 22318 28254 22370
rect 28306 22318 28308 22370
rect 27804 22148 27860 22158
rect 27580 22146 27860 22148
rect 27580 22094 27806 22146
rect 27858 22094 27860 22146
rect 27580 22092 27860 22094
rect 27804 22082 27860 22092
rect 27468 21588 27524 21598
rect 27524 21532 27972 21588
rect 27468 21494 27524 21532
rect 27692 21364 27748 21374
rect 27580 21362 27748 21364
rect 27580 21310 27694 21362
rect 27746 21310 27748 21362
rect 27580 21308 27748 21310
rect 27468 21028 27524 21038
rect 27580 21028 27636 21308
rect 27692 21298 27748 21308
rect 27468 21026 27636 21028
rect 27468 20974 27470 21026
rect 27522 20974 27636 21026
rect 27468 20972 27636 20974
rect 27468 20962 27524 20972
rect 27692 20916 27748 20926
rect 27692 20822 27748 20860
rect 27356 20638 27358 20690
rect 27410 20638 27412 20690
rect 27356 20626 27412 20638
rect 27916 20690 27972 21532
rect 28028 21364 28084 21374
rect 28028 21270 28084 21308
rect 27916 20638 27918 20690
rect 27970 20638 27972 20690
rect 27916 20626 27972 20638
rect 28028 20914 28084 20926
rect 28028 20862 28030 20914
rect 28082 20862 28084 20914
rect 27132 20580 27188 20590
rect 27132 20578 27300 20580
rect 27132 20526 27134 20578
rect 27186 20526 27300 20578
rect 27132 20524 27300 20526
rect 27132 20514 27188 20524
rect 27020 20300 27188 20356
rect 25228 20020 25284 20030
rect 25228 19926 25284 19964
rect 26124 19908 26180 19918
rect 25004 19234 25172 19236
rect 25004 19182 25006 19234
rect 25058 19182 25172 19234
rect 25004 19180 25172 19182
rect 26012 19236 26068 19246
rect 24556 18676 24612 18686
rect 24556 18582 24612 18620
rect 24444 18564 24500 18574
rect 24444 18470 24500 18508
rect 24780 18452 24836 18462
rect 24780 18358 24836 18396
rect 24332 17668 24388 17678
rect 24332 16994 24388 17612
rect 24332 16942 24334 16994
rect 24386 16942 24388 16994
rect 24332 16930 24388 16942
rect 24444 17666 24500 17678
rect 24444 17614 24446 17666
rect 24498 17614 24500 17666
rect 24444 16996 24500 17614
rect 25004 17668 25060 19180
rect 26012 19142 26068 19180
rect 26124 19234 26180 19852
rect 26124 19182 26126 19234
rect 26178 19182 26180 19234
rect 26124 19170 26180 19182
rect 25228 19124 25284 19134
rect 25564 19124 25620 19134
rect 25228 19122 25620 19124
rect 25228 19070 25230 19122
rect 25282 19070 25566 19122
rect 25618 19070 25620 19122
rect 25228 19068 25620 19070
rect 25228 19058 25284 19068
rect 25564 19058 25620 19068
rect 25788 19122 25844 19134
rect 25788 19070 25790 19122
rect 25842 19070 25844 19122
rect 25452 18900 25508 18910
rect 25004 17602 25060 17612
rect 25228 18676 25284 18686
rect 24444 16930 24500 16940
rect 24220 16380 24388 16436
rect 24220 16100 24276 16110
rect 24220 16006 24276 16044
rect 24108 15934 24110 15986
rect 24162 15934 24164 15986
rect 23884 15876 23940 15886
rect 23884 15782 23940 15820
rect 24108 15148 24164 15934
rect 23996 15092 24164 15148
rect 23660 13806 23662 13858
rect 23714 13806 23716 13858
rect 23660 13794 23716 13806
rect 23884 14644 23940 14654
rect 23884 13858 23940 14588
rect 23884 13806 23886 13858
rect 23938 13806 23940 13858
rect 23436 13570 23492 13580
rect 23548 13634 23604 13646
rect 23548 13582 23550 13634
rect 23602 13582 23604 13634
rect 21980 12348 22260 12404
rect 22540 13524 22596 13534
rect 21868 11732 21924 11742
rect 21756 11676 21868 11732
rect 21532 11396 21588 11406
rect 21532 11302 21588 11340
rect 21868 11282 21924 11676
rect 21868 11230 21870 11282
rect 21922 11230 21924 11282
rect 21868 11218 21924 11230
rect 21420 9884 21812 9940
rect 21420 9714 21476 9884
rect 21420 9662 21422 9714
rect 21474 9662 21476 9714
rect 21420 9650 21476 9662
rect 21532 9714 21588 9726
rect 21532 9662 21534 9714
rect 21586 9662 21588 9714
rect 21196 9602 21252 9614
rect 21196 9550 21198 9602
rect 21250 9550 21252 9602
rect 20636 9156 20692 9166
rect 21196 9156 21252 9550
rect 21532 9268 21588 9662
rect 21532 9202 21588 9212
rect 20636 9154 21252 9156
rect 20636 9102 20638 9154
rect 20690 9102 21252 9154
rect 20636 9100 21252 9102
rect 20636 9090 20692 9100
rect 21196 9044 21252 9100
rect 21196 8988 21476 9044
rect 20076 8930 20244 8932
rect 20076 8878 20078 8930
rect 20130 8878 20244 8930
rect 20076 8876 20244 8878
rect 20076 8484 20132 8876
rect 19180 8418 19236 8428
rect 20076 8258 20132 8428
rect 20076 8206 20078 8258
rect 20130 8206 20132 8258
rect 20076 8194 20132 8206
rect 20524 8260 20580 8270
rect 20748 8260 20804 8270
rect 21308 8260 21364 8270
rect 20524 8258 20692 8260
rect 20524 8206 20526 8258
rect 20578 8206 20692 8258
rect 20524 8204 20692 8206
rect 20524 8194 20580 8204
rect 18284 7970 18340 7980
rect 20524 8036 20580 8046
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19404 7588 19460 7598
rect 19404 7494 19460 7532
rect 20300 7588 20356 7598
rect 16380 7422 16382 7474
rect 16434 7422 16436 7474
rect 16380 7410 16436 7422
rect 16604 7476 16660 7486
rect 18172 7476 18228 7486
rect 16604 7382 16660 7420
rect 17948 7420 18172 7476
rect 18228 7420 18452 7476
rect 15708 6748 16436 6804
rect 15260 6290 15316 6300
rect 16156 6580 16212 6590
rect 13804 6018 13972 6020
rect 13804 5966 13806 6018
rect 13858 5966 13972 6018
rect 13804 5964 13972 5966
rect 16156 6018 16212 6524
rect 16268 6130 16324 6748
rect 16380 6690 16436 6748
rect 16380 6638 16382 6690
rect 16434 6638 16436 6690
rect 16380 6626 16436 6638
rect 16492 6802 16548 6814
rect 16492 6750 16494 6802
rect 16546 6750 16548 6802
rect 16492 6692 16548 6750
rect 16492 6626 16548 6636
rect 17276 6692 17332 6702
rect 17948 6692 18004 7420
rect 18172 7382 18228 7420
rect 18060 6804 18116 6842
rect 18060 6738 18116 6748
rect 17276 6598 17332 6636
rect 17836 6690 18004 6692
rect 17836 6638 17950 6690
rect 18002 6638 18004 6690
rect 17836 6636 18004 6638
rect 18396 6692 18452 7420
rect 18620 7474 18676 7486
rect 18620 7422 18622 7474
rect 18674 7422 18676 7474
rect 18508 6692 18564 6702
rect 18396 6690 18564 6692
rect 18396 6638 18510 6690
rect 18562 6638 18564 6690
rect 18396 6636 18564 6638
rect 16268 6078 16270 6130
rect 16322 6078 16324 6130
rect 16268 6066 16324 6078
rect 16492 6468 16548 6478
rect 16492 6130 16548 6412
rect 17724 6468 17780 6478
rect 17724 6374 17780 6412
rect 16492 6078 16494 6130
rect 16546 6078 16548 6130
rect 16492 6066 16548 6078
rect 16156 5966 16158 6018
rect 16210 5966 16212 6018
rect 13804 5954 13860 5964
rect 16156 5954 16212 5966
rect 13132 5854 13134 5906
rect 13186 5854 13188 5906
rect 13132 5842 13188 5854
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 17836 5236 17892 6636
rect 17948 6626 18004 6636
rect 18508 6626 18564 6636
rect 18620 6692 18676 7422
rect 19964 7476 20020 7486
rect 19964 7382 20020 7420
rect 20300 7474 20356 7532
rect 20300 7422 20302 7474
rect 20354 7422 20356 7474
rect 20300 7410 20356 7422
rect 20524 7586 20580 7980
rect 20524 7534 20526 7586
rect 20578 7534 20580 7586
rect 18732 7364 18788 7374
rect 18732 7362 19236 7364
rect 18732 7310 18734 7362
rect 18786 7310 19236 7362
rect 18732 7308 19236 7310
rect 18732 7298 18788 7308
rect 18732 6692 18788 6702
rect 18620 6636 18732 6692
rect 18172 6468 18228 6478
rect 18620 6468 18676 6636
rect 18732 6598 18788 6636
rect 18172 6466 18676 6468
rect 18172 6414 18174 6466
rect 18226 6414 18676 6466
rect 18172 6412 18676 6414
rect 19068 6466 19124 6478
rect 19068 6414 19070 6466
rect 19122 6414 19124 6466
rect 18172 6402 18228 6412
rect 19068 5906 19124 6414
rect 19068 5854 19070 5906
rect 19122 5854 19124 5906
rect 19068 5842 19124 5854
rect 18396 5796 18452 5806
rect 17948 5236 18004 5246
rect 17836 5234 18004 5236
rect 17836 5182 17950 5234
rect 18002 5182 18004 5234
rect 17836 5180 18004 5182
rect 17948 5170 18004 5180
rect 18396 5010 18452 5740
rect 19180 5794 19236 7308
rect 20524 7252 20580 7534
rect 20300 7196 20580 7252
rect 19180 5742 19182 5794
rect 19234 5742 19236 5794
rect 19180 5730 19236 5742
rect 19404 6692 19460 6702
rect 19404 5122 19460 6636
rect 19852 6580 19908 6590
rect 20188 6580 20244 6590
rect 19852 6578 20244 6580
rect 19852 6526 19854 6578
rect 19906 6526 20190 6578
rect 20242 6526 20244 6578
rect 19852 6524 20244 6526
rect 19852 6514 19908 6524
rect 20188 6468 20244 6524
rect 20300 6578 20356 7196
rect 20300 6526 20302 6578
rect 20354 6526 20356 6578
rect 20300 6514 20356 6526
rect 20524 6692 20580 6702
rect 20188 6402 20244 6412
rect 20524 6466 20580 6636
rect 20524 6414 20526 6466
rect 20578 6414 20580 6466
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 20524 5572 20580 6414
rect 20636 5908 20692 8204
rect 20748 8258 21364 8260
rect 20748 8206 20750 8258
rect 20802 8206 21310 8258
rect 21362 8206 21364 8258
rect 20748 8204 21364 8206
rect 21420 8260 21476 8988
rect 21644 9042 21700 9054
rect 21644 8990 21646 9042
rect 21698 8990 21700 9042
rect 21532 8260 21588 8270
rect 21420 8258 21588 8260
rect 21420 8206 21534 8258
rect 21586 8206 21588 8258
rect 21420 8204 21588 8206
rect 20748 8194 20804 8204
rect 21308 8194 21364 8204
rect 21532 8194 21588 8204
rect 20860 7362 20916 7374
rect 20860 7310 20862 7362
rect 20914 7310 20916 7362
rect 20748 5908 20804 5918
rect 20636 5852 20748 5908
rect 20524 5506 20580 5516
rect 20748 5346 20804 5852
rect 20860 5906 20916 7310
rect 20860 5854 20862 5906
rect 20914 5854 20916 5906
rect 20860 5796 20916 5854
rect 21644 5908 21700 8990
rect 21756 8260 21812 9884
rect 21756 8194 21812 8204
rect 21868 8484 21924 8494
rect 21644 5814 21700 5852
rect 20860 5730 20916 5740
rect 21868 5794 21924 8428
rect 21868 5742 21870 5794
rect 21922 5742 21924 5794
rect 21868 5730 21924 5742
rect 20748 5294 20750 5346
rect 20802 5294 20804 5346
rect 20748 5282 20804 5294
rect 21868 5572 21924 5582
rect 21868 5234 21924 5516
rect 21868 5182 21870 5234
rect 21922 5182 21924 5234
rect 21868 5170 21924 5182
rect 19404 5070 19406 5122
rect 19458 5070 19460 5122
rect 19404 5058 19460 5070
rect 18396 4958 18398 5010
rect 18450 4958 18452 5010
rect 18396 4946 18452 4958
rect 21980 4900 22036 12348
rect 22092 12178 22148 12190
rect 22092 12126 22094 12178
rect 22146 12126 22148 12178
rect 22092 11170 22148 12126
rect 22540 12178 22596 13468
rect 23548 13076 23604 13582
rect 23884 13524 23940 13806
rect 23884 13458 23940 13468
rect 23996 13188 24052 15092
rect 24108 13748 24164 13758
rect 24108 13654 24164 13692
rect 24052 13132 24164 13188
rect 23996 13122 24052 13132
rect 23548 13020 23940 13076
rect 23324 12964 23380 12974
rect 23324 12962 23828 12964
rect 23324 12910 23326 12962
rect 23378 12910 23828 12962
rect 23324 12908 23828 12910
rect 23324 12898 23380 12908
rect 23100 12850 23156 12862
rect 23100 12798 23102 12850
rect 23154 12798 23156 12850
rect 23100 12740 23156 12798
rect 22540 12126 22542 12178
rect 22594 12126 22596 12178
rect 22540 11844 22596 12126
rect 22988 12178 23044 12190
rect 22988 12126 22990 12178
rect 23042 12126 23044 12178
rect 22988 12068 23044 12126
rect 22540 11788 22932 11844
rect 22428 11284 22484 11294
rect 22428 11282 22820 11284
rect 22428 11230 22430 11282
rect 22482 11230 22820 11282
rect 22428 11228 22820 11230
rect 22428 11218 22484 11228
rect 22092 11118 22094 11170
rect 22146 11118 22148 11170
rect 22092 11060 22148 11118
rect 22092 11004 22708 11060
rect 22652 10610 22708 11004
rect 22652 10558 22654 10610
rect 22706 10558 22708 10610
rect 22652 10546 22708 10558
rect 22092 9044 22148 9054
rect 22092 8370 22148 8988
rect 22092 8318 22094 8370
rect 22146 8318 22148 8370
rect 22092 8306 22148 8318
rect 22764 8372 22820 11228
rect 22876 10610 22932 11788
rect 22876 10558 22878 10610
rect 22930 10558 22932 10610
rect 22876 10546 22932 10558
rect 22876 9156 22932 9166
rect 22988 9156 23044 12012
rect 23100 11956 23156 12684
rect 23324 12292 23380 12302
rect 23324 12198 23380 12236
rect 23100 11890 23156 11900
rect 23772 12178 23828 12908
rect 23772 12126 23774 12178
rect 23826 12126 23828 12178
rect 23772 11508 23828 12126
rect 23884 11732 23940 13020
rect 23996 12962 24052 12974
rect 23996 12910 23998 12962
rect 24050 12910 24052 12962
rect 23996 12068 24052 12910
rect 23996 11974 24052 12012
rect 23884 11676 24052 11732
rect 23884 11508 23940 11518
rect 23212 11506 23940 11508
rect 23212 11454 23886 11506
rect 23938 11454 23940 11506
rect 23212 11452 23940 11454
rect 23212 10834 23268 11452
rect 23884 11442 23940 11452
rect 23212 10782 23214 10834
rect 23266 10782 23268 10834
rect 23212 10770 23268 10782
rect 23996 10724 24052 11676
rect 23660 10668 24052 10724
rect 23436 9940 23492 9950
rect 23436 9826 23492 9884
rect 23436 9774 23438 9826
rect 23490 9774 23492 9826
rect 23436 9762 23492 9774
rect 23660 9828 23716 10668
rect 23660 9714 23716 9772
rect 23660 9662 23662 9714
rect 23714 9662 23716 9714
rect 23660 9650 23716 9662
rect 23996 10052 24052 10062
rect 22876 9154 23044 9156
rect 22876 9102 22878 9154
rect 22930 9102 23044 9154
rect 22876 9100 23044 9102
rect 22876 9090 22932 9100
rect 23660 9044 23716 9054
rect 23660 8950 23716 8988
rect 23996 8930 24052 9996
rect 24108 9940 24164 13132
rect 24332 12404 24388 16380
rect 25116 16100 25172 16110
rect 25116 16006 25172 16044
rect 25228 15986 25284 18620
rect 25340 18452 25396 18462
rect 25340 17444 25396 18396
rect 25452 17666 25508 18844
rect 25676 18450 25732 18462
rect 25676 18398 25678 18450
rect 25730 18398 25732 18450
rect 25676 17892 25732 18398
rect 25788 18340 25844 19070
rect 26572 18676 26628 20076
rect 26572 18582 26628 18620
rect 26684 19122 26740 19134
rect 26684 19070 26686 19122
rect 26738 19070 26740 19122
rect 25788 18274 25844 18284
rect 26012 18450 26068 18462
rect 26012 18398 26014 18450
rect 26066 18398 26068 18450
rect 26012 17892 26068 18398
rect 26236 18452 26292 18462
rect 26684 18452 26740 19070
rect 26236 18450 26740 18452
rect 26236 18398 26238 18450
rect 26290 18398 26740 18450
rect 26236 18396 26740 18398
rect 26796 19010 26852 19022
rect 26796 18958 26798 19010
rect 26850 18958 26852 19010
rect 26796 18452 26852 18958
rect 27020 19012 27076 19022
rect 27020 18918 27076 18956
rect 26236 18386 26292 18396
rect 26796 18386 26852 18396
rect 26908 18562 26964 18574
rect 26908 18510 26910 18562
rect 26962 18510 26964 18562
rect 26908 18340 26964 18510
rect 25676 17836 25956 17892
rect 25452 17614 25454 17666
rect 25506 17614 25508 17666
rect 25452 17602 25508 17614
rect 25788 17668 25844 17678
rect 25900 17668 25956 17836
rect 26012 17826 26068 17836
rect 26124 17890 26180 17902
rect 26124 17838 26126 17890
rect 26178 17838 26180 17890
rect 26124 17668 26180 17838
rect 25900 17612 26180 17668
rect 25788 17574 25844 17612
rect 25340 17388 25620 17444
rect 25564 16994 25620 17388
rect 25564 16942 25566 16994
rect 25618 16942 25620 16994
rect 25564 16930 25620 16942
rect 26124 16882 26180 17612
rect 26796 17892 26852 17902
rect 26572 16884 26628 16894
rect 26124 16830 26126 16882
rect 26178 16830 26180 16882
rect 25788 16100 25844 16110
rect 25228 15934 25230 15986
rect 25282 15934 25284 15986
rect 25228 15922 25284 15934
rect 25340 16098 25844 16100
rect 25340 16046 25790 16098
rect 25842 16046 25844 16098
rect 25340 16044 25844 16046
rect 24668 15204 24724 15242
rect 24668 15138 24724 15148
rect 25340 15148 25396 16044
rect 25788 16034 25844 16044
rect 26012 16098 26068 16110
rect 26012 16046 26014 16098
rect 26066 16046 26068 16098
rect 25452 15874 25508 15886
rect 25452 15822 25454 15874
rect 25506 15822 25508 15874
rect 25452 15540 25508 15822
rect 26012 15764 26068 16046
rect 26012 15698 26068 15708
rect 25452 15474 25508 15484
rect 26012 15540 26068 15550
rect 26012 15426 26068 15484
rect 26012 15374 26014 15426
rect 26066 15374 26068 15426
rect 26012 15362 26068 15374
rect 25564 15316 25620 15326
rect 25564 15148 25620 15260
rect 25340 15092 25620 15148
rect 25004 14532 25060 14542
rect 24556 14530 25060 14532
rect 24556 14478 25006 14530
rect 25058 14478 25060 14530
rect 24556 14476 25060 14478
rect 24556 13970 24612 14476
rect 25004 14466 25060 14476
rect 24556 13918 24558 13970
rect 24610 13918 24612 13970
rect 24556 13906 24612 13918
rect 24668 12850 24724 12862
rect 24668 12798 24670 12850
rect 24722 12798 24724 12850
rect 24668 12740 24724 12798
rect 24668 12674 24724 12684
rect 24332 12348 24500 12404
rect 24332 12180 24388 12190
rect 24332 12086 24388 12124
rect 24332 11956 24388 11966
rect 24332 11394 24388 11900
rect 24332 11342 24334 11394
rect 24386 11342 24388 11394
rect 24332 11330 24388 11342
rect 24444 10388 24500 12348
rect 25452 12180 25508 12190
rect 25452 12086 25508 12124
rect 25340 12068 25396 12078
rect 25340 11394 25396 12012
rect 25564 11618 25620 15092
rect 25900 15204 25956 15214
rect 25900 14530 25956 15148
rect 25900 14478 25902 14530
rect 25954 14478 25956 14530
rect 25900 14466 25956 14478
rect 26124 14532 26180 16830
rect 26460 16828 26572 16884
rect 26460 15876 26516 16828
rect 26572 16818 26628 16828
rect 26796 16882 26852 17836
rect 26796 16830 26798 16882
rect 26850 16830 26852 16882
rect 26796 16436 26852 16830
rect 26908 16884 26964 18284
rect 27132 18004 27188 20300
rect 27244 18788 27300 20524
rect 27468 20018 27524 20030
rect 27468 19966 27470 20018
rect 27522 19966 27524 20018
rect 27468 19236 27524 19966
rect 28028 19906 28084 20862
rect 28252 20132 28308 22318
rect 28252 20038 28308 20076
rect 28364 21362 28420 21374
rect 28364 21310 28366 21362
rect 28418 21310 28420 21362
rect 28028 19854 28030 19906
rect 28082 19854 28084 19906
rect 27804 19460 27860 19470
rect 28028 19460 28084 19854
rect 27804 19458 28084 19460
rect 27804 19406 27806 19458
rect 27858 19406 28084 19458
rect 27804 19404 28084 19406
rect 28140 20018 28196 20030
rect 28140 19966 28142 20018
rect 28194 19966 28196 20018
rect 27804 19394 27860 19404
rect 27580 19236 27636 19246
rect 27468 19234 27636 19236
rect 27468 19182 27582 19234
rect 27634 19182 27636 19234
rect 27468 19180 27636 19182
rect 27244 18732 27412 18788
rect 27356 18452 27412 18732
rect 27468 18676 27524 19180
rect 27580 19170 27636 19180
rect 28028 19236 28084 19246
rect 28140 19236 28196 19966
rect 28084 19180 28196 19236
rect 28028 19142 28084 19180
rect 27692 19012 27748 19022
rect 28364 19012 28420 21310
rect 27692 19010 28420 19012
rect 27692 18958 27694 19010
rect 27746 18958 28420 19010
rect 27692 18956 28420 18958
rect 27692 18946 27748 18956
rect 27468 18620 27636 18676
rect 27356 18386 27412 18396
rect 27468 18450 27524 18462
rect 27468 18398 27470 18450
rect 27522 18398 27524 18450
rect 27468 18340 27524 18398
rect 27468 18274 27524 18284
rect 27356 18228 27412 18238
rect 27244 18004 27300 18014
rect 27132 17948 27244 18004
rect 27244 17938 27300 17948
rect 26908 16818 26964 16828
rect 26236 15820 26516 15876
rect 26572 16380 26852 16436
rect 26236 14756 26292 15820
rect 26348 15652 26404 15662
rect 26348 15314 26404 15596
rect 26348 15262 26350 15314
rect 26402 15262 26404 15314
rect 26348 14868 26404 15262
rect 26460 15204 26516 15214
rect 26572 15204 26628 16380
rect 26684 16100 26740 16110
rect 27020 16100 27076 16110
rect 26684 16098 27076 16100
rect 26684 16046 26686 16098
rect 26738 16046 27022 16098
rect 27074 16046 27076 16098
rect 26684 16044 27076 16046
rect 26684 16034 26740 16044
rect 27020 16034 27076 16044
rect 27244 15316 27300 15326
rect 27244 15222 27300 15260
rect 26516 15148 26628 15204
rect 26460 15138 26516 15148
rect 26348 14812 26628 14868
rect 26236 14700 26516 14756
rect 26348 14532 26404 14542
rect 26124 14530 26404 14532
rect 26124 14478 26350 14530
rect 26402 14478 26404 14530
rect 26124 14476 26404 14478
rect 26348 14466 26404 14476
rect 26348 13972 26404 13982
rect 26460 13972 26516 14700
rect 26572 14644 26628 14812
rect 26908 14644 26964 14654
rect 26572 14642 26964 14644
rect 26572 14590 26910 14642
rect 26962 14590 26964 14642
rect 26572 14588 26964 14590
rect 25900 13970 26516 13972
rect 25900 13918 26350 13970
rect 26402 13918 26516 13970
rect 25900 13916 26516 13918
rect 25788 12850 25844 12862
rect 25788 12798 25790 12850
rect 25842 12798 25844 12850
rect 25788 12516 25844 12798
rect 25900 12850 25956 13916
rect 26348 13906 26404 13916
rect 26572 13860 26628 13870
rect 26628 13804 26740 13860
rect 26572 13766 26628 13804
rect 26236 13746 26292 13758
rect 26236 13694 26238 13746
rect 26290 13694 26292 13746
rect 25900 12798 25902 12850
rect 25954 12798 25956 12850
rect 25900 12786 25956 12798
rect 26124 12852 26180 12862
rect 26124 12758 26180 12796
rect 25788 12460 26068 12516
rect 25564 11566 25566 11618
rect 25618 11566 25620 11618
rect 25564 11554 25620 11566
rect 25900 12292 25956 12302
rect 25900 12066 25956 12236
rect 25900 12014 25902 12066
rect 25954 12014 25956 12066
rect 25340 11342 25342 11394
rect 25394 11342 25396 11394
rect 25340 11330 25396 11342
rect 24444 10332 24724 10388
rect 24108 9874 24164 9884
rect 24332 9716 24388 9726
rect 23996 8878 23998 8930
rect 24050 8878 24052 8930
rect 23996 8866 24052 8878
rect 24108 9602 24164 9614
rect 24108 9550 24110 9602
rect 24162 9550 24164 9602
rect 22876 8372 22932 8382
rect 22764 8316 22876 8372
rect 22876 8278 22932 8316
rect 24108 8370 24164 9550
rect 24220 9602 24276 9614
rect 24220 9550 24222 9602
rect 24274 9550 24276 9602
rect 24220 9044 24276 9550
rect 24220 8978 24276 8988
rect 24332 8930 24388 9660
rect 24556 9602 24612 9614
rect 24556 9550 24558 9602
rect 24610 9550 24612 9602
rect 24332 8878 24334 8930
rect 24386 8878 24388 8930
rect 24332 8866 24388 8878
rect 24444 9042 24500 9054
rect 24444 8990 24446 9042
rect 24498 8990 24500 9042
rect 24108 8318 24110 8370
rect 24162 8318 24164 8370
rect 24108 8306 24164 8318
rect 22428 8260 22484 8270
rect 22428 8166 22484 8204
rect 23436 8260 23492 8270
rect 23436 8146 23492 8204
rect 24444 8260 24500 8990
rect 23436 8094 23438 8146
rect 23490 8094 23492 8146
rect 23436 8082 23492 8094
rect 23548 8146 23604 8158
rect 23548 8094 23550 8146
rect 23602 8094 23604 8146
rect 23212 8036 23268 8046
rect 22764 8034 23268 8036
rect 22764 7982 23214 8034
rect 23266 7982 23268 8034
rect 22764 7980 23268 7982
rect 22764 7474 22820 7980
rect 23212 7970 23268 7980
rect 22764 7422 22766 7474
rect 22818 7422 22820 7474
rect 22764 7410 22820 7422
rect 23548 7476 23604 8094
rect 24444 7586 24500 8204
rect 24556 8146 24612 9550
rect 24556 8094 24558 8146
rect 24610 8094 24612 8146
rect 24556 8082 24612 8094
rect 24444 7534 24446 7586
rect 24498 7534 24500 7586
rect 24444 7522 24500 7534
rect 23548 7410 23604 7420
rect 24108 7474 24164 7486
rect 24108 7422 24110 7474
rect 24162 7422 24164 7474
rect 22428 7362 22484 7374
rect 22428 7310 22430 7362
rect 22482 7310 22484 7362
rect 22204 6804 22260 6842
rect 22092 6692 22148 6702
rect 22092 6598 22148 6636
rect 22092 5348 22148 5358
rect 22204 5348 22260 6748
rect 22428 6580 22484 7310
rect 23996 6804 24052 6814
rect 23996 6710 24052 6748
rect 22540 6692 22596 6702
rect 22988 6692 23044 6702
rect 22540 6598 22596 6636
rect 22652 6690 23044 6692
rect 22652 6638 22990 6690
rect 23042 6638 23044 6690
rect 22652 6636 23044 6638
rect 22428 6356 22484 6524
rect 22316 6300 22484 6356
rect 22316 5682 22372 6300
rect 22652 5796 22708 6636
rect 22988 6626 23044 6636
rect 24108 6692 24164 7422
rect 24556 6692 24612 6702
rect 24164 6690 24612 6692
rect 24164 6638 24558 6690
rect 24610 6638 24612 6690
rect 24164 6636 24612 6638
rect 24108 6598 24164 6636
rect 24556 6626 24612 6636
rect 23660 6580 23716 6590
rect 23660 6486 23716 6524
rect 22316 5630 22318 5682
rect 22370 5630 22372 5682
rect 22316 5618 22372 5630
rect 22428 5740 22708 5796
rect 22092 5346 22260 5348
rect 22092 5294 22094 5346
rect 22146 5294 22260 5346
rect 22092 5292 22260 5294
rect 22428 5346 22484 5740
rect 22428 5294 22430 5346
rect 22482 5294 22484 5346
rect 22092 5282 22148 5292
rect 22428 5282 22484 5294
rect 21980 4844 22596 4900
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 22204 3444 22260 3482
rect 22428 3444 22484 3454
rect 22204 3442 22484 3444
rect 22204 3390 22206 3442
rect 22258 3390 22430 3442
rect 22482 3390 22484 3442
rect 22204 3388 22484 3390
rect 22540 3444 22596 4844
rect 22764 3444 22820 3454
rect 22540 3442 22820 3444
rect 22540 3390 22766 3442
rect 22818 3390 22820 3442
rect 22540 3388 22820 3390
rect 19740 3332 19796 3342
rect 19516 3330 19796 3332
rect 19516 3278 19742 3330
rect 19794 3278 19796 3330
rect 19516 3276 19796 3278
rect 19516 800 19572 3276
rect 19740 3266 19796 3276
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 22204 800 22260 3388
rect 22428 3378 22484 3388
rect 22764 3378 22820 3388
rect 24556 3444 24612 3454
rect 24668 3444 24724 10332
rect 25452 10052 25508 10062
rect 24780 9940 24836 9950
rect 24780 9714 24836 9884
rect 24780 9662 24782 9714
rect 24834 9662 24836 9714
rect 24780 9650 24836 9662
rect 24892 9714 24948 9726
rect 24892 9662 24894 9714
rect 24946 9662 24948 9714
rect 24892 9268 24948 9662
rect 24892 9202 24948 9212
rect 25228 9044 25284 9054
rect 25228 8950 25284 8988
rect 25452 9042 25508 9996
rect 25900 10052 25956 12014
rect 25900 9986 25956 9996
rect 25900 9828 25956 9838
rect 25900 9734 25956 9772
rect 26012 9714 26068 12460
rect 26236 11732 26292 13694
rect 26684 12850 26740 13804
rect 26684 12798 26686 12850
rect 26738 12798 26740 12850
rect 26684 12786 26740 12798
rect 26908 12292 26964 14588
rect 27244 14532 27300 14542
rect 26908 12226 26964 12236
rect 27132 14476 27244 14532
rect 27020 12180 27076 12190
rect 27020 12086 27076 12124
rect 26236 11666 26292 11676
rect 27020 11394 27076 11406
rect 27020 11342 27022 11394
rect 27074 11342 27076 11394
rect 26908 10052 26964 10062
rect 27020 10052 27076 11342
rect 26908 10050 27076 10052
rect 26908 9998 26910 10050
rect 26962 9998 27076 10050
rect 26908 9996 27076 9998
rect 26908 9986 26964 9996
rect 26460 9828 26516 9838
rect 26348 9826 26516 9828
rect 26348 9774 26462 9826
rect 26514 9774 26516 9826
rect 26348 9772 26516 9774
rect 26012 9662 26014 9714
rect 26066 9662 26068 9714
rect 26012 9268 26068 9662
rect 26236 9716 26292 9726
rect 26236 9622 26292 9660
rect 26348 9380 26404 9772
rect 26460 9762 26516 9772
rect 26908 9828 26964 9838
rect 26012 9202 26068 9212
rect 26124 9324 26404 9380
rect 26124 9266 26180 9324
rect 26124 9214 26126 9266
rect 26178 9214 26180 9266
rect 26124 9202 26180 9214
rect 25452 8990 25454 9042
rect 25506 8990 25508 9042
rect 25452 8978 25508 8990
rect 25676 8818 25732 8830
rect 25676 8766 25678 8818
rect 25730 8766 25732 8818
rect 25564 8260 25620 8270
rect 25676 8260 25732 8766
rect 26908 8482 26964 9772
rect 26908 8430 26910 8482
rect 26962 8430 26964 8482
rect 26908 8418 26964 8430
rect 25620 8204 25732 8260
rect 26572 8372 26628 8382
rect 25564 8166 25620 8204
rect 25340 7700 25396 7710
rect 25676 7700 25732 7710
rect 25340 7698 25732 7700
rect 25340 7646 25342 7698
rect 25394 7646 25678 7698
rect 25730 7646 25732 7698
rect 25340 7644 25732 7646
rect 24780 6690 24836 6702
rect 24780 6638 24782 6690
rect 24834 6638 24836 6690
rect 24780 6580 24836 6638
rect 24780 6514 24836 6524
rect 25340 6468 25396 7644
rect 25676 7634 25732 7644
rect 26012 7586 26068 7598
rect 26012 7534 26014 7586
rect 26066 7534 26068 7586
rect 25452 7476 25508 7486
rect 25452 6690 25508 7420
rect 26012 7364 26068 7534
rect 26572 7588 26628 8316
rect 26796 8148 26852 8158
rect 26796 7698 26852 8092
rect 26796 7646 26798 7698
rect 26850 7646 26852 7698
rect 26796 7634 26852 7646
rect 26572 7494 26628 7532
rect 26012 7298 26068 7308
rect 26348 7474 26404 7486
rect 26348 7422 26350 7474
rect 26402 7422 26404 7474
rect 26348 6804 26404 7422
rect 27020 7476 27076 7486
rect 27132 7476 27188 14476
rect 27244 14466 27300 14476
rect 27356 14196 27412 18172
rect 27468 16996 27524 17006
rect 27580 16996 27636 18620
rect 27692 18562 27748 18574
rect 27692 18510 27694 18562
rect 27746 18510 27748 18562
rect 27692 18452 27748 18510
rect 28252 18564 28308 18574
rect 27748 18396 28196 18452
rect 27692 18386 27748 18396
rect 27468 16994 27636 16996
rect 27468 16942 27470 16994
rect 27522 16942 27636 16994
rect 27468 16940 27636 16942
rect 28140 17108 28196 18396
rect 27468 16930 27524 16940
rect 28028 16884 28084 16922
rect 28028 16818 28084 16828
rect 28028 16660 28084 16670
rect 28028 16210 28084 16604
rect 28028 16158 28030 16210
rect 28082 16158 28084 16210
rect 28028 16146 28084 16158
rect 27580 16100 27636 16110
rect 27580 16006 27636 16044
rect 28140 15986 28196 17052
rect 28140 15934 28142 15986
rect 28194 15934 28196 15986
rect 28140 15922 28196 15934
rect 28252 18450 28308 18508
rect 28252 18398 28254 18450
rect 28306 18398 28308 18450
rect 27916 15428 27972 15438
rect 28252 15428 28308 18398
rect 28364 18228 28420 18238
rect 28476 18228 28532 23996
rect 28700 22484 28756 27916
rect 28924 27748 28980 28364
rect 28700 22418 28756 22428
rect 28812 27746 28980 27748
rect 28812 27694 28926 27746
rect 28978 27694 28980 27746
rect 28812 27692 28980 27694
rect 28812 26180 28868 27692
rect 28924 27682 28980 27692
rect 29148 26908 29204 29260
rect 29484 29204 29540 29708
rect 29372 29148 29540 29204
rect 29260 28756 29316 28766
rect 29372 28756 29428 29148
rect 29260 28754 29428 28756
rect 29260 28702 29262 28754
rect 29314 28702 29428 28754
rect 29260 28700 29428 28702
rect 29260 27748 29316 28700
rect 29484 28644 29540 28654
rect 29372 27972 29428 27982
rect 29372 27878 29428 27916
rect 29484 27860 29540 28588
rect 29596 28644 29652 30270
rect 29708 29764 29764 31724
rect 29820 31714 29876 31724
rect 29820 29988 29876 29998
rect 30268 29988 30324 35756
rect 30380 35588 30436 38612
rect 30492 37828 30548 40684
rect 31052 39844 31108 41356
rect 32172 41300 32228 41310
rect 32060 41298 32228 41300
rect 32060 41246 32174 41298
rect 32226 41246 32228 41298
rect 32060 41244 32228 41246
rect 31948 41188 32004 41198
rect 31948 41094 32004 41132
rect 31164 41076 31220 41086
rect 31164 41074 31668 41076
rect 31164 41022 31166 41074
rect 31218 41022 31668 41074
rect 31164 41020 31668 41022
rect 31164 41010 31220 41020
rect 31052 39778 31108 39788
rect 31612 39842 31668 41020
rect 31836 40964 31892 40974
rect 31836 40870 31892 40908
rect 32060 40404 32116 41244
rect 32172 41234 32228 41244
rect 32284 41188 32340 42140
rect 32396 41972 32452 42702
rect 32396 41906 32452 41916
rect 32956 43372 33236 43428
rect 32284 41094 32340 41132
rect 32508 40964 32564 40974
rect 32564 40908 32900 40964
rect 32508 40870 32564 40908
rect 31612 39790 31614 39842
rect 31666 39790 31668 39842
rect 31612 39778 31668 39790
rect 31836 40348 32116 40404
rect 30828 39618 30884 39630
rect 30828 39566 30830 39618
rect 30882 39566 30884 39618
rect 30828 39060 30884 39566
rect 30828 38994 30884 39004
rect 30940 39506 30996 39518
rect 30940 39454 30942 39506
rect 30994 39454 30996 39506
rect 30940 38668 30996 39454
rect 31164 39060 31220 39070
rect 31164 38966 31220 39004
rect 30940 38612 31108 38668
rect 30492 37156 30548 37772
rect 30492 37090 30548 37100
rect 30940 37492 30996 37502
rect 30940 36482 30996 37436
rect 30940 36430 30942 36482
rect 30994 36430 30996 36482
rect 30940 35700 30996 36430
rect 30716 35644 30996 35700
rect 30492 35588 30548 35598
rect 30380 35586 30548 35588
rect 30380 35534 30494 35586
rect 30546 35534 30548 35586
rect 30380 35532 30548 35534
rect 30380 35028 30436 35532
rect 30492 35522 30548 35532
rect 30380 34962 30436 34972
rect 30492 35028 30548 35038
rect 30716 35028 30772 35644
rect 31052 35588 31108 38612
rect 31612 37492 31668 37502
rect 31612 37398 31668 37436
rect 31164 37156 31220 37166
rect 31164 37062 31220 37100
rect 31612 36372 31668 36382
rect 31612 36278 31668 36316
rect 30492 35026 30772 35028
rect 30492 34974 30494 35026
rect 30546 34974 30772 35026
rect 30492 34972 30772 34974
rect 30492 34962 30548 34972
rect 30604 34804 30660 34814
rect 30604 33570 30660 34748
rect 30716 34130 30772 34972
rect 30940 35532 31108 35588
rect 30940 35026 30996 35532
rect 30940 34974 30942 35026
rect 30994 34974 30996 35026
rect 30940 34962 30996 34974
rect 31052 35028 31108 35038
rect 30828 34804 30884 34814
rect 31052 34804 31108 34972
rect 30828 34802 31108 34804
rect 30828 34750 30830 34802
rect 30882 34750 31108 34802
rect 30828 34748 31108 34750
rect 31164 34802 31220 34814
rect 31164 34750 31166 34802
rect 31218 34750 31220 34802
rect 30828 34738 30884 34748
rect 31164 34244 31220 34750
rect 31388 34802 31444 34814
rect 31388 34750 31390 34802
rect 31442 34750 31444 34802
rect 31276 34244 31332 34254
rect 30716 34078 30718 34130
rect 30770 34078 30772 34130
rect 30716 34066 30772 34078
rect 31052 34242 31332 34244
rect 31052 34190 31278 34242
rect 31330 34190 31332 34242
rect 31052 34188 31332 34190
rect 30604 33518 30606 33570
rect 30658 33518 30660 33570
rect 30604 33506 30660 33518
rect 30492 33234 30548 33246
rect 30492 33182 30494 33234
rect 30546 33182 30548 33234
rect 30492 32900 30548 33182
rect 30604 33236 30660 33246
rect 31052 33236 31108 34188
rect 31276 34132 31332 34188
rect 31276 34066 31332 34076
rect 31388 33796 31444 34750
rect 31612 34244 31668 34254
rect 31612 34150 31668 34188
rect 31388 33730 31444 33740
rect 31388 33348 31444 33358
rect 31612 33348 31668 33358
rect 31388 33346 31668 33348
rect 31388 33294 31390 33346
rect 31442 33294 31614 33346
rect 31666 33294 31668 33346
rect 31388 33292 31668 33294
rect 31388 33282 31444 33292
rect 31612 33282 31668 33292
rect 30604 33234 31108 33236
rect 30604 33182 30606 33234
rect 30658 33182 31054 33234
rect 31106 33182 31108 33234
rect 30604 33180 31108 33182
rect 30604 33170 30660 33180
rect 31052 33170 31108 33180
rect 31164 33236 31220 33246
rect 31164 33142 31220 33180
rect 30492 32834 30548 32844
rect 31052 32674 31108 32686
rect 31052 32622 31054 32674
rect 31106 32622 31108 32674
rect 30716 32562 30772 32574
rect 30716 32510 30718 32562
rect 30770 32510 30772 32562
rect 29820 29986 30324 29988
rect 29820 29934 29822 29986
rect 29874 29934 30324 29986
rect 29820 29932 30324 29934
rect 30380 32450 30436 32462
rect 30380 32398 30382 32450
rect 30434 32398 30436 32450
rect 29820 29922 29876 29932
rect 30380 29876 30436 32398
rect 30716 32004 30772 32510
rect 30716 31938 30772 31948
rect 31052 31778 31108 32622
rect 31500 32452 31556 32462
rect 31500 32358 31556 32396
rect 31836 31892 31892 40348
rect 32508 40292 32564 40302
rect 31948 40236 32508 40292
rect 31948 39842 32004 40236
rect 32508 40198 32564 40236
rect 31948 39790 31950 39842
rect 32002 39790 32004 39842
rect 31948 39778 32004 39790
rect 32732 39618 32788 39630
rect 32732 39566 32734 39618
rect 32786 39566 32788 39618
rect 32508 39508 32564 39518
rect 32284 39506 32564 39508
rect 32284 39454 32510 39506
rect 32562 39454 32564 39506
rect 32284 39452 32564 39454
rect 32172 36372 32228 36382
rect 32172 35922 32228 36316
rect 32172 35870 32174 35922
rect 32226 35870 32228 35922
rect 32172 35858 32228 35870
rect 31948 35586 32004 35598
rect 31948 35534 31950 35586
rect 32002 35534 32004 35586
rect 31948 35252 32004 35534
rect 32284 35364 32340 39452
rect 32508 39442 32564 39452
rect 32732 39060 32788 39566
rect 32396 38612 32452 38622
rect 32396 38050 32452 38556
rect 32396 37998 32398 38050
rect 32450 37998 32452 38050
rect 32396 37492 32452 37998
rect 32396 37426 32452 37436
rect 32732 37492 32788 39004
rect 32732 37426 32788 37436
rect 32844 36148 32900 40908
rect 32956 36820 33012 43372
rect 33180 43204 33236 43214
rect 33180 39956 33236 43148
rect 33292 42868 33348 44940
rect 33404 44940 33516 44996
rect 33404 44322 33460 44940
rect 33516 44902 33572 44940
rect 34524 44994 34580 45006
rect 34524 44942 34526 44994
rect 34578 44942 34580 44994
rect 33404 44270 33406 44322
rect 33458 44270 33460 44322
rect 33404 44258 33460 44270
rect 33516 44212 33572 44222
rect 33292 42802 33348 42812
rect 33404 43650 33460 43662
rect 33404 43598 33406 43650
rect 33458 43598 33460 43650
rect 33404 42196 33460 43598
rect 33516 42754 33572 44156
rect 34412 44212 34468 44222
rect 34524 44212 34580 44942
rect 34468 44156 34580 44212
rect 34412 44118 34468 44156
rect 33516 42702 33518 42754
rect 33570 42702 33572 42754
rect 33516 42690 33572 42702
rect 33628 43764 33684 43774
rect 33404 42140 33572 42196
rect 33404 41972 33460 41982
rect 33292 41860 33348 41870
rect 33292 41766 33348 41804
rect 33404 41298 33460 41916
rect 33404 41246 33406 41298
rect 33458 41246 33460 41298
rect 33404 41234 33460 41246
rect 33292 41188 33348 41198
rect 33292 41094 33348 41132
rect 33516 41076 33572 42140
rect 33628 41188 33684 43708
rect 34076 43652 34132 43662
rect 33852 43596 34076 43652
rect 33740 43540 33796 43550
rect 33740 42866 33796 43484
rect 33740 42814 33742 42866
rect 33794 42814 33796 42866
rect 33740 41860 33796 42814
rect 33852 42194 33908 43596
rect 34076 43558 34132 43596
rect 34748 43316 34804 45164
rect 34860 45220 34916 45230
rect 34860 45106 34916 45164
rect 34860 45054 34862 45106
rect 34914 45054 34916 45106
rect 34860 45042 34916 45054
rect 34972 45108 35028 46510
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 35308 46116 35364 46126
rect 35308 45890 35364 46060
rect 35308 45838 35310 45890
rect 35362 45838 35364 45890
rect 35308 45220 35364 45838
rect 35308 45154 35364 45164
rect 35532 45778 35588 47068
rect 35532 45726 35534 45778
rect 35586 45726 35588 45778
rect 34972 44436 35028 45052
rect 35532 44884 35588 45726
rect 35532 44818 35588 44828
rect 35644 44996 35700 47404
rect 35868 47348 35924 49196
rect 35980 48914 36036 49420
rect 36092 49028 36148 49038
rect 36316 49028 36372 49758
rect 36148 48972 36372 49028
rect 36652 49586 36708 49598
rect 36652 49534 36654 49586
rect 36706 49534 36708 49586
rect 36092 48934 36148 48972
rect 35980 48862 35982 48914
rect 36034 48862 36036 48914
rect 35980 48850 36036 48862
rect 36092 48804 36148 48814
rect 36540 48804 36596 48814
rect 36092 48356 36148 48748
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 35644 44548 35700 44940
rect 35756 47346 35924 47348
rect 35756 47294 35870 47346
rect 35922 47294 35924 47346
rect 35756 47292 35924 47294
rect 35756 44994 35812 47292
rect 35868 47282 35924 47292
rect 35980 48354 36148 48356
rect 35980 48302 36094 48354
rect 36146 48302 36148 48354
rect 35980 48300 36148 48302
rect 35756 44942 35758 44994
rect 35810 44942 35812 44994
rect 35756 44930 35812 44942
rect 35868 45890 35924 45902
rect 35868 45838 35870 45890
rect 35922 45838 35924 45890
rect 35756 44548 35812 44558
rect 35644 44546 35812 44548
rect 35644 44494 35758 44546
rect 35810 44494 35812 44546
rect 35644 44492 35812 44494
rect 35756 44482 35812 44492
rect 34972 44342 35028 44380
rect 35420 44434 35476 44446
rect 35420 44382 35422 44434
rect 35474 44382 35476 44434
rect 35420 43708 35476 44382
rect 35532 44436 35588 44446
rect 35532 44210 35588 44380
rect 35532 44158 35534 44210
rect 35586 44158 35588 44210
rect 35532 44146 35588 44158
rect 35868 43876 35924 45838
rect 35980 45668 36036 48300
rect 36092 48290 36148 48300
rect 36316 48802 36596 48804
rect 36316 48750 36542 48802
rect 36594 48750 36596 48802
rect 36316 48748 36596 48750
rect 36316 47458 36372 48748
rect 36540 48738 36596 48748
rect 36652 48242 36708 49534
rect 36764 49476 36820 50372
rect 36876 49924 36932 49934
rect 36876 49810 36932 49868
rect 36876 49758 36878 49810
rect 36930 49758 36932 49810
rect 36876 49746 36932 49758
rect 36764 49410 36820 49420
rect 36988 49028 37044 49038
rect 36988 48934 37044 48972
rect 36652 48190 36654 48242
rect 36706 48190 36708 48242
rect 36652 48178 36708 48190
rect 36764 48916 36820 48926
rect 36316 47406 36318 47458
rect 36370 47406 36372 47458
rect 36316 47394 36372 47406
rect 36540 46676 36596 46686
rect 36764 46676 36820 48860
rect 37100 48580 37156 50764
rect 37324 50594 37380 50606
rect 37324 50542 37326 50594
rect 37378 50542 37380 50594
rect 37324 49700 37380 50542
rect 37436 50484 37492 50764
rect 37548 50754 37604 50764
rect 37772 50708 37828 50718
rect 37884 50708 37940 51660
rect 37772 50706 37940 50708
rect 37772 50654 37774 50706
rect 37826 50654 37940 50706
rect 37772 50652 37940 50654
rect 37772 50596 37828 50652
rect 37772 50530 37828 50540
rect 37548 50484 37604 50494
rect 37436 50482 37604 50484
rect 37436 50430 37550 50482
rect 37602 50430 37604 50482
rect 37436 50428 37604 50430
rect 38108 50428 38164 55412
rect 38780 55076 38836 55086
rect 38780 54626 38836 55020
rect 38780 54574 38782 54626
rect 38834 54574 38836 54626
rect 38780 53730 38836 54574
rect 38780 53678 38782 53730
rect 38834 53678 38836 53730
rect 38780 53666 38836 53678
rect 38556 53508 38612 53518
rect 38444 52836 38500 52846
rect 38556 52836 38612 53452
rect 38780 53060 38836 53070
rect 38780 52966 38836 53004
rect 38892 52948 38948 56142
rect 39228 56084 39284 56094
rect 39228 55300 39284 56028
rect 40236 56082 40292 56702
rect 40236 56030 40238 56082
rect 40290 56030 40292 56082
rect 39788 55970 39844 55982
rect 39788 55918 39790 55970
rect 39842 55918 39844 55970
rect 39228 55234 39284 55244
rect 39452 55298 39508 55310
rect 39452 55246 39454 55298
rect 39506 55246 39508 55298
rect 39452 55188 39508 55246
rect 39228 54290 39284 54302
rect 39228 54238 39230 54290
rect 39282 54238 39284 54290
rect 38892 52882 38948 52892
rect 39116 53506 39172 53518
rect 39116 53454 39118 53506
rect 39170 53454 39172 53506
rect 38444 52834 38612 52836
rect 38444 52782 38446 52834
rect 38498 52782 38612 52834
rect 38444 52780 38612 52782
rect 38444 52770 38500 52780
rect 38332 52162 38388 52174
rect 38332 52110 38334 52162
rect 38386 52110 38388 52162
rect 38332 51492 38388 52110
rect 38444 51940 38500 51950
rect 38444 51846 38500 51884
rect 38556 51716 38612 52780
rect 39004 52722 39060 52734
rect 39004 52670 39006 52722
rect 39058 52670 39060 52722
rect 38780 52276 38836 52286
rect 39004 52276 39060 52670
rect 38780 52274 39060 52276
rect 38780 52222 38782 52274
rect 38834 52222 39060 52274
rect 38780 52220 39060 52222
rect 38780 52210 38836 52220
rect 38668 52162 38724 52174
rect 38668 52110 38670 52162
rect 38722 52110 38724 52162
rect 38668 51828 38724 52110
rect 39116 52052 39172 53454
rect 39004 51996 39172 52052
rect 38668 51762 38724 51772
rect 38780 51938 38836 51950
rect 38780 51886 38782 51938
rect 38834 51886 38836 51938
rect 38332 51426 38388 51436
rect 38444 51660 38612 51716
rect 37548 50418 37604 50428
rect 37884 50372 38164 50428
rect 38220 51154 38276 51166
rect 38220 51102 38222 51154
rect 38274 51102 38276 51154
rect 37660 49922 37716 49934
rect 37660 49870 37662 49922
rect 37714 49870 37716 49922
rect 37548 49812 37604 49822
rect 37324 49634 37380 49644
rect 37436 49810 37604 49812
rect 37436 49758 37550 49810
rect 37602 49758 37604 49810
rect 37436 49756 37604 49758
rect 37212 49476 37268 49486
rect 37212 49026 37268 49420
rect 37212 48974 37214 49026
rect 37266 48974 37268 49026
rect 37212 48962 37268 48974
rect 37100 48514 37156 48524
rect 37324 48802 37380 48814
rect 37324 48750 37326 48802
rect 37378 48750 37380 48802
rect 37100 48244 37156 48254
rect 37100 48150 37156 48188
rect 37324 48130 37380 48750
rect 37436 48804 37492 49756
rect 37548 49746 37604 49756
rect 37660 49476 37716 49870
rect 37660 49410 37716 49420
rect 37772 49924 37828 49934
rect 37436 48710 37492 48748
rect 37548 49140 37604 49150
rect 37324 48078 37326 48130
rect 37378 48078 37380 48130
rect 37324 48066 37380 48078
rect 36540 46674 36820 46676
rect 36540 46622 36542 46674
rect 36594 46622 36820 46674
rect 36540 46620 36820 46622
rect 36988 46676 37044 46686
rect 36540 46610 36596 46620
rect 36988 46582 37044 46620
rect 37548 46562 37604 49084
rect 37660 49028 37716 49038
rect 37772 49028 37828 49868
rect 37660 49026 37828 49028
rect 37660 48974 37662 49026
rect 37714 48974 37828 49026
rect 37660 48972 37828 48974
rect 37660 48962 37716 48972
rect 37772 48916 37828 48972
rect 37772 48850 37828 48860
rect 37884 48580 37940 50372
rect 38108 49924 38164 49934
rect 37996 48916 38052 48926
rect 37996 48822 38052 48860
rect 38108 48580 38164 49868
rect 38220 49810 38276 51102
rect 38332 51154 38388 51166
rect 38332 51102 38334 51154
rect 38386 51102 38388 51154
rect 38332 50596 38388 51102
rect 38332 50530 38388 50540
rect 38220 49758 38222 49810
rect 38274 49758 38276 49810
rect 38220 49746 38276 49758
rect 38332 49700 38388 49710
rect 38332 49028 38388 49644
rect 38332 48934 38388 48972
rect 37548 46510 37550 46562
rect 37602 46510 37604 46562
rect 37548 46498 37604 46510
rect 37660 48524 37940 48580
rect 37996 48524 38164 48580
rect 36316 46116 36372 46126
rect 36092 45892 36148 45902
rect 36092 45890 36260 45892
rect 36092 45838 36094 45890
rect 36146 45838 36260 45890
rect 36092 45836 36260 45838
rect 36092 45826 36148 45836
rect 36092 45668 36148 45678
rect 35980 45612 36092 45668
rect 36092 44212 36148 45612
rect 36204 45444 36260 45836
rect 36204 45378 36260 45388
rect 36204 45218 36260 45230
rect 36204 45166 36206 45218
rect 36258 45166 36260 45218
rect 36204 44546 36260 45166
rect 36204 44494 36206 44546
rect 36258 44494 36260 44546
rect 36204 44482 36260 44494
rect 36316 44322 36372 46060
rect 37660 45892 37716 48524
rect 37772 48356 37828 48366
rect 37996 48356 38052 48524
rect 37772 48354 38388 48356
rect 37772 48302 37774 48354
rect 37826 48302 38388 48354
rect 37772 48300 38388 48302
rect 37772 48290 37828 48300
rect 37212 45836 37716 45892
rect 38108 47460 38164 47470
rect 36428 45780 36484 45790
rect 36428 45686 36484 45724
rect 37100 45668 37156 45678
rect 37100 45574 37156 45612
rect 36316 44270 36318 44322
rect 36370 44270 36372 44322
rect 36316 44258 36372 44270
rect 36764 45332 36820 45342
rect 36204 44212 36260 44222
rect 36092 44210 36260 44212
rect 36092 44158 36206 44210
rect 36258 44158 36260 44210
rect 36092 44156 36260 44158
rect 36204 44146 36260 44156
rect 36764 44212 36820 45276
rect 36988 44212 37044 44222
rect 36764 44210 37044 44212
rect 36764 44158 36990 44210
rect 37042 44158 37044 44210
rect 36764 44156 37044 44158
rect 35868 43820 36260 43876
rect 34748 43250 34804 43260
rect 35084 43652 35476 43708
rect 36204 43764 36260 43820
rect 36092 43652 36148 43662
rect 34524 42868 34580 42878
rect 34524 42774 34580 42812
rect 34748 42868 34804 42878
rect 33852 42142 33854 42194
rect 33906 42142 33908 42194
rect 33852 42130 33908 42142
rect 34300 41860 34356 41870
rect 33740 41858 34356 41860
rect 33740 41806 34302 41858
rect 34354 41806 34356 41858
rect 33740 41804 34356 41806
rect 34300 41794 34356 41804
rect 34748 41860 34804 42812
rect 35084 42754 35140 43652
rect 35980 43316 36036 43326
rect 35868 43204 35924 43214
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 35084 42702 35086 42754
rect 35138 42702 35140 42754
rect 35084 42690 35140 42702
rect 34860 42644 34916 42654
rect 34860 42082 34916 42588
rect 35756 42644 35812 42654
rect 35756 42550 35812 42588
rect 35868 42420 35924 43148
rect 35980 42532 36036 43260
rect 36092 42754 36148 43596
rect 36204 43540 36260 43708
rect 36204 43446 36260 43484
rect 36092 42702 36094 42754
rect 36146 42702 36148 42754
rect 36092 42690 36148 42702
rect 36428 43428 36484 43438
rect 36764 43428 36820 44156
rect 36988 44146 37044 44156
rect 37100 44098 37156 44110
rect 37100 44046 37102 44098
rect 37154 44046 37156 44098
rect 37100 43764 37156 44046
rect 37100 43698 37156 43708
rect 36428 43426 36820 43428
rect 36428 43374 36430 43426
rect 36482 43374 36820 43426
rect 36428 43372 36820 43374
rect 36876 43428 36932 43438
rect 35980 42530 36260 42532
rect 35980 42478 35982 42530
rect 36034 42478 36260 42530
rect 35980 42476 36260 42478
rect 35980 42466 36036 42476
rect 34860 42030 34862 42082
rect 34914 42030 34916 42082
rect 34860 42018 34916 42030
rect 35756 42364 35924 42420
rect 34076 41298 34132 41310
rect 34076 41246 34078 41298
rect 34130 41246 34132 41298
rect 33628 41132 34020 41188
rect 33516 41010 33572 41020
rect 33852 40964 33908 40974
rect 33404 40628 33460 40638
rect 33852 40628 33908 40908
rect 33404 40626 33908 40628
rect 33404 40574 33406 40626
rect 33458 40574 33908 40626
rect 33404 40572 33908 40574
rect 33404 40562 33460 40572
rect 33852 40514 33908 40572
rect 33852 40462 33854 40514
rect 33906 40462 33908 40514
rect 33852 40450 33908 40462
rect 33292 40404 33348 40414
rect 33292 40310 33348 40348
rect 33404 40180 33460 40190
rect 33404 40178 33796 40180
rect 33404 40126 33406 40178
rect 33458 40126 33796 40178
rect 33404 40124 33796 40126
rect 33404 40114 33460 40124
rect 33180 39900 33460 39956
rect 33292 39396 33348 39406
rect 33180 39394 33348 39396
rect 33180 39342 33294 39394
rect 33346 39342 33348 39394
rect 33180 39340 33348 39342
rect 33180 38612 33236 39340
rect 33292 39330 33348 39340
rect 33180 38546 33236 38556
rect 33292 38946 33348 38958
rect 33292 38894 33294 38946
rect 33346 38894 33348 38946
rect 33292 38276 33348 38894
rect 33068 38220 33348 38276
rect 33068 38162 33124 38220
rect 33068 38110 33070 38162
rect 33122 38110 33124 38162
rect 33068 38098 33124 38110
rect 32956 36754 33012 36764
rect 33180 36596 33236 36606
rect 32844 36092 33124 36148
rect 32396 35924 32452 35934
rect 32956 35924 33012 35934
rect 32396 35922 33012 35924
rect 32396 35870 32398 35922
rect 32450 35870 32958 35922
rect 33010 35870 33012 35922
rect 32396 35868 33012 35870
rect 32396 35858 32452 35868
rect 32956 35858 33012 35868
rect 32508 35698 32564 35710
rect 32508 35646 32510 35698
rect 32562 35646 32564 35698
rect 32284 35308 32452 35364
rect 31948 33908 32004 35196
rect 32060 34804 32116 34814
rect 32060 34710 32116 34748
rect 32284 34690 32340 34702
rect 32284 34638 32286 34690
rect 32338 34638 32340 34690
rect 32172 34356 32228 34366
rect 32060 34300 32172 34356
rect 32060 34130 32116 34300
rect 32172 34290 32228 34300
rect 32060 34078 32062 34130
rect 32114 34078 32116 34130
rect 32060 34066 32116 34078
rect 32172 34132 32228 34142
rect 32172 34038 32228 34076
rect 31948 33842 32004 33852
rect 31948 33684 32004 33694
rect 31948 33458 32004 33628
rect 31948 33406 31950 33458
rect 32002 33406 32004 33458
rect 31948 33394 32004 33406
rect 31948 33124 32004 33134
rect 31948 33030 32004 33068
rect 32172 33122 32228 33134
rect 32172 33070 32174 33122
rect 32226 33070 32228 33122
rect 32172 32676 32228 33070
rect 32172 32610 32228 32620
rect 31836 31826 31892 31836
rect 31052 31726 31054 31778
rect 31106 31726 31108 31778
rect 30716 30996 30772 31006
rect 30492 30212 30548 30222
rect 30492 30118 30548 30156
rect 30380 29810 30436 29820
rect 30604 29988 30660 29998
rect 30156 29764 30212 29774
rect 29708 29708 30100 29764
rect 30044 29650 30100 29708
rect 30044 29598 30046 29650
rect 30098 29598 30100 29650
rect 30044 29586 30100 29598
rect 30044 28644 30100 28654
rect 29596 28642 30100 28644
rect 29596 28590 29598 28642
rect 29650 28590 30046 28642
rect 30098 28590 30100 28642
rect 29596 28588 30100 28590
rect 29596 28578 29652 28588
rect 30044 28578 30100 28588
rect 30156 28420 30212 29708
rect 30380 29538 30436 29550
rect 30380 29486 30382 29538
rect 30434 29486 30436 29538
rect 30380 28644 30436 29486
rect 30604 29426 30660 29932
rect 30604 29374 30606 29426
rect 30658 29374 30660 29426
rect 30604 29362 30660 29374
rect 30716 29652 30772 30940
rect 30828 30548 30884 30558
rect 30828 30098 30884 30492
rect 30828 30046 30830 30098
rect 30882 30046 30884 30098
rect 30828 30034 30884 30046
rect 30716 29204 30772 29596
rect 31052 29652 31108 31726
rect 31948 31778 32004 31790
rect 31948 31726 31950 31778
rect 32002 31726 32004 31778
rect 31164 31666 31220 31678
rect 31164 31614 31166 31666
rect 31218 31614 31220 31666
rect 31164 30100 31220 31614
rect 31500 31666 31556 31678
rect 31500 31614 31502 31666
rect 31554 31614 31556 31666
rect 31500 31220 31556 31614
rect 31500 30772 31556 31164
rect 31836 30884 31892 30894
rect 31836 30790 31892 30828
rect 31500 30706 31556 30716
rect 31500 30548 31556 30558
rect 31948 30548 32004 31726
rect 32284 30772 32340 34638
rect 32396 34130 32452 35308
rect 32508 35026 32564 35646
rect 32508 34974 32510 35026
rect 32562 34974 32564 35026
rect 32508 34962 32564 34974
rect 32396 34078 32398 34130
rect 32450 34078 32452 34130
rect 32396 34066 32452 34078
rect 32508 34690 32564 34702
rect 32508 34638 32510 34690
rect 32562 34638 32564 34690
rect 32396 33908 32452 33918
rect 32396 31890 32452 33852
rect 32508 32676 32564 34638
rect 32956 34356 33012 34366
rect 33068 34356 33124 36092
rect 33180 35922 33236 36540
rect 33180 35870 33182 35922
rect 33234 35870 33236 35922
rect 33180 35858 33236 35870
rect 33292 35698 33348 35710
rect 33292 35646 33294 35698
rect 33346 35646 33348 35698
rect 33292 35364 33348 35646
rect 33292 35298 33348 35308
rect 33180 35140 33236 35150
rect 33404 35140 33460 39900
rect 33740 39620 33796 40124
rect 33852 39620 33908 39630
rect 33740 39618 33908 39620
rect 33740 39566 33854 39618
rect 33906 39566 33908 39618
rect 33740 39564 33908 39566
rect 33852 39554 33908 39564
rect 33516 38834 33572 38846
rect 33516 38782 33518 38834
rect 33570 38782 33572 38834
rect 33516 38668 33572 38782
rect 33964 38724 34020 41132
rect 34076 40404 34132 41246
rect 34748 41186 34804 41804
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 35420 41188 35476 41198
rect 34748 41134 34750 41186
rect 34802 41134 34804 41186
rect 34748 41122 34804 41134
rect 35308 41186 35476 41188
rect 35308 41134 35422 41186
rect 35474 41134 35476 41186
rect 35308 41132 35476 41134
rect 34636 41076 34692 41086
rect 34636 40982 34692 41020
rect 34412 40964 34468 40974
rect 34412 40870 34468 40908
rect 34076 40310 34132 40348
rect 35308 40626 35364 41132
rect 35420 41122 35476 41132
rect 35308 40574 35310 40626
rect 35362 40574 35364 40626
rect 34412 40292 34468 40302
rect 34188 40236 34412 40292
rect 34188 39618 34244 40236
rect 34412 40198 34468 40236
rect 35308 40292 35364 40574
rect 35420 40628 35476 40638
rect 35420 40534 35476 40572
rect 35644 40514 35700 40526
rect 35644 40462 35646 40514
rect 35698 40462 35700 40514
rect 35532 40404 35588 40414
rect 35644 40404 35700 40462
rect 35532 40402 35700 40404
rect 35532 40350 35534 40402
rect 35586 40350 35700 40402
rect 35532 40348 35700 40350
rect 35532 40338 35588 40348
rect 35308 40180 35364 40236
rect 35308 40124 35588 40180
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 34188 39566 34190 39618
rect 34242 39566 34244 39618
rect 34188 39554 34244 39566
rect 35532 39618 35588 40124
rect 35532 39566 35534 39618
rect 35586 39566 35588 39618
rect 35532 39554 35588 39566
rect 34412 39394 34468 39406
rect 34412 39342 34414 39394
rect 34466 39342 34468 39394
rect 33516 38612 33908 38668
rect 33964 38658 34020 38668
rect 34076 38722 34132 38734
rect 34076 38670 34078 38722
rect 34130 38670 34132 38722
rect 34076 38668 34132 38670
rect 34412 38668 34468 39342
rect 34524 39396 34580 39406
rect 34524 39394 35140 39396
rect 34524 39342 34526 39394
rect 34578 39342 35140 39394
rect 34524 39340 35140 39342
rect 34524 39330 34580 39340
rect 34076 38612 34468 38668
rect 34748 38724 34804 38734
rect 34748 38612 35028 38668
rect 33516 37492 33572 37502
rect 33852 37492 33908 38612
rect 34300 38164 34356 38174
rect 33964 37492 34020 37502
rect 33852 37490 34020 37492
rect 33852 37438 33966 37490
rect 34018 37438 34020 37490
rect 33852 37436 34020 37438
rect 33516 37398 33572 37436
rect 33964 37426 34020 37436
rect 34300 37266 34356 38108
rect 34300 37214 34302 37266
rect 34354 37214 34356 37266
rect 34300 37202 34356 37214
rect 34412 37156 34468 38612
rect 34524 37492 34580 37502
rect 34524 37378 34580 37436
rect 34860 37380 34916 37390
rect 34524 37326 34526 37378
rect 34578 37326 34580 37378
rect 34524 37314 34580 37326
rect 34748 37378 34916 37380
rect 34748 37326 34862 37378
rect 34914 37326 34916 37378
rect 34748 37324 34916 37326
rect 34412 37100 34580 37156
rect 34188 36820 34244 36830
rect 34244 36764 34356 36820
rect 34188 36754 34244 36764
rect 33852 36596 33908 36606
rect 33852 36502 33908 36540
rect 33852 35588 33908 35598
rect 34188 35588 34244 35598
rect 33852 35586 34244 35588
rect 33852 35534 33854 35586
rect 33906 35534 34190 35586
rect 34242 35534 34244 35586
rect 33852 35532 34244 35534
rect 33852 35522 33908 35532
rect 33180 35138 33460 35140
rect 33180 35086 33182 35138
rect 33234 35086 33460 35138
rect 33180 35084 33460 35086
rect 33180 35074 33236 35084
rect 33964 35028 34020 35532
rect 34188 35522 34244 35532
rect 34300 35140 34356 36764
rect 34412 36596 34468 36606
rect 34412 36502 34468 36540
rect 34412 35140 34468 35150
rect 34300 35138 34468 35140
rect 34300 35086 34414 35138
rect 34466 35086 34468 35138
rect 34300 35084 34468 35086
rect 34412 35074 34468 35084
rect 33740 34972 34020 35028
rect 33516 34916 33572 34926
rect 33740 34916 33796 34972
rect 33516 34914 33796 34916
rect 33516 34862 33518 34914
rect 33570 34862 33796 34914
rect 33516 34860 33796 34862
rect 33964 34914 34020 34972
rect 33964 34862 33966 34914
rect 34018 34862 34020 34914
rect 33516 34850 33572 34860
rect 33292 34692 33348 34702
rect 33292 34598 33348 34636
rect 33068 34300 33236 34356
rect 32956 34262 33012 34300
rect 32620 34132 32676 34142
rect 32620 34038 32676 34076
rect 33068 34130 33124 34142
rect 33068 34078 33070 34130
rect 33122 34078 33124 34130
rect 32508 32610 32564 32620
rect 32732 33124 32788 33134
rect 32396 31838 32398 31890
rect 32450 31838 32452 31890
rect 32396 31108 32452 31838
rect 32396 31042 32452 31052
rect 32284 30716 32676 30772
rect 31500 30434 31556 30492
rect 31500 30382 31502 30434
rect 31554 30382 31556 30434
rect 31500 30370 31556 30382
rect 31724 30492 32004 30548
rect 31276 30100 31332 30110
rect 31164 30098 31332 30100
rect 31164 30046 31278 30098
rect 31330 30046 31332 30098
rect 31164 30044 31332 30046
rect 31276 29876 31332 30044
rect 31612 29988 31668 29998
rect 31724 29988 31780 30492
rect 31836 30322 31892 30334
rect 31836 30270 31838 30322
rect 31890 30270 31892 30322
rect 31836 30212 31892 30270
rect 32284 30212 32340 30222
rect 32508 30212 32564 30222
rect 31836 30210 32452 30212
rect 31836 30158 32286 30210
rect 32338 30158 32452 30210
rect 31836 30156 32452 30158
rect 32284 30146 32340 30156
rect 31668 29932 31780 29988
rect 31612 29922 31668 29932
rect 31276 29810 31332 29820
rect 31052 29586 31108 29596
rect 31164 29764 31220 29774
rect 31164 29540 31220 29708
rect 31948 29652 32004 29662
rect 32284 29652 32340 29662
rect 31948 29558 32004 29596
rect 32060 29596 32284 29652
rect 31164 29314 31220 29484
rect 31164 29262 31166 29314
rect 31218 29262 31220 29314
rect 31164 29250 31220 29262
rect 31612 29426 31668 29438
rect 31612 29374 31614 29426
rect 31666 29374 31668 29426
rect 30380 28578 30436 28588
rect 30492 29148 30772 29204
rect 29932 28364 30212 28420
rect 30380 28418 30436 28430
rect 30380 28366 30382 28418
rect 30434 28366 30436 28418
rect 29596 27860 29652 27870
rect 29484 27858 29652 27860
rect 29484 27806 29598 27858
rect 29650 27806 29652 27858
rect 29484 27804 29652 27806
rect 29596 27794 29652 27804
rect 29260 27692 29540 27748
rect 28924 26852 29204 26908
rect 29260 27186 29316 27198
rect 29260 27134 29262 27186
rect 29314 27134 29316 27186
rect 29260 26964 29316 27134
rect 29260 26898 29316 26908
rect 28924 26514 28980 26852
rect 28924 26462 28926 26514
rect 28978 26462 28980 26514
rect 28924 26450 28980 26462
rect 29260 26180 29316 26190
rect 28812 26178 29316 26180
rect 28812 26126 29262 26178
rect 29314 26126 29316 26178
rect 28812 26124 29316 26126
rect 28588 22260 28644 22270
rect 28588 22258 28756 22260
rect 28588 22206 28590 22258
rect 28642 22206 28756 22258
rect 28588 22204 28756 22206
rect 28588 22194 28644 22204
rect 28588 21698 28644 21710
rect 28588 21646 28590 21698
rect 28642 21646 28644 21698
rect 28588 21476 28644 21646
rect 28588 21410 28644 21420
rect 28700 21474 28756 22204
rect 28700 21422 28702 21474
rect 28754 21422 28756 21474
rect 28700 21410 28756 21422
rect 28812 21252 28868 26124
rect 29260 26114 29316 26124
rect 29484 25956 29540 27692
rect 29708 27076 29764 27086
rect 29708 26982 29764 27020
rect 29932 26514 29988 28364
rect 30044 27860 30100 27870
rect 30380 27860 30436 28366
rect 30044 27858 30436 27860
rect 30044 27806 30046 27858
rect 30098 27806 30436 27858
rect 30044 27804 30436 27806
rect 30044 27076 30100 27804
rect 30380 27300 30436 27310
rect 30380 27186 30436 27244
rect 30380 27134 30382 27186
rect 30434 27134 30436 27186
rect 30380 27122 30436 27134
rect 30044 27010 30100 27020
rect 29932 26462 29934 26514
rect 29986 26462 29988 26514
rect 29932 26450 29988 26462
rect 29708 26404 29764 26414
rect 29708 26310 29764 26348
rect 30156 26292 30212 26302
rect 30380 26292 30436 26302
rect 30156 26290 30436 26292
rect 30156 26238 30158 26290
rect 30210 26238 30382 26290
rect 30434 26238 30436 26290
rect 30156 26236 30436 26238
rect 30156 26226 30212 26236
rect 30380 26226 30436 26236
rect 29484 25890 29540 25900
rect 30044 26178 30100 26190
rect 30044 26126 30046 26178
rect 30098 26126 30100 26178
rect 29932 25620 29988 25630
rect 30044 25620 30100 26126
rect 29932 25618 30100 25620
rect 29932 25566 29934 25618
rect 29986 25566 30100 25618
rect 29932 25564 30100 25566
rect 29932 25554 29988 25564
rect 29260 25506 29316 25518
rect 29260 25454 29262 25506
rect 29314 25454 29316 25506
rect 29260 24948 29316 25454
rect 30492 25060 30548 29148
rect 30604 28868 30660 28878
rect 30604 27746 30660 28812
rect 31164 28756 31220 28766
rect 31164 28662 31220 28700
rect 30828 28644 30884 28654
rect 30828 28550 30884 28588
rect 31612 28644 31668 29374
rect 31612 28550 31668 28588
rect 31724 28420 31780 28430
rect 30940 27860 30996 27870
rect 30604 27694 30606 27746
rect 30658 27694 30660 27746
rect 30604 26740 30660 27694
rect 30828 27858 30996 27860
rect 30828 27806 30942 27858
rect 30994 27806 30996 27858
rect 30828 27804 30996 27806
rect 30828 27076 30884 27804
rect 30940 27794 30996 27804
rect 30828 26982 30884 27020
rect 31388 27746 31444 27758
rect 31388 27694 31390 27746
rect 31442 27694 31444 27746
rect 31388 27076 31444 27694
rect 30604 26674 30660 26684
rect 30492 24994 30548 25004
rect 30604 26402 30660 26414
rect 30604 26350 30606 26402
rect 30658 26350 30660 26402
rect 29316 24892 29540 24948
rect 29260 24882 29316 24892
rect 29260 23828 29316 23838
rect 28700 21196 28868 21252
rect 29036 23826 29316 23828
rect 29036 23774 29262 23826
rect 29314 23774 29316 23826
rect 29036 23772 29316 23774
rect 28588 20132 28644 20142
rect 28588 19236 28644 20076
rect 28588 18674 28644 19180
rect 28588 18622 28590 18674
rect 28642 18622 28644 18674
rect 28588 18610 28644 18622
rect 28420 18172 28532 18228
rect 28364 18162 28420 18172
rect 28476 18004 28532 18014
rect 28364 17556 28420 17566
rect 28364 17106 28420 17500
rect 28364 17054 28366 17106
rect 28418 17054 28420 17106
rect 28364 17042 28420 17054
rect 27916 15426 28308 15428
rect 27916 15374 27918 15426
rect 27970 15374 28308 15426
rect 27916 15372 28308 15374
rect 27916 15362 27972 15372
rect 27580 14980 27636 14990
rect 27356 14130 27412 14140
rect 27468 14924 27580 14980
rect 27244 13746 27300 13758
rect 27244 13694 27246 13746
rect 27298 13694 27300 13746
rect 27244 12962 27300 13694
rect 27244 12910 27246 12962
rect 27298 12910 27300 12962
rect 27244 12066 27300 12910
rect 27244 12014 27246 12066
rect 27298 12014 27300 12066
rect 27244 11284 27300 12014
rect 27244 11218 27300 11228
rect 27468 9940 27524 14924
rect 27580 14914 27636 14924
rect 28476 14980 28532 17948
rect 28700 17780 28756 21196
rect 28924 19794 28980 19806
rect 28924 19742 28926 19794
rect 28978 19742 28980 19794
rect 28812 19012 28868 19022
rect 28812 18674 28868 18956
rect 28812 18622 28814 18674
rect 28866 18622 28868 18674
rect 28812 18610 28868 18622
rect 28924 18450 28980 19742
rect 29036 18788 29092 23772
rect 29260 23762 29316 23772
rect 29372 23714 29428 23726
rect 29372 23662 29374 23714
rect 29426 23662 29428 23714
rect 29372 23380 29428 23662
rect 29372 23314 29428 23324
rect 29260 22484 29316 22494
rect 29148 21476 29204 21486
rect 29148 20692 29204 21420
rect 29260 20916 29316 22428
rect 29484 21812 29540 24892
rect 30268 24834 30324 24846
rect 30268 24782 30270 24834
rect 30322 24782 30324 24834
rect 30044 24724 30100 24734
rect 29596 24722 30100 24724
rect 29596 24670 30046 24722
rect 30098 24670 30100 24722
rect 29596 24668 30100 24670
rect 29596 23938 29652 24668
rect 30044 24658 30100 24668
rect 30268 24388 30324 24782
rect 30380 24836 30436 24846
rect 30380 24742 30436 24780
rect 30380 24612 30436 24622
rect 30604 24612 30660 26350
rect 30940 26404 30996 26414
rect 30940 26310 30996 26348
rect 31164 26404 31220 26414
rect 30716 26292 30772 26302
rect 30716 26198 30772 26236
rect 30828 25396 30884 25406
rect 30828 24722 30884 25340
rect 31164 25284 31220 26348
rect 31276 26290 31332 26302
rect 31276 26238 31278 26290
rect 31330 26238 31332 26290
rect 31276 25508 31332 26238
rect 31276 25442 31332 25452
rect 31164 25218 31220 25228
rect 30828 24670 30830 24722
rect 30882 24670 30884 24722
rect 30828 24658 30884 24670
rect 30380 24610 30660 24612
rect 30380 24558 30382 24610
rect 30434 24558 30660 24610
rect 30380 24556 30660 24558
rect 30380 24546 30436 24556
rect 30268 24332 30660 24388
rect 30156 24276 30212 24286
rect 30044 24220 30156 24276
rect 30044 24050 30100 24220
rect 30156 24210 30212 24220
rect 30268 24164 30324 24174
rect 30268 24052 30324 24108
rect 30044 23998 30046 24050
rect 30098 23998 30100 24050
rect 30044 23986 30100 23998
rect 30156 23996 30324 24052
rect 29596 23886 29598 23938
rect 29650 23886 29652 23938
rect 29596 23874 29652 23886
rect 30156 23826 30212 23996
rect 30492 23940 30548 23950
rect 30492 23846 30548 23884
rect 30156 23774 30158 23826
rect 30210 23774 30212 23826
rect 30156 23762 30212 23774
rect 29820 23714 29876 23726
rect 29820 23662 29822 23714
rect 29874 23662 29876 23714
rect 29820 23492 29876 23662
rect 30044 23714 30100 23726
rect 30044 23662 30046 23714
rect 30098 23662 30100 23714
rect 30044 23604 30100 23662
rect 30044 23548 30212 23604
rect 29820 23436 30100 23492
rect 29708 23380 29764 23390
rect 29764 23324 29876 23380
rect 29708 23314 29764 23324
rect 29820 23266 29876 23324
rect 30044 23378 30100 23436
rect 30044 23326 30046 23378
rect 30098 23326 30100 23378
rect 30044 23314 30100 23326
rect 29820 23214 29822 23266
rect 29874 23214 29876 23266
rect 29820 23202 29876 23214
rect 29708 23156 29764 23166
rect 29484 21586 29540 21756
rect 29484 21534 29486 21586
rect 29538 21534 29540 21586
rect 29484 21522 29540 21534
rect 29596 23154 29764 23156
rect 29596 23102 29710 23154
rect 29762 23102 29764 23154
rect 29596 23100 29764 23102
rect 29596 20916 29652 23100
rect 29708 23090 29764 23100
rect 30156 20916 30212 23548
rect 30492 22148 30548 22158
rect 30268 22092 30492 22148
rect 30268 21698 30324 22092
rect 30492 22082 30548 22092
rect 30268 21646 30270 21698
rect 30322 21646 30324 21698
rect 30268 21634 30324 21646
rect 29260 20860 29428 20916
rect 29260 20692 29316 20702
rect 29148 20690 29316 20692
rect 29148 20638 29262 20690
rect 29314 20638 29316 20690
rect 29148 20636 29316 20638
rect 29260 20580 29316 20636
rect 29260 20514 29316 20524
rect 29372 20130 29428 20860
rect 29372 20078 29374 20130
rect 29426 20078 29428 20130
rect 29372 19460 29428 20078
rect 29484 20860 29652 20916
rect 29708 20860 30212 20916
rect 29484 19794 29540 20860
rect 29708 20804 29764 20860
rect 29484 19742 29486 19794
rect 29538 19742 29540 19794
rect 29484 19730 29540 19742
rect 29596 20748 29764 20804
rect 29372 19394 29428 19404
rect 29596 19348 29652 20748
rect 29932 20692 29988 20702
rect 29932 20690 30212 20692
rect 29932 20638 29934 20690
rect 29986 20638 30212 20690
rect 29932 20636 30212 20638
rect 29932 20626 29988 20636
rect 29708 20580 29764 20590
rect 29708 20486 29764 20524
rect 29820 20578 29876 20590
rect 29820 20526 29822 20578
rect 29874 20526 29876 20578
rect 29820 20356 29876 20526
rect 30156 20468 30212 20636
rect 30156 20412 30436 20468
rect 29820 20300 30212 20356
rect 29820 20130 29876 20142
rect 29820 20078 29822 20130
rect 29874 20078 29876 20130
rect 29708 20018 29764 20030
rect 29708 19966 29710 20018
rect 29762 19966 29764 20018
rect 29708 19684 29764 19966
rect 29708 19618 29764 19628
rect 29820 19572 29876 20078
rect 30156 20132 30212 20300
rect 30268 20132 30324 20142
rect 30156 20130 30324 20132
rect 30156 20078 30270 20130
rect 30322 20078 30324 20130
rect 30156 20076 30324 20078
rect 30268 20066 30324 20076
rect 30380 20132 30436 20412
rect 30380 20066 30436 20076
rect 30044 20020 30100 20030
rect 30044 19926 30100 19964
rect 30492 20020 30548 20030
rect 30492 19926 30548 19964
rect 29820 19506 29876 19516
rect 29596 19346 29764 19348
rect 29596 19294 29598 19346
rect 29650 19294 29764 19346
rect 29596 19292 29764 19294
rect 29596 19282 29652 19292
rect 29148 19236 29204 19246
rect 29148 19142 29204 19180
rect 29260 19122 29316 19134
rect 29260 19070 29262 19122
rect 29314 19070 29316 19122
rect 29260 19012 29316 19070
rect 29260 18946 29316 18956
rect 29036 18732 29316 18788
rect 28924 18398 28926 18450
rect 28978 18398 28980 18450
rect 28924 18386 28980 18398
rect 29260 17892 29316 18732
rect 29148 17890 29316 17892
rect 29148 17838 29262 17890
rect 29314 17838 29316 17890
rect 29148 17836 29316 17838
rect 28812 17780 28868 17790
rect 28700 17724 28812 17780
rect 28812 17714 28868 17724
rect 28700 17108 28756 17118
rect 28700 17014 28756 17052
rect 28924 17108 28980 17118
rect 28924 17014 28980 17052
rect 28476 14914 28532 14924
rect 28588 16882 28644 16894
rect 28588 16830 28590 16882
rect 28642 16830 28644 16882
rect 28588 14756 28644 16830
rect 29148 15652 29204 17836
rect 29260 17826 29316 17836
rect 29708 17780 29764 19292
rect 30044 19234 30100 19246
rect 30044 19182 30046 19234
rect 30098 19182 30100 19234
rect 30044 18564 30100 19182
rect 30604 18788 30660 24332
rect 31276 23828 31332 23838
rect 31276 23734 31332 23772
rect 30940 23714 30996 23726
rect 30940 23662 30942 23714
rect 30994 23662 30996 23714
rect 30828 23380 30884 23390
rect 30940 23380 30996 23662
rect 31164 23714 31220 23726
rect 31164 23662 31166 23714
rect 31218 23662 31220 23714
rect 31052 23380 31108 23390
rect 30940 23378 31108 23380
rect 30940 23326 31054 23378
rect 31106 23326 31108 23378
rect 30940 23324 31108 23326
rect 30828 23286 30884 23324
rect 31052 23314 31108 23324
rect 30716 23154 30772 23166
rect 30716 23102 30718 23154
rect 30770 23102 30772 23154
rect 30716 22036 30772 23102
rect 30716 21970 30772 21980
rect 30828 23156 30884 23166
rect 30716 20804 30772 20814
rect 30828 20804 30884 23100
rect 30940 23044 30996 23054
rect 30940 22370 30996 22988
rect 30940 22318 30942 22370
rect 30994 22318 30996 22370
rect 30940 22306 30996 22318
rect 31164 22372 31220 23662
rect 31276 23156 31332 23166
rect 31388 23156 31444 27020
rect 31724 27412 31780 28364
rect 31612 26850 31668 26862
rect 31612 26798 31614 26850
rect 31666 26798 31668 26850
rect 31612 26404 31668 26798
rect 31724 26514 31780 27356
rect 31724 26462 31726 26514
rect 31778 26462 31780 26514
rect 31724 26450 31780 26462
rect 31612 26338 31668 26348
rect 31500 26292 31556 26302
rect 31500 26198 31556 26236
rect 31836 26292 31892 26302
rect 31836 26198 31892 26236
rect 31836 25508 31892 25518
rect 31332 23100 31444 23156
rect 31500 25060 31556 25070
rect 31724 25060 31780 25070
rect 31276 23090 31332 23100
rect 31500 22596 31556 25004
rect 31612 25004 31724 25060
rect 31612 23940 31668 25004
rect 31724 24994 31780 25004
rect 31724 24724 31780 24734
rect 31724 24050 31780 24668
rect 31836 24612 31892 25452
rect 31836 24546 31892 24556
rect 31948 25284 32004 25294
rect 31724 23998 31726 24050
rect 31778 23998 31780 24050
rect 31724 23986 31780 23998
rect 31612 23846 31668 23884
rect 31500 22540 31668 22596
rect 31500 22372 31556 22382
rect 31164 22316 31444 22372
rect 31052 22148 31108 22158
rect 31052 22054 31108 22092
rect 31164 22146 31220 22158
rect 31164 22094 31166 22146
rect 31218 22094 31220 22146
rect 31164 21812 31220 22094
rect 30716 20802 30884 20804
rect 30716 20750 30718 20802
rect 30770 20750 30884 20802
rect 30716 20748 30884 20750
rect 31052 21756 31220 21812
rect 30716 20738 30772 20748
rect 31052 20242 31108 21756
rect 31276 21364 31332 21374
rect 31276 20802 31332 21308
rect 31276 20750 31278 20802
rect 31330 20750 31332 20802
rect 31276 20738 31332 20750
rect 31052 20190 31054 20242
rect 31106 20190 31108 20242
rect 31052 20178 31108 20190
rect 30716 20020 30772 20030
rect 30716 19926 30772 19964
rect 30828 20018 30884 20030
rect 30828 19966 30830 20018
rect 30882 19966 30884 20018
rect 30828 19460 30884 19966
rect 31388 19460 31444 22316
rect 31500 22278 31556 22316
rect 31612 20356 31668 22540
rect 31724 22372 31780 22382
rect 31948 22372 32004 25228
rect 32060 23380 32116 29596
rect 32284 29558 32340 29596
rect 32172 28642 32228 28654
rect 32172 28590 32174 28642
rect 32226 28590 32228 28642
rect 32172 28420 32228 28590
rect 32396 28644 32452 30156
rect 32508 30098 32564 30156
rect 32508 30046 32510 30098
rect 32562 30046 32564 30098
rect 32508 30034 32564 30046
rect 32508 28644 32564 28654
rect 32396 28642 32564 28644
rect 32396 28590 32510 28642
rect 32562 28590 32564 28642
rect 32396 28588 32564 28590
rect 32508 28578 32564 28588
rect 32620 28420 32676 30716
rect 32172 28354 32228 28364
rect 32396 28364 32676 28420
rect 32172 28196 32228 28206
rect 32172 27524 32228 28140
rect 32172 27186 32228 27468
rect 32172 27134 32174 27186
rect 32226 27134 32228 27186
rect 32172 27122 32228 27134
rect 32396 27076 32452 28364
rect 32508 27748 32564 27758
rect 32732 27748 32788 33068
rect 33068 32788 33124 34078
rect 33068 32722 33124 32732
rect 33180 32452 33236 34300
rect 33516 34244 33572 34254
rect 33516 34130 33572 34188
rect 33516 34078 33518 34130
rect 33570 34078 33572 34130
rect 33516 34066 33572 34078
rect 33292 34020 33348 34030
rect 33292 33926 33348 33964
rect 33068 32450 33236 32452
rect 33068 32398 33182 32450
rect 33234 32398 33236 32450
rect 33068 32396 33236 32398
rect 32956 32004 33012 32014
rect 32844 31554 32900 31566
rect 32844 31502 32846 31554
rect 32898 31502 32900 31554
rect 32844 30996 32900 31502
rect 32956 31218 33012 31948
rect 32956 31166 32958 31218
rect 33010 31166 33012 31218
rect 32956 31154 33012 31166
rect 33068 30996 33124 32396
rect 33180 32386 33236 32396
rect 33180 31780 33236 31790
rect 33180 31686 33236 31724
rect 33516 31668 33572 31678
rect 33516 31574 33572 31612
rect 32844 30994 33124 30996
rect 32844 30942 33070 30994
rect 33122 30942 33124 30994
rect 32844 30940 33124 30942
rect 32956 30324 33012 30940
rect 33068 30930 33124 30940
rect 33404 31554 33460 31566
rect 33404 31502 33406 31554
rect 33458 31502 33460 31554
rect 32956 30268 33348 30324
rect 33292 30210 33348 30268
rect 33292 30158 33294 30210
rect 33346 30158 33348 30210
rect 33292 30100 33348 30158
rect 33180 30044 33348 30100
rect 32844 29428 32900 29438
rect 32844 28418 32900 29372
rect 33180 28868 33236 30044
rect 33404 29652 33460 31502
rect 33628 31444 33684 34860
rect 33964 34850 34020 34862
rect 33852 34804 33908 34814
rect 33740 34244 33796 34254
rect 33740 34150 33796 34188
rect 33852 34020 33908 34748
rect 33404 29586 33460 29596
rect 33516 31388 33684 31444
rect 33740 33964 33908 34020
rect 33964 34132 34020 34142
rect 34524 34132 34580 37100
rect 34636 35588 34692 35598
rect 34636 35138 34692 35532
rect 34748 35476 34804 37324
rect 34860 37314 34916 37324
rect 34860 37044 34916 37054
rect 34860 36258 34916 36988
rect 34860 36206 34862 36258
rect 34914 36206 34916 36258
rect 34860 35698 34916 36206
rect 34860 35646 34862 35698
rect 34914 35646 34916 35698
rect 34860 35634 34916 35646
rect 34860 35476 34916 35486
rect 34748 35420 34860 35476
rect 34860 35410 34916 35420
rect 34636 35086 34638 35138
rect 34690 35086 34692 35138
rect 34636 35074 34692 35086
rect 34972 34916 35028 38612
rect 34860 34860 35028 34916
rect 35084 34914 35140 39340
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 35308 38164 35364 38174
rect 35308 38070 35364 38108
rect 35644 38164 35700 38174
rect 35644 37490 35700 38108
rect 35644 37438 35646 37490
rect 35698 37438 35700 37490
rect 35644 37426 35700 37438
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35756 36596 35812 42364
rect 36204 42308 36260 42476
rect 36204 42242 36260 42252
rect 36092 42196 36148 42206
rect 35868 42194 36148 42196
rect 35868 42142 36094 42194
rect 36146 42142 36148 42194
rect 35868 42140 36148 42142
rect 35868 41298 35924 42140
rect 36092 42130 36148 42140
rect 36204 42084 36260 42094
rect 36428 42084 36484 43372
rect 36876 43334 36932 43372
rect 37212 43204 37268 45836
rect 37436 45668 37492 45678
rect 37436 45574 37492 45612
rect 37324 45444 37380 45454
rect 37324 44322 37380 45388
rect 37436 45108 37492 45118
rect 38108 45108 38164 47404
rect 38332 47458 38388 48300
rect 38332 47406 38334 47458
rect 38386 47406 38388 47458
rect 38332 47394 38388 47406
rect 38332 46564 38388 46574
rect 38332 45668 38388 46508
rect 38332 45602 38388 45612
rect 38220 45332 38276 45342
rect 38220 45218 38276 45276
rect 38220 45166 38222 45218
rect 38274 45166 38276 45218
rect 38220 45154 38276 45166
rect 37436 45106 38164 45108
rect 37436 45054 37438 45106
rect 37490 45054 38164 45106
rect 37436 45052 38164 45054
rect 37436 45042 37492 45052
rect 38444 44436 38500 51660
rect 38780 51604 38836 51886
rect 38892 51604 38948 51614
rect 38780 51548 38892 51604
rect 38892 51538 38948 51548
rect 38780 51378 38836 51390
rect 38780 51326 38782 51378
rect 38834 51326 38836 51378
rect 38556 51268 38612 51278
rect 38556 51174 38612 51212
rect 38780 51156 38836 51326
rect 38780 51090 38836 51100
rect 38668 50818 38724 50830
rect 38668 50766 38670 50818
rect 38722 50766 38724 50818
rect 38556 49140 38612 49150
rect 38556 47460 38612 49084
rect 38668 48132 38724 50766
rect 38780 50596 38836 50606
rect 39004 50596 39060 51996
rect 39116 51604 39172 51614
rect 39116 51510 39172 51548
rect 38780 50594 39060 50596
rect 38780 50542 38782 50594
rect 38834 50542 39060 50594
rect 38780 50540 39060 50542
rect 38780 50530 38836 50540
rect 39228 50036 39284 54238
rect 39340 53620 39396 53630
rect 39340 53170 39396 53564
rect 39340 53118 39342 53170
rect 39394 53118 39396 53170
rect 39340 53106 39396 53118
rect 39116 49980 39284 50036
rect 39340 52948 39396 52958
rect 39452 52948 39508 55132
rect 39788 54180 39844 55918
rect 40236 55524 40292 56030
rect 40236 55458 40292 55468
rect 40684 56194 40740 56206
rect 40684 56142 40686 56194
rect 40738 56142 40740 56194
rect 39900 55300 39956 55310
rect 40124 55300 40180 55310
rect 39900 55298 40068 55300
rect 39900 55246 39902 55298
rect 39954 55246 40068 55298
rect 39900 55244 40068 55246
rect 39900 55234 39956 55244
rect 39788 54114 39844 54124
rect 39900 54626 39956 54638
rect 39900 54574 39902 54626
rect 39954 54574 39956 54626
rect 39900 53956 39956 54574
rect 39788 53900 39956 53956
rect 39564 53620 39620 53630
rect 39564 53526 39620 53564
rect 39452 52892 39620 52948
rect 38892 49924 38948 49934
rect 38892 49830 38948 49868
rect 39116 49810 39172 49980
rect 39116 49758 39118 49810
rect 39170 49758 39172 49810
rect 39116 49140 39172 49758
rect 39228 49812 39284 49822
rect 39228 49698 39284 49756
rect 39228 49646 39230 49698
rect 39282 49646 39284 49698
rect 39228 49634 39284 49646
rect 39116 49074 39172 49084
rect 39116 48916 39172 48926
rect 38780 48914 39284 48916
rect 38780 48862 39118 48914
rect 39170 48862 39284 48914
rect 38780 48860 39284 48862
rect 38780 48354 38836 48860
rect 39116 48850 39172 48860
rect 38780 48302 38782 48354
rect 38834 48302 38836 48354
rect 38780 48290 38836 48302
rect 38892 48244 38948 48254
rect 38892 48132 38948 48188
rect 38668 48076 38948 48132
rect 38556 47394 38612 47404
rect 39228 47458 39284 48860
rect 39228 47406 39230 47458
rect 39282 47406 39284 47458
rect 39228 47394 39284 47406
rect 39004 47346 39060 47358
rect 39004 47294 39006 47346
rect 39058 47294 39060 47346
rect 39004 46788 39060 47294
rect 39004 46722 39060 46732
rect 38556 45892 38612 45902
rect 38556 45798 38612 45836
rect 38780 45890 38836 45902
rect 38780 45838 38782 45890
rect 38834 45838 38836 45890
rect 38780 45780 38836 45838
rect 38780 45714 38836 45724
rect 38892 45892 38948 45902
rect 37324 44270 37326 44322
rect 37378 44270 37380 44322
rect 37324 44258 37380 44270
rect 38220 44380 38500 44436
rect 38556 45668 38612 45678
rect 37324 43652 37380 43662
rect 37324 43558 37380 43596
rect 37212 43138 37268 43148
rect 37884 43428 37940 43438
rect 37100 42756 37156 42766
rect 37100 42754 37828 42756
rect 37100 42702 37102 42754
rect 37154 42702 37828 42754
rect 37100 42700 37828 42702
rect 37100 42690 37156 42700
rect 36988 42644 37044 42654
rect 36988 42550 37044 42588
rect 37772 42642 37828 42700
rect 37772 42590 37774 42642
rect 37826 42590 37828 42642
rect 36204 42082 36484 42084
rect 36204 42030 36206 42082
rect 36258 42030 36484 42082
rect 36204 42028 36484 42030
rect 36540 42532 36596 42542
rect 36204 42018 36260 42028
rect 35868 41246 35870 41298
rect 35922 41246 35924 41298
rect 35868 40514 35924 41246
rect 36316 41300 36372 41310
rect 36316 41206 36372 41244
rect 36540 41186 36596 42476
rect 37548 42532 37604 42542
rect 37548 42438 37604 42476
rect 37548 42308 37604 42318
rect 36988 42196 37044 42206
rect 36988 42102 37044 42140
rect 36540 41134 36542 41186
rect 36594 41134 36596 41186
rect 36540 41122 36596 41134
rect 36764 41970 36820 41982
rect 36764 41918 36766 41970
rect 36818 41918 36820 41970
rect 36764 40628 36820 41918
rect 36764 40562 36820 40572
rect 37100 41076 37156 41086
rect 35868 40462 35870 40514
rect 35922 40462 35924 40514
rect 35868 39730 35924 40462
rect 35868 39678 35870 39730
rect 35922 39678 35924 39730
rect 35868 39666 35924 39678
rect 36316 40290 36372 40302
rect 36316 40238 36318 40290
rect 36370 40238 36372 40290
rect 35980 38722 36036 38734
rect 35980 38670 35982 38722
rect 36034 38670 36036 38722
rect 35868 38612 35924 38622
rect 35868 37826 35924 38556
rect 35868 37774 35870 37826
rect 35922 37774 35924 37826
rect 35868 37044 35924 37774
rect 35980 37828 36036 38670
rect 36316 38668 36372 40238
rect 36428 39508 36484 39518
rect 36428 39506 36820 39508
rect 36428 39454 36430 39506
rect 36482 39454 36820 39506
rect 36428 39452 36820 39454
rect 36428 39442 36484 39452
rect 36764 38948 36820 39452
rect 37100 39506 37156 41020
rect 37324 41074 37380 41086
rect 37324 41022 37326 41074
rect 37378 41022 37380 41074
rect 37212 40404 37268 40414
rect 37324 40404 37380 41022
rect 37212 40402 37380 40404
rect 37212 40350 37214 40402
rect 37266 40350 37380 40402
rect 37212 40348 37380 40350
rect 37212 40338 37268 40348
rect 37100 39454 37102 39506
rect 37154 39454 37156 39506
rect 36876 39396 36932 39406
rect 36876 39394 37044 39396
rect 36876 39342 36878 39394
rect 36930 39342 37044 39394
rect 36876 39340 37044 39342
rect 36876 39330 36932 39340
rect 36988 38948 37044 39340
rect 37100 39172 37156 39454
rect 37212 39508 37268 39518
rect 37212 39414 37268 39452
rect 37324 39172 37380 40348
rect 37548 39396 37604 42252
rect 37772 42082 37828 42590
rect 37772 42030 37774 42082
rect 37826 42030 37828 42082
rect 37772 42018 37828 42030
rect 37884 42754 37940 43372
rect 37884 42702 37886 42754
rect 37938 42702 37940 42754
rect 37884 41970 37940 42702
rect 37884 41918 37886 41970
rect 37938 41918 37940 41970
rect 37884 41906 37940 41918
rect 38108 41972 38164 41982
rect 38108 41186 38164 41916
rect 38108 41134 38110 41186
rect 38162 41134 38164 41186
rect 38108 41122 38164 41134
rect 37660 40404 37716 40414
rect 37660 39842 37716 40348
rect 38220 39956 38276 44380
rect 38444 44210 38500 44222
rect 38444 44158 38446 44210
rect 38498 44158 38500 44210
rect 38444 43876 38500 44158
rect 38444 43810 38500 43820
rect 38332 42644 38388 42654
rect 38556 42644 38612 45612
rect 38892 45330 38948 45836
rect 38892 45278 38894 45330
rect 38946 45278 38948 45330
rect 38892 45266 38948 45278
rect 39116 45780 39172 45790
rect 39116 45218 39172 45724
rect 39116 45166 39118 45218
rect 39170 45166 39172 45218
rect 39116 45154 39172 45166
rect 38780 44882 38836 44894
rect 38780 44830 38782 44882
rect 38834 44830 38836 44882
rect 38668 44436 38724 44446
rect 38780 44436 38836 44830
rect 38724 44380 38836 44436
rect 38668 44322 38724 44380
rect 38668 44270 38670 44322
rect 38722 44270 38724 44322
rect 38668 44258 38724 44270
rect 38332 42642 38612 42644
rect 38332 42590 38334 42642
rect 38386 42590 38612 42642
rect 38332 42588 38612 42590
rect 38780 43988 38836 43998
rect 38332 41748 38388 42588
rect 38556 41972 38612 41982
rect 38556 41878 38612 41916
rect 38332 41692 38612 41748
rect 38332 41076 38388 41086
rect 38332 40404 38388 41020
rect 38556 40628 38612 41692
rect 38556 40562 38612 40572
rect 38332 40310 38388 40348
rect 38556 40292 38612 40302
rect 38556 40198 38612 40236
rect 38220 39900 38388 39956
rect 37660 39790 37662 39842
rect 37714 39790 37716 39842
rect 37660 39778 37716 39790
rect 38220 39732 38276 39742
rect 37772 39676 38220 39732
rect 37772 39618 37828 39676
rect 38220 39638 38276 39676
rect 37772 39566 37774 39618
rect 37826 39566 37828 39618
rect 37772 39554 37828 39566
rect 37660 39396 37716 39406
rect 37548 39394 37940 39396
rect 37548 39342 37662 39394
rect 37714 39342 37940 39394
rect 37548 39340 37940 39342
rect 37660 39330 37716 39340
rect 37100 39116 37268 39172
rect 37324 39116 37828 39172
rect 37212 39060 37268 39116
rect 37212 39004 37604 39060
rect 37100 38948 37156 38958
rect 36764 38892 36932 38948
rect 36988 38946 37156 38948
rect 36988 38894 37102 38946
rect 37154 38894 37156 38946
rect 36988 38892 37156 38894
rect 36540 38836 36596 38846
rect 36540 38722 36596 38780
rect 36540 38670 36542 38722
rect 36594 38670 36596 38722
rect 36540 38668 36596 38670
rect 36316 38612 36596 38668
rect 36876 38834 36932 38892
rect 36876 38782 36878 38834
rect 36930 38782 36932 38834
rect 36876 38668 36932 38782
rect 36876 38612 37044 38668
rect 36092 38052 36148 38062
rect 36092 37958 36148 37996
rect 36428 38050 36484 38612
rect 36428 37998 36430 38050
rect 36482 37998 36484 38050
rect 36428 37986 36484 37998
rect 36988 38050 37044 38612
rect 36988 37998 36990 38050
rect 37042 37998 37044 38050
rect 36988 37986 37044 37998
rect 37100 38052 37156 38892
rect 37212 38052 37268 38062
rect 37100 38050 37268 38052
rect 37100 37998 37214 38050
rect 37266 37998 37268 38050
rect 37100 37996 37268 37998
rect 37212 37986 37268 37996
rect 37436 38052 37492 38062
rect 37436 37958 37492 37996
rect 36316 37828 36372 37838
rect 37100 37828 37156 37838
rect 35980 37826 36372 37828
rect 35980 37774 36318 37826
rect 36370 37774 36372 37826
rect 35980 37772 36372 37774
rect 35868 36978 35924 36988
rect 35756 36530 35812 36540
rect 36316 36260 36372 37772
rect 36316 35700 36372 36204
rect 36316 35634 36372 35644
rect 36988 37826 37156 37828
rect 36988 37774 37102 37826
rect 37154 37774 37156 37826
rect 36988 37772 37156 37774
rect 35532 35588 35588 35598
rect 35532 35586 36036 35588
rect 35532 35534 35534 35586
rect 35586 35534 36036 35586
rect 35532 35532 36036 35534
rect 35532 35522 35588 35532
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35980 35138 36036 35532
rect 35980 35086 35982 35138
rect 36034 35086 36036 35138
rect 35980 35074 36036 35086
rect 36428 35476 36484 35486
rect 35084 34862 35086 34914
rect 35138 34862 35140 34914
rect 33964 34130 34580 34132
rect 33964 34078 33966 34130
rect 34018 34078 34580 34130
rect 33964 34076 34580 34078
rect 34748 34690 34804 34702
rect 34748 34638 34750 34690
rect 34802 34638 34804 34690
rect 33404 29426 33460 29438
rect 33404 29374 33406 29426
rect 33458 29374 33460 29426
rect 33180 28802 33236 28812
rect 33292 28980 33348 28990
rect 32844 28366 32846 28418
rect 32898 28366 32900 28418
rect 32844 28196 32900 28366
rect 33292 28644 33348 28924
rect 32844 28130 32900 28140
rect 33180 28196 33236 28206
rect 32508 27746 32788 27748
rect 32508 27694 32510 27746
rect 32562 27694 32788 27746
rect 32508 27692 32788 27694
rect 32508 27682 32564 27692
rect 32732 27300 32788 27692
rect 32732 27234 32788 27244
rect 33068 27524 33124 27534
rect 32508 27186 32564 27198
rect 32508 27134 32510 27186
rect 32562 27134 32564 27186
rect 32508 27076 32564 27134
rect 32396 27020 32564 27076
rect 32620 27188 32676 27198
rect 32620 27074 32676 27132
rect 32620 27022 32622 27074
rect 32674 27022 32676 27074
rect 32620 27010 32676 27022
rect 32844 27188 32900 27198
rect 32844 27074 32900 27132
rect 32844 27022 32846 27074
rect 32898 27022 32900 27074
rect 32844 27010 32900 27022
rect 32172 26964 32228 26974
rect 32228 26908 32340 26964
rect 32172 26898 32228 26908
rect 32172 26404 32228 26414
rect 32172 25508 32228 26348
rect 32172 25442 32228 25452
rect 32172 25284 32228 25294
rect 32172 25190 32228 25228
rect 32172 24948 32228 24958
rect 32284 24948 32340 26908
rect 33068 26962 33124 27468
rect 33068 26910 33070 26962
rect 33122 26910 33124 26962
rect 33068 26898 33124 26910
rect 33068 26628 33124 26638
rect 32508 26290 32564 26302
rect 32508 26238 32510 26290
rect 32562 26238 32564 26290
rect 32508 25620 32564 26238
rect 33068 26180 33124 26572
rect 33180 26404 33236 28140
rect 33292 28082 33348 28588
rect 33292 28030 33294 28082
rect 33346 28030 33348 28082
rect 33292 28018 33348 28030
rect 33404 27300 33460 29374
rect 33516 27524 33572 31388
rect 33740 29316 33796 33964
rect 33964 33124 34020 34076
rect 34300 33796 34356 33806
rect 34300 33236 34356 33740
rect 34412 33460 34468 33470
rect 34748 33460 34804 34638
rect 34860 34020 34916 34860
rect 35084 34850 35140 34862
rect 35196 34804 35252 34814
rect 35196 34710 35252 34748
rect 35868 34802 35924 34814
rect 35868 34750 35870 34802
rect 35922 34750 35924 34802
rect 34972 34692 35028 34702
rect 34972 34242 35028 34636
rect 35420 34692 35476 34702
rect 35420 34690 35812 34692
rect 35420 34638 35422 34690
rect 35474 34638 35812 34690
rect 35420 34636 35812 34638
rect 35420 34626 35476 34636
rect 35420 34356 35476 34366
rect 35420 34262 35476 34300
rect 34972 34190 34974 34242
rect 35026 34190 35028 34242
rect 34972 34178 35028 34190
rect 35196 34130 35252 34142
rect 35196 34078 35198 34130
rect 35250 34078 35252 34130
rect 35196 34020 35252 34078
rect 35644 34130 35700 34142
rect 35644 34078 35646 34130
rect 35698 34078 35700 34130
rect 34860 33964 35252 34020
rect 35308 34018 35364 34030
rect 35308 33966 35310 34018
rect 35362 33966 35364 34018
rect 35308 33908 35364 33966
rect 35308 33852 35588 33908
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 34748 33404 35140 33460
rect 34412 33366 34468 33404
rect 34524 33346 34580 33358
rect 34524 33294 34526 33346
rect 34578 33294 34580 33346
rect 34300 33180 34468 33236
rect 33964 33058 34020 33068
rect 34188 31892 34244 31902
rect 33852 31780 33908 31790
rect 34076 31780 34132 31790
rect 33852 31686 33908 31724
rect 33964 31724 34076 31780
rect 33964 31444 34020 31724
rect 34076 31714 34132 31724
rect 34188 31666 34244 31836
rect 34188 31614 34190 31666
rect 34242 31614 34244 31666
rect 34188 31602 34244 31614
rect 34300 31666 34356 31678
rect 34300 31614 34302 31666
rect 34354 31614 34356 31666
rect 34076 31556 34132 31566
rect 34076 31462 34132 31500
rect 33852 31388 34020 31444
rect 33852 30996 33908 31388
rect 34300 31332 34356 31614
rect 34412 31668 34468 33180
rect 34524 31892 34580 33294
rect 34860 33234 34916 33246
rect 34860 33182 34862 33234
rect 34914 33182 34916 33234
rect 34860 32900 34916 33182
rect 34972 33124 35028 33134
rect 34972 33030 35028 33068
rect 34524 31826 34580 31836
rect 34636 32844 34916 32900
rect 34636 31890 34692 32844
rect 34636 31838 34638 31890
rect 34690 31838 34692 31890
rect 34636 31826 34692 31838
rect 34748 32562 34804 32574
rect 34748 32510 34750 32562
rect 34802 32510 34804 32562
rect 34412 31612 34692 31668
rect 33852 30930 33908 30940
rect 33964 31276 34300 31332
rect 33740 29250 33796 29260
rect 33852 30772 33908 30782
rect 33852 28644 33908 30716
rect 33964 30436 34020 31276
rect 34300 31238 34356 31276
rect 34188 31108 34244 31118
rect 34244 31052 34468 31108
rect 34188 31014 34244 31052
rect 34076 30996 34132 31006
rect 34076 30902 34132 30940
rect 33964 30370 34020 30380
rect 34412 30098 34468 31052
rect 34412 30046 34414 30098
rect 34466 30046 34468 30098
rect 34412 30034 34468 30046
rect 34524 30210 34580 30222
rect 34524 30158 34526 30210
rect 34578 30158 34580 30210
rect 34300 29988 34356 29998
rect 34300 29894 34356 29932
rect 33628 28588 33908 28644
rect 33628 28530 33684 28588
rect 33628 28478 33630 28530
rect 33682 28478 33684 28530
rect 33628 28466 33684 28478
rect 33516 27458 33572 27468
rect 33628 28084 33684 28094
rect 33852 28084 33908 28588
rect 33964 29540 34020 29550
rect 33964 28418 34020 29484
rect 34524 29204 34580 30158
rect 34636 29650 34692 31612
rect 34748 30884 34804 32510
rect 34748 30324 34804 30828
rect 34860 32452 34916 32462
rect 34860 30436 34916 32396
rect 35084 32228 35140 33404
rect 35532 33346 35588 33852
rect 35644 33572 35700 34078
rect 35644 33506 35700 33516
rect 35532 33294 35534 33346
rect 35586 33294 35588 33346
rect 35532 33282 35588 33294
rect 35756 33348 35812 34636
rect 35868 33460 35924 34750
rect 35980 34692 36036 34702
rect 35980 34598 36036 34636
rect 35868 33404 36036 33460
rect 35756 33282 35812 33292
rect 35868 33236 35924 33274
rect 35868 33170 35924 33180
rect 35196 33122 35252 33134
rect 35196 33070 35198 33122
rect 35250 33070 35252 33122
rect 35196 32452 35252 33070
rect 35756 33124 35812 33134
rect 35756 33030 35812 33068
rect 35196 32386 35252 32396
rect 35868 33012 35924 33022
rect 34972 32172 35140 32228
rect 35196 32172 35460 32182
rect 34972 32002 35028 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 34972 31950 34974 32002
rect 35026 31950 35028 32002
rect 34972 31938 35028 31950
rect 35308 32004 35364 32014
rect 35084 31892 35140 31902
rect 35308 31892 35364 31948
rect 35084 31890 35364 31892
rect 35084 31838 35086 31890
rect 35138 31838 35364 31890
rect 35084 31836 35364 31838
rect 35532 31892 35588 31902
rect 35084 31826 35140 31836
rect 35532 31780 35588 31836
rect 35308 31724 35588 31780
rect 35308 31666 35364 31724
rect 35644 31668 35700 31678
rect 35308 31614 35310 31666
rect 35362 31614 35364 31666
rect 35196 31108 35252 31118
rect 35196 31014 35252 31052
rect 35084 30994 35140 31006
rect 35084 30942 35086 30994
rect 35138 30942 35140 30994
rect 35084 30436 35140 30942
rect 35308 30772 35364 31614
rect 35532 31666 35700 31668
rect 35532 31614 35646 31666
rect 35698 31614 35700 31666
rect 35532 31612 35700 31614
rect 35532 31108 35588 31612
rect 35644 31602 35700 31612
rect 35868 31666 35924 32956
rect 35980 31890 36036 33404
rect 36092 33236 36148 33246
rect 36092 33234 36372 33236
rect 36092 33182 36094 33234
rect 36146 33182 36372 33234
rect 36092 33180 36372 33182
rect 36092 33170 36148 33180
rect 35980 31838 35982 31890
rect 36034 31838 36036 31890
rect 35980 31826 36036 31838
rect 35868 31614 35870 31666
rect 35922 31614 35924 31666
rect 35532 31042 35588 31052
rect 35644 31108 35700 31118
rect 35868 31108 35924 31614
rect 35980 31332 36036 31342
rect 35980 31218 36036 31276
rect 35980 31166 35982 31218
rect 36034 31166 36036 31218
rect 35980 31154 36036 31166
rect 35644 31106 35924 31108
rect 35644 31054 35646 31106
rect 35698 31054 35924 31106
rect 35644 31052 35924 31054
rect 36204 31108 36260 31118
rect 35308 30706 35364 30716
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 34860 30380 35028 30436
rect 35084 30380 35252 30436
rect 34972 30324 35028 30380
rect 34748 30268 34916 30324
rect 34972 30268 35140 30324
rect 34636 29598 34638 29650
rect 34690 29598 34692 29650
rect 34636 29586 34692 29598
rect 34748 29538 34804 29550
rect 34748 29486 34750 29538
rect 34802 29486 34804 29538
rect 34524 29138 34580 29148
rect 34636 29426 34692 29438
rect 34636 29374 34638 29426
rect 34690 29374 34692 29426
rect 34524 28642 34580 28654
rect 34524 28590 34526 28642
rect 34578 28590 34580 28642
rect 34524 28532 34580 28590
rect 34524 28466 34580 28476
rect 33964 28366 33966 28418
rect 34018 28366 34020 28418
rect 33964 28354 34020 28366
rect 33852 28028 34356 28084
rect 33404 27234 33460 27244
rect 33292 26962 33348 26974
rect 33292 26910 33294 26962
rect 33346 26910 33348 26962
rect 33292 26908 33348 26910
rect 33628 26908 33684 28028
rect 33964 27858 34020 27870
rect 33964 27806 33966 27858
rect 34018 27806 34020 27858
rect 33964 27076 34020 27806
rect 33964 26908 34020 27020
rect 33292 26852 33460 26908
rect 33628 26852 33796 26908
rect 33180 26348 33348 26404
rect 33180 26180 33236 26190
rect 33068 26178 33236 26180
rect 33068 26126 33182 26178
rect 33234 26126 33236 26178
rect 33068 26124 33236 26126
rect 32508 25554 32564 25564
rect 33068 25956 33124 25966
rect 33068 25618 33124 25900
rect 33068 25566 33070 25618
rect 33122 25566 33124 25618
rect 33068 25554 33124 25566
rect 32620 25506 32676 25518
rect 32620 25454 32622 25506
rect 32674 25454 32676 25506
rect 32620 25396 32676 25454
rect 32620 25330 32676 25340
rect 32844 25396 32900 25406
rect 32172 24946 32340 24948
rect 32172 24894 32174 24946
rect 32226 24894 32340 24946
rect 32172 24892 32340 24894
rect 32172 24882 32228 24892
rect 32284 24836 32340 24892
rect 32508 24948 32564 24958
rect 32508 24854 32564 24892
rect 32284 24770 32340 24780
rect 32060 23314 32116 23324
rect 32172 24612 32228 24622
rect 31724 22278 31780 22316
rect 31836 22316 32004 22372
rect 32060 22372 32116 22382
rect 32172 22372 32228 24556
rect 32844 23548 32900 25340
rect 33068 25394 33124 25406
rect 33068 25342 33070 25394
rect 33122 25342 33124 25394
rect 32956 24836 33012 24846
rect 32956 24722 33012 24780
rect 32956 24670 32958 24722
rect 33010 24670 33012 24722
rect 32956 24658 33012 24670
rect 33068 24612 33124 25342
rect 33180 25396 33236 26124
rect 33292 25620 33348 26348
rect 33404 26292 33460 26852
rect 33740 26516 33796 26852
rect 33852 26852 33908 26862
rect 33964 26852 34244 26908
rect 33852 26758 33908 26796
rect 33740 26460 33908 26516
rect 33516 26404 33572 26414
rect 33516 26310 33572 26348
rect 33740 26292 33796 26302
rect 33404 26180 33460 26236
rect 33628 26290 33796 26292
rect 33628 26238 33742 26290
rect 33794 26238 33796 26290
rect 33628 26236 33796 26238
rect 33404 26124 33572 26180
rect 33292 25554 33348 25564
rect 33404 25508 33460 25518
rect 33404 25414 33460 25452
rect 33180 25302 33236 25340
rect 33516 25060 33572 26124
rect 33404 25004 33572 25060
rect 33292 24722 33348 24734
rect 33292 24670 33294 24722
rect 33346 24670 33348 24722
rect 33180 24612 33236 24622
rect 33068 24610 33236 24612
rect 33068 24558 33182 24610
rect 33234 24558 33236 24610
rect 33068 24556 33236 24558
rect 33180 24546 33236 24556
rect 33292 23716 33348 24670
rect 33292 23622 33348 23660
rect 32060 22370 32228 22372
rect 32060 22318 32062 22370
rect 32114 22318 32228 22370
rect 32060 22316 32228 22318
rect 31836 21364 31892 22316
rect 32060 22306 32116 22316
rect 31948 22146 32004 22158
rect 31948 22094 31950 22146
rect 32002 22094 32004 22146
rect 31948 21476 32004 22094
rect 32172 21700 32228 22316
rect 32732 23492 32900 23548
rect 33180 23604 33236 23614
rect 32172 21634 32228 21644
rect 32620 21700 32676 21710
rect 32396 21476 32452 21486
rect 31948 21474 32452 21476
rect 31948 21422 32398 21474
rect 32450 21422 32452 21474
rect 31948 21420 32452 21422
rect 31836 21308 32004 21364
rect 31724 20692 31780 20702
rect 31724 20598 31780 20636
rect 31612 20300 31892 20356
rect 30828 19394 30884 19404
rect 30940 19404 31444 19460
rect 31500 20130 31556 20142
rect 31500 20078 31502 20130
rect 31554 20078 31556 20130
rect 31500 19572 31556 20078
rect 31612 20132 31668 20142
rect 31612 20038 31668 20076
rect 30044 18498 30100 18508
rect 30268 18732 30660 18788
rect 30268 18116 30324 18732
rect 30492 18564 30548 18574
rect 29484 17778 29764 17780
rect 29484 17726 29710 17778
rect 29762 17726 29764 17778
rect 29484 17724 29764 17726
rect 29260 17666 29316 17678
rect 29260 17614 29262 17666
rect 29314 17614 29316 17666
rect 29260 16882 29316 17614
rect 29260 16830 29262 16882
rect 29314 16830 29316 16882
rect 29260 16324 29316 16830
rect 29484 16882 29540 17724
rect 29708 17714 29764 17724
rect 29932 18060 30324 18116
rect 30380 18562 30548 18564
rect 30380 18510 30494 18562
rect 30546 18510 30548 18562
rect 30380 18508 30548 18510
rect 29820 17666 29876 17678
rect 29820 17614 29822 17666
rect 29874 17614 29876 17666
rect 29820 16884 29876 17614
rect 29484 16830 29486 16882
rect 29538 16830 29540 16882
rect 29484 16818 29540 16830
rect 29708 16828 29876 16884
rect 29708 16660 29764 16828
rect 29708 16566 29764 16604
rect 29820 16660 29876 16670
rect 29932 16660 29988 18060
rect 30380 17556 30436 18508
rect 30492 18498 30548 18508
rect 30604 18452 30660 18462
rect 30828 18452 30884 18462
rect 30604 18358 30660 18396
rect 30716 18450 30884 18452
rect 30716 18398 30830 18450
rect 30882 18398 30884 18450
rect 30716 18396 30884 18398
rect 30492 18228 30548 18238
rect 30716 18228 30772 18396
rect 30828 18386 30884 18396
rect 30940 18228 30996 19404
rect 31500 19348 31556 19516
rect 31276 19292 31556 19348
rect 31724 19794 31780 19806
rect 31724 19742 31726 19794
rect 31778 19742 31780 19794
rect 31724 19684 31780 19742
rect 31276 18562 31332 19292
rect 31612 19236 31668 19246
rect 31500 19124 31556 19134
rect 31388 19068 31500 19124
rect 31388 18674 31444 19068
rect 31500 19030 31556 19068
rect 31388 18622 31390 18674
rect 31442 18622 31444 18674
rect 31388 18610 31444 18622
rect 31500 18676 31556 18686
rect 31276 18510 31278 18562
rect 31330 18510 31332 18562
rect 31052 18340 31108 18350
rect 31108 18284 31220 18340
rect 31052 18274 31108 18284
rect 30492 18226 30772 18228
rect 30492 18174 30494 18226
rect 30546 18174 30772 18226
rect 30492 18172 30772 18174
rect 30828 18172 30996 18228
rect 30492 18162 30548 18172
rect 30380 17490 30436 17500
rect 30604 17780 30660 17790
rect 29820 16658 29988 16660
rect 29820 16606 29822 16658
rect 29874 16606 29988 16658
rect 29820 16604 29988 16606
rect 30156 16772 30212 16782
rect 29820 16594 29876 16604
rect 29260 16258 29316 16268
rect 29820 16098 29876 16110
rect 30044 16100 30100 16110
rect 29820 16046 29822 16098
rect 29874 16046 29876 16098
rect 29820 15652 29876 16046
rect 29148 15586 29204 15596
rect 29260 15596 29876 15652
rect 29932 16098 30100 16100
rect 29932 16046 30046 16098
rect 30098 16046 30100 16098
rect 29932 16044 30100 16046
rect 29260 15316 29316 15596
rect 29932 15540 29988 16044
rect 30044 16034 30100 16044
rect 28364 14700 28644 14756
rect 28700 15314 29316 15316
rect 28700 15262 29262 15314
rect 29314 15262 29316 15314
rect 28700 15260 29316 15262
rect 28364 14532 28420 14700
rect 28364 14438 28420 14476
rect 28700 14530 28756 15260
rect 29260 15250 29316 15260
rect 29596 15484 29988 15540
rect 29596 15314 29652 15484
rect 29596 15262 29598 15314
rect 29650 15262 29652 15314
rect 28700 14478 28702 14530
rect 28754 14478 28756 14530
rect 28700 14466 28756 14478
rect 28476 14308 28532 14318
rect 28700 14308 28756 14318
rect 28364 14306 28532 14308
rect 28364 14254 28478 14306
rect 28530 14254 28532 14306
rect 28364 14252 28532 14254
rect 28252 13860 28308 13870
rect 28252 13766 28308 13804
rect 27692 13746 27748 13758
rect 27692 13694 27694 13746
rect 27746 13694 27748 13746
rect 27692 12964 27748 13694
rect 27804 13748 27860 13758
rect 28140 13748 28196 13758
rect 27804 13746 28196 13748
rect 27804 13694 27806 13746
rect 27858 13694 28142 13746
rect 28194 13694 28196 13746
rect 27804 13692 28196 13694
rect 27804 13682 27860 13692
rect 28140 13682 28196 13692
rect 28028 13524 28084 13534
rect 28084 13468 28196 13524
rect 28028 13458 28084 13468
rect 27916 12964 27972 12974
rect 27692 12962 27972 12964
rect 27692 12910 27918 12962
rect 27970 12910 27972 12962
rect 27692 12908 27972 12910
rect 27244 9884 27524 9940
rect 27580 11396 27636 11406
rect 27916 11396 27972 12908
rect 28028 12180 28084 12190
rect 28028 12086 28084 12124
rect 28028 11732 28084 11742
rect 28028 11506 28084 11676
rect 28028 11454 28030 11506
rect 28082 11454 28084 11506
rect 28028 11442 28084 11454
rect 27580 11394 27972 11396
rect 27580 11342 27582 11394
rect 27634 11342 27972 11394
rect 27580 11340 27972 11342
rect 27244 7700 27300 9884
rect 27580 9828 27636 11340
rect 28028 11284 28084 11294
rect 28028 11190 28084 11228
rect 28140 11060 28196 13468
rect 28028 11004 28196 11060
rect 28028 10778 28084 11004
rect 28364 10948 28420 14252
rect 28476 14242 28532 14252
rect 28588 14252 28700 14308
rect 28476 13972 28532 13982
rect 28588 13972 28644 14252
rect 28700 14242 28756 14252
rect 29484 14308 29540 14318
rect 29484 14214 29540 14252
rect 28924 14196 28980 14206
rect 28980 14140 29092 14196
rect 28924 14130 28980 14140
rect 28476 13970 28644 13972
rect 28476 13918 28478 13970
rect 28530 13918 28644 13970
rect 28476 13916 28644 13918
rect 28476 13906 28532 13916
rect 28588 13076 28644 13086
rect 28588 12982 28644 13020
rect 28588 12740 28644 12750
rect 28588 12178 28644 12684
rect 28588 12126 28590 12178
rect 28642 12126 28644 12178
rect 28588 12114 28644 12126
rect 28028 10726 28030 10778
rect 28082 10726 28084 10778
rect 28028 10724 28084 10726
rect 27580 9762 27636 9772
rect 27804 10668 28084 10724
rect 28140 10892 28420 10948
rect 28140 10834 28196 10892
rect 28140 10782 28142 10834
rect 28194 10782 28196 10834
rect 27356 9716 27412 9726
rect 27804 9716 27860 10668
rect 28140 10612 28196 10782
rect 28924 10612 28980 10622
rect 27916 10556 28196 10612
rect 28476 10610 28980 10612
rect 28476 10558 28926 10610
rect 28978 10558 28980 10610
rect 28476 10556 28980 10558
rect 27916 9940 27972 10556
rect 28140 10388 28196 10398
rect 28196 10332 28308 10388
rect 28140 10294 28196 10332
rect 27916 9874 27972 9884
rect 27804 9660 28084 9716
rect 27356 9042 27412 9660
rect 27692 9268 27748 9278
rect 27692 9174 27748 9212
rect 27468 9156 27524 9166
rect 27468 9154 27636 9156
rect 27468 9102 27470 9154
rect 27522 9102 27636 9154
rect 27468 9100 27636 9102
rect 27468 9090 27524 9100
rect 27356 8990 27358 9042
rect 27410 8990 27412 9042
rect 27356 8260 27412 8990
rect 27468 8260 27524 8270
rect 27356 8258 27524 8260
rect 27356 8206 27470 8258
rect 27522 8206 27524 8258
rect 27356 8204 27524 8206
rect 27468 8194 27524 8204
rect 27580 8146 27636 9100
rect 27580 8094 27582 8146
rect 27634 8094 27636 8146
rect 27244 7644 27524 7700
rect 27020 7474 27188 7476
rect 27020 7422 27022 7474
rect 27074 7422 27188 7474
rect 27020 7420 27188 7422
rect 27244 7476 27300 7486
rect 27020 7364 27076 7420
rect 27244 7382 27300 7420
rect 27020 7298 27076 7308
rect 26348 6738 26404 6748
rect 25452 6638 25454 6690
rect 25506 6638 25508 6690
rect 25452 6626 25508 6638
rect 25340 6402 25396 6412
rect 27468 4564 27524 7644
rect 27580 7698 27636 8094
rect 27580 7646 27582 7698
rect 27634 7646 27636 7698
rect 27580 7634 27636 7646
rect 28028 7700 28084 9660
rect 28252 9154 28308 10332
rect 28364 9940 28420 9950
rect 28364 9716 28420 9884
rect 28476 9938 28532 10556
rect 28924 10546 28980 10556
rect 28476 9886 28478 9938
rect 28530 9886 28532 9938
rect 28476 9874 28532 9886
rect 29036 9828 29092 14140
rect 29260 13074 29316 13086
rect 29260 13022 29262 13074
rect 29314 13022 29316 13074
rect 29260 11844 29316 13022
rect 29484 12852 29540 12862
rect 29484 12758 29540 12796
rect 29260 11778 29316 11788
rect 29372 10610 29428 10622
rect 29372 10558 29374 10610
rect 29426 10558 29428 10610
rect 29372 10388 29428 10558
rect 29260 9940 29316 9950
rect 29372 9940 29428 10332
rect 29372 9884 29540 9940
rect 29260 9846 29316 9884
rect 28924 9772 29092 9828
rect 28588 9716 28644 9726
rect 28364 9714 28532 9716
rect 28364 9662 28366 9714
rect 28418 9662 28532 9714
rect 28364 9660 28532 9662
rect 28364 9650 28420 9660
rect 28252 9102 28254 9154
rect 28306 9102 28308 9154
rect 28252 9090 28308 9102
rect 28476 9268 28532 9660
rect 28588 9622 28644 9660
rect 28476 9044 28532 9212
rect 28588 9044 28644 9054
rect 28476 9042 28644 9044
rect 28476 8990 28590 9042
rect 28642 8990 28644 9042
rect 28476 8988 28644 8990
rect 28588 8978 28644 8988
rect 28476 8372 28532 8382
rect 28364 8260 28420 8270
rect 28364 8166 28420 8204
rect 28476 8034 28532 8316
rect 28924 8148 28980 9772
rect 29148 9716 29204 9726
rect 29204 9660 29428 9716
rect 29148 9650 29204 9660
rect 29372 9044 29428 9660
rect 29484 9714 29540 9884
rect 29484 9662 29486 9714
rect 29538 9662 29540 9714
rect 29484 9650 29540 9662
rect 29484 9044 29540 9054
rect 29260 9042 29540 9044
rect 29260 8990 29486 9042
rect 29538 8990 29540 9042
rect 29260 8988 29540 8990
rect 28476 7982 28478 8034
rect 28530 7982 28532 8034
rect 28476 7970 28532 7982
rect 28812 8092 28980 8148
rect 29148 8148 29204 8158
rect 27804 7588 27860 7598
rect 27692 7364 27748 7374
rect 27692 6692 27748 7308
rect 27804 6804 27860 7532
rect 28028 7586 28084 7644
rect 28028 7534 28030 7586
rect 28082 7534 28084 7586
rect 28028 7522 28084 7534
rect 28140 7476 28196 7486
rect 27804 6748 27972 6804
rect 27692 6636 27860 6692
rect 27804 6578 27860 6636
rect 27804 6526 27806 6578
rect 27858 6526 27860 6578
rect 27804 6514 27860 6526
rect 27916 6578 27972 6748
rect 28140 6690 28196 7420
rect 28140 6638 28142 6690
rect 28194 6638 28196 6690
rect 28140 6626 28196 6638
rect 27916 6526 27918 6578
rect 27970 6526 27972 6578
rect 27916 6514 27972 6526
rect 28588 5236 28644 5246
rect 28364 5124 28420 5134
rect 28364 5030 28420 5068
rect 28588 5010 28644 5180
rect 28588 4958 28590 5010
rect 28642 4958 28644 5010
rect 28588 4946 28644 4958
rect 28700 4900 28756 4910
rect 27692 4564 27748 4574
rect 27468 4562 27748 4564
rect 27468 4510 27694 4562
rect 27746 4510 27748 4562
rect 27468 4508 27748 4510
rect 25340 4228 25396 4238
rect 24556 3442 24724 3444
rect 24556 3390 24558 3442
rect 24610 3390 24724 3442
rect 24556 3388 24724 3390
rect 24892 4226 25396 4228
rect 24892 4174 25342 4226
rect 25394 4174 25396 4226
rect 24892 4172 25396 4174
rect 24892 3554 24948 4172
rect 25340 4162 25396 4172
rect 26796 3668 26852 3678
rect 26796 3666 26964 3668
rect 26796 3614 26798 3666
rect 26850 3614 26964 3666
rect 26796 3612 26964 3614
rect 26796 3602 26852 3612
rect 24892 3502 24894 3554
rect 24946 3502 24948 3554
rect 24556 3378 24612 3388
rect 24892 800 24948 3502
rect 26908 800 26964 3612
rect 27692 3554 27748 4508
rect 28252 4228 28308 4238
rect 28252 4226 28420 4228
rect 28252 4174 28254 4226
rect 28306 4174 28420 4226
rect 28252 4172 28420 4174
rect 28252 4162 28308 4172
rect 27692 3502 27694 3554
rect 27746 3502 27748 3554
rect 27692 3490 27748 3502
rect 28364 3444 28420 4172
rect 28364 3378 28420 3388
rect 28476 4116 28532 4126
rect 28476 2100 28532 4060
rect 28700 3442 28756 4844
rect 28812 4564 28868 8092
rect 29148 8054 29204 8092
rect 29148 7476 29204 7486
rect 29148 7382 29204 7420
rect 28924 7364 28980 7374
rect 28924 6804 28980 7308
rect 29260 7250 29316 8988
rect 29484 8978 29540 8988
rect 29484 8708 29540 8718
rect 29372 8372 29428 8382
rect 29372 8278 29428 8316
rect 29260 7198 29262 7250
rect 29314 7198 29316 7250
rect 29260 7186 29316 7198
rect 28924 6738 28980 6748
rect 29484 5906 29540 8652
rect 29596 8372 29652 15262
rect 29708 15316 29764 15326
rect 29708 15222 29764 15260
rect 30156 15148 30212 16716
rect 30380 15876 30436 15886
rect 30380 15782 30436 15820
rect 30380 15314 30436 15326
rect 30380 15262 30382 15314
rect 30434 15262 30436 15314
rect 30380 15204 30436 15262
rect 30492 15204 30548 15214
rect 30380 15148 30492 15204
rect 29708 15092 29764 15102
rect 29708 14532 29764 15036
rect 29820 15092 30212 15148
rect 29820 14754 29876 15092
rect 29820 14702 29822 14754
rect 29874 14702 29876 14754
rect 29820 14690 29876 14702
rect 29708 14438 29764 14476
rect 30044 14530 30100 14542
rect 30044 14478 30046 14530
rect 30098 14478 30100 14530
rect 30044 14420 30100 14478
rect 30268 14532 30324 14542
rect 30268 14438 30324 14476
rect 30044 14354 30100 14364
rect 30380 14418 30436 14430
rect 30380 14366 30382 14418
rect 30434 14366 30436 14418
rect 30380 14308 30436 14366
rect 30380 14242 30436 14252
rect 30268 13858 30324 13870
rect 30268 13806 30270 13858
rect 30322 13806 30324 13858
rect 30268 12852 30324 13806
rect 30268 12786 30324 12796
rect 30492 12628 30548 15148
rect 30156 12572 30548 12628
rect 30156 10722 30212 12572
rect 30604 12292 30660 17724
rect 30716 17668 30772 17678
rect 30716 13972 30772 17612
rect 30828 14642 30884 18172
rect 31164 17778 31220 18284
rect 31164 17726 31166 17778
rect 31218 17726 31220 17778
rect 31052 17666 31108 17678
rect 31052 17614 31054 17666
rect 31106 17614 31108 17666
rect 31052 17556 31108 17614
rect 31052 17490 31108 17500
rect 31052 15428 31108 15438
rect 31164 15428 31220 17726
rect 31276 16660 31332 18510
rect 31388 18340 31444 18350
rect 31388 17108 31444 18284
rect 31500 17890 31556 18620
rect 31500 17838 31502 17890
rect 31554 17838 31556 17890
rect 31500 17826 31556 17838
rect 31388 16882 31444 17052
rect 31388 16830 31390 16882
rect 31442 16830 31444 16882
rect 31388 16818 31444 16830
rect 31500 16884 31556 16894
rect 31612 16884 31668 19180
rect 31724 18676 31780 19628
rect 31836 19012 31892 20300
rect 31836 18946 31892 18956
rect 31724 18610 31780 18620
rect 31948 18452 32004 21308
rect 32060 20690 32116 20702
rect 32060 20638 32062 20690
rect 32114 20638 32116 20690
rect 32060 20020 32116 20638
rect 32060 19010 32116 19964
rect 32060 18958 32062 19010
rect 32114 18958 32116 19010
rect 32060 18946 32116 18958
rect 32172 19234 32228 19246
rect 32172 19182 32174 19234
rect 32226 19182 32228 19234
rect 32172 18676 32228 19182
rect 32172 18610 32228 18620
rect 31948 18396 32228 18452
rect 31836 18340 31892 18350
rect 31836 18246 31892 18284
rect 32060 18226 32116 18238
rect 32060 18174 32062 18226
rect 32114 18174 32116 18226
rect 32060 16884 32116 18174
rect 31612 16828 31892 16884
rect 31500 16770 31556 16828
rect 31500 16718 31502 16770
rect 31554 16718 31556 16770
rect 31276 16604 31444 16660
rect 31052 15426 31220 15428
rect 31052 15374 31054 15426
rect 31106 15374 31220 15426
rect 31052 15372 31220 15374
rect 31052 15362 31108 15372
rect 30940 15316 30996 15326
rect 30940 15222 30996 15260
rect 31276 15316 31332 15326
rect 31276 15222 31332 15260
rect 30828 14590 30830 14642
rect 30882 14590 30884 14642
rect 30828 14420 30884 14590
rect 31276 14532 31332 14542
rect 31276 14438 31332 14476
rect 30828 14364 31220 14420
rect 30716 13916 31108 13972
rect 30716 13746 30772 13758
rect 30716 13694 30718 13746
rect 30770 13694 30772 13746
rect 30716 12740 30772 13694
rect 30716 12684 30996 12740
rect 30940 12292 30996 12684
rect 31052 12516 31108 13916
rect 31164 13746 31220 14364
rect 31276 13972 31332 13982
rect 31388 13972 31444 16604
rect 31500 15538 31556 16718
rect 31836 16770 31892 16828
rect 32060 16818 32116 16828
rect 31836 16718 31838 16770
rect 31890 16718 31892 16770
rect 31836 16706 31892 16718
rect 31500 15486 31502 15538
rect 31554 15486 31556 15538
rect 31500 15474 31556 15486
rect 31836 15876 31892 15886
rect 31612 15314 31668 15326
rect 31612 15262 31614 15314
rect 31666 15262 31668 15314
rect 31612 15204 31668 15262
rect 31836 15314 31892 15820
rect 31836 15262 31838 15314
rect 31890 15262 31892 15314
rect 31836 15250 31892 15262
rect 31612 15138 31668 15148
rect 31276 13970 31444 13972
rect 31276 13918 31278 13970
rect 31330 13918 31444 13970
rect 31276 13916 31444 13918
rect 31500 14532 31556 14542
rect 31276 13906 31332 13916
rect 31164 13694 31166 13746
rect 31218 13694 31220 13746
rect 31164 13682 31220 13694
rect 31388 13076 31444 13086
rect 31500 13076 31556 14476
rect 31388 13074 31556 13076
rect 31388 13022 31390 13074
rect 31442 13022 31556 13074
rect 31388 13020 31556 13022
rect 31388 13010 31444 13020
rect 31164 12852 31220 12862
rect 31164 12850 31444 12852
rect 31164 12798 31166 12850
rect 31218 12798 31444 12850
rect 31164 12796 31444 12798
rect 31164 12786 31220 12796
rect 31052 12460 31220 12516
rect 31052 12292 31108 12302
rect 30604 12236 30884 12292
rect 30940 12290 31108 12292
rect 30940 12238 31054 12290
rect 31106 12238 31108 12290
rect 30940 12236 31108 12238
rect 30156 10670 30158 10722
rect 30210 10670 30212 10722
rect 30156 10658 30212 10670
rect 30380 12178 30436 12190
rect 30380 12126 30382 12178
rect 30434 12126 30436 12178
rect 30380 11844 30436 12126
rect 29820 10610 29876 10622
rect 29820 10558 29822 10610
rect 29874 10558 29876 10610
rect 29708 8372 29764 8382
rect 29596 8370 29764 8372
rect 29596 8318 29710 8370
rect 29762 8318 29764 8370
rect 29596 8316 29764 8318
rect 29708 8306 29764 8316
rect 29820 8372 29876 10558
rect 30380 10498 30436 11788
rect 30604 12066 30660 12078
rect 30604 12014 30606 12066
rect 30658 12014 30660 12066
rect 30604 10612 30660 12014
rect 30380 10446 30382 10498
rect 30434 10446 30436 10498
rect 30380 10434 30436 10446
rect 30492 10610 30660 10612
rect 30492 10558 30606 10610
rect 30658 10558 30660 10610
rect 30492 10556 30660 10558
rect 30492 10276 30548 10556
rect 30604 10546 30660 10556
rect 30156 10220 30548 10276
rect 30156 9154 30212 10220
rect 30716 9828 30772 9838
rect 30156 9102 30158 9154
rect 30210 9102 30212 9154
rect 30156 9090 30212 9102
rect 30268 9826 30772 9828
rect 30268 9774 30718 9826
rect 30770 9774 30772 9826
rect 30268 9772 30772 9774
rect 29820 8306 29876 8316
rect 30268 8260 30324 9772
rect 30716 9762 30772 9772
rect 30828 9716 30884 12236
rect 31052 12226 31108 12236
rect 30828 9660 30996 9716
rect 30716 9492 30772 9502
rect 30604 9436 30716 9492
rect 30604 9266 30660 9436
rect 30716 9426 30772 9436
rect 30604 9214 30606 9266
rect 30658 9214 30660 9266
rect 30492 9042 30548 9054
rect 30492 8990 30494 9042
rect 30546 8990 30548 9042
rect 30492 8372 30548 8990
rect 30492 8306 30548 8316
rect 30268 7700 30324 8204
rect 30604 8260 30660 9214
rect 30828 9268 30884 9278
rect 30828 9174 30884 9212
rect 30604 8194 30660 8204
rect 30156 7644 30324 7700
rect 30156 7586 30212 7644
rect 30156 7534 30158 7586
rect 30210 7534 30212 7586
rect 30156 7522 30212 7534
rect 30268 7474 30324 7486
rect 30268 7422 30270 7474
rect 30322 7422 30324 7474
rect 30268 7364 30324 7422
rect 30604 7476 30660 7486
rect 30604 7382 30660 7420
rect 30268 7298 30324 7308
rect 30940 6692 30996 9660
rect 31164 9492 31220 12460
rect 31388 9938 31444 12796
rect 32172 11844 32228 18396
rect 32172 11778 32228 11788
rect 31948 10500 32004 10510
rect 31948 10406 32004 10444
rect 31388 9886 31390 9938
rect 31442 9886 31444 9938
rect 31388 9874 31444 9886
rect 32172 10386 32228 10398
rect 32172 10334 32174 10386
rect 32226 10334 32228 10386
rect 32172 9716 32228 10334
rect 32284 10164 32340 21420
rect 32396 21410 32452 21420
rect 32508 20916 32564 20926
rect 32508 20822 32564 20860
rect 32396 20802 32452 20814
rect 32396 20750 32398 20802
rect 32450 20750 32452 20802
rect 32396 18674 32452 20750
rect 32620 20692 32676 21644
rect 32732 21476 32788 23492
rect 32732 21410 32788 21420
rect 32844 21812 32900 21822
rect 32620 20130 32676 20636
rect 32844 20802 32900 21756
rect 33180 21812 33236 23548
rect 33180 21718 33236 21756
rect 32844 20750 32846 20802
rect 32898 20750 32900 20802
rect 32844 20244 32900 20750
rect 32844 20178 32900 20188
rect 32620 20078 32622 20130
rect 32674 20078 32676 20130
rect 32620 20066 32676 20078
rect 33068 20018 33124 20030
rect 33068 19966 33070 20018
rect 33122 19966 33124 20018
rect 33068 19458 33124 19966
rect 33292 20020 33348 20030
rect 33292 19926 33348 19964
rect 33068 19406 33070 19458
rect 33122 19406 33124 19458
rect 33068 19394 33124 19406
rect 32732 19236 32788 19246
rect 32732 19142 32788 19180
rect 32508 19124 32564 19134
rect 32508 19030 32564 19068
rect 32396 18622 32398 18674
rect 32450 18622 32452 18674
rect 32396 18610 32452 18622
rect 32732 19012 32788 19022
rect 32732 17778 32788 18956
rect 33292 18676 33348 18686
rect 33292 18582 33348 18620
rect 33404 18452 33460 25004
rect 33516 24836 33572 24846
rect 33628 24836 33684 26236
rect 33740 26226 33796 26236
rect 33516 24834 33684 24836
rect 33516 24782 33518 24834
rect 33570 24782 33684 24834
rect 33516 24780 33684 24782
rect 33516 24770 33572 24780
rect 33628 24052 33684 24780
rect 33628 23986 33684 23996
rect 33740 25396 33796 25406
rect 33740 24050 33796 25340
rect 33740 23998 33742 24050
rect 33794 23998 33796 24050
rect 33740 23548 33796 23998
rect 33628 23492 33796 23548
rect 33852 23548 33908 26460
rect 34076 26292 34132 26302
rect 34076 26198 34132 26236
rect 33964 26178 34020 26190
rect 33964 26126 33966 26178
rect 34018 26126 34020 26178
rect 33964 25732 34020 26126
rect 33964 25666 34020 25676
rect 34076 26068 34132 26078
rect 33852 23492 34020 23548
rect 33628 21812 33684 23492
rect 33964 23156 34020 23492
rect 33852 23154 34020 23156
rect 33852 23102 33966 23154
rect 34018 23102 34020 23154
rect 33852 23100 34020 23102
rect 33852 22258 33908 23100
rect 33964 23090 34020 23100
rect 34076 22820 34132 26012
rect 34188 25506 34244 26852
rect 34188 25454 34190 25506
rect 34242 25454 34244 25506
rect 34188 25442 34244 25454
rect 34300 24948 34356 28028
rect 34524 27748 34580 27758
rect 34524 27412 34580 27692
rect 34636 27524 34692 29374
rect 34748 28756 34804 29486
rect 34748 28690 34804 28700
rect 34748 28420 34804 28430
rect 34748 28326 34804 28364
rect 34636 27458 34692 27468
rect 34748 27860 34804 27870
rect 34524 27346 34580 27356
rect 34748 27300 34804 27804
rect 34748 27234 34804 27244
rect 34860 27076 34916 30268
rect 34972 30100 35028 30110
rect 34972 30006 35028 30044
rect 35084 28642 35140 30268
rect 35196 30212 35252 30380
rect 35308 30212 35364 30222
rect 35196 30156 35308 30212
rect 35308 29426 35364 30156
rect 35308 29374 35310 29426
rect 35362 29374 35364 29426
rect 35308 29362 35364 29374
rect 35532 29538 35588 29550
rect 35532 29486 35534 29538
rect 35586 29486 35588 29538
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35420 28868 35476 28878
rect 35532 28868 35588 29486
rect 35476 28812 35588 28868
rect 35420 28802 35476 28812
rect 35084 28590 35086 28642
rect 35138 28590 35140 28642
rect 34972 28532 35028 28542
rect 34972 28196 35028 28476
rect 34972 28130 35028 28140
rect 34972 27858 35028 27870
rect 34972 27806 34974 27858
rect 35026 27806 35028 27858
rect 34972 27412 35028 27806
rect 35084 27860 35140 28590
rect 35084 27794 35140 27804
rect 35196 28756 35252 28766
rect 35644 28756 35700 31052
rect 35756 29986 35812 29998
rect 35756 29934 35758 29986
rect 35810 29934 35812 29986
rect 35756 29540 35812 29934
rect 36204 29988 36260 31052
rect 36316 30882 36372 33180
rect 36428 33124 36484 35420
rect 36876 34692 36932 34702
rect 36876 34598 36932 34636
rect 36652 34018 36708 34030
rect 36652 33966 36654 34018
rect 36706 33966 36708 34018
rect 36652 33684 36708 33966
rect 36652 33618 36708 33628
rect 36428 33058 36484 33068
rect 36540 33236 36596 33246
rect 36428 31780 36484 31790
rect 36428 31686 36484 31724
rect 36428 31332 36484 31342
rect 36428 31218 36484 31276
rect 36428 31166 36430 31218
rect 36482 31166 36484 31218
rect 36428 31154 36484 31166
rect 36316 30830 36318 30882
rect 36370 30830 36372 30882
rect 36316 30818 36372 30830
rect 36540 30548 36596 33180
rect 36988 31556 37044 37772
rect 37100 37762 37156 37772
rect 37548 37492 37604 39004
rect 37660 38836 37716 38846
rect 37660 38742 37716 38780
rect 37772 38722 37828 39116
rect 37772 38670 37774 38722
rect 37826 38670 37828 38722
rect 37772 38658 37828 38670
rect 37884 38050 37940 39340
rect 38332 38668 38388 39900
rect 37884 37998 37886 38050
rect 37938 37998 37940 38050
rect 37884 37986 37940 37998
rect 37996 38612 38388 38668
rect 38556 38834 38612 38846
rect 38556 38782 38558 38834
rect 38610 38782 38612 38834
rect 37324 37490 37604 37492
rect 37324 37438 37550 37490
rect 37602 37438 37604 37490
rect 37324 37436 37604 37438
rect 37212 37268 37268 37278
rect 37212 37174 37268 37212
rect 37324 36482 37380 37436
rect 37548 37426 37604 37436
rect 37436 37268 37492 37278
rect 37436 37174 37492 37212
rect 37772 37266 37828 37278
rect 37772 37214 37774 37266
rect 37826 37214 37828 37266
rect 37772 37156 37828 37214
rect 37772 37090 37828 37100
rect 37660 37044 37716 37054
rect 37660 36932 37716 36988
rect 37660 36876 37828 36932
rect 37324 36430 37326 36482
rect 37378 36430 37380 36482
rect 37324 36418 37380 36430
rect 37548 36258 37604 36270
rect 37548 36206 37550 36258
rect 37602 36206 37604 36258
rect 37548 35700 37604 36206
rect 37548 35634 37604 35644
rect 37660 35586 37716 35598
rect 37660 35534 37662 35586
rect 37714 35534 37716 35586
rect 37100 35476 37156 35486
rect 37660 35476 37716 35534
rect 37100 34802 37156 35420
rect 37548 35420 37660 35476
rect 37100 34750 37102 34802
rect 37154 34750 37156 34802
rect 37100 34738 37156 34750
rect 37212 35140 37268 35150
rect 37212 34802 37268 35084
rect 37212 34750 37214 34802
rect 37266 34750 37268 34802
rect 37212 33684 37268 34750
rect 37548 34354 37604 35420
rect 37660 35410 37716 35420
rect 37772 35028 37828 36876
rect 37996 35924 38052 38612
rect 38220 37828 38276 37838
rect 38220 37734 38276 37772
rect 38556 37380 38612 38782
rect 38780 38164 38836 43932
rect 39004 43876 39060 43886
rect 39004 43204 39060 43820
rect 39340 43652 39396 52892
rect 39452 52724 39508 52734
rect 39452 52164 39508 52668
rect 39564 52388 39620 52892
rect 39676 52834 39732 52846
rect 39676 52782 39678 52834
rect 39730 52782 39732 52834
rect 39676 52500 39732 52782
rect 39788 52724 39844 53900
rect 40012 53844 40068 55244
rect 40124 55298 40292 55300
rect 40124 55246 40126 55298
rect 40178 55246 40292 55298
rect 40124 55244 40292 55246
rect 40124 55234 40180 55244
rect 40124 54628 40180 54638
rect 40124 54514 40180 54572
rect 40124 54462 40126 54514
rect 40178 54462 40180 54514
rect 40124 54450 40180 54462
rect 39900 53732 39956 53742
rect 40012 53732 40068 53788
rect 39900 53730 40068 53732
rect 39900 53678 39902 53730
rect 39954 53678 40068 53730
rect 39900 53676 40068 53678
rect 40236 53956 40292 55244
rect 40460 55076 40516 55086
rect 40460 54982 40516 55020
rect 40236 53730 40292 53900
rect 40236 53678 40238 53730
rect 40290 53678 40292 53730
rect 39900 53666 39956 53676
rect 40236 53666 40292 53678
rect 39788 52658 39844 52668
rect 39900 53508 39956 53518
rect 39676 52444 39844 52500
rect 39564 52332 39732 52388
rect 39452 51602 39508 52108
rect 39564 52052 39620 52062
rect 39564 51958 39620 51996
rect 39452 51550 39454 51602
rect 39506 51550 39508 51602
rect 39452 51538 39508 51550
rect 39452 50706 39508 50718
rect 39452 50654 39454 50706
rect 39506 50654 39508 50706
rect 39452 49252 39508 50654
rect 39452 49186 39508 49196
rect 39564 49812 39620 49822
rect 39564 49026 39620 49756
rect 39564 48974 39566 49026
rect 39618 48974 39620 49026
rect 39564 48962 39620 48974
rect 39452 48580 39508 48590
rect 39452 47460 39508 48524
rect 39452 47346 39508 47404
rect 39452 47294 39454 47346
rect 39506 47294 39508 47346
rect 39452 47282 39508 47294
rect 39564 47346 39620 47358
rect 39564 47294 39566 47346
rect 39618 47294 39620 47346
rect 39564 47124 39620 47294
rect 39564 47058 39620 47068
rect 39564 46450 39620 46462
rect 39564 46398 39566 46450
rect 39618 46398 39620 46450
rect 39564 45892 39620 46398
rect 39564 45826 39620 45836
rect 39676 45668 39732 52332
rect 39788 51268 39844 52444
rect 39900 51604 39956 53452
rect 40012 53506 40068 53518
rect 40012 53454 40014 53506
rect 40066 53454 40068 53506
rect 40012 52948 40068 53454
rect 40124 52948 40180 52958
rect 40012 52892 40124 52948
rect 40124 52854 40180 52892
rect 40012 52276 40068 52286
rect 40012 52162 40068 52220
rect 40012 52110 40014 52162
rect 40066 52110 40068 52162
rect 40012 52098 40068 52110
rect 39900 51538 39956 51548
rect 39788 51202 39844 51212
rect 40348 50596 40404 50606
rect 40348 50502 40404 50540
rect 40684 50428 40740 56142
rect 40908 55300 40964 59276
rect 49728 59200 49840 60000
rect 50400 59200 50512 60000
rect 41020 56308 41076 56318
rect 41020 56214 41076 56252
rect 43036 56308 43092 56318
rect 43036 56214 43092 56252
rect 49756 56308 49812 59200
rect 50428 56754 50484 59200
rect 50428 56702 50430 56754
rect 50482 56702 50484 56754
rect 50428 56690 50484 56702
rect 51212 56754 51268 56766
rect 51212 56702 51214 56754
rect 51266 56702 51268 56754
rect 50556 56476 50820 56486
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50556 56410 50820 56420
rect 49756 56306 50036 56308
rect 49756 56254 49758 56306
rect 49810 56254 50036 56306
rect 49756 56252 50036 56254
rect 49756 56242 49812 56252
rect 41356 56194 41412 56206
rect 41356 56142 41358 56194
rect 41410 56142 41412 56194
rect 41020 55300 41076 55310
rect 40908 55244 41020 55300
rect 41020 55206 41076 55244
rect 40796 55074 40852 55086
rect 40796 55022 40798 55074
rect 40850 55022 40852 55074
rect 40796 52388 40852 55022
rect 41020 54628 41076 54638
rect 41020 54534 41076 54572
rect 41356 54068 41412 56142
rect 41580 56196 41636 56206
rect 41580 56082 41636 56140
rect 43708 56196 43764 56206
rect 43708 56102 43764 56140
rect 49980 56194 50036 56252
rect 51212 56306 51268 56702
rect 51212 56254 51214 56306
rect 51266 56254 51268 56306
rect 49980 56142 49982 56194
rect 50034 56142 50036 56194
rect 49980 56130 50036 56142
rect 50316 56194 50372 56206
rect 50316 56142 50318 56194
rect 50370 56142 50372 56194
rect 41580 56030 41582 56082
rect 41634 56030 41636 56082
rect 41580 56018 41636 56030
rect 42588 56084 42644 56094
rect 42588 55990 42644 56028
rect 42140 55972 42196 55982
rect 42140 55878 42196 55916
rect 42028 55412 42084 55422
rect 42028 55318 42084 55356
rect 42476 55300 42532 55310
rect 42476 55206 42532 55244
rect 41580 55188 41636 55198
rect 41580 55094 41636 55132
rect 41356 54002 41412 54012
rect 42588 53620 42644 53630
rect 42364 53508 42420 53518
rect 42588 53508 42644 53564
rect 43372 53618 43428 53630
rect 43372 53566 43374 53618
rect 43426 53566 43428 53618
rect 42364 53506 42644 53508
rect 42364 53454 42366 53506
rect 42418 53454 42644 53506
rect 42364 53452 42644 53454
rect 42700 53508 42756 53518
rect 42924 53508 42980 53518
rect 42364 53396 42420 53452
rect 42700 53414 42756 53452
rect 42812 53506 42980 53508
rect 42812 53454 42926 53506
rect 42978 53454 42980 53506
rect 42812 53452 42980 53454
rect 42364 53330 42420 53340
rect 41020 53172 41076 53182
rect 41020 53078 41076 53116
rect 41132 53060 41188 53070
rect 40908 52948 40964 52958
rect 40908 52854 40964 52892
rect 41132 52388 41188 53004
rect 40796 52332 40964 52388
rect 40908 51940 40964 52332
rect 40572 50372 40740 50428
rect 40796 51884 40964 51940
rect 41020 52332 41132 52388
rect 40124 48692 40180 48702
rect 40124 48354 40180 48636
rect 40124 48302 40126 48354
rect 40178 48302 40180 48354
rect 40124 48290 40180 48302
rect 40236 48466 40292 48478
rect 40236 48414 40238 48466
rect 40290 48414 40292 48466
rect 40124 47012 40180 47022
rect 40012 46788 40068 46798
rect 40012 46694 40068 46732
rect 40124 46786 40180 46956
rect 40236 46900 40292 48414
rect 40236 46834 40292 46844
rect 40124 46734 40126 46786
rect 40178 46734 40180 46786
rect 40124 46722 40180 46734
rect 40348 46674 40404 46686
rect 40348 46622 40350 46674
rect 40402 46622 40404 46674
rect 40348 46564 40404 46622
rect 40348 46498 40404 46508
rect 40572 46116 40628 50372
rect 40684 49026 40740 49038
rect 40684 48974 40686 49026
rect 40738 48974 40740 49026
rect 40684 48692 40740 48974
rect 40684 48626 40740 48636
rect 40796 46676 40852 51884
rect 40908 51380 40964 51390
rect 41020 51380 41076 52332
rect 41132 52294 41188 52332
rect 41356 53058 41412 53070
rect 41356 53006 41358 53058
rect 41410 53006 41412 53058
rect 41356 52836 41412 53006
rect 42700 52948 42756 52958
rect 42812 52948 42868 53452
rect 42924 53442 42980 53452
rect 43036 53506 43092 53518
rect 43036 53454 43038 53506
rect 43090 53454 43092 53506
rect 43036 53284 43092 53454
rect 42700 52946 42812 52948
rect 42700 52894 42702 52946
rect 42754 52894 42812 52946
rect 42700 52892 42812 52894
rect 42700 52882 42756 52892
rect 42812 52854 42868 52892
rect 42924 53228 43092 53284
rect 43260 53506 43316 53518
rect 43260 53454 43262 53506
rect 43314 53454 43316 53506
rect 42924 52946 42980 53228
rect 42924 52894 42926 52946
rect 42978 52894 42980 52946
rect 41356 52276 41412 52780
rect 42028 52836 42084 52846
rect 42028 52742 42084 52780
rect 42924 52836 42980 52894
rect 42924 52770 42980 52780
rect 42700 52388 42756 52398
rect 42756 52332 42868 52388
rect 42700 52322 42756 52332
rect 41132 52164 41188 52174
rect 41132 52070 41188 52108
rect 40908 51378 41076 51380
rect 40908 51326 40910 51378
rect 40962 51326 41076 51378
rect 40908 51324 41076 51326
rect 41356 51378 41412 52220
rect 42476 52164 42532 52174
rect 41916 52162 42532 52164
rect 41916 52110 42478 52162
rect 42530 52110 42532 52162
rect 41916 52108 42532 52110
rect 41804 52052 41860 52062
rect 41356 51326 41358 51378
rect 41410 51326 41412 51378
rect 40908 51314 40964 51324
rect 41356 51314 41412 51326
rect 41692 52050 41860 52052
rect 41692 51998 41806 52050
rect 41858 51998 41860 52050
rect 41692 51996 41860 51998
rect 41132 51268 41188 51278
rect 41132 51174 41188 51212
rect 41244 51156 41300 51166
rect 41244 50594 41300 51100
rect 41244 50542 41246 50594
rect 41298 50542 41300 50594
rect 41244 50530 41300 50542
rect 41468 49810 41524 49822
rect 41468 49758 41470 49810
rect 41522 49758 41524 49810
rect 41468 49028 41524 49758
rect 41468 48962 41524 48972
rect 41356 48914 41412 48926
rect 41356 48862 41358 48914
rect 41410 48862 41412 48914
rect 41132 47234 41188 47246
rect 41132 47182 41134 47234
rect 41186 47182 41188 47234
rect 41132 47012 41188 47182
rect 41020 46956 41132 47012
rect 40796 46620 40964 46676
rect 40908 46116 40964 46620
rect 41020 46674 41076 46956
rect 41132 46946 41188 46956
rect 41020 46622 41022 46674
rect 41074 46622 41076 46674
rect 41020 46610 41076 46622
rect 41244 46786 41300 46798
rect 41244 46734 41246 46786
rect 41298 46734 41300 46786
rect 41244 46676 41300 46734
rect 41244 46610 41300 46620
rect 40908 46060 41300 46116
rect 40572 46050 40628 46060
rect 39564 45612 39732 45668
rect 39788 46004 39844 46014
rect 39788 45778 39844 45948
rect 40908 45892 40964 45902
rect 40908 45798 40964 45836
rect 39788 45726 39790 45778
rect 39842 45726 39844 45778
rect 39452 43988 39508 43998
rect 39564 43988 39620 45612
rect 39788 44210 39844 45726
rect 40572 45780 40628 45790
rect 40796 45780 40852 45790
rect 40628 45724 40740 45780
rect 40572 45714 40628 45724
rect 39788 44158 39790 44210
rect 39842 44158 39844 44210
rect 39788 44146 39844 44158
rect 40236 45666 40292 45678
rect 40236 45614 40238 45666
rect 40290 45614 40292 45666
rect 39508 43932 39620 43988
rect 39676 44098 39732 44110
rect 39676 44046 39678 44098
rect 39730 44046 39732 44098
rect 39452 43922 39508 43932
rect 39676 43708 39732 44046
rect 39340 43586 39396 43596
rect 39564 43652 39732 43708
rect 38892 42868 38948 42878
rect 38892 42754 38948 42812
rect 39004 42866 39060 43148
rect 39004 42814 39006 42866
rect 39058 42814 39060 42866
rect 39004 42802 39060 42814
rect 38892 42702 38894 42754
rect 38946 42702 38948 42754
rect 38892 42690 38948 42702
rect 39228 42082 39284 42094
rect 39228 42030 39230 42082
rect 39282 42030 39284 42082
rect 38892 41972 38948 41982
rect 39228 41972 39284 42030
rect 38892 41970 39284 41972
rect 38892 41918 38894 41970
rect 38946 41918 39284 41970
rect 38892 41916 39284 41918
rect 38892 41906 38948 41916
rect 38892 41746 38948 41758
rect 38892 41694 38894 41746
rect 38946 41694 38948 41746
rect 38892 40402 38948 41694
rect 39228 41300 39284 41916
rect 39564 41972 39620 43652
rect 40236 43540 40292 45614
rect 40684 45666 40740 45724
rect 40796 45686 40852 45724
rect 40684 45614 40686 45666
rect 40738 45614 40740 45666
rect 40684 45602 40740 45614
rect 40460 44436 40516 44446
rect 40460 44342 40516 44380
rect 40796 44210 40852 44222
rect 40796 44158 40798 44210
rect 40850 44158 40852 44210
rect 40796 43764 40852 44158
rect 40796 43708 41076 43764
rect 41244 43708 41300 46060
rect 41356 46004 41412 48862
rect 41692 48692 41748 51996
rect 41804 51986 41860 51996
rect 41804 51380 41860 51390
rect 41804 51286 41860 51324
rect 41916 51268 41972 52108
rect 42476 52098 42532 52108
rect 42588 52164 42644 52174
rect 42588 52070 42644 52108
rect 42812 52162 42868 52332
rect 42812 52110 42814 52162
rect 42866 52110 42868 52162
rect 42812 52098 42868 52110
rect 43260 52162 43316 53454
rect 43372 53396 43428 53566
rect 44828 53618 44884 53630
rect 44828 53566 44830 53618
rect 44882 53566 44884 53618
rect 43372 53330 43428 53340
rect 44380 53508 44436 53518
rect 44268 53060 44324 53070
rect 43820 53058 44324 53060
rect 43820 53006 44270 53058
rect 44322 53006 44324 53058
rect 43820 53004 44324 53006
rect 43372 52948 43428 52958
rect 43372 52854 43428 52892
rect 43596 52836 43652 52846
rect 43596 52742 43652 52780
rect 43260 52110 43262 52162
rect 43314 52110 43316 52162
rect 43260 51828 43316 52110
rect 43260 51762 43316 51772
rect 43596 52388 43652 52398
rect 43596 52274 43652 52332
rect 43596 52222 43598 52274
rect 43650 52222 43652 52274
rect 42588 51604 42644 51614
rect 42924 51604 42980 51614
rect 42644 51548 42756 51604
rect 42476 51492 42532 51502
rect 42476 51380 42532 51436
rect 41916 50706 41972 51212
rect 41916 50654 41918 50706
rect 41970 50654 41972 50706
rect 41916 50642 41972 50654
rect 42140 51378 42532 51380
rect 42140 51326 42478 51378
rect 42530 51326 42532 51378
rect 42140 51324 42532 51326
rect 42140 50428 42196 51324
rect 42476 51314 42532 51324
rect 42588 51044 42644 51548
rect 42700 51490 42756 51548
rect 42924 51510 42980 51548
rect 42700 51438 42702 51490
rect 42754 51438 42756 51490
rect 42700 51426 42756 51438
rect 43036 51380 43092 51390
rect 43484 51380 43540 51390
rect 43092 51324 43204 51380
rect 43036 51286 43092 51324
rect 41916 50372 42196 50428
rect 42252 50988 42644 51044
rect 42812 51266 42868 51278
rect 42812 51214 42814 51266
rect 42866 51214 42868 51266
rect 41804 50036 41860 50046
rect 41916 50036 41972 50372
rect 41804 50034 41972 50036
rect 41804 49982 41806 50034
rect 41858 49982 41972 50034
rect 41804 49980 41972 49982
rect 42252 50034 42308 50988
rect 42252 49982 42254 50034
rect 42306 49982 42308 50034
rect 41804 49970 41860 49980
rect 42252 49970 42308 49982
rect 42476 50820 42532 50830
rect 42812 50820 42868 51214
rect 42812 50764 43092 50820
rect 41692 48356 41748 48636
rect 41692 48354 41972 48356
rect 41692 48302 41694 48354
rect 41746 48302 41972 48354
rect 41692 48300 41972 48302
rect 41692 48290 41748 48300
rect 41916 47570 41972 48300
rect 41916 47518 41918 47570
rect 41970 47518 41972 47570
rect 41916 47506 41972 47518
rect 42028 48244 42084 48254
rect 42028 47460 42084 48188
rect 42140 47460 42196 47470
rect 42028 47458 42196 47460
rect 42028 47406 42142 47458
rect 42194 47406 42196 47458
rect 42028 47404 42196 47406
rect 42140 47394 42196 47404
rect 41468 47234 41524 47246
rect 41468 47182 41470 47234
rect 41522 47182 41524 47234
rect 41468 47124 41524 47182
rect 41468 47058 41524 47068
rect 42140 46900 42196 46910
rect 41468 46788 41524 46798
rect 41468 46674 41524 46732
rect 42028 46786 42084 46798
rect 42028 46734 42030 46786
rect 42082 46734 42084 46786
rect 41468 46622 41470 46674
rect 41522 46622 41524 46674
rect 41468 46610 41524 46622
rect 41804 46676 41860 46686
rect 41804 46582 41860 46620
rect 41356 45890 41412 45948
rect 41916 46562 41972 46574
rect 41916 46510 41918 46562
rect 41970 46510 41972 46562
rect 41356 45838 41358 45890
rect 41410 45838 41412 45890
rect 41356 45826 41412 45838
rect 41468 45890 41524 45902
rect 41468 45838 41470 45890
rect 41522 45838 41524 45890
rect 41468 45444 41524 45838
rect 41916 45890 41972 46510
rect 42028 46564 42084 46734
rect 42028 46498 42084 46508
rect 41916 45838 41918 45890
rect 41970 45838 41972 45890
rect 41916 45826 41972 45838
rect 42140 45890 42196 46844
rect 42140 45838 42142 45890
rect 42194 45838 42196 45890
rect 41468 45378 41524 45388
rect 41692 45666 41748 45678
rect 41692 45614 41694 45666
rect 41746 45614 41748 45666
rect 41692 45108 41748 45614
rect 41580 45106 41748 45108
rect 41580 45054 41694 45106
rect 41746 45054 41748 45106
rect 41580 45052 41748 45054
rect 41580 43708 41636 45052
rect 41692 45042 41748 45052
rect 42140 44322 42196 45838
rect 42140 44270 42142 44322
rect 42194 44270 42196 44322
rect 42140 44258 42196 44270
rect 42252 44994 42308 45006
rect 42252 44942 42254 44994
rect 42306 44942 42308 44994
rect 42252 44772 42308 44942
rect 39676 43484 40292 43540
rect 40572 43652 40628 43662
rect 39676 43314 39732 43484
rect 39676 43262 39678 43314
rect 39730 43262 39732 43314
rect 39676 42756 39732 43262
rect 39788 43316 39844 43326
rect 39788 43222 39844 43260
rect 40012 43314 40068 43326
rect 40012 43262 40014 43314
rect 40066 43262 40068 43314
rect 40012 43204 40068 43262
rect 40124 43316 40180 43326
rect 40572 43316 40628 43596
rect 40124 43314 40292 43316
rect 40124 43262 40126 43314
rect 40178 43262 40292 43314
rect 40124 43260 40292 43262
rect 40124 43250 40180 43260
rect 40012 43138 40068 43148
rect 39788 42756 39844 42766
rect 39676 42754 39844 42756
rect 39676 42702 39790 42754
rect 39842 42702 39844 42754
rect 39676 42700 39844 42702
rect 39788 42690 39844 42700
rect 39788 42308 39844 42318
rect 39844 42252 39956 42308
rect 39788 42242 39844 42252
rect 39564 41878 39620 41916
rect 39228 41186 39284 41244
rect 39228 41134 39230 41186
rect 39282 41134 39284 41186
rect 39228 41122 39284 41134
rect 39340 41076 39396 41086
rect 39340 40982 39396 41020
rect 38892 40350 38894 40402
rect 38946 40350 38948 40402
rect 38892 40338 38948 40350
rect 39676 40292 39732 40302
rect 39676 40290 39844 40292
rect 39676 40238 39678 40290
rect 39730 40238 39844 40290
rect 39676 40236 39844 40238
rect 39676 40226 39732 40236
rect 39788 39842 39844 40236
rect 39788 39790 39790 39842
rect 39842 39790 39844 39842
rect 39788 39778 39844 39790
rect 39452 39732 39508 39742
rect 39452 39618 39508 39676
rect 39452 39566 39454 39618
rect 39506 39566 39508 39618
rect 39452 39554 39508 39566
rect 39900 39506 39956 42252
rect 40124 42196 40180 42206
rect 40124 42102 40180 42140
rect 40124 41972 40180 41982
rect 40124 39842 40180 41916
rect 40236 41970 40292 43260
rect 40572 42866 40628 43260
rect 40572 42814 40574 42866
rect 40626 42814 40628 42866
rect 40572 42802 40628 42814
rect 40908 43314 40964 43326
rect 40908 43262 40910 43314
rect 40962 43262 40964 43314
rect 40908 42084 40964 43262
rect 41020 43204 41076 43708
rect 41132 43652 41300 43708
rect 41468 43652 41636 43708
rect 41692 43764 41748 43802
rect 41692 43698 41748 43708
rect 42252 43652 42308 44716
rect 42476 43708 42532 50764
rect 42924 50370 42980 50382
rect 42924 50318 42926 50370
rect 42978 50318 42980 50370
rect 42588 50036 42644 50046
rect 42588 49942 42644 49980
rect 42924 49252 42980 50318
rect 43036 49810 43092 50764
rect 43148 50594 43204 51324
rect 43484 51286 43540 51324
rect 43484 50820 43540 50830
rect 43596 50820 43652 52222
rect 43820 51604 43876 53004
rect 44268 52994 44324 53004
rect 43932 52722 43988 52734
rect 43932 52670 43934 52722
rect 43986 52670 43988 52722
rect 43932 52052 43988 52670
rect 43932 51986 43988 51996
rect 43540 50764 43652 50820
rect 43708 51492 43764 51502
rect 43820 51492 43876 51548
rect 43708 51490 43876 51492
rect 43708 51438 43710 51490
rect 43762 51438 43876 51490
rect 43708 51436 43876 51438
rect 44156 51492 44212 51502
rect 43484 50754 43540 50764
rect 43148 50542 43150 50594
rect 43202 50542 43204 50594
rect 43148 50530 43204 50542
rect 43596 50596 43652 50606
rect 43708 50596 43764 51436
rect 44156 51378 44212 51436
rect 44156 51326 44158 51378
rect 44210 51326 44212 51378
rect 44156 51314 44212 51326
rect 44156 51154 44212 51166
rect 44156 51102 44158 51154
rect 44210 51102 44212 51154
rect 43596 50594 43764 50596
rect 43596 50542 43598 50594
rect 43650 50542 43764 50594
rect 43596 50540 43764 50542
rect 43932 50594 43988 50606
rect 43932 50542 43934 50594
rect 43986 50542 43988 50594
rect 43596 50530 43652 50540
rect 43820 50482 43876 50494
rect 43820 50430 43822 50482
rect 43874 50430 43876 50482
rect 43820 50148 43876 50430
rect 43820 50082 43876 50092
rect 43932 50036 43988 50542
rect 43036 49758 43038 49810
rect 43090 49758 43092 49810
rect 43036 49746 43092 49758
rect 43260 49812 43316 49822
rect 43260 49718 43316 49756
rect 42924 49196 43316 49252
rect 43260 48242 43316 49196
rect 43260 48190 43262 48242
rect 43314 48190 43316 48242
rect 43260 48178 43316 48190
rect 43708 48580 43764 48590
rect 43708 48466 43764 48524
rect 43708 48414 43710 48466
rect 43762 48414 43764 48466
rect 43148 47460 43204 47470
rect 42812 47346 42868 47358
rect 42812 47294 42814 47346
rect 42866 47294 42868 47346
rect 42700 46676 42756 46686
rect 42812 46676 42868 47294
rect 43148 46898 43204 47404
rect 43148 46846 43150 46898
rect 43202 46846 43204 46898
rect 43148 46834 43204 46846
rect 43484 47234 43540 47246
rect 43484 47182 43486 47234
rect 43538 47182 43540 47234
rect 42700 46674 42868 46676
rect 42700 46622 42702 46674
rect 42754 46622 42868 46674
rect 42700 46620 42868 46622
rect 42924 46676 42980 46686
rect 42700 45892 42756 46620
rect 42924 46228 42980 46620
rect 43260 46452 43316 46462
rect 43260 46358 43316 46396
rect 43484 46340 43540 47182
rect 43708 46562 43764 48414
rect 43820 47348 43876 47358
rect 43820 47254 43876 47292
rect 43932 47234 43988 49980
rect 44156 49810 44212 51102
rect 44380 50428 44436 53452
rect 44492 53172 44548 53182
rect 44828 53172 44884 53566
rect 47852 53620 47908 53630
rect 47908 53564 48132 53620
rect 47852 53526 47908 53564
rect 44548 53116 44884 53172
rect 44940 53506 44996 53518
rect 44940 53454 44942 53506
rect 44994 53454 44996 53506
rect 44492 52946 44548 53116
rect 44492 52894 44494 52946
rect 44546 52894 44548 52946
rect 44492 52882 44548 52894
rect 44940 52052 44996 53454
rect 45164 53506 45220 53518
rect 45164 53454 45166 53506
rect 45218 53454 45220 53506
rect 45164 52836 45220 53454
rect 46284 53172 46340 53182
rect 45724 53058 45780 53070
rect 45724 53006 45726 53058
rect 45778 53006 45780 53058
rect 45164 52834 45444 52836
rect 45164 52782 45166 52834
rect 45218 52782 45444 52834
rect 45164 52780 45444 52782
rect 45164 52770 45220 52780
rect 45388 52274 45444 52780
rect 45388 52222 45390 52274
rect 45442 52222 45444 52274
rect 45388 52210 45444 52222
rect 44828 51492 44884 51502
rect 44716 51380 44772 51390
rect 44604 51378 44772 51380
rect 44604 51326 44718 51378
rect 44770 51326 44772 51378
rect 44604 51324 44772 51326
rect 44380 50372 44548 50428
rect 44492 50306 44548 50316
rect 44492 50036 44548 50046
rect 44604 50036 44660 51324
rect 44716 51314 44772 51324
rect 44828 50596 44884 51436
rect 44940 51380 44996 51996
rect 45724 52162 45780 53006
rect 45724 52110 45726 52162
rect 45778 52110 45780 52162
rect 45500 51604 45556 51614
rect 45500 51490 45556 51548
rect 45500 51438 45502 51490
rect 45554 51438 45556 51490
rect 45500 51426 45556 51438
rect 45612 51492 45668 51502
rect 45612 51398 45668 51436
rect 45388 51380 45444 51390
rect 44940 51378 45444 51380
rect 44940 51326 45390 51378
rect 45442 51326 45444 51378
rect 44940 51324 45444 51326
rect 45388 51268 45444 51324
rect 45388 51202 45444 51212
rect 44940 50596 44996 50606
rect 44828 50594 44996 50596
rect 44828 50542 44942 50594
rect 44994 50542 44996 50594
rect 44828 50540 44996 50542
rect 44828 50428 44884 50540
rect 44940 50530 44996 50540
rect 44548 49980 44660 50036
rect 44716 50372 44884 50428
rect 45164 50482 45220 50494
rect 45164 50430 45166 50482
rect 45218 50430 45220 50482
rect 45164 50372 45220 50430
rect 45612 50484 45668 50522
rect 45724 50484 45780 52110
rect 46284 51378 46340 53116
rect 46956 52946 47012 52958
rect 46956 52894 46958 52946
rect 47010 52894 47012 52946
rect 46956 52162 47012 52894
rect 47628 52836 47684 52846
rect 46956 52110 46958 52162
rect 47010 52110 47012 52162
rect 46956 52052 47012 52110
rect 46956 51492 47012 51996
rect 46956 51398 47012 51436
rect 47404 52834 47684 52836
rect 47404 52782 47630 52834
rect 47682 52782 47684 52834
rect 47404 52780 47684 52782
rect 46284 51326 46286 51378
rect 46338 51326 46340 51378
rect 46284 51314 46340 51326
rect 46508 51380 46564 51390
rect 46508 51286 46564 51324
rect 46620 51378 46676 51390
rect 46620 51326 46622 51378
rect 46674 51326 46676 51378
rect 46620 51268 46676 51326
rect 47292 51268 47348 51278
rect 46620 51202 46676 51212
rect 47180 51266 47348 51268
rect 47180 51214 47294 51266
rect 47346 51214 47348 51266
rect 47180 51212 47348 51214
rect 46060 51154 46116 51166
rect 46060 51102 46062 51154
rect 46114 51102 46116 51154
rect 46060 50596 46116 51102
rect 47180 51156 47236 51212
rect 47292 51202 47348 51212
rect 47180 50820 47236 51100
rect 47404 50820 47460 52780
rect 47628 52770 47684 52780
rect 48076 52162 48132 53564
rect 48076 52110 48078 52162
rect 48130 52110 48132 52162
rect 46844 50764 47236 50820
rect 47292 50764 47460 50820
rect 47628 52050 47684 52062
rect 47628 51998 47630 52050
rect 47682 51998 47684 52050
rect 46060 50530 46116 50540
rect 46620 50596 46676 50606
rect 45668 50428 45780 50484
rect 45612 50418 45668 50428
rect 44492 49970 44548 49980
rect 44156 49758 44158 49810
rect 44210 49758 44212 49810
rect 44156 49746 44212 49758
rect 44716 49810 44772 50372
rect 45164 50306 45220 50316
rect 44716 49758 44718 49810
rect 44770 49758 44772 49810
rect 44716 49746 44772 49758
rect 44940 50148 44996 50158
rect 44940 50034 44996 50092
rect 44940 49982 44942 50034
rect 44994 49982 44996 50034
rect 44044 49698 44100 49710
rect 44044 49646 44046 49698
rect 44098 49646 44100 49698
rect 44044 48916 44100 49646
rect 44044 48132 44100 48860
rect 44940 48804 44996 49982
rect 46620 49810 46676 50540
rect 46844 50428 46900 50764
rect 46620 49758 46622 49810
rect 46674 49758 46676 49810
rect 46620 49746 46676 49758
rect 46732 50372 46900 50428
rect 46956 50484 47012 50494
rect 46732 49810 46788 50372
rect 46732 49758 46734 49810
rect 46786 49758 46788 49810
rect 46732 49746 46788 49758
rect 46956 49810 47012 50428
rect 46956 49758 46958 49810
rect 47010 49758 47012 49810
rect 46956 49746 47012 49758
rect 47068 49586 47124 49598
rect 47068 49534 47070 49586
rect 47122 49534 47124 49586
rect 47068 49252 47124 49534
rect 46732 49196 47124 49252
rect 46732 49026 46788 49196
rect 46732 48974 46734 49026
rect 46786 48974 46788 49026
rect 46732 48962 46788 48974
rect 47292 49026 47348 50764
rect 47628 50594 47684 51998
rect 47852 51380 47908 51390
rect 47852 51286 47908 51324
rect 48076 51044 48132 52110
rect 48188 53396 48244 53406
rect 48188 52276 48244 53340
rect 49084 53058 49140 53070
rect 49084 53006 49086 53058
rect 49138 53006 49140 53058
rect 48188 52050 48244 52220
rect 48860 52946 48916 52958
rect 48860 52894 48862 52946
rect 48914 52894 48916 52946
rect 48412 52164 48468 52174
rect 48412 52070 48468 52108
rect 48860 52162 48916 52894
rect 49084 52388 49140 53006
rect 49084 52322 49140 52332
rect 49196 52946 49252 52958
rect 49196 52894 49198 52946
rect 49250 52894 49252 52946
rect 48860 52110 48862 52162
rect 48914 52110 48916 52162
rect 48860 52098 48916 52110
rect 48188 51998 48190 52050
rect 48242 51998 48244 52050
rect 48188 51986 48244 51998
rect 48636 52052 48692 52062
rect 48636 51958 48692 51996
rect 49196 52052 49252 52894
rect 49644 52834 49700 52846
rect 49644 52782 49646 52834
rect 49698 52782 49700 52834
rect 49644 52388 49700 52782
rect 49644 52322 49700 52332
rect 50316 52276 50372 56142
rect 51212 55468 51268 56254
rect 50988 55412 51268 55468
rect 51548 56194 51604 56206
rect 51548 56142 51550 56194
rect 51602 56142 51604 56194
rect 50988 55410 51044 55412
rect 50988 55358 50990 55410
rect 51042 55358 51044 55410
rect 50988 55346 51044 55358
rect 50556 54908 50820 54918
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50556 54842 50820 54852
rect 50556 53340 50820 53350
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50556 53274 50820 53284
rect 49308 52164 49364 52174
rect 49308 52070 49364 52108
rect 50204 52164 50260 52174
rect 50316 52164 50372 52220
rect 50876 52388 50932 52398
rect 50932 52332 51156 52388
rect 50876 52274 50932 52332
rect 50876 52222 50878 52274
rect 50930 52222 50932 52274
rect 50876 52210 50932 52222
rect 50204 52162 50372 52164
rect 50204 52110 50206 52162
rect 50258 52110 50372 52162
rect 50204 52108 50372 52110
rect 50988 52164 51044 52174
rect 50204 52098 50260 52108
rect 48748 51380 48804 51390
rect 48748 51286 48804 51324
rect 49084 51378 49140 51390
rect 49084 51326 49086 51378
rect 49138 51326 49140 51378
rect 48076 50978 48132 50988
rect 48972 51266 49028 51278
rect 48972 51214 48974 51266
rect 49026 51214 49028 51266
rect 47628 50542 47630 50594
rect 47682 50542 47684 50594
rect 47628 50530 47684 50542
rect 47852 50706 47908 50718
rect 47852 50654 47854 50706
rect 47906 50654 47908 50706
rect 47404 50372 47460 50382
rect 47404 50034 47460 50316
rect 47404 49982 47406 50034
rect 47458 49982 47460 50034
rect 47404 49970 47460 49982
rect 47292 48974 47294 49026
rect 47346 48974 47348 49026
rect 46844 48916 46900 48926
rect 46900 48860 47012 48916
rect 46844 48822 46900 48860
rect 44940 48738 44996 48748
rect 45276 48692 45332 48702
rect 44492 48356 44548 48366
rect 44044 48066 44100 48076
rect 44156 48354 44548 48356
rect 44156 48302 44494 48354
rect 44546 48302 44548 48354
rect 44156 48300 44548 48302
rect 43932 47182 43934 47234
rect 43986 47182 43988 47234
rect 43932 46900 43988 47182
rect 43932 46834 43988 46844
rect 44156 47458 44212 48300
rect 44492 48290 44548 48300
rect 44268 48132 44324 48142
rect 44268 48038 44324 48076
rect 44156 47406 44158 47458
rect 44210 47406 44212 47458
rect 44156 46786 44212 47406
rect 44156 46734 44158 46786
rect 44210 46734 44212 46786
rect 44156 46722 44212 46734
rect 45276 46674 45332 48636
rect 46172 48692 46228 48702
rect 46060 48468 46116 48478
rect 45276 46622 45278 46674
rect 45330 46622 45332 46674
rect 45276 46610 45332 46622
rect 45388 48466 46116 48468
rect 45388 48414 46062 48466
rect 46114 48414 46116 48466
rect 45388 48412 46116 48414
rect 43708 46510 43710 46562
rect 43762 46510 43764 46562
rect 43708 46498 43764 46510
rect 45052 46452 45108 46462
rect 43484 46284 43876 46340
rect 42924 46172 43652 46228
rect 43484 45892 43540 45902
rect 42700 45890 43540 45892
rect 42700 45838 43486 45890
rect 43538 45838 43540 45890
rect 42700 45836 43540 45838
rect 43484 45826 43540 45836
rect 43596 45778 43652 46172
rect 43596 45726 43598 45778
rect 43650 45726 43652 45778
rect 43036 45666 43092 45678
rect 43036 45614 43038 45666
rect 43090 45614 43092 45666
rect 43036 45108 43092 45614
rect 43596 45668 43652 45726
rect 43596 45602 43652 45612
rect 43820 45890 43876 46284
rect 43820 45838 43822 45890
rect 43874 45838 43876 45890
rect 42924 44210 42980 44222
rect 42924 44158 42926 44210
rect 42978 44158 42980 44210
rect 42924 43708 42980 44158
rect 41132 43650 41188 43652
rect 41132 43598 41134 43650
rect 41186 43598 41188 43650
rect 41132 43314 41188 43598
rect 41468 43650 41524 43652
rect 41468 43598 41470 43650
rect 41522 43598 41524 43650
rect 41468 43586 41524 43598
rect 42252 43586 42308 43596
rect 42364 43652 42532 43708
rect 41804 43428 41860 43438
rect 42252 43428 42308 43438
rect 41132 43262 41134 43314
rect 41186 43262 41188 43314
rect 41132 43250 41188 43262
rect 41692 43426 42308 43428
rect 41692 43374 41806 43426
rect 41858 43374 42254 43426
rect 42306 43374 42308 43426
rect 41692 43372 42308 43374
rect 41020 42756 41076 43148
rect 41356 42756 41412 42766
rect 41020 42754 41412 42756
rect 41020 42702 41358 42754
rect 41410 42702 41412 42754
rect 41020 42700 41412 42702
rect 41356 42690 41412 42700
rect 41468 42196 41524 42206
rect 40236 41918 40238 41970
rect 40290 41918 40292 41970
rect 40236 41906 40292 41918
rect 40572 42082 40964 42084
rect 40572 42030 40910 42082
rect 40962 42030 40964 42082
rect 40572 42028 40964 42030
rect 40124 39790 40126 39842
rect 40178 39790 40180 39842
rect 40124 39778 40180 39790
rect 40348 40292 40404 40302
rect 39900 39454 39902 39506
rect 39954 39454 39956 39506
rect 39900 39442 39956 39454
rect 39116 39394 39172 39406
rect 39116 39342 39118 39394
rect 39170 39342 39172 39394
rect 39116 39284 39172 39342
rect 39116 39218 39172 39228
rect 38780 38098 38836 38108
rect 40348 38836 40404 40236
rect 40572 39732 40628 42028
rect 40908 42018 40964 42028
rect 41020 42084 41076 42094
rect 41020 42082 41188 42084
rect 41020 42030 41022 42082
rect 41074 42030 41188 42082
rect 41020 42028 41188 42030
rect 41020 42018 41076 42028
rect 41020 41746 41076 41758
rect 41020 41694 41022 41746
rect 41074 41694 41076 41746
rect 41020 41074 41076 41694
rect 41020 41022 41022 41074
rect 41074 41022 41076 41074
rect 41020 41010 41076 41022
rect 40908 40628 40964 40638
rect 40908 40534 40964 40572
rect 40572 39638 40628 39676
rect 40684 40516 40740 40526
rect 40348 38162 40404 38780
rect 40348 38110 40350 38162
rect 40402 38110 40404 38162
rect 40348 38098 40404 38110
rect 40236 38052 40292 38062
rect 39788 37828 39844 37838
rect 38556 37378 39172 37380
rect 38556 37326 38558 37378
rect 38610 37326 39172 37378
rect 38556 37324 39172 37326
rect 38556 37286 38612 37324
rect 38108 37266 38164 37278
rect 38108 37214 38110 37266
rect 38162 37214 38164 37266
rect 38108 36706 38164 37214
rect 38220 37268 38276 37278
rect 38220 37044 38276 37212
rect 38332 37266 38388 37278
rect 38332 37214 38334 37266
rect 38386 37214 38388 37266
rect 38332 37156 38388 37214
rect 39116 37266 39172 37324
rect 39116 37214 39118 37266
rect 39170 37214 39172 37266
rect 39116 37202 39172 37214
rect 38332 37090 38388 37100
rect 38444 37154 38500 37166
rect 38892 37156 38948 37166
rect 38444 37102 38446 37154
rect 38498 37102 38500 37154
rect 38444 37044 38500 37102
rect 38556 37100 38836 37156
rect 38556 37044 38612 37100
rect 38444 36988 38612 37044
rect 38220 36978 38276 36988
rect 38108 36654 38110 36706
rect 38162 36654 38164 36706
rect 38108 36642 38164 36654
rect 38220 36484 38276 36494
rect 38220 36390 38276 36428
rect 38108 36260 38164 36270
rect 38108 36166 38164 36204
rect 38668 36260 38724 36270
rect 38668 36166 38724 36204
rect 38780 36036 38836 37100
rect 38892 37062 38948 37100
rect 39788 37154 39844 37772
rect 40236 37492 40292 37996
rect 40348 37492 40404 37502
rect 40236 37490 40404 37492
rect 40236 37438 40350 37490
rect 40402 37438 40404 37490
rect 40236 37436 40404 37438
rect 40348 37426 40404 37436
rect 40460 37492 40516 37502
rect 39788 37102 39790 37154
rect 39842 37102 39844 37154
rect 39452 37042 39508 37054
rect 39452 36990 39454 37042
rect 39506 36990 39508 37042
rect 39452 36484 39508 36990
rect 39452 36418 39508 36428
rect 38780 35980 38948 36036
rect 37996 35858 38052 35868
rect 38332 35924 38388 35934
rect 37884 35812 37940 35822
rect 37884 35140 37940 35756
rect 38220 35812 38276 35822
rect 38220 35718 38276 35756
rect 38108 35698 38164 35710
rect 38108 35646 38110 35698
rect 38162 35646 38164 35698
rect 37996 35140 38052 35150
rect 37884 35138 38052 35140
rect 37884 35086 37998 35138
rect 38050 35086 38052 35138
rect 37884 35084 38052 35086
rect 37996 35074 38052 35084
rect 38108 35140 38164 35646
rect 38332 35700 38388 35868
rect 38780 35812 38836 35822
rect 38444 35700 38500 35710
rect 38332 35698 38500 35700
rect 38332 35646 38446 35698
rect 38498 35646 38500 35698
rect 38332 35644 38500 35646
rect 38444 35634 38500 35644
rect 38556 35700 38612 35710
rect 38220 35588 38276 35598
rect 38220 35494 38276 35532
rect 38108 35074 38164 35084
rect 37772 34962 37828 34972
rect 38444 35028 38500 35038
rect 38220 34914 38276 34926
rect 38220 34862 38222 34914
rect 38274 34862 38276 34914
rect 37548 34302 37550 34354
rect 37602 34302 37604 34354
rect 37548 34290 37604 34302
rect 37660 34690 37716 34702
rect 37660 34638 37662 34690
rect 37714 34638 37716 34690
rect 37660 34244 37716 34638
rect 37660 34178 37716 34188
rect 38220 34244 38276 34862
rect 38220 34178 38276 34188
rect 37212 33618 37268 33628
rect 37996 33684 38052 33694
rect 37100 33572 37156 33582
rect 37100 33458 37156 33516
rect 37100 33406 37102 33458
rect 37154 33406 37156 33458
rect 37100 33394 37156 33406
rect 37884 33348 37940 33358
rect 37548 33346 37940 33348
rect 37548 33294 37886 33346
rect 37938 33294 37940 33346
rect 37548 33292 37940 33294
rect 37324 33234 37380 33246
rect 37324 33182 37326 33234
rect 37378 33182 37380 33234
rect 37100 33124 37156 33134
rect 37100 33122 37268 33124
rect 37100 33070 37102 33122
rect 37154 33070 37268 33122
rect 37100 33068 37268 33070
rect 37100 33058 37156 33068
rect 37100 31780 37156 31790
rect 37100 31686 37156 31724
rect 36988 31500 37156 31556
rect 36988 30996 37044 31006
rect 36540 30482 36596 30492
rect 36652 30770 36708 30782
rect 36652 30718 36654 30770
rect 36706 30718 36708 30770
rect 36316 30212 36372 30222
rect 36316 30118 36372 30156
rect 36652 30100 36708 30718
rect 36204 29932 36372 29988
rect 35756 29474 35812 29484
rect 35980 29538 36036 29550
rect 35980 29486 35982 29538
rect 36034 29486 36036 29538
rect 35980 29316 36036 29486
rect 36204 29428 36260 29438
rect 36204 29334 36260 29372
rect 35980 29250 36036 29260
rect 35196 27970 35252 28700
rect 35532 28700 35700 28756
rect 35980 28868 36036 28878
rect 35308 28642 35364 28654
rect 35308 28590 35310 28642
rect 35362 28590 35364 28642
rect 35308 28084 35364 28590
rect 35308 28018 35364 28028
rect 35420 28308 35476 28318
rect 35420 28082 35476 28252
rect 35420 28030 35422 28082
rect 35474 28030 35476 28082
rect 35420 28018 35476 28030
rect 35196 27918 35198 27970
rect 35250 27918 35252 27970
rect 35196 27748 35252 27918
rect 35196 27682 35252 27692
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 34972 27356 35140 27412
rect 35196 27402 35460 27412
rect 34860 27020 35028 27076
rect 34524 26292 34580 26302
rect 34524 26178 34580 26236
rect 34972 26290 35028 27020
rect 34972 26238 34974 26290
rect 35026 26238 35028 26290
rect 34972 26226 35028 26238
rect 34524 26126 34526 26178
rect 34578 26126 34580 26178
rect 34524 25956 34580 26126
rect 34524 25890 34580 25900
rect 35084 25732 35140 27356
rect 35196 27188 35252 27198
rect 35196 26962 35252 27132
rect 35196 26910 35198 26962
rect 35250 26910 35252 26962
rect 35196 26898 35252 26910
rect 35308 27074 35364 27086
rect 35308 27022 35310 27074
rect 35362 27022 35364 27074
rect 35308 26740 35364 27022
rect 35196 26684 35364 26740
rect 35196 26068 35252 26684
rect 35196 26002 35252 26012
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 34972 25676 35140 25732
rect 34300 24834 34356 24892
rect 34300 24782 34302 24834
rect 34354 24782 34356 24834
rect 34300 24770 34356 24782
rect 34524 25620 34580 25630
rect 34412 24722 34468 24734
rect 34412 24670 34414 24722
rect 34466 24670 34468 24722
rect 34188 24612 34244 24622
rect 34188 23156 34244 24556
rect 34412 24276 34468 24670
rect 34412 24210 34468 24220
rect 34524 23940 34580 25564
rect 34860 25060 34916 25070
rect 34636 24948 34692 24958
rect 34636 24834 34692 24892
rect 34636 24782 34638 24834
rect 34690 24782 34692 24834
rect 34636 24770 34692 24782
rect 34860 24722 34916 25004
rect 34860 24670 34862 24722
rect 34914 24670 34916 24722
rect 34748 24610 34804 24622
rect 34748 24558 34750 24610
rect 34802 24558 34804 24610
rect 34748 24500 34804 24558
rect 34748 24434 34804 24444
rect 34860 24164 34916 24670
rect 34972 24724 35028 25676
rect 35084 25506 35140 25518
rect 35532 25508 35588 28700
rect 35980 28642 36036 28812
rect 35980 28590 35982 28642
rect 36034 28590 36036 28642
rect 35980 28578 36036 28590
rect 35756 28420 35812 28430
rect 35084 25454 35086 25506
rect 35138 25454 35140 25506
rect 35084 25172 35140 25454
rect 35420 25452 35588 25508
rect 35644 28418 35812 28420
rect 35644 28366 35758 28418
rect 35810 28366 35812 28418
rect 35644 28364 35812 28366
rect 35196 25396 35252 25406
rect 35196 25302 35252 25340
rect 35084 25106 35140 25116
rect 35420 24948 35476 25452
rect 35644 24948 35700 28364
rect 35756 28354 35812 28364
rect 35868 28420 35924 28430
rect 35868 28326 35924 28364
rect 36092 28308 36148 28318
rect 35980 28196 36036 28206
rect 35868 28084 35924 28094
rect 35868 27970 35924 28028
rect 35868 27918 35870 27970
rect 35922 27918 35924 27970
rect 35868 27906 35924 27918
rect 35980 27858 36036 28140
rect 35980 27806 35982 27858
rect 36034 27806 36036 27858
rect 35980 27074 36036 27806
rect 35980 27022 35982 27074
rect 36034 27022 36036 27074
rect 35756 26516 35812 26526
rect 35756 25618 35812 26460
rect 35756 25566 35758 25618
rect 35810 25566 35812 25618
rect 35756 25554 35812 25566
rect 35980 25506 36036 27022
rect 36092 26962 36148 28252
rect 36092 26910 36094 26962
rect 36146 26910 36148 26962
rect 36092 26898 36148 26910
rect 36316 26964 36372 29932
rect 36652 29428 36708 30044
rect 36988 29986 37044 30940
rect 36988 29934 36990 29986
rect 37042 29934 37044 29986
rect 36988 29540 37044 29934
rect 36876 29484 37044 29540
rect 36652 29362 36708 29372
rect 36764 29426 36820 29438
rect 36764 29374 36766 29426
rect 36818 29374 36820 29426
rect 36428 29204 36484 29214
rect 36428 28754 36484 29148
rect 36428 28702 36430 28754
rect 36482 28702 36484 28754
rect 36428 28690 36484 28702
rect 36652 28084 36708 28094
rect 36764 28084 36820 29374
rect 36876 28420 36932 29484
rect 37100 29426 37156 31500
rect 37212 30548 37268 33068
rect 37324 32900 37380 33182
rect 37324 32834 37380 32844
rect 37548 31218 37604 33292
rect 37884 33282 37940 33292
rect 37996 33124 38052 33628
rect 38332 33236 38388 33246
rect 38332 33142 38388 33180
rect 37884 33068 38052 33124
rect 38220 33122 38276 33134
rect 38220 33070 38222 33122
rect 38274 33070 38276 33122
rect 37548 31166 37550 31218
rect 37602 31166 37604 31218
rect 37548 31154 37604 31166
rect 37772 31666 37828 31678
rect 37772 31614 37774 31666
rect 37826 31614 37828 31666
rect 37772 31220 37828 31614
rect 37772 31154 37828 31164
rect 37324 30996 37380 31006
rect 37324 30902 37380 30940
rect 37660 30772 37716 30782
rect 37660 30678 37716 30716
rect 37212 30492 37828 30548
rect 37212 30436 37268 30492
rect 37212 30210 37268 30380
rect 37212 30158 37214 30210
rect 37266 30158 37268 30210
rect 37212 30146 37268 30158
rect 37436 30324 37492 30334
rect 37436 29764 37492 30268
rect 37100 29374 37102 29426
rect 37154 29374 37156 29426
rect 37100 29362 37156 29374
rect 37212 29708 37492 29764
rect 37660 30322 37716 30334
rect 37660 30270 37662 30322
rect 37714 30270 37716 30322
rect 36988 29316 37044 29326
rect 36988 28642 37044 29260
rect 36988 28590 36990 28642
rect 37042 28590 37044 28642
rect 36988 28578 37044 28590
rect 37212 28532 37268 29708
rect 37324 29540 37380 29550
rect 37324 29446 37380 29484
rect 37548 29540 37604 29550
rect 37660 29540 37716 30270
rect 37772 30098 37828 30492
rect 37772 30046 37774 30098
rect 37826 30046 37828 30098
rect 37772 30034 37828 30046
rect 37884 29876 37940 33068
rect 38220 30994 38276 33070
rect 38332 32452 38388 32462
rect 38444 32452 38500 34972
rect 38556 34244 38612 35644
rect 38780 35026 38836 35756
rect 38780 34974 38782 35026
rect 38834 34974 38836 35026
rect 38780 34962 38836 34974
rect 38556 34178 38612 34188
rect 38556 33348 38612 33358
rect 38556 33254 38612 33292
rect 38892 32788 38948 35980
rect 39676 35924 39732 35934
rect 39676 35830 39732 35868
rect 39788 35700 39844 37102
rect 40012 37044 40068 37054
rect 39900 36596 39956 36606
rect 40012 36596 40068 36988
rect 39900 36594 40012 36596
rect 39900 36542 39902 36594
rect 39954 36542 40012 36594
rect 39900 36540 40012 36542
rect 39900 36530 39956 36540
rect 40012 36530 40068 36540
rect 40460 36594 40516 37436
rect 40572 37044 40628 37054
rect 40572 36706 40628 36988
rect 40572 36654 40574 36706
rect 40626 36654 40628 36706
rect 40572 36642 40628 36654
rect 40460 36542 40462 36594
rect 40514 36542 40516 36594
rect 40460 36530 40516 36542
rect 40236 36484 40292 36494
rect 40236 36390 40292 36428
rect 40012 35924 40068 35934
rect 40012 35830 40068 35868
rect 40684 35924 40740 40460
rect 41132 40404 41188 42028
rect 41468 41186 41524 42140
rect 41692 41858 41748 43372
rect 41804 43362 41860 43372
rect 42252 43362 42308 43372
rect 42364 42980 42420 43652
rect 41692 41806 41694 41858
rect 41746 41806 41748 41858
rect 41692 41794 41748 41806
rect 42028 42924 42420 42980
rect 42588 43650 42644 43662
rect 42588 43598 42590 43650
rect 42642 43598 42644 43650
rect 42588 43316 42644 43598
rect 41468 41134 41470 41186
rect 41522 41134 41524 41186
rect 41468 41122 41524 41134
rect 42028 40516 42084 42924
rect 42364 42754 42420 42766
rect 42364 42702 42366 42754
rect 42418 42702 42420 42754
rect 42364 42308 42420 42702
rect 42364 42242 42420 42252
rect 42140 42084 42196 42094
rect 42588 42084 42644 43260
rect 42140 42082 42644 42084
rect 42140 42030 42142 42082
rect 42194 42030 42644 42082
rect 42140 42028 42644 42030
rect 42700 43652 42980 43708
rect 43036 43764 43092 45052
rect 43036 43698 43092 43708
rect 43372 45444 43428 45454
rect 43820 45444 43876 45838
rect 44940 45892 44996 45902
rect 44828 45780 44884 45790
rect 44828 45686 44884 45724
rect 44940 45444 44996 45836
rect 45052 45890 45108 46396
rect 45052 45838 45054 45890
rect 45106 45838 45108 45890
rect 45052 45826 45108 45838
rect 45388 45890 45444 48412
rect 46060 48402 46116 48412
rect 46172 48354 46228 48636
rect 46172 48302 46174 48354
rect 46226 48302 46228 48354
rect 46172 48290 46228 48302
rect 46844 48692 46900 48702
rect 46844 48242 46900 48636
rect 46956 48356 47012 48860
rect 47068 48802 47124 48814
rect 47068 48750 47070 48802
rect 47122 48750 47124 48802
rect 47068 48468 47124 48750
rect 47292 48692 47348 48974
rect 47292 48626 47348 48636
rect 47740 49922 47796 49934
rect 47740 49870 47742 49922
rect 47794 49870 47796 49922
rect 47068 48412 47572 48468
rect 46956 48300 47124 48356
rect 46844 48190 46846 48242
rect 46898 48190 46900 48242
rect 46844 48178 46900 48190
rect 47068 48242 47124 48300
rect 47068 48190 47070 48242
rect 47122 48190 47124 48242
rect 47068 48178 47124 48190
rect 47516 47570 47572 48412
rect 47740 48356 47796 49870
rect 47852 48580 47908 50654
rect 48636 50706 48692 50718
rect 48636 50654 48638 50706
rect 48690 50654 48692 50706
rect 48636 49028 48692 50654
rect 48748 50594 48804 50606
rect 48748 50542 48750 50594
rect 48802 50542 48804 50594
rect 48748 50484 48804 50542
rect 48748 50418 48804 50428
rect 48972 49698 49028 51214
rect 49084 51268 49140 51326
rect 49084 51202 49140 51212
rect 48972 49646 48974 49698
rect 49026 49646 49028 49698
rect 48972 49634 49028 49646
rect 49084 51044 49140 51054
rect 48636 48962 48692 48972
rect 49084 49138 49140 50988
rect 49084 49086 49086 49138
rect 49138 49086 49140 49138
rect 49084 48804 49140 49086
rect 49196 49028 49252 51996
rect 50428 51938 50484 51950
rect 50428 51886 50430 51938
rect 50482 51886 50484 51938
rect 50428 51380 50484 51886
rect 50556 51772 50820 51782
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50556 51706 50820 51716
rect 50988 51604 51044 52108
rect 50764 51548 51044 51604
rect 50428 51324 50708 51380
rect 49532 51268 49588 51278
rect 49532 51174 49588 51212
rect 49756 51156 49812 51166
rect 49756 51062 49812 51100
rect 49980 51154 50036 51166
rect 49980 51102 49982 51154
rect 50034 51102 50036 51154
rect 49532 50596 49588 50606
rect 49532 50502 49588 50540
rect 49980 50372 50036 51102
rect 50092 51156 50148 51166
rect 50092 50708 50148 51100
rect 50092 50614 50148 50652
rect 50428 51154 50484 51166
rect 50428 51102 50430 51154
rect 50482 51102 50484 51154
rect 49532 49922 49588 49934
rect 49532 49870 49534 49922
rect 49586 49870 49588 49922
rect 49532 49476 49588 49870
rect 49980 49812 50036 50316
rect 50428 50036 50484 51102
rect 50652 50372 50708 51324
rect 50764 51378 50820 51548
rect 51100 51492 51156 52332
rect 51548 52052 51604 56142
rect 51548 51604 51604 51996
rect 50764 51326 50766 51378
rect 50818 51326 50820 51378
rect 50764 51314 50820 51326
rect 50988 51436 51156 51492
rect 51324 51602 51604 51604
rect 51324 51550 51550 51602
rect 51602 51550 51604 51602
rect 51324 51548 51604 51550
rect 50988 51378 51044 51436
rect 50988 51326 50990 51378
rect 51042 51326 51044 51378
rect 50988 51314 51044 51326
rect 51324 51378 51380 51548
rect 51548 51538 51604 51548
rect 51884 51492 51940 51502
rect 51884 51398 51940 51436
rect 52668 51492 52724 51502
rect 51324 51326 51326 51378
rect 51378 51326 51380 51378
rect 51324 51314 51380 51326
rect 51100 51268 51156 51278
rect 51100 50596 51156 51212
rect 51884 50708 51940 50718
rect 51660 50596 51716 50606
rect 51100 50594 51716 50596
rect 51100 50542 51662 50594
rect 51714 50542 51716 50594
rect 51100 50540 51716 50542
rect 51660 50530 51716 50540
rect 51884 50594 51940 50652
rect 51884 50542 51886 50594
rect 51938 50542 51940 50594
rect 51884 50530 51940 50542
rect 52668 50482 52724 51436
rect 52668 50430 52670 50482
rect 52722 50430 52724 50482
rect 51436 50372 51492 50382
rect 50652 50316 50932 50372
rect 50556 50204 50820 50214
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50556 50138 50820 50148
rect 50428 49970 50484 49980
rect 50428 49812 50484 49822
rect 49980 49810 50484 49812
rect 49980 49758 50430 49810
rect 50482 49758 50484 49810
rect 49980 49756 50484 49758
rect 49532 49410 49588 49420
rect 50316 49476 50372 49486
rect 49532 49252 49588 49262
rect 49532 49158 49588 49196
rect 49420 49028 49476 49038
rect 49196 49026 49476 49028
rect 49196 48974 49422 49026
rect 49474 48974 49476 49026
rect 49196 48972 49476 48974
rect 49420 48962 49476 48972
rect 49532 48804 49588 48814
rect 49084 48802 49588 48804
rect 49084 48750 49534 48802
rect 49586 48750 49588 48802
rect 49084 48748 49588 48750
rect 50316 48804 50372 49420
rect 50428 49252 50484 49756
rect 50428 49186 50484 49196
rect 50428 49028 50484 49038
rect 50484 48972 50596 49028
rect 50428 48962 50484 48972
rect 50540 48914 50596 48972
rect 50540 48862 50542 48914
rect 50594 48862 50596 48914
rect 50540 48850 50596 48862
rect 50316 48748 50484 48804
rect 49532 48738 49588 48748
rect 47852 48514 47908 48524
rect 50428 48468 50484 48748
rect 50556 48636 50820 48646
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50556 48570 50820 48580
rect 50876 48580 50932 50316
rect 51436 50278 51492 50316
rect 51772 50370 51828 50382
rect 51772 50318 51774 50370
rect 51826 50318 51828 50370
rect 51772 49810 51828 50318
rect 52444 50372 52500 50382
rect 51772 49758 51774 49810
rect 51826 49758 51828 49810
rect 51772 49746 51828 49758
rect 52108 50036 52164 50046
rect 52108 49810 52164 49980
rect 52108 49758 52110 49810
rect 52162 49758 52164 49810
rect 52108 49746 52164 49758
rect 52332 49810 52388 49822
rect 52332 49758 52334 49810
rect 52386 49758 52388 49810
rect 51996 49698 52052 49710
rect 51996 49646 51998 49698
rect 52050 49646 52052 49698
rect 51212 49588 51268 49598
rect 50988 49586 51268 49588
rect 50988 49534 51214 49586
rect 51266 49534 51268 49586
rect 50988 49532 51268 49534
rect 50988 49026 51044 49532
rect 50988 48974 50990 49026
rect 51042 48974 51044 49026
rect 50988 48962 51044 48974
rect 51100 49028 51156 49038
rect 50876 48524 51044 48580
rect 50652 48468 50708 48478
rect 50428 48466 50708 48468
rect 50428 48414 50654 48466
rect 50706 48414 50708 48466
rect 50428 48412 50708 48414
rect 50652 48402 50708 48412
rect 50764 48468 50820 48478
rect 50764 48356 50820 48412
rect 50876 48356 50932 48366
rect 47740 48300 47908 48356
rect 50764 48354 50932 48356
rect 50764 48302 50878 48354
rect 50930 48302 50932 48354
rect 50764 48300 50932 48302
rect 47740 48132 47796 48142
rect 47516 47518 47518 47570
rect 47570 47518 47572 47570
rect 47516 47506 47572 47518
rect 47628 48130 47796 48132
rect 47628 48078 47742 48130
rect 47794 48078 47796 48130
rect 47628 48076 47796 48078
rect 45388 45838 45390 45890
rect 45442 45838 45444 45890
rect 43820 45388 44324 45444
rect 42700 42754 42756 43652
rect 42700 42702 42702 42754
rect 42754 42702 42756 42754
rect 42140 42018 42196 42028
rect 42700 41972 42756 42702
rect 43372 42082 43428 45388
rect 43708 45276 44212 45332
rect 43708 45106 43764 45276
rect 43708 45054 43710 45106
rect 43762 45054 43764 45106
rect 43708 45042 43764 45054
rect 43932 45106 43988 45118
rect 43932 45054 43934 45106
rect 43986 45054 43988 45106
rect 43820 44994 43876 45006
rect 43820 44942 43822 44994
rect 43874 44942 43876 44994
rect 43820 44436 43876 44942
rect 43932 44996 43988 45054
rect 43932 44930 43988 44940
rect 44044 44882 44100 44894
rect 44044 44830 44046 44882
rect 44098 44830 44100 44882
rect 43932 44436 43988 44446
rect 43820 44380 43932 44436
rect 43932 44370 43988 44380
rect 43708 44324 43764 44334
rect 43708 44322 43876 44324
rect 43708 44270 43710 44322
rect 43762 44270 43876 44322
rect 43708 44268 43876 44270
rect 43708 44258 43764 44268
rect 43820 43876 43876 44268
rect 43708 43820 43876 43876
rect 43932 44212 43988 44222
rect 43708 43652 43764 43820
rect 43596 42980 43652 42990
rect 43372 42030 43374 42082
rect 43426 42030 43428 42082
rect 43372 42018 43428 42030
rect 43484 42978 43652 42980
rect 43484 42926 43598 42978
rect 43650 42926 43652 42978
rect 43484 42924 43652 42926
rect 42700 41906 42756 41916
rect 43484 41972 43540 42924
rect 43596 42914 43652 42924
rect 43708 42868 43764 43596
rect 43932 43538 43988 44156
rect 43932 43486 43934 43538
rect 43986 43486 43988 43538
rect 43932 43474 43988 43486
rect 43708 42802 43764 42812
rect 43596 42756 43652 42766
rect 43596 42194 43652 42700
rect 43596 42142 43598 42194
rect 43650 42142 43652 42194
rect 43596 42130 43652 42142
rect 43484 41906 43540 41916
rect 44044 41970 44100 44830
rect 44156 44434 44212 45276
rect 44156 44382 44158 44434
rect 44210 44382 44212 44434
rect 44156 43316 44212 44382
rect 44156 43250 44212 43260
rect 44268 44210 44324 45388
rect 44828 45388 44996 45444
rect 45052 45666 45108 45678
rect 45052 45614 45054 45666
rect 45106 45614 45108 45666
rect 44268 44158 44270 44210
rect 44322 44158 44324 44210
rect 44268 42084 44324 44158
rect 44492 45106 44548 45118
rect 44492 45054 44494 45106
rect 44546 45054 44548 45106
rect 44492 44212 44548 45054
rect 44828 44884 44884 45388
rect 45052 45332 45108 45614
rect 45388 45444 45444 45838
rect 45388 45378 45444 45388
rect 45612 46898 45668 46910
rect 45612 46846 45614 46898
rect 45666 46846 45668 46898
rect 45052 45266 45108 45276
rect 45164 45220 45220 45230
rect 45164 45218 45332 45220
rect 45164 45166 45166 45218
rect 45218 45166 45332 45218
rect 45164 45164 45332 45166
rect 45164 45154 45220 45164
rect 44940 45108 44996 45118
rect 44940 45014 44996 45052
rect 45052 44994 45108 45006
rect 45052 44942 45054 44994
rect 45106 44942 45108 44994
rect 45052 44884 45108 44942
rect 44828 44828 45108 44884
rect 45276 44772 45332 45164
rect 44492 44146 44548 44156
rect 45052 44434 45108 44446
rect 45052 44382 45054 44434
rect 45106 44382 45108 44434
rect 45052 44212 45108 44382
rect 45164 44324 45220 44334
rect 45276 44324 45332 44716
rect 45164 44322 45332 44324
rect 45164 44270 45166 44322
rect 45218 44270 45332 44322
rect 45164 44268 45332 44270
rect 45500 45108 45556 45118
rect 45500 44322 45556 45052
rect 45500 44270 45502 44322
rect 45554 44270 45556 44322
rect 45164 44258 45220 44268
rect 45500 44258 45556 44270
rect 45052 44146 45108 44156
rect 45612 44212 45668 46846
rect 46060 46900 46116 46910
rect 46060 46806 46116 46844
rect 46396 46786 46452 46798
rect 46396 46734 46398 46786
rect 46450 46734 46452 46786
rect 46396 46004 46452 46734
rect 47628 46340 47684 48076
rect 47740 48066 47796 48076
rect 47852 46786 47908 48300
rect 50876 48290 50932 48300
rect 50988 48356 51044 48524
rect 50988 48262 51044 48300
rect 49308 47572 49364 47582
rect 49308 47460 49364 47516
rect 51100 47460 51156 48972
rect 51212 47572 51268 49532
rect 51996 49364 52052 49646
rect 52332 49476 52388 49758
rect 52332 49410 52388 49420
rect 51548 49308 52052 49364
rect 51548 49026 51604 49308
rect 51548 48974 51550 49026
rect 51602 48974 51604 49026
rect 51548 48962 51604 48974
rect 51436 48802 51492 48814
rect 51436 48750 51438 48802
rect 51490 48750 51492 48802
rect 51436 48468 51492 48750
rect 52444 48804 52500 50316
rect 52444 48738 52500 48748
rect 51436 48402 51492 48412
rect 51212 47478 51268 47516
rect 51324 48356 51380 48366
rect 48972 47458 49364 47460
rect 48972 47406 49310 47458
rect 49362 47406 49364 47458
rect 48972 47404 49364 47406
rect 48076 47346 48132 47358
rect 48076 47294 48078 47346
rect 48130 47294 48132 47346
rect 47964 47012 48020 47022
rect 47964 46898 48020 46956
rect 47964 46846 47966 46898
rect 48018 46846 48020 46898
rect 47964 46834 48020 46846
rect 47852 46734 47854 46786
rect 47906 46734 47908 46786
rect 47852 46564 47908 46734
rect 48076 46788 48132 47294
rect 48188 46788 48244 46798
rect 48076 46732 48188 46788
rect 48188 46694 48244 46732
rect 48972 46786 49028 47404
rect 49308 47394 49364 47404
rect 50876 47458 51156 47460
rect 50876 47406 51102 47458
rect 51154 47406 51156 47458
rect 50876 47404 51156 47406
rect 49980 47346 50036 47358
rect 49980 47294 49982 47346
rect 50034 47294 50036 47346
rect 49084 46900 49140 46910
rect 49084 46898 49700 46900
rect 49084 46846 49086 46898
rect 49138 46846 49700 46898
rect 49084 46844 49700 46846
rect 49084 46834 49140 46844
rect 48972 46734 48974 46786
rect 49026 46734 49028 46786
rect 48972 46722 49028 46734
rect 47852 46498 47908 46508
rect 46396 45938 46452 45948
rect 47404 46284 47796 46340
rect 47404 45890 47460 46284
rect 47404 45838 47406 45890
rect 47458 45838 47460 45890
rect 47404 45826 47460 45838
rect 47628 46004 47684 46014
rect 47628 45890 47684 45948
rect 47628 45838 47630 45890
rect 47682 45838 47684 45890
rect 46172 45780 46228 45790
rect 46172 45686 46228 45724
rect 47516 45780 47572 45790
rect 47516 45686 47572 45724
rect 45836 45668 45892 45678
rect 45836 45574 45892 45612
rect 46956 45666 47012 45678
rect 46956 45614 46958 45666
rect 47010 45614 47012 45666
rect 45836 45332 45892 45342
rect 45836 45238 45892 45276
rect 46732 45332 46788 45342
rect 46284 44996 46340 45006
rect 46284 44902 46340 44940
rect 46732 44546 46788 45276
rect 46732 44494 46734 44546
rect 46786 44494 46788 44546
rect 46732 44482 46788 44494
rect 46844 44996 46900 45006
rect 45612 44146 45668 44156
rect 46060 44436 46116 44446
rect 46060 44100 46116 44380
rect 46060 44098 46228 44100
rect 46060 44046 46062 44098
rect 46114 44046 46228 44098
rect 46060 44044 46228 44046
rect 46060 44034 46116 44044
rect 45052 43314 45108 43326
rect 45052 43262 45054 43314
rect 45106 43262 45108 43314
rect 44940 42754 44996 42766
rect 44940 42702 44942 42754
rect 44994 42702 44996 42754
rect 44940 42196 44996 42702
rect 44940 42130 44996 42140
rect 44268 42018 44324 42028
rect 44044 41918 44046 41970
rect 44098 41918 44100 41970
rect 44044 41906 44100 41918
rect 44940 41972 44996 41982
rect 45052 41972 45108 43262
rect 46172 42866 46228 44044
rect 46732 43652 46788 43662
rect 46732 43558 46788 43596
rect 46172 42814 46174 42866
rect 46226 42814 46228 42866
rect 46172 42802 46228 42814
rect 46396 43316 46452 43326
rect 45388 42756 45444 42766
rect 45388 42662 45444 42700
rect 46396 42754 46452 43260
rect 46396 42702 46398 42754
rect 46450 42702 46452 42754
rect 46396 42690 46452 42702
rect 46508 42978 46564 42990
rect 46508 42926 46510 42978
rect 46562 42926 46564 42978
rect 45500 42084 45556 42094
rect 44940 41970 45108 41972
rect 44940 41918 44942 41970
rect 44994 41918 45108 41970
rect 44940 41916 45108 41918
rect 45388 41972 45444 41982
rect 44044 41412 44100 41422
rect 44044 41410 44436 41412
rect 44044 41358 44046 41410
rect 44098 41358 44436 41410
rect 44044 41356 44436 41358
rect 44044 41346 44100 41356
rect 42588 41188 42644 41198
rect 42588 41094 42644 41132
rect 43484 41074 43540 41086
rect 43484 41022 43486 41074
rect 43538 41022 43540 41074
rect 43260 40740 43316 40750
rect 42028 40450 42084 40460
rect 42476 40516 42532 40526
rect 42476 40422 42532 40460
rect 43036 40514 43092 40526
rect 43036 40462 43038 40514
rect 43090 40462 43092 40514
rect 41468 40404 41524 40414
rect 41132 40348 41468 40404
rect 41468 40310 41524 40348
rect 43036 40404 43092 40462
rect 40908 39618 40964 39630
rect 40908 39566 40910 39618
rect 40962 39566 40964 39618
rect 40908 38052 40964 39566
rect 41804 39620 41860 39630
rect 42140 39620 42196 39630
rect 41244 38836 41300 38846
rect 41804 38836 41860 39564
rect 41916 39618 42196 39620
rect 41916 39566 42142 39618
rect 42194 39566 42196 39618
rect 41916 39564 42196 39566
rect 41916 38946 41972 39564
rect 42140 39554 42196 39564
rect 42812 39618 42868 39630
rect 42812 39566 42814 39618
rect 42866 39566 42868 39618
rect 41916 38894 41918 38946
rect 41970 38894 41972 38946
rect 41916 38882 41972 38894
rect 42700 39394 42756 39406
rect 42700 39342 42702 39394
rect 42754 39342 42756 39394
rect 41244 38742 41300 38780
rect 41580 38834 41860 38836
rect 41580 38782 41806 38834
rect 41858 38782 41860 38834
rect 41580 38780 41860 38782
rect 40908 37986 40964 37996
rect 41580 38050 41636 38780
rect 41804 38770 41860 38780
rect 42588 38722 42644 38734
rect 42588 38670 42590 38722
rect 42642 38670 42644 38722
rect 41580 37998 41582 38050
rect 41634 37998 41636 38050
rect 41580 37986 41636 37998
rect 41692 38274 41748 38286
rect 41692 38222 41694 38274
rect 41746 38222 41748 38274
rect 41692 37044 41748 38222
rect 41692 36594 41748 36988
rect 41692 36542 41694 36594
rect 41746 36542 41748 36594
rect 41692 36530 41748 36542
rect 42588 37266 42644 38670
rect 42588 37214 42590 37266
rect 42642 37214 42644 37266
rect 41356 36484 41412 36494
rect 41356 36390 41412 36428
rect 40684 35858 40740 35868
rect 40908 36370 40964 36382
rect 40908 36318 40910 36370
rect 40962 36318 40964 36370
rect 39676 35644 39844 35700
rect 39900 35700 39956 35710
rect 39116 35586 39172 35598
rect 39116 35534 39118 35586
rect 39170 35534 39172 35586
rect 39116 35140 39172 35534
rect 39116 35074 39172 35084
rect 39676 35252 39732 35644
rect 39452 35028 39508 35038
rect 39452 34934 39508 34972
rect 39676 34802 39732 35196
rect 39788 35140 39844 35150
rect 39900 35140 39956 35644
rect 39788 35138 39956 35140
rect 39788 35086 39790 35138
rect 39842 35086 39956 35138
rect 39788 35084 39956 35086
rect 39788 35074 39844 35084
rect 40012 35028 40068 35038
rect 39900 34972 40012 35028
rect 39676 34750 39678 34802
rect 39730 34750 39732 34802
rect 39676 34580 39732 34750
rect 39788 34804 39844 34814
rect 39900 34804 39956 34972
rect 40012 34962 40068 34972
rect 40348 35026 40404 35038
rect 40348 34974 40350 35026
rect 40402 34974 40404 35026
rect 39788 34802 39956 34804
rect 39788 34750 39790 34802
rect 39842 34750 39956 34802
rect 39788 34748 39956 34750
rect 39788 34738 39844 34748
rect 39676 34514 39732 34524
rect 40236 34690 40292 34702
rect 40236 34638 40238 34690
rect 40290 34638 40292 34690
rect 40236 34244 40292 34638
rect 40236 34178 40292 34188
rect 39900 34130 39956 34142
rect 39900 34078 39902 34130
rect 39954 34078 39956 34130
rect 39228 34020 39284 34030
rect 39228 33926 39284 33964
rect 39900 33572 39956 34078
rect 40124 34020 40180 34030
rect 40124 33926 40180 33964
rect 40124 33572 40180 33582
rect 39900 33516 40124 33572
rect 40124 33458 40180 33516
rect 40348 33570 40404 34974
rect 40796 34916 40852 34926
rect 40908 34916 40964 36318
rect 41132 35700 41188 35710
rect 41132 35606 41188 35644
rect 41804 35700 41860 35710
rect 41804 35606 41860 35644
rect 42588 35698 42644 37214
rect 42588 35646 42590 35698
rect 42642 35646 42644 35698
rect 40796 34914 40964 34916
rect 40796 34862 40798 34914
rect 40850 34862 40964 34914
rect 40796 34860 40964 34862
rect 40796 34850 40852 34860
rect 40348 33518 40350 33570
rect 40402 33518 40404 33570
rect 40348 33506 40404 33518
rect 40460 34690 40516 34702
rect 40460 34638 40462 34690
rect 40514 34638 40516 34690
rect 40124 33406 40126 33458
rect 40178 33406 40180 33458
rect 40124 33394 40180 33406
rect 40460 33236 40516 34638
rect 40908 34242 40964 34860
rect 41132 35028 41188 35038
rect 41132 34914 41188 34972
rect 41804 35028 41860 35038
rect 41804 34934 41860 34972
rect 42588 35026 42644 35646
rect 42588 34974 42590 35026
rect 42642 34974 42644 35026
rect 42588 34962 42644 34974
rect 42700 37154 42756 39342
rect 42812 37492 42868 39566
rect 42812 37426 42868 37436
rect 42700 37102 42702 37154
rect 42754 37102 42756 37154
rect 42700 35700 42756 37102
rect 41132 34862 41134 34914
rect 41186 34862 41188 34914
rect 41132 34850 41188 34862
rect 42700 34914 42756 35644
rect 43036 36482 43092 40348
rect 43260 40402 43316 40684
rect 43260 40350 43262 40402
rect 43314 40350 43316 40402
rect 43260 40338 43316 40350
rect 43372 40404 43428 40414
rect 43372 40310 43428 40348
rect 43484 39620 43540 41022
rect 44156 41074 44212 41086
rect 44156 41022 44158 41074
rect 44210 41022 44212 41074
rect 44044 40964 44100 40974
rect 43932 40962 44100 40964
rect 43932 40910 44046 40962
rect 44098 40910 44100 40962
rect 43932 40908 44100 40910
rect 43596 40404 43652 40414
rect 43932 40404 43988 40908
rect 44044 40898 44100 40908
rect 43652 40348 43988 40404
rect 44044 40516 44100 40526
rect 44156 40516 44212 41022
rect 44044 40514 44212 40516
rect 44044 40462 44046 40514
rect 44098 40462 44212 40514
rect 44044 40460 44212 40462
rect 43596 40310 43652 40348
rect 44044 39730 44100 40460
rect 44044 39678 44046 39730
rect 44098 39678 44100 39730
rect 44044 39666 44100 39678
rect 43596 39620 43652 39630
rect 43540 39618 43652 39620
rect 43540 39566 43598 39618
rect 43650 39566 43652 39618
rect 43540 39564 43652 39566
rect 43484 39526 43540 39564
rect 43596 39554 43652 39564
rect 43708 39506 43764 39518
rect 43708 39454 43710 39506
rect 43762 39454 43764 39506
rect 43708 39060 43764 39454
rect 43708 38994 43764 39004
rect 43484 38948 43540 38958
rect 43484 37266 43540 38892
rect 43596 38836 43652 38846
rect 44380 38836 44436 41356
rect 44940 41188 44996 41916
rect 44940 41094 44996 41132
rect 45388 41186 45444 41916
rect 45388 41134 45390 41186
rect 45442 41134 45444 41186
rect 45388 41122 45444 41134
rect 44828 41074 44884 41086
rect 44828 41022 44830 41074
rect 44882 41022 44884 41074
rect 44828 40740 44884 41022
rect 44828 40674 44884 40684
rect 45388 40402 45444 40414
rect 45388 40350 45390 40402
rect 45442 40350 45444 40402
rect 45164 40290 45220 40302
rect 45164 40238 45166 40290
rect 45218 40238 45220 40290
rect 44492 38948 44548 38958
rect 44492 38854 44548 38892
rect 43652 38780 43764 38836
rect 43596 38742 43652 38780
rect 43708 38274 43764 38780
rect 43708 38222 43710 38274
rect 43762 38222 43764 38274
rect 43708 38210 43764 38222
rect 43932 38834 44436 38836
rect 43932 38782 44382 38834
rect 44434 38782 44436 38834
rect 43932 38780 44436 38782
rect 43932 37938 43988 38780
rect 44380 38770 44436 38780
rect 45164 38668 45220 40238
rect 45388 39394 45444 40350
rect 45388 39342 45390 39394
rect 45442 39342 45444 39394
rect 45388 39330 45444 39342
rect 45500 38948 45556 42028
rect 46172 41860 46228 41870
rect 46172 41766 46228 41804
rect 45948 40292 46004 40302
rect 45948 39618 46004 40236
rect 46284 40292 46340 40302
rect 46284 40290 46452 40292
rect 46284 40238 46286 40290
rect 46338 40238 46452 40290
rect 46284 40236 46452 40238
rect 46284 40226 46340 40236
rect 45948 39566 45950 39618
rect 46002 39566 46004 39618
rect 45948 39554 46004 39566
rect 45612 39284 45668 39294
rect 45612 39058 45668 39228
rect 45612 39006 45614 39058
rect 45666 39006 45668 39058
rect 45612 38994 45668 39006
rect 45836 39060 45892 39070
rect 45836 38966 45892 39004
rect 44940 38612 45220 38668
rect 45388 38946 45556 38948
rect 45388 38894 45502 38946
rect 45554 38894 45556 38946
rect 45388 38892 45556 38894
rect 43932 37886 43934 37938
rect 43986 37886 43988 37938
rect 43932 37874 43988 37886
rect 44044 38162 44100 38174
rect 44044 38110 44046 38162
rect 44098 38110 44100 38162
rect 43484 37214 43486 37266
rect 43538 37214 43540 37266
rect 43484 36706 43540 37214
rect 44044 37268 44100 38110
rect 44940 38164 44996 38612
rect 44268 37268 44324 37278
rect 44044 37266 44324 37268
rect 44044 37214 44270 37266
rect 44322 37214 44324 37266
rect 44044 37212 44324 37214
rect 44268 37202 44324 37212
rect 44940 37266 44996 38108
rect 45388 38050 45444 38892
rect 45500 38882 45556 38892
rect 46284 38836 46340 38846
rect 46284 38742 46340 38780
rect 46396 38834 46452 40236
rect 46508 39620 46564 42926
rect 46844 42754 46900 44940
rect 46956 44212 47012 45614
rect 47068 44436 47124 44446
rect 47516 44436 47572 44446
rect 47068 44434 47572 44436
rect 47068 44382 47070 44434
rect 47122 44382 47518 44434
rect 47570 44382 47572 44434
rect 47068 44380 47572 44382
rect 47068 44370 47124 44380
rect 46956 44118 47012 44156
rect 46844 42702 46846 42754
rect 46898 42702 46900 42754
rect 46844 42690 46900 42702
rect 47292 43426 47348 43438
rect 47292 43374 47294 43426
rect 47346 43374 47348 43426
rect 47292 42532 47348 43374
rect 47404 42532 47460 42542
rect 47292 42476 47404 42532
rect 47404 42082 47460 42476
rect 47404 42030 47406 42082
rect 47458 42030 47460 42082
rect 47404 42018 47460 42030
rect 46956 41860 47012 41870
rect 46956 40402 47012 41804
rect 47404 41858 47460 41870
rect 47404 41806 47406 41858
rect 47458 41806 47460 41858
rect 47404 41636 47460 41806
rect 47404 41074 47460 41580
rect 47516 41186 47572 44380
rect 47628 43708 47684 45838
rect 47740 45218 47796 46284
rect 48188 46004 48244 46014
rect 47964 45780 48020 45790
rect 47964 45330 48020 45724
rect 47964 45278 47966 45330
rect 48018 45278 48020 45330
rect 47964 45266 48020 45278
rect 48188 45330 48244 45948
rect 48972 46002 49028 46014
rect 48972 45950 48974 46002
rect 49026 45950 49028 46002
rect 48748 45892 48804 45902
rect 48748 45798 48804 45836
rect 48860 45778 48916 45790
rect 48860 45726 48862 45778
rect 48914 45726 48916 45778
rect 48860 45556 48916 45726
rect 48188 45278 48190 45330
rect 48242 45278 48244 45330
rect 48188 45266 48244 45278
rect 48300 45500 48916 45556
rect 48300 45330 48356 45500
rect 48300 45278 48302 45330
rect 48354 45278 48356 45330
rect 48300 45266 48356 45278
rect 47740 45166 47742 45218
rect 47794 45166 47796 45218
rect 47740 45154 47796 45166
rect 47964 44210 48020 44222
rect 47964 44158 47966 44210
rect 48018 44158 48020 44210
rect 47628 43652 47796 43708
rect 47516 41134 47518 41186
rect 47570 41134 47572 41186
rect 47516 41122 47572 41134
rect 47628 41972 47684 41982
rect 47740 41972 47796 43652
rect 47628 41970 47796 41972
rect 47628 41918 47630 41970
rect 47682 41918 47796 41970
rect 47628 41916 47796 41918
rect 47404 41022 47406 41074
rect 47458 41022 47460 41074
rect 47404 41010 47460 41022
rect 47628 40626 47684 41916
rect 47964 41636 48020 44158
rect 48188 44212 48244 44222
rect 48188 42866 48244 44156
rect 48860 43314 48916 43326
rect 48860 43262 48862 43314
rect 48914 43262 48916 43314
rect 48860 42980 48916 43262
rect 48972 43314 49028 45950
rect 49644 45892 49700 46844
rect 49420 45890 49700 45892
rect 49420 45838 49646 45890
rect 49698 45838 49700 45890
rect 49420 45836 49700 45838
rect 49196 45106 49252 45118
rect 49196 45054 49198 45106
rect 49250 45054 49252 45106
rect 49084 44996 49140 45006
rect 49084 44902 49140 44940
rect 49196 44212 49252 45054
rect 49196 44146 49252 44156
rect 49420 44210 49476 45836
rect 49644 45826 49700 45836
rect 49980 45106 50036 47294
rect 50556 47068 50820 47078
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50556 47002 50820 47012
rect 50428 46788 50484 46798
rect 50428 46694 50484 46732
rect 49980 45054 49982 45106
rect 50034 45054 50036 45106
rect 49756 44996 49812 45006
rect 49420 44158 49422 44210
rect 49474 44158 49476 44210
rect 49420 44146 49476 44158
rect 49644 44210 49700 44222
rect 49644 44158 49646 44210
rect 49698 44158 49700 44210
rect 48972 43262 48974 43314
rect 49026 43262 49028 43314
rect 48972 43092 49028 43262
rect 49196 43316 49252 43326
rect 49196 43222 49252 43260
rect 49308 43316 49364 43326
rect 49308 43314 49476 43316
rect 49308 43262 49310 43314
rect 49362 43262 49476 43314
rect 49308 43260 49476 43262
rect 49308 43250 49364 43260
rect 48972 43036 49252 43092
rect 48860 42924 49140 42980
rect 48188 42814 48190 42866
rect 48242 42814 48244 42866
rect 48188 42802 48244 42814
rect 48972 42756 49028 42766
rect 48972 42644 49028 42700
rect 47964 41570 48020 41580
rect 48636 42642 49028 42644
rect 48636 42590 48974 42642
rect 49026 42590 49028 42642
rect 48636 42588 49028 42590
rect 48636 41186 48692 42588
rect 48972 42578 49028 42588
rect 49084 42420 49140 42924
rect 48972 42364 49140 42420
rect 48636 41134 48638 41186
rect 48690 41134 48692 41186
rect 48636 41122 48692 41134
rect 48860 41970 48916 41982
rect 48860 41918 48862 41970
rect 48914 41918 48916 41970
rect 48748 40962 48804 40974
rect 48748 40910 48750 40962
rect 48802 40910 48804 40962
rect 47628 40574 47630 40626
rect 47682 40574 47684 40626
rect 47628 40562 47684 40574
rect 48300 40628 48356 40638
rect 46956 40350 46958 40402
rect 47010 40350 47012 40402
rect 46956 40338 47012 40350
rect 48188 40402 48244 40414
rect 48188 40350 48190 40402
rect 48242 40350 48244 40402
rect 47180 40292 47236 40302
rect 47180 40198 47236 40236
rect 48188 39732 48244 40350
rect 48300 39844 48356 40572
rect 48748 40292 48804 40910
rect 48300 39842 48692 39844
rect 48300 39790 48302 39842
rect 48354 39790 48692 39842
rect 48300 39788 48692 39790
rect 48300 39778 48356 39788
rect 48188 39666 48244 39676
rect 46620 39620 46676 39630
rect 46508 39564 46620 39620
rect 46620 39526 46676 39564
rect 47852 39618 47908 39630
rect 48076 39620 48132 39630
rect 47852 39566 47854 39618
rect 47906 39566 47908 39618
rect 46396 38782 46398 38834
rect 46450 38782 46452 38834
rect 45388 37998 45390 38050
rect 45442 37998 45444 38050
rect 45388 37986 45444 37998
rect 46396 38050 46452 38782
rect 46396 37998 46398 38050
rect 46450 37998 46452 38050
rect 46396 37986 46452 37998
rect 46844 39506 46900 39518
rect 46844 39454 46846 39506
rect 46898 39454 46900 39506
rect 46844 39060 46900 39454
rect 46844 38834 46900 39004
rect 46844 38782 46846 38834
rect 46898 38782 46900 38834
rect 46844 38050 46900 38782
rect 47740 38948 47796 38958
rect 47852 38948 47908 39566
rect 47740 38946 47908 38948
rect 47740 38894 47742 38946
rect 47794 38894 47908 38946
rect 47740 38892 47908 38894
rect 47964 39618 48132 39620
rect 47964 39566 48078 39618
rect 48130 39566 48132 39618
rect 47964 39564 48132 39566
rect 47628 38610 47684 38622
rect 47628 38558 47630 38610
rect 47682 38558 47684 38610
rect 47628 38164 47684 38558
rect 47404 38108 47684 38164
rect 46844 37998 46846 38050
rect 46898 37998 46900 38050
rect 46844 37986 46900 37998
rect 47180 38052 47236 38062
rect 47180 37958 47236 37996
rect 44940 37214 44942 37266
rect 44994 37214 44996 37266
rect 44940 37202 44996 37214
rect 45612 37826 45668 37838
rect 45612 37774 45614 37826
rect 45666 37774 45668 37826
rect 45612 37268 45668 37774
rect 46844 37380 46900 37390
rect 46844 37378 47012 37380
rect 46844 37326 46846 37378
rect 46898 37326 47012 37378
rect 46844 37324 47012 37326
rect 46844 37314 46900 37324
rect 45612 37202 45668 37212
rect 46732 37268 46788 37278
rect 43484 36654 43486 36706
rect 43538 36654 43540 36706
rect 43484 36642 43540 36654
rect 43596 37154 43652 37166
rect 43596 37102 43598 37154
rect 43650 37102 43652 37154
rect 43036 36430 43038 36482
rect 43090 36430 43092 36482
rect 42700 34862 42702 34914
rect 42754 34862 42756 34914
rect 42700 34850 42756 34862
rect 42812 35474 42868 35486
rect 42812 35422 42814 35474
rect 42866 35422 42868 35474
rect 41356 34692 41412 34702
rect 41580 34692 41636 34702
rect 41356 34690 41580 34692
rect 41356 34638 41358 34690
rect 41410 34638 41580 34690
rect 41356 34636 41580 34638
rect 41356 34626 41412 34636
rect 41244 34354 41300 34366
rect 41244 34302 41246 34354
rect 41298 34302 41300 34354
rect 40908 34190 40910 34242
rect 40962 34190 40964 34242
rect 40908 34178 40964 34190
rect 41132 34244 41188 34254
rect 41132 34150 41188 34188
rect 41020 34132 41076 34142
rect 41020 33572 41076 34076
rect 41020 33478 41076 33516
rect 41132 33460 41188 33470
rect 41244 33460 41300 34302
rect 41580 34130 41636 34636
rect 42588 34580 42644 34590
rect 42140 34244 42196 34254
rect 42140 34150 42196 34188
rect 41580 34078 41582 34130
rect 41634 34078 41636 34130
rect 41580 34066 41636 34078
rect 41804 34132 41860 34142
rect 41804 34038 41860 34076
rect 42588 34130 42644 34524
rect 42812 34244 42868 35422
rect 43036 34916 43092 36430
rect 43372 36596 43428 36606
rect 43372 36370 43428 36540
rect 43372 36318 43374 36370
rect 43426 36318 43428 36370
rect 43372 36306 43428 36318
rect 43596 35252 43652 37102
rect 46172 37156 46228 37166
rect 46172 37062 46228 37100
rect 45612 37044 45668 37054
rect 44044 36596 44100 36606
rect 44044 36502 44100 36540
rect 45612 36596 45668 36988
rect 45612 36482 45668 36540
rect 45612 36430 45614 36482
rect 45666 36430 45668 36482
rect 45612 36418 45668 36430
rect 45948 36932 46004 36942
rect 45948 36370 46004 36876
rect 45948 36318 45950 36370
rect 46002 36318 46004 36370
rect 45948 36306 46004 36318
rect 46732 36148 46788 37212
rect 46844 37042 46900 37054
rect 46844 36990 46846 37042
rect 46898 36990 46900 37042
rect 46844 36370 46900 36990
rect 46956 36932 47012 37324
rect 47292 37156 47348 37166
rect 46956 36866 47012 36876
rect 47180 37154 47348 37156
rect 47180 37102 47294 37154
rect 47346 37102 47348 37154
rect 47180 37100 47348 37102
rect 46844 36318 46846 36370
rect 46898 36318 46900 36370
rect 46844 36306 46900 36318
rect 47180 36260 47236 37100
rect 47292 37090 47348 37100
rect 47292 36484 47348 36494
rect 47404 36484 47460 38108
rect 47740 38052 47796 38892
rect 47964 38722 48020 39564
rect 48076 39554 48132 39564
rect 47964 38670 47966 38722
rect 48018 38670 48020 38722
rect 47964 38276 48020 38670
rect 47964 38210 48020 38220
rect 48076 39396 48132 39406
rect 47964 38052 48020 38062
rect 47740 37996 47964 38052
rect 47964 37958 48020 37996
rect 47628 37940 47684 37950
rect 47628 37378 47684 37884
rect 47628 37326 47630 37378
rect 47682 37326 47684 37378
rect 47628 37314 47684 37326
rect 47516 37268 47572 37278
rect 47516 37174 47572 37212
rect 48076 37266 48132 39340
rect 48188 38164 48244 38174
rect 48188 38070 48244 38108
rect 48636 38052 48692 39788
rect 48748 39620 48804 40236
rect 48860 39844 48916 41918
rect 48972 41972 49028 42364
rect 48972 41906 49028 41916
rect 49084 42082 49140 42094
rect 49084 42030 49086 42082
rect 49138 42030 49140 42082
rect 49084 40516 49140 42030
rect 49196 41748 49252 43036
rect 49308 41748 49364 41758
rect 49196 41692 49308 41748
rect 49308 41682 49364 41692
rect 49084 40450 49140 40460
rect 49196 40514 49252 40526
rect 49196 40462 49198 40514
rect 49250 40462 49252 40514
rect 48972 40292 49028 40302
rect 48972 40290 49140 40292
rect 48972 40238 48974 40290
rect 49026 40238 49140 40290
rect 48972 40236 49140 40238
rect 48972 40226 49028 40236
rect 48860 39778 48916 39788
rect 48972 39732 49028 39742
rect 48860 39620 48916 39630
rect 48748 39618 48916 39620
rect 48748 39566 48862 39618
rect 48914 39566 48916 39618
rect 48748 39564 48916 39566
rect 48860 39554 48916 39564
rect 48748 39396 48804 39406
rect 48748 39302 48804 39340
rect 48860 39284 48916 39294
rect 48860 39058 48916 39228
rect 48860 39006 48862 39058
rect 48914 39006 48916 39058
rect 48860 38994 48916 39006
rect 48748 38834 48804 38846
rect 48748 38782 48750 38834
rect 48802 38782 48804 38834
rect 48748 38724 48804 38782
rect 48972 38724 49028 39676
rect 49084 39730 49140 40236
rect 49084 39678 49086 39730
rect 49138 39678 49140 39730
rect 49084 39666 49140 39678
rect 49084 39060 49140 39070
rect 49196 39060 49252 40462
rect 49308 39620 49364 39630
rect 49308 39526 49364 39564
rect 49420 39618 49476 43260
rect 49644 41970 49700 44158
rect 49756 43708 49812 44940
rect 49756 43652 49924 43708
rect 49644 41918 49646 41970
rect 49698 41918 49700 41970
rect 49644 41906 49700 41918
rect 49756 43316 49812 43326
rect 49532 41860 49588 41870
rect 49532 41766 49588 41804
rect 49756 41860 49812 43260
rect 49868 42754 49924 43652
rect 49868 42702 49870 42754
rect 49922 42702 49924 42754
rect 49868 42690 49924 42702
rect 49980 42756 50036 45054
rect 50316 46564 50372 46574
rect 50092 44884 50148 44894
rect 50092 44790 50148 44828
rect 49980 42690 50036 42700
rect 50316 42642 50372 46508
rect 50876 46562 50932 47404
rect 51100 47394 51156 47404
rect 51324 46788 51380 48300
rect 52668 47908 52724 50430
rect 52780 50482 52836 50494
rect 52780 50430 52782 50482
rect 52834 50430 52836 50482
rect 52780 50372 52836 50430
rect 53228 50482 53284 50494
rect 53228 50430 53230 50482
rect 53282 50430 53284 50482
rect 52780 50306 52836 50316
rect 53004 50370 53060 50382
rect 53004 50318 53006 50370
rect 53058 50318 53060 50370
rect 52780 50036 52836 50046
rect 52780 49810 52836 49980
rect 52780 49758 52782 49810
rect 52834 49758 52836 49810
rect 52780 49746 52836 49758
rect 53004 49810 53060 50318
rect 53228 50372 53284 50430
rect 53228 50306 53284 50316
rect 53340 50372 53396 50382
rect 53340 50370 53956 50372
rect 53340 50318 53342 50370
rect 53394 50318 53956 50370
rect 53340 50316 53956 50318
rect 53340 50306 53396 50316
rect 53676 50036 53732 50046
rect 53676 49922 53732 49980
rect 53900 50034 53956 50316
rect 53900 49982 53902 50034
rect 53954 49982 53956 50034
rect 53900 49970 53956 49982
rect 53676 49870 53678 49922
rect 53730 49870 53732 49922
rect 53676 49858 53732 49870
rect 53004 49758 53006 49810
rect 53058 49758 53060 49810
rect 53004 49746 53060 49758
rect 53900 49698 53956 49710
rect 53900 49646 53902 49698
rect 53954 49646 53956 49698
rect 53340 49588 53396 49598
rect 52892 49586 53620 49588
rect 52892 49534 53342 49586
rect 53394 49534 53620 49586
rect 52892 49532 53620 49534
rect 52332 47852 52724 47908
rect 52780 49138 52836 49150
rect 52780 49086 52782 49138
rect 52834 49086 52836 49138
rect 51660 47346 51716 47358
rect 51660 47294 51662 47346
rect 51714 47294 51716 47346
rect 51436 46900 51492 46910
rect 51436 46806 51492 46844
rect 50876 46510 50878 46562
rect 50930 46510 50932 46562
rect 50876 46498 50932 46510
rect 51100 46786 51380 46788
rect 51100 46734 51326 46786
rect 51378 46734 51380 46786
rect 51100 46732 51380 46734
rect 50988 45780 51044 45790
rect 50988 45686 51044 45724
rect 50556 45500 50820 45510
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50556 45434 50820 45444
rect 50652 44884 50708 44894
rect 50652 44322 50708 44828
rect 50652 44270 50654 44322
rect 50706 44270 50708 44322
rect 50652 44258 50708 44270
rect 50764 44212 50820 44222
rect 50764 44118 50820 44156
rect 50988 44098 51044 44110
rect 50988 44046 50990 44098
rect 51042 44046 51044 44098
rect 50556 43932 50820 43942
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50556 43866 50820 43876
rect 50988 43708 51044 44046
rect 50876 43652 51044 43708
rect 51100 43764 51156 46732
rect 51324 46722 51380 46732
rect 51548 46564 51604 46574
rect 51436 46452 51492 46462
rect 51436 46358 51492 46396
rect 51548 45778 51604 46508
rect 51660 45892 51716 47294
rect 51772 45892 51828 45902
rect 51660 45890 51828 45892
rect 51660 45838 51774 45890
rect 51826 45838 51828 45890
rect 51660 45836 51828 45838
rect 51772 45826 51828 45836
rect 51548 45726 51550 45778
rect 51602 45726 51604 45778
rect 51548 45714 51604 45726
rect 52332 45780 52388 47852
rect 52780 47572 52836 49086
rect 52892 48914 52948 49532
rect 53340 49522 53396 49532
rect 53116 49252 53172 49262
rect 53564 49252 53620 49532
rect 53900 49252 53956 49646
rect 53172 49196 53396 49252
rect 53564 49196 53844 49252
rect 53116 49158 53172 49196
rect 52892 48862 52894 48914
rect 52946 48862 52948 48914
rect 52892 48850 52948 48862
rect 52668 46676 52724 46686
rect 52780 46676 52836 47516
rect 53116 48468 53172 48478
rect 53116 47460 53172 48412
rect 53340 48466 53396 49196
rect 53788 49138 53844 49196
rect 53900 49186 53956 49196
rect 53788 49086 53790 49138
rect 53842 49086 53844 49138
rect 53788 49074 53844 49086
rect 53340 48414 53342 48466
rect 53394 48414 53396 48466
rect 53340 48402 53396 48414
rect 53676 48802 53732 48814
rect 53676 48750 53678 48802
rect 53730 48750 53732 48802
rect 53676 48242 53732 48750
rect 53676 48190 53678 48242
rect 53730 48190 53732 48242
rect 53676 48178 53732 48190
rect 53004 47458 53172 47460
rect 53004 47406 53118 47458
rect 53170 47406 53172 47458
rect 53004 47404 53172 47406
rect 52668 46674 52836 46676
rect 52668 46622 52670 46674
rect 52722 46622 52836 46674
rect 52668 46620 52836 46622
rect 52892 47346 52948 47358
rect 52892 47294 52894 47346
rect 52946 47294 52948 47346
rect 52668 46610 52724 46620
rect 52780 46116 52836 46126
rect 52780 46022 52836 46060
rect 52668 45780 52724 45790
rect 52332 45778 52724 45780
rect 52332 45726 52670 45778
rect 52722 45726 52724 45778
rect 52332 45724 52724 45726
rect 51324 45668 51380 45678
rect 51324 45666 51492 45668
rect 51324 45614 51326 45666
rect 51378 45614 51492 45666
rect 51324 45612 51492 45614
rect 51324 45602 51380 45612
rect 51436 45332 51492 45612
rect 51436 45276 51716 45332
rect 51660 45220 51716 45276
rect 52556 45330 52612 45342
rect 52556 45278 52558 45330
rect 52610 45278 52612 45330
rect 52444 45220 52500 45230
rect 51660 45218 51940 45220
rect 51660 45166 51662 45218
rect 51714 45166 51940 45218
rect 51660 45164 51940 45166
rect 51660 45154 51716 45164
rect 51548 45106 51604 45118
rect 51548 45054 51550 45106
rect 51602 45054 51604 45106
rect 51548 44884 51604 45054
rect 51604 44828 51828 44884
rect 51548 44818 51604 44828
rect 51660 44324 51716 44334
rect 51660 44230 51716 44268
rect 51772 44322 51828 44828
rect 51772 44270 51774 44322
rect 51826 44270 51828 44322
rect 51772 44258 51828 44270
rect 51884 44212 51940 45164
rect 51884 44118 51940 44156
rect 51996 45108 52052 45118
rect 51100 43698 51156 43708
rect 51212 44098 51268 44110
rect 51212 44046 51214 44098
rect 51266 44046 51268 44098
rect 50876 43426 50932 43652
rect 50876 43374 50878 43426
rect 50930 43374 50932 43426
rect 50876 43362 50932 43374
rect 51212 42866 51268 44046
rect 51996 43988 52052 45052
rect 51884 43932 52052 43988
rect 52444 45106 52500 45164
rect 52444 45054 52446 45106
rect 52498 45054 52500 45106
rect 52444 44324 52500 45054
rect 52556 45108 52612 45278
rect 52556 45042 52612 45052
rect 51324 43652 51380 43662
rect 51324 43650 51492 43652
rect 51324 43598 51326 43650
rect 51378 43598 51492 43650
rect 51324 43596 51492 43598
rect 51324 43586 51380 43596
rect 51212 42814 51214 42866
rect 51266 42814 51268 42866
rect 51212 42802 51268 42814
rect 51436 42756 51492 43596
rect 51324 42754 51492 42756
rect 51324 42702 51438 42754
rect 51490 42702 51492 42754
rect 51324 42700 51492 42702
rect 50316 42590 50318 42642
rect 50370 42590 50372 42642
rect 49868 42530 49924 42542
rect 49868 42478 49870 42530
rect 49922 42478 49924 42530
rect 49868 41972 49924 42478
rect 49868 41906 49924 41916
rect 49756 41636 49812 41804
rect 49756 41570 49812 41580
rect 50316 41524 50372 42590
rect 50652 42644 50708 42654
rect 51324 42644 51380 42700
rect 51436 42690 51492 42700
rect 51548 43428 51604 43438
rect 50652 42642 51380 42644
rect 50652 42590 50654 42642
rect 50706 42590 51380 42642
rect 50652 42588 51380 42590
rect 50652 42578 50708 42588
rect 50428 42532 50484 42542
rect 50428 42438 50484 42476
rect 50556 42364 50820 42374
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50556 42298 50820 42308
rect 51436 41970 51492 41982
rect 51436 41918 51438 41970
rect 51490 41918 51492 41970
rect 51436 41860 51492 41918
rect 51436 41794 51492 41804
rect 50316 41458 50372 41468
rect 50428 41746 50484 41758
rect 50428 41694 50430 41746
rect 50482 41694 50484 41746
rect 50428 41188 50484 41694
rect 51212 41188 51268 41198
rect 51548 41188 51604 43372
rect 51884 42754 51940 43932
rect 51884 42702 51886 42754
rect 51938 42702 51940 42754
rect 51884 42690 51940 42702
rect 51996 43764 52052 43774
rect 50428 41094 50484 41132
rect 50876 41186 51604 41188
rect 50876 41134 51214 41186
rect 51266 41134 51604 41186
rect 50876 41132 51604 41134
rect 50556 40796 50820 40806
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50556 40730 50820 40740
rect 50652 40628 50708 40638
rect 50652 40534 50708 40572
rect 50764 40516 50820 40526
rect 50876 40516 50932 41132
rect 51212 41122 51268 41132
rect 50764 40514 50932 40516
rect 50764 40462 50766 40514
rect 50818 40462 50932 40514
rect 50764 40460 50932 40462
rect 50764 40450 50820 40460
rect 51548 40402 51604 41132
rect 51660 42530 51716 42542
rect 51660 42478 51662 42530
rect 51714 42478 51716 42530
rect 51660 41186 51716 42478
rect 51996 41860 52052 43708
rect 52444 43538 52500 44268
rect 52444 43486 52446 43538
rect 52498 43486 52500 43538
rect 52444 43474 52500 43486
rect 52668 42642 52724 45724
rect 52780 45780 52836 45790
rect 52780 45686 52836 45724
rect 52892 45220 52948 47294
rect 53004 46674 53060 47404
rect 53116 47394 53172 47404
rect 53228 48130 53284 48142
rect 53228 48078 53230 48130
rect 53282 48078 53284 48130
rect 53228 46900 53284 48078
rect 54124 47572 54180 47582
rect 54124 47458 54180 47516
rect 54124 47406 54126 47458
rect 54178 47406 54180 47458
rect 54124 47394 54180 47406
rect 54460 47458 54516 47470
rect 54460 47406 54462 47458
rect 54514 47406 54516 47458
rect 53228 46834 53284 46844
rect 54124 46900 54180 46910
rect 54124 46786 54180 46844
rect 54124 46734 54126 46786
rect 54178 46734 54180 46786
rect 53004 46622 53006 46674
rect 53058 46622 53060 46674
rect 53004 46610 53060 46622
rect 53788 46674 53844 46686
rect 53788 46622 53790 46674
rect 53842 46622 53844 46674
rect 53116 46564 53172 46574
rect 53452 46564 53508 46574
rect 53116 46562 53508 46564
rect 53116 46510 53118 46562
rect 53170 46510 53454 46562
rect 53506 46510 53508 46562
rect 53116 46508 53508 46510
rect 53116 46498 53172 46508
rect 53452 46498 53508 46508
rect 53564 46562 53620 46574
rect 53564 46510 53566 46562
rect 53618 46510 53620 46562
rect 52892 45154 52948 45164
rect 53004 45108 53060 45118
rect 53004 45014 53060 45052
rect 53452 45108 53508 45118
rect 53564 45108 53620 46510
rect 53788 46452 53844 46622
rect 53788 46386 53844 46396
rect 54124 46002 54180 46734
rect 54236 46788 54292 46798
rect 54236 46786 54404 46788
rect 54236 46734 54238 46786
rect 54290 46734 54404 46786
rect 54236 46732 54404 46734
rect 54236 46722 54292 46732
rect 54124 45950 54126 46002
rect 54178 45950 54180 46002
rect 54124 45938 54180 45950
rect 54236 46450 54292 46462
rect 54236 46398 54238 46450
rect 54290 46398 54292 46450
rect 53452 45106 53620 45108
rect 53452 45054 53454 45106
rect 53506 45054 53620 45106
rect 53452 45052 53620 45054
rect 53788 45108 53844 45118
rect 53452 45042 53508 45052
rect 53788 45014 53844 45052
rect 54124 45108 54180 45118
rect 53900 44210 53956 44222
rect 53900 44158 53902 44210
rect 53954 44158 53956 44210
rect 53228 43428 53284 43438
rect 53228 43334 53284 43372
rect 53900 42756 53956 44158
rect 54124 43764 54180 45052
rect 54236 45106 54292 46398
rect 54348 46116 54404 46732
rect 54460 46452 54516 47406
rect 54460 46386 54516 46396
rect 54348 45890 54404 46060
rect 54348 45838 54350 45890
rect 54402 45838 54404 45890
rect 54348 45826 54404 45838
rect 54796 46002 54852 46014
rect 54796 45950 54798 46002
rect 54850 45950 54852 46002
rect 54796 45330 54852 45950
rect 54796 45278 54798 45330
rect 54850 45278 54852 45330
rect 54236 45054 54238 45106
rect 54290 45054 54292 45106
rect 54236 45042 54292 45054
rect 54572 45108 54628 45118
rect 54572 45014 54628 45052
rect 54684 44994 54740 45006
rect 54684 44942 54686 44994
rect 54738 44942 54740 44994
rect 54684 44548 54740 44942
rect 54124 43538 54180 43708
rect 54124 43486 54126 43538
rect 54178 43486 54180 43538
rect 54124 43474 54180 43486
rect 54236 44492 54740 44548
rect 54236 43204 54292 44492
rect 54796 44322 54852 45278
rect 55692 44324 55748 44334
rect 54796 44270 54798 44322
rect 54850 44270 54852 44322
rect 54796 43708 54852 44270
rect 55468 44322 55748 44324
rect 55468 44270 55694 44322
rect 55746 44270 55748 44322
rect 55468 44268 55748 44270
rect 55244 43764 55300 43802
rect 55468 43764 55524 44268
rect 55692 44258 55748 44268
rect 55300 43708 55524 43764
rect 55804 44210 55860 44222
rect 55804 44158 55806 44210
rect 55858 44158 55860 44210
rect 55804 43708 55860 44158
rect 54348 43652 55076 43708
rect 55244 43698 55300 43708
rect 54348 43538 54404 43652
rect 55020 43650 55076 43652
rect 55020 43598 55022 43650
rect 55074 43598 55076 43650
rect 55020 43586 55076 43598
rect 55692 43652 55860 43708
rect 54348 43486 54350 43538
rect 54402 43486 54404 43538
rect 54348 43474 54404 43486
rect 54684 43314 54740 43326
rect 54684 43262 54686 43314
rect 54738 43262 54740 43314
rect 54236 43148 54628 43204
rect 54348 42980 54404 42990
rect 54348 42978 54516 42980
rect 54348 42926 54350 42978
rect 54402 42926 54516 42978
rect 54348 42924 54516 42926
rect 54348 42914 54404 42924
rect 54124 42756 54180 42766
rect 53900 42754 54180 42756
rect 53900 42702 54126 42754
rect 54178 42702 54180 42754
rect 53900 42700 54180 42702
rect 52668 42590 52670 42642
rect 52722 42590 52724 42642
rect 52444 41972 52500 41982
rect 52444 41878 52500 41916
rect 51996 41748 52052 41804
rect 51884 41692 52052 41748
rect 52668 41748 52724 42590
rect 52780 42532 52836 42542
rect 52780 42084 52836 42476
rect 52780 42018 52836 42028
rect 53004 42530 53060 42542
rect 53004 42478 53006 42530
rect 53058 42478 53060 42530
rect 52892 41858 52948 41870
rect 52892 41806 52894 41858
rect 52946 41806 52948 41858
rect 52892 41748 52948 41806
rect 52668 41692 52836 41748
rect 51660 41134 51662 41186
rect 51714 41134 51716 41186
rect 51660 41122 51716 41134
rect 51772 41188 51828 41198
rect 51548 40350 51550 40402
rect 51602 40350 51604 40402
rect 51548 40338 51604 40350
rect 51772 40402 51828 41132
rect 51772 40350 51774 40402
rect 51826 40350 51828 40402
rect 51772 40338 51828 40350
rect 51324 40290 51380 40302
rect 51324 40238 51326 40290
rect 51378 40238 51380 40290
rect 51100 39730 51156 39742
rect 51100 39678 51102 39730
rect 51154 39678 51156 39730
rect 49420 39566 49422 39618
rect 49474 39566 49476 39618
rect 49420 39554 49476 39566
rect 49980 39618 50036 39630
rect 49980 39566 49982 39618
rect 50034 39566 50036 39618
rect 49084 39058 49252 39060
rect 49084 39006 49086 39058
rect 49138 39006 49252 39058
rect 49084 39004 49252 39006
rect 49084 38994 49140 39004
rect 49644 38946 49700 38958
rect 49644 38894 49646 38946
rect 49698 38894 49700 38946
rect 49308 38836 49364 38846
rect 49196 38780 49308 38836
rect 49196 38724 49252 38780
rect 49308 38742 49364 38780
rect 48748 38668 49252 38724
rect 48748 38052 48804 38062
rect 48636 38050 48804 38052
rect 48636 37998 48750 38050
rect 48802 37998 48804 38050
rect 48636 37996 48804 37998
rect 48300 37940 48356 37950
rect 48300 37846 48356 37884
rect 48076 37214 48078 37266
rect 48130 37214 48132 37266
rect 48076 37202 48132 37214
rect 47292 36482 47460 36484
rect 47292 36430 47294 36482
rect 47346 36430 47460 36482
rect 47292 36428 47460 36430
rect 48300 37042 48356 37054
rect 48300 36990 48302 37042
rect 48354 36990 48356 37042
rect 47292 36418 47348 36428
rect 47180 36204 47348 36260
rect 46396 36092 46788 36148
rect 44044 35810 44100 35822
rect 44044 35758 44046 35810
rect 44098 35758 44100 35810
rect 43596 35186 43652 35196
rect 43708 35586 43764 35598
rect 43708 35534 43710 35586
rect 43762 35534 43764 35586
rect 43036 34850 43092 34860
rect 43148 35138 43204 35150
rect 43148 35086 43150 35138
rect 43202 35086 43204 35138
rect 42812 34178 42868 34188
rect 42924 34354 42980 34366
rect 42924 34302 42926 34354
rect 42978 34302 42980 34354
rect 42588 34078 42590 34130
rect 42642 34078 42644 34130
rect 42588 34066 42644 34078
rect 41916 34018 41972 34030
rect 41916 33966 41918 34018
rect 41970 33966 41972 34018
rect 41804 33572 41860 33582
rect 41804 33478 41860 33516
rect 41132 33458 41300 33460
rect 41132 33406 41134 33458
rect 41186 33406 41300 33458
rect 41132 33404 41300 33406
rect 41132 33394 41188 33404
rect 41916 33348 41972 33966
rect 42140 33572 42196 33582
rect 42924 33572 42980 34302
rect 43036 34244 43092 34254
rect 43036 34150 43092 34188
rect 43148 34130 43204 35086
rect 43484 34356 43540 34366
rect 43708 34356 43764 35534
rect 43820 34916 43876 34926
rect 43820 34822 43876 34860
rect 44044 34916 44100 35758
rect 44268 35812 44324 35822
rect 44044 34850 44100 34860
rect 44156 34916 44212 34926
rect 44268 34916 44324 35756
rect 45276 35812 45332 35822
rect 45276 35718 45332 35756
rect 45724 35586 45780 35598
rect 45724 35534 45726 35586
rect 45778 35534 45780 35586
rect 45276 35252 45332 35262
rect 44156 34914 44548 34916
rect 44156 34862 44158 34914
rect 44210 34862 44548 34914
rect 44156 34860 44548 34862
rect 44156 34850 44212 34860
rect 43932 34692 43988 34702
rect 43932 34598 43988 34636
rect 43708 34300 43988 34356
rect 43484 34262 43540 34300
rect 43596 34244 43652 34254
rect 43596 34242 43764 34244
rect 43596 34190 43598 34242
rect 43650 34190 43764 34242
rect 43596 34188 43764 34190
rect 43596 34178 43652 34188
rect 43148 34078 43150 34130
rect 43202 34078 43204 34130
rect 43148 34066 43204 34078
rect 42140 33570 42980 33572
rect 42140 33518 42142 33570
rect 42194 33518 42980 33570
rect 42140 33516 42980 33518
rect 42140 33506 42196 33516
rect 41916 33254 41972 33292
rect 42700 33348 42756 33358
rect 42700 33254 42756 33292
rect 42924 33346 42980 33516
rect 42924 33294 42926 33346
rect 42978 33294 42980 33346
rect 42924 33282 42980 33294
rect 43708 34020 43764 34188
rect 40460 33170 40516 33180
rect 42252 33234 42308 33246
rect 42252 33182 42254 33234
rect 42306 33182 42308 33234
rect 40684 33124 40740 33134
rect 40684 33122 40964 33124
rect 40684 33070 40686 33122
rect 40738 33070 40964 33122
rect 40684 33068 40964 33070
rect 40684 33058 40740 33068
rect 38892 32722 38948 32732
rect 40684 32788 40740 32798
rect 38332 32450 38500 32452
rect 38332 32398 38334 32450
rect 38386 32398 38500 32450
rect 38332 32396 38500 32398
rect 38556 32676 38612 32686
rect 38332 31780 38388 32396
rect 38556 31948 38612 32620
rect 38556 31892 38724 31948
rect 38332 31714 38388 31724
rect 38332 31220 38388 31230
rect 38556 31220 38612 31230
rect 38388 31218 38612 31220
rect 38388 31166 38558 31218
rect 38610 31166 38612 31218
rect 38388 31164 38612 31166
rect 38332 31154 38388 31164
rect 38556 31154 38612 31164
rect 38668 31218 38724 31892
rect 39900 31890 39956 31902
rect 39900 31838 39902 31890
rect 39954 31838 39956 31890
rect 39564 31780 39620 31790
rect 38668 31166 38670 31218
rect 38722 31166 38724 31218
rect 38220 30942 38222 30994
rect 38274 30942 38276 30994
rect 38220 30930 38276 30942
rect 38444 30996 38500 31006
rect 38444 30902 38500 30940
rect 37996 30772 38052 30782
rect 37996 30770 38164 30772
rect 37996 30718 37998 30770
rect 38050 30718 38164 30770
rect 37996 30716 38164 30718
rect 37996 30706 38052 30716
rect 37996 30324 38052 30334
rect 37996 30230 38052 30268
rect 37548 29538 37716 29540
rect 37548 29486 37550 29538
rect 37602 29486 37716 29538
rect 37548 29484 37716 29486
rect 37772 29820 37940 29876
rect 37548 29474 37604 29484
rect 37436 29314 37492 29326
rect 37436 29262 37438 29314
rect 37490 29262 37492 29314
rect 37324 28532 37380 28542
rect 37212 28476 37324 28532
rect 37324 28438 37380 28476
rect 37100 28420 37156 28430
rect 36876 28364 37044 28420
rect 36652 28082 36820 28084
rect 36652 28030 36654 28082
rect 36706 28030 36820 28082
rect 36652 28028 36820 28030
rect 36652 27972 36708 28028
rect 36652 27906 36708 27916
rect 36988 27860 37044 28364
rect 37100 28082 37156 28364
rect 37100 28030 37102 28082
rect 37154 28030 37156 28082
rect 37100 28018 37156 28030
rect 37324 28084 37380 28094
rect 37436 28084 37492 29262
rect 37660 28644 37716 28654
rect 37660 28550 37716 28588
rect 37772 28420 37828 29820
rect 37996 29652 38052 29662
rect 38108 29652 38164 30716
rect 37996 29650 38164 29652
rect 37996 29598 37998 29650
rect 38050 29598 38164 29650
rect 37996 29596 38164 29598
rect 38220 30548 38276 30558
rect 37996 29586 38052 29596
rect 37324 28082 37492 28084
rect 37324 28030 37326 28082
rect 37378 28030 37492 28082
rect 37324 28028 37492 28030
rect 37660 28364 37828 28420
rect 37884 29426 37940 29438
rect 37884 29374 37886 29426
rect 37938 29374 37940 29426
rect 37884 28532 37940 29374
rect 38108 29428 38164 29438
rect 38220 29428 38276 30492
rect 38556 30436 38612 30446
rect 38668 30436 38724 31166
rect 39228 31444 39284 31454
rect 39228 31106 39284 31388
rect 39228 31054 39230 31106
rect 39282 31054 39284 31106
rect 39228 31042 39284 31054
rect 39116 30996 39172 31006
rect 39116 30902 39172 30940
rect 38612 30380 38724 30436
rect 38556 30098 38612 30380
rect 39564 30212 39620 31724
rect 39900 31444 39956 31838
rect 40348 31780 40404 31790
rect 40348 31686 40404 31724
rect 39900 31378 39956 31388
rect 39676 30884 39732 30894
rect 39676 30790 39732 30828
rect 40572 30436 40628 30446
rect 39788 30212 39844 30222
rect 39564 30210 39844 30212
rect 39564 30158 39566 30210
rect 39618 30158 39790 30210
rect 39842 30158 39844 30210
rect 39564 30156 39844 30158
rect 39564 30146 39620 30156
rect 39788 30146 39844 30156
rect 40572 30210 40628 30380
rect 40572 30158 40574 30210
rect 40626 30158 40628 30210
rect 40572 30146 40628 30158
rect 38556 30046 38558 30098
rect 38610 30046 38612 30098
rect 38556 30034 38612 30046
rect 38892 29986 38948 29998
rect 38892 29934 38894 29986
rect 38946 29934 38948 29986
rect 38108 29426 38276 29428
rect 38108 29374 38110 29426
rect 38162 29374 38276 29426
rect 38108 29372 38276 29374
rect 38556 29428 38612 29438
rect 38892 29428 38948 29934
rect 40348 29876 40404 29886
rect 38556 29426 38948 29428
rect 38556 29374 38558 29426
rect 38610 29374 38948 29426
rect 38556 29372 38948 29374
rect 40012 29652 40068 29662
rect 38108 29362 38164 29372
rect 38556 29362 38612 29372
rect 38668 28644 38724 29372
rect 39900 29316 39956 29326
rect 37324 28018 37380 28028
rect 36988 27804 37156 27860
rect 36316 26898 36372 26908
rect 36988 27074 37044 27086
rect 36988 27022 36990 27074
rect 37042 27022 37044 27074
rect 36988 26180 37044 27022
rect 37100 26628 37156 27804
rect 37212 27746 37268 27758
rect 37212 27694 37214 27746
rect 37266 27694 37268 27746
rect 37212 27300 37268 27694
rect 37660 27636 37716 28364
rect 37884 28084 37940 28476
rect 37996 28642 38724 28644
rect 37996 28590 38670 28642
rect 38722 28590 38724 28642
rect 37996 28588 38724 28590
rect 37996 28530 38052 28588
rect 37996 28478 37998 28530
rect 38050 28478 38052 28530
rect 37996 28466 38052 28478
rect 37884 28018 37940 28028
rect 38556 28418 38612 28430
rect 38556 28366 38558 28418
rect 38610 28366 38612 28418
rect 38444 27972 38500 27982
rect 38444 27878 38500 27916
rect 37772 27860 37828 27870
rect 38220 27860 38276 27870
rect 37772 27858 38276 27860
rect 37772 27806 37774 27858
rect 37826 27806 38222 27858
rect 38274 27806 38276 27858
rect 37772 27804 38276 27806
rect 37772 27794 37828 27804
rect 38220 27794 38276 27804
rect 38556 27858 38612 28366
rect 38556 27806 38558 27858
rect 38610 27806 38612 27858
rect 38556 27636 38612 27806
rect 38668 27860 38724 28588
rect 38892 28756 38948 28766
rect 38780 28532 38836 28542
rect 38780 28196 38836 28476
rect 38780 28130 38836 28140
rect 38780 27860 38836 27870
rect 38668 27858 38836 27860
rect 38668 27806 38782 27858
rect 38834 27806 38836 27858
rect 38668 27804 38836 27806
rect 38780 27794 38836 27804
rect 37660 27580 37940 27636
rect 37212 27244 37828 27300
rect 37772 27186 37828 27244
rect 37772 27134 37774 27186
rect 37826 27134 37828 27186
rect 37772 27122 37828 27134
rect 37884 26908 37940 27580
rect 38556 27570 38612 27580
rect 38892 27076 38948 28700
rect 39900 28756 39956 29260
rect 39900 28690 39956 28700
rect 39004 28532 39060 28542
rect 39004 28308 39060 28476
rect 39340 28532 39396 28542
rect 39340 28438 39396 28476
rect 39004 28242 39060 28252
rect 39116 28420 39172 28430
rect 39116 28084 39172 28364
rect 39228 28418 39284 28430
rect 39228 28366 39230 28418
rect 39282 28366 39284 28418
rect 39228 28308 39284 28366
rect 39228 28242 39284 28252
rect 39900 28418 39956 28430
rect 39900 28366 39902 28418
rect 39954 28366 39956 28418
rect 39340 28140 39844 28196
rect 39228 28084 39284 28094
rect 39116 28082 39284 28084
rect 39116 28030 39230 28082
rect 39282 28030 39284 28082
rect 39116 28028 39284 28030
rect 39228 28018 39284 28028
rect 39340 28082 39396 28140
rect 39340 28030 39342 28082
rect 39394 28030 39396 28082
rect 39340 28018 39396 28030
rect 39788 28082 39844 28140
rect 39788 28030 39790 28082
rect 39842 28030 39844 28082
rect 39788 28018 39844 28030
rect 39900 27972 39956 28366
rect 40012 28082 40068 29596
rect 40348 29650 40404 29820
rect 40348 29598 40350 29650
rect 40402 29598 40404 29650
rect 40348 29586 40404 29598
rect 40684 29092 40740 32732
rect 40908 31220 40964 33068
rect 42140 32788 42196 32798
rect 42252 32788 42308 33182
rect 42140 32786 42308 32788
rect 42140 32734 42142 32786
rect 42194 32734 42308 32786
rect 42140 32732 42308 32734
rect 42700 32788 42756 32798
rect 42140 32722 42196 32732
rect 42364 32564 42420 32574
rect 42588 32564 42644 32574
rect 42364 32562 42644 32564
rect 42364 32510 42366 32562
rect 42418 32510 42590 32562
rect 42642 32510 42644 32562
rect 42364 32508 42644 32510
rect 42364 32498 42420 32508
rect 42588 32498 42644 32508
rect 42028 32338 42084 32350
rect 42028 32286 42030 32338
rect 42082 32286 42084 32338
rect 42028 32004 42084 32286
rect 42028 31938 42084 31948
rect 40908 31164 41860 31220
rect 41356 30994 41412 31006
rect 41356 30942 41358 30994
rect 41410 30942 41412 30994
rect 41020 30884 41076 30894
rect 41356 30884 41412 30942
rect 41020 30882 41412 30884
rect 41020 30830 41022 30882
rect 41074 30830 41412 30882
rect 41020 30828 41412 30830
rect 41020 30548 41076 30828
rect 41020 30482 41076 30492
rect 41580 29988 41636 29998
rect 40796 29652 40852 29662
rect 40796 29558 40852 29596
rect 40908 29426 40964 29438
rect 40908 29374 40910 29426
rect 40962 29374 40964 29426
rect 40908 29316 40964 29374
rect 40908 29250 40964 29260
rect 40684 29036 41300 29092
rect 41244 28866 41300 29036
rect 41244 28814 41246 28866
rect 41298 28814 41300 28866
rect 41244 28802 41300 28814
rect 40012 28030 40014 28082
rect 40066 28030 40068 28082
rect 40012 28018 40068 28030
rect 40348 28642 40404 28654
rect 40348 28590 40350 28642
rect 40402 28590 40404 28642
rect 39900 27906 39956 27916
rect 40124 27972 40180 27982
rect 38892 27010 38948 27020
rect 39452 27860 39508 27870
rect 37884 26852 38500 26908
rect 37100 26562 37156 26572
rect 37100 26180 37156 26190
rect 36988 26178 37156 26180
rect 36988 26126 37102 26178
rect 37154 26126 37156 26178
rect 36988 26124 37156 26126
rect 35980 25454 35982 25506
rect 36034 25454 36036 25506
rect 35980 25442 36036 25454
rect 36204 25508 36260 25518
rect 36204 25394 36260 25452
rect 36204 25342 36206 25394
rect 36258 25342 36260 25394
rect 36204 25330 36260 25342
rect 35420 24854 35476 24892
rect 35532 24892 35700 24948
rect 37100 25284 37156 26124
rect 37772 25732 37828 25742
rect 37548 25730 37828 25732
rect 37548 25678 37774 25730
rect 37826 25678 37828 25730
rect 37548 25676 37828 25678
rect 37548 25506 37604 25676
rect 37772 25666 37828 25676
rect 38220 25730 38276 25742
rect 38220 25678 38222 25730
rect 38274 25678 38276 25730
rect 37548 25454 37550 25506
rect 37602 25454 37604 25506
rect 37548 25442 37604 25454
rect 37996 25508 38052 25518
rect 37996 25414 38052 25452
rect 37436 25396 37492 25406
rect 37436 25302 37492 25340
rect 35196 24724 35252 24734
rect 34972 24722 35252 24724
rect 34972 24670 35198 24722
rect 35250 24670 35252 24722
rect 34972 24668 35252 24670
rect 34972 24164 35028 24174
rect 34860 24162 35028 24164
rect 34860 24110 34974 24162
rect 35026 24110 35028 24162
rect 34860 24108 35028 24110
rect 34972 24098 35028 24108
rect 34636 23940 34692 23950
rect 34524 23938 34692 23940
rect 34524 23886 34638 23938
rect 34690 23886 34692 23938
rect 34524 23884 34692 23886
rect 34636 23874 34692 23884
rect 34748 23940 34804 23950
rect 34412 23828 34468 23838
rect 34300 23156 34356 23166
rect 34188 23100 34300 23156
rect 34300 23090 34356 23100
rect 34412 23154 34468 23772
rect 34748 23268 34804 23884
rect 34748 23202 34804 23212
rect 34412 23102 34414 23154
rect 34466 23102 34468 23154
rect 34076 22754 34132 22764
rect 34412 22484 34468 23102
rect 34636 23156 34692 23166
rect 34636 23062 34692 23100
rect 34524 23044 34580 23054
rect 34524 22950 34580 22988
rect 35084 22484 35140 24668
rect 35196 24658 35252 24668
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 35196 24162 35252 24174
rect 35196 24110 35198 24162
rect 35250 24110 35252 24162
rect 35196 23714 35252 24110
rect 35532 23828 35588 24892
rect 35756 24836 35812 24846
rect 35756 24742 35812 24780
rect 36316 24836 36372 24846
rect 35644 24724 35700 24734
rect 35644 24630 35700 24668
rect 36316 24722 36372 24780
rect 37100 24836 37156 25228
rect 37100 24770 37156 24780
rect 37212 25282 37268 25294
rect 37212 25230 37214 25282
rect 37266 25230 37268 25282
rect 36316 24670 36318 24722
rect 36370 24670 36372 24722
rect 35980 24610 36036 24622
rect 35980 24558 35982 24610
rect 36034 24558 36036 24610
rect 35868 23940 35924 23950
rect 35980 23940 36036 24558
rect 35868 23938 36036 23940
rect 35868 23886 35870 23938
rect 35922 23886 36036 23938
rect 35868 23884 36036 23886
rect 35868 23874 35924 23884
rect 35532 23762 35588 23772
rect 35196 23662 35198 23714
rect 35250 23662 35252 23714
rect 35196 22932 35252 23662
rect 35980 23716 36036 23726
rect 36204 23716 36260 23726
rect 35980 23622 36036 23660
rect 36092 23714 36260 23716
rect 36092 23662 36206 23714
rect 36258 23662 36260 23714
rect 36092 23660 36260 23662
rect 35308 23604 35364 23614
rect 35308 23154 35364 23548
rect 35980 23268 36036 23278
rect 36092 23268 36148 23660
rect 36204 23650 36260 23660
rect 36316 23604 36372 24670
rect 37100 24610 37156 24622
rect 37100 24558 37102 24610
rect 37154 24558 37156 24610
rect 36988 24500 37044 24510
rect 36316 23538 36372 23548
rect 36428 24052 36484 24062
rect 35980 23266 36148 23268
rect 35980 23214 35982 23266
rect 36034 23214 36148 23266
rect 35980 23212 36148 23214
rect 35980 23202 36036 23212
rect 35308 23102 35310 23154
rect 35362 23102 35364 23154
rect 35308 23090 35364 23102
rect 35196 22866 35252 22876
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 34076 22428 34468 22484
rect 34076 22370 34132 22428
rect 34076 22318 34078 22370
rect 34130 22318 34132 22370
rect 34076 22306 34132 22318
rect 33852 22206 33854 22258
rect 33906 22206 33908 22258
rect 33852 22148 33908 22206
rect 33852 22082 33908 22092
rect 34188 22258 34244 22270
rect 34188 22206 34190 22258
rect 34242 22206 34244 22258
rect 34188 21924 34244 22206
rect 34412 22260 34468 22428
rect 34748 22428 35140 22484
rect 36204 22596 36260 22606
rect 34412 22194 34468 22204
rect 34524 22370 34580 22382
rect 34524 22318 34526 22370
rect 34578 22318 34580 22370
rect 34300 22148 34356 22158
rect 34300 22054 34356 22092
rect 34524 22036 34580 22318
rect 34524 21970 34580 21980
rect 33516 21756 33684 21812
rect 33740 21868 34244 21924
rect 33740 21810 33796 21868
rect 33740 21758 33742 21810
rect 33794 21758 33796 21810
rect 33516 21700 33572 21756
rect 33740 21746 33796 21758
rect 33516 21634 33572 21644
rect 33964 21586 34020 21598
rect 33964 21534 33966 21586
rect 34018 21534 34020 21586
rect 33852 21474 33908 21486
rect 33852 21422 33854 21474
rect 33906 21422 33908 21474
rect 33852 21028 33908 21422
rect 33628 20972 33908 21028
rect 33628 20914 33684 20972
rect 33628 20862 33630 20914
rect 33682 20862 33684 20914
rect 33628 20850 33684 20862
rect 33852 20244 33908 20254
rect 33964 20244 34020 21534
rect 34412 21588 34468 21598
rect 34412 21494 34468 21532
rect 33852 20242 34020 20244
rect 33852 20190 33854 20242
rect 33906 20190 34020 20242
rect 33852 20188 34020 20190
rect 33852 20178 33908 20188
rect 34412 20132 34468 20142
rect 33852 20018 33908 20030
rect 33852 19966 33854 20018
rect 33906 19966 33908 20018
rect 33628 19796 33684 19806
rect 33628 19702 33684 19740
rect 33852 19460 33908 19966
rect 34412 20018 34468 20076
rect 34412 19966 34414 20018
rect 34466 19966 34468 20018
rect 34412 19954 34468 19966
rect 33628 19404 33852 19460
rect 33628 19346 33684 19404
rect 33852 19394 33908 19404
rect 33628 19294 33630 19346
rect 33682 19294 33684 19346
rect 33628 19282 33684 19294
rect 32732 17726 32734 17778
rect 32786 17726 32788 17778
rect 32732 17714 32788 17726
rect 33292 18396 33460 18452
rect 33068 17668 33124 17678
rect 33068 17574 33124 17612
rect 33292 16322 33348 18396
rect 34524 18228 34580 18238
rect 34300 17778 34356 17790
rect 34300 17726 34302 17778
rect 34354 17726 34356 17778
rect 33516 17668 33572 17678
rect 33516 17574 33572 17612
rect 33292 16270 33294 16322
rect 33346 16270 33348 16322
rect 33292 16258 33348 16270
rect 34300 16100 34356 17726
rect 34524 17666 34580 18172
rect 34748 17892 34804 22428
rect 35196 22372 35252 22382
rect 35196 22278 35252 22316
rect 35980 22372 36036 22382
rect 36204 22372 36260 22540
rect 35980 22370 36260 22372
rect 35980 22318 35982 22370
rect 36034 22318 36206 22370
rect 36258 22318 36260 22370
rect 35980 22316 36260 22318
rect 35980 22306 36036 22316
rect 36204 22306 36260 22316
rect 34972 22260 35028 22270
rect 34972 22166 35028 22204
rect 36316 22260 36372 22270
rect 36428 22260 36484 23996
rect 36988 23938 37044 24444
rect 37100 24162 37156 24558
rect 37100 24110 37102 24162
rect 37154 24110 37156 24162
rect 37100 24098 37156 24110
rect 36988 23886 36990 23938
rect 37042 23886 37044 23938
rect 36988 23874 37044 23886
rect 37100 23828 37156 23838
rect 37212 23828 37268 25230
rect 38220 24164 38276 25678
rect 38332 25732 38388 25742
rect 38332 25508 38388 25676
rect 38444 25730 38500 26852
rect 38444 25678 38446 25730
rect 38498 25678 38500 25730
rect 38444 25618 38500 25678
rect 38444 25566 38446 25618
rect 38498 25566 38500 25618
rect 38444 25554 38500 25566
rect 39452 25620 39508 27804
rect 39900 27748 39956 27758
rect 39900 27654 39956 27692
rect 39900 27188 39956 27198
rect 40124 27188 40180 27916
rect 40348 27972 40404 28590
rect 41020 28644 41076 28654
rect 41020 28550 41076 28588
rect 41580 28642 41636 29932
rect 41804 29428 41860 31164
rect 42476 31108 42532 31118
rect 42476 31014 42532 31052
rect 42252 30994 42308 31006
rect 42252 30942 42254 30994
rect 42306 30942 42308 30994
rect 42252 30212 42308 30942
rect 42700 30996 42756 32732
rect 42812 32674 42868 32686
rect 42812 32622 42814 32674
rect 42866 32622 42868 32674
rect 42812 31220 42868 32622
rect 42924 32676 42980 32686
rect 42924 32582 42980 32620
rect 43708 32674 43764 33964
rect 43708 32622 43710 32674
rect 43762 32622 43764 32674
rect 43708 32610 43764 32622
rect 43820 34130 43876 34142
rect 43820 34078 43822 34130
rect 43874 34078 43876 34130
rect 43820 33570 43876 34078
rect 43820 33518 43822 33570
rect 43874 33518 43876 33570
rect 43820 32676 43876 33518
rect 43932 33572 43988 34300
rect 44492 34354 44548 34860
rect 45276 34914 45332 35196
rect 45724 35252 45780 35534
rect 45724 35186 45780 35196
rect 45276 34862 45278 34914
rect 45330 34862 45332 34914
rect 45276 34850 45332 34862
rect 45724 34916 45780 34926
rect 45724 34822 45780 34860
rect 44828 34804 44884 34814
rect 44492 34302 44494 34354
rect 44546 34302 44548 34354
rect 44492 34290 44548 34302
rect 44604 34802 44884 34804
rect 44604 34750 44830 34802
rect 44882 34750 44884 34802
rect 44604 34748 44884 34750
rect 44604 34242 44660 34748
rect 44828 34738 44884 34748
rect 46172 34802 46228 34814
rect 46172 34750 46174 34802
rect 46226 34750 46228 34802
rect 45388 34692 45444 34702
rect 44604 34190 44606 34242
rect 44658 34190 44660 34242
rect 44604 34178 44660 34190
rect 45164 34356 45220 34366
rect 44156 34132 44212 34142
rect 44156 34038 44212 34076
rect 44268 34130 44324 34142
rect 44268 34078 44270 34130
rect 44322 34078 44324 34130
rect 44268 34020 44324 34078
rect 44268 33954 44324 33964
rect 44716 34132 44772 34142
rect 43932 33346 43988 33516
rect 43932 33294 43934 33346
rect 43986 33294 43988 33346
rect 43932 33282 43988 33294
rect 43820 32562 43876 32620
rect 43820 32510 43822 32562
rect 43874 32510 43876 32562
rect 43820 32498 43876 32510
rect 43932 32900 43988 32910
rect 43932 32450 43988 32844
rect 44716 32562 44772 34076
rect 45164 33346 45220 34300
rect 45388 34130 45444 34636
rect 46172 34468 46228 34750
rect 46284 34692 46340 34702
rect 46284 34598 46340 34636
rect 46396 34468 46452 36092
rect 47292 35812 47348 36204
rect 48300 35924 48356 36990
rect 48412 36484 48468 36494
rect 48636 36484 48692 37996
rect 48748 37986 48804 37996
rect 48412 36482 48692 36484
rect 48412 36430 48414 36482
rect 48466 36430 48692 36482
rect 48412 36428 48692 36430
rect 48972 37154 49028 37166
rect 48972 37102 48974 37154
rect 49026 37102 49028 37154
rect 48412 36418 48468 36428
rect 48300 35868 48804 35924
rect 47180 35700 47236 35710
rect 47068 35252 47124 35262
rect 47068 34914 47124 35196
rect 47180 35028 47236 35644
rect 47180 34962 47236 34972
rect 47068 34862 47070 34914
rect 47122 34862 47124 34914
rect 47068 34850 47124 34862
rect 46508 34692 46564 34702
rect 47292 34692 47348 35756
rect 48076 35364 48132 35374
rect 46508 34598 46564 34636
rect 47068 34636 47348 34692
rect 47516 34692 47572 34702
rect 46172 34412 46452 34468
rect 46620 34580 46676 34590
rect 45612 34356 45668 34366
rect 45612 34262 45668 34300
rect 45388 34078 45390 34130
rect 45442 34078 45444 34130
rect 45388 34066 45444 34078
rect 45948 34132 46004 34142
rect 45948 34038 46004 34076
rect 45164 33294 45166 33346
rect 45218 33294 45220 33346
rect 45164 33282 45220 33294
rect 45836 33516 46228 33572
rect 44828 33236 44884 33246
rect 44828 33142 44884 33180
rect 45276 32900 45332 32910
rect 45164 32674 45220 32686
rect 45164 32622 45166 32674
rect 45218 32622 45220 32674
rect 44716 32510 44718 32562
rect 44770 32510 44772 32562
rect 44716 32498 44772 32510
rect 45052 32564 45108 32574
rect 43932 32398 43934 32450
rect 43986 32398 43988 32450
rect 43932 32386 43988 32398
rect 45052 31890 45108 32508
rect 45052 31838 45054 31890
rect 45106 31838 45108 31890
rect 45052 31826 45108 31838
rect 44940 31666 44996 31678
rect 44940 31614 44942 31666
rect 44994 31614 44996 31666
rect 44940 31332 44996 31614
rect 45164 31668 45220 32622
rect 45276 32562 45332 32844
rect 45276 32510 45278 32562
rect 45330 32510 45332 32562
rect 45276 32002 45332 32510
rect 45836 32564 45892 33516
rect 46172 33458 46228 33516
rect 46172 33406 46174 33458
rect 46226 33406 46228 33458
rect 46172 33394 46228 33406
rect 46284 33346 46340 34412
rect 46620 34130 46676 34524
rect 46620 34078 46622 34130
rect 46674 34078 46676 34130
rect 46620 34066 46676 34078
rect 46284 33294 46286 33346
rect 46338 33294 46340 33346
rect 46284 33282 46340 33294
rect 46060 33236 46116 33246
rect 45836 32470 45892 32508
rect 45948 33180 46060 33236
rect 45276 31950 45278 32002
rect 45330 31950 45332 32002
rect 45276 31938 45332 31950
rect 45500 32004 45556 32014
rect 45500 31778 45556 31948
rect 45500 31726 45502 31778
rect 45554 31726 45556 31778
rect 45500 31714 45556 31726
rect 45948 31892 46004 33180
rect 46060 33142 46116 33180
rect 46620 33124 46676 33134
rect 47068 33124 47124 34636
rect 47516 34242 47572 34636
rect 47516 34190 47518 34242
rect 47570 34190 47572 34242
rect 47516 34178 47572 34190
rect 48076 34018 48132 35308
rect 48524 34916 48580 34926
rect 48748 34916 48804 35868
rect 48972 35364 49028 37102
rect 48860 34916 48916 34926
rect 48748 34914 48916 34916
rect 48748 34862 48862 34914
rect 48914 34862 48916 34914
rect 48748 34860 48916 34862
rect 48524 34822 48580 34860
rect 48860 34850 48916 34860
rect 48972 34802 49028 35308
rect 49084 36370 49140 36382
rect 49084 36318 49086 36370
rect 49138 36318 49140 36370
rect 49084 34916 49140 36318
rect 49084 34850 49140 34860
rect 48972 34750 48974 34802
rect 49026 34750 49028 34802
rect 48972 34738 49028 34750
rect 48076 33966 48078 34018
rect 48130 33966 48132 34018
rect 47180 33348 47236 33358
rect 47516 33348 47572 33358
rect 47180 33346 47572 33348
rect 47180 33294 47182 33346
rect 47234 33294 47518 33346
rect 47570 33294 47572 33346
rect 47180 33292 47572 33294
rect 47180 33282 47236 33292
rect 47516 33282 47572 33292
rect 48076 33346 48132 33966
rect 48412 34580 48468 34590
rect 48412 33458 48468 34524
rect 49196 34242 49252 38668
rect 49644 36932 49700 38894
rect 49868 38722 49924 38734
rect 49868 38670 49870 38722
rect 49922 38670 49924 38722
rect 49868 37268 49924 38670
rect 49980 38724 50036 39566
rect 50204 39620 50260 39630
rect 51100 39620 51156 39678
rect 50204 39618 50372 39620
rect 50204 39566 50206 39618
rect 50258 39566 50372 39618
rect 50204 39564 50372 39566
rect 50204 39554 50260 39564
rect 50204 38724 50260 38734
rect 49980 38722 50260 38724
rect 49980 38670 50206 38722
rect 50258 38670 50260 38722
rect 49980 38668 50260 38670
rect 50204 38050 50260 38668
rect 50204 37998 50206 38050
rect 50258 37998 50260 38050
rect 50204 37986 50260 37998
rect 50092 37940 50148 37950
rect 50092 37828 50148 37884
rect 50316 37828 50372 39564
rect 51100 39554 51156 39564
rect 50540 39396 50596 39406
rect 50540 39394 51268 39396
rect 50540 39342 50542 39394
rect 50594 39342 51268 39394
rect 50540 39340 51268 39342
rect 50540 39330 50596 39340
rect 50556 39228 50820 39238
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50556 39162 50820 39172
rect 50876 38946 50932 38958
rect 50876 38894 50878 38946
rect 50930 38894 50932 38946
rect 50876 38612 50932 38894
rect 51100 38946 51156 38958
rect 51100 38894 51102 38946
rect 51154 38894 51156 38946
rect 51100 38836 51156 38894
rect 51100 38770 51156 38780
rect 50876 38546 50932 38556
rect 50092 37772 50372 37828
rect 50556 37660 50820 37670
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50556 37594 50820 37604
rect 49868 37202 49924 37212
rect 50092 37268 50148 37278
rect 50764 37268 50820 37278
rect 50092 37266 50260 37268
rect 50092 37214 50094 37266
rect 50146 37214 50260 37266
rect 50092 37212 50260 37214
rect 50092 37202 50148 37212
rect 49644 35698 49700 36876
rect 49644 35646 49646 35698
rect 49698 35646 49700 35698
rect 49644 35476 49700 35646
rect 49644 35410 49700 35420
rect 49756 36370 49812 36382
rect 49756 36318 49758 36370
rect 49810 36318 49812 36370
rect 49308 34692 49364 34702
rect 49308 34356 49364 34636
rect 49644 34690 49700 34702
rect 49644 34638 49646 34690
rect 49698 34638 49700 34690
rect 49644 34356 49700 34638
rect 49756 34580 49812 36318
rect 49868 35812 49924 35822
rect 49868 35028 49924 35756
rect 50204 35810 50260 37212
rect 50764 37174 50820 37212
rect 50204 35758 50206 35810
rect 50258 35758 50260 35810
rect 50204 35746 50260 35758
rect 50316 37042 50372 37054
rect 50316 36990 50318 37042
rect 50370 36990 50372 37042
rect 49868 34962 49924 34972
rect 49980 34916 50036 34926
rect 49980 34822 50036 34860
rect 49868 34692 49924 34702
rect 49868 34598 49924 34636
rect 49756 34514 49812 34524
rect 49644 34300 50036 34356
rect 49308 34262 49364 34300
rect 49196 34190 49198 34242
rect 49250 34190 49252 34242
rect 49196 34178 49252 34190
rect 48412 33406 48414 33458
rect 48466 33406 48468 33458
rect 48412 33394 48468 33406
rect 49532 34130 49588 34142
rect 49532 34078 49534 34130
rect 49586 34078 49588 34130
rect 48076 33294 48078 33346
rect 48130 33294 48132 33346
rect 48076 33282 48132 33294
rect 49532 33236 49588 34078
rect 49868 34132 49924 34142
rect 49308 33124 49364 33134
rect 47068 33068 47236 33124
rect 46620 32562 46676 33068
rect 46620 32510 46622 32562
rect 46674 32510 46676 32562
rect 46620 32004 46676 32510
rect 46620 31938 46676 31948
rect 46732 32676 46788 32686
rect 45948 31836 46564 31892
rect 45164 31602 45220 31612
rect 45948 31666 46004 31836
rect 45948 31614 45950 31666
rect 46002 31614 46004 31666
rect 45948 31602 46004 31614
rect 46060 31668 46116 31678
rect 46060 31574 46116 31612
rect 46508 31666 46564 31836
rect 46620 31780 46676 31790
rect 46732 31780 46788 32620
rect 46620 31778 46788 31780
rect 46620 31726 46622 31778
rect 46674 31726 46788 31778
rect 46620 31724 46788 31726
rect 46620 31714 46676 31724
rect 46508 31614 46510 31666
rect 46562 31614 46564 31666
rect 46508 31602 46564 31614
rect 47068 31668 47124 31678
rect 47068 31574 47124 31612
rect 47180 31666 47236 33068
rect 49308 33030 49364 33068
rect 49308 32900 49364 32910
rect 47964 31892 48020 31902
rect 47964 31798 48020 31836
rect 48300 31892 48356 31902
rect 48972 31892 49252 31948
rect 47180 31614 47182 31666
rect 47234 31614 47236 31666
rect 47180 31602 47236 31614
rect 48188 31778 48244 31790
rect 48188 31726 48190 31778
rect 48242 31726 48244 31778
rect 44940 31266 44996 31276
rect 45724 31554 45780 31566
rect 46284 31556 46340 31566
rect 45724 31502 45726 31554
rect 45778 31502 45780 31554
rect 42812 31164 42980 31220
rect 42812 30996 42868 31006
rect 42700 30994 42868 30996
rect 42700 30942 42814 30994
rect 42866 30942 42868 30994
rect 42700 30940 42868 30942
rect 42252 30146 42308 30156
rect 42364 30882 42420 30894
rect 42364 30830 42366 30882
rect 42418 30830 42420 30882
rect 41916 29876 41972 29886
rect 41916 29652 41972 29820
rect 42364 29652 42420 30830
rect 42700 30322 42756 30940
rect 42812 30930 42868 30940
rect 42700 30270 42702 30322
rect 42754 30270 42756 30322
rect 42700 30258 42756 30270
rect 42812 30772 42868 30782
rect 41916 29596 42084 29652
rect 42028 29538 42084 29596
rect 42028 29486 42030 29538
rect 42082 29486 42084 29538
rect 42028 29474 42084 29486
rect 42140 29596 42756 29652
rect 41916 29428 41972 29438
rect 41804 29426 41972 29428
rect 41804 29374 41918 29426
rect 41970 29374 41972 29426
rect 41804 29372 41972 29374
rect 41916 29362 41972 29372
rect 42140 29204 42196 29596
rect 42700 29538 42756 29596
rect 42700 29486 42702 29538
rect 42754 29486 42756 29538
rect 42700 29474 42756 29486
rect 42812 29426 42868 30716
rect 42924 30100 42980 31164
rect 42924 30034 42980 30044
rect 43148 31106 43204 31118
rect 43148 31054 43150 31106
rect 43202 31054 43204 31106
rect 43036 29988 43092 29998
rect 43036 29894 43092 29932
rect 43148 29876 43204 31054
rect 43596 31108 43652 31118
rect 43372 30322 43428 30334
rect 43372 30270 43374 30322
rect 43426 30270 43428 30322
rect 43372 30212 43428 30270
rect 43596 30322 43652 31052
rect 44492 31108 44548 31118
rect 45724 31108 45780 31502
rect 46172 31554 46340 31556
rect 46172 31502 46286 31554
rect 46338 31502 46340 31554
rect 46172 31500 46340 31502
rect 45836 31108 45892 31118
rect 44492 31014 44548 31052
rect 45388 31106 45892 31108
rect 45388 31054 45838 31106
rect 45890 31054 45892 31106
rect 45388 31052 45892 31054
rect 44380 30996 44436 31006
rect 44268 30994 44436 30996
rect 44268 30942 44382 30994
rect 44434 30942 44436 30994
rect 44268 30940 44436 30942
rect 43596 30270 43598 30322
rect 43650 30270 43652 30322
rect 43596 30258 43652 30270
rect 43932 30324 43988 30334
rect 43932 30230 43988 30268
rect 43372 30146 43428 30156
rect 44268 30212 44324 30940
rect 44380 30930 44436 30940
rect 44604 30996 44660 31006
rect 44604 30994 44772 30996
rect 44604 30942 44606 30994
rect 44658 30942 44772 30994
rect 44604 30940 44772 30942
rect 44604 30930 44660 30940
rect 44268 30118 44324 30156
rect 44604 30100 44660 30110
rect 44044 29988 44100 29998
rect 44044 29894 44100 29932
rect 43148 29810 43204 29820
rect 44604 29538 44660 30044
rect 44716 29988 44772 30940
rect 44716 29922 44772 29932
rect 45052 30994 45108 31006
rect 45052 30942 45054 30994
rect 45106 30942 45108 30994
rect 45052 29652 45108 30942
rect 45276 30772 45332 30782
rect 45276 30678 45332 30716
rect 45388 30548 45444 31052
rect 45836 31042 45892 31052
rect 45612 30772 45668 30782
rect 45276 30492 45444 30548
rect 45500 30716 45612 30772
rect 45164 30434 45220 30446
rect 45164 30382 45166 30434
rect 45218 30382 45220 30434
rect 45164 30212 45220 30382
rect 45164 30146 45220 30156
rect 45052 29586 45108 29596
rect 44604 29486 44606 29538
rect 44658 29486 44660 29538
rect 44604 29474 44660 29486
rect 42812 29374 42814 29426
rect 42866 29374 42868 29426
rect 42812 29362 42868 29374
rect 44492 29428 44548 29438
rect 41580 28590 41582 28642
rect 41634 28590 41636 28642
rect 41580 28578 41636 28590
rect 41804 29148 42196 29204
rect 41804 28530 41860 29148
rect 42252 28644 42308 28654
rect 41804 28478 41806 28530
rect 41858 28478 41860 28530
rect 41804 28466 41860 28478
rect 41916 28642 42308 28644
rect 41916 28590 42254 28642
rect 42306 28590 42308 28642
rect 41916 28588 42308 28590
rect 40796 28420 40852 28430
rect 41692 28420 41748 28430
rect 40796 28418 40964 28420
rect 40796 28366 40798 28418
rect 40850 28366 40964 28418
rect 40796 28364 40964 28366
rect 40796 28354 40852 28364
rect 40348 27906 40404 27916
rect 39900 27186 40180 27188
rect 39900 27134 39902 27186
rect 39954 27134 40180 27186
rect 39900 27132 40180 27134
rect 40460 27858 40516 27870
rect 40460 27806 40462 27858
rect 40514 27806 40516 27858
rect 39900 25844 39956 27132
rect 40348 27074 40404 27086
rect 40348 27022 40350 27074
rect 40402 27022 40404 27074
rect 40348 26740 40404 27022
rect 40460 26908 40516 27806
rect 40908 27858 40964 28364
rect 41692 28326 41748 28364
rect 41916 28084 41972 28588
rect 42252 28578 42308 28588
rect 42700 28644 42756 28654
rect 42924 28644 42980 28654
rect 42700 28642 42980 28644
rect 42700 28590 42702 28642
rect 42754 28590 42926 28642
rect 42978 28590 42980 28642
rect 42700 28588 42980 28590
rect 42700 28578 42756 28588
rect 42924 28578 42980 28588
rect 43708 28642 43764 28654
rect 43708 28590 43710 28642
rect 43762 28590 43764 28642
rect 43148 28532 43204 28542
rect 43148 28438 43204 28476
rect 43260 28532 43316 28542
rect 43708 28532 43764 28590
rect 43260 28530 43764 28532
rect 43260 28478 43262 28530
rect 43314 28478 43764 28530
rect 43260 28476 43764 28478
rect 43820 28532 43876 28542
rect 42140 28418 42196 28430
rect 42140 28366 42142 28418
rect 42194 28366 42196 28418
rect 42140 28308 42196 28366
rect 42364 28420 42420 28430
rect 42364 28326 42420 28364
rect 42140 28242 42196 28252
rect 41692 28028 41972 28084
rect 41692 27970 41748 28028
rect 41692 27918 41694 27970
rect 41746 27918 41748 27970
rect 41692 27906 41748 27918
rect 40908 27806 40910 27858
rect 40962 27806 40964 27858
rect 40908 26908 40964 27806
rect 41020 27748 41076 27758
rect 41020 27186 41076 27692
rect 41020 27134 41022 27186
rect 41074 27134 41076 27186
rect 41020 27122 41076 27134
rect 41916 27636 41972 27646
rect 40460 26852 40852 26908
rect 40908 26852 41076 26908
rect 40348 26674 40404 26684
rect 40796 26066 40852 26852
rect 40796 26014 40798 26066
rect 40850 26014 40852 26066
rect 40796 26002 40852 26014
rect 41020 26740 41076 26852
rect 41020 26178 41076 26684
rect 41804 26516 41860 26526
rect 41804 26422 41860 26460
rect 41916 26516 41972 27580
rect 43260 27636 43316 28476
rect 43820 27746 43876 28476
rect 44492 27970 44548 29372
rect 45276 29426 45332 30492
rect 45276 29374 45278 29426
rect 45330 29374 45332 29426
rect 45276 29362 45332 29374
rect 45500 29426 45556 30716
rect 45612 30678 45668 30716
rect 46172 30436 46228 31500
rect 46284 31490 46340 31500
rect 46844 31556 46900 31566
rect 46844 31106 46900 31500
rect 47404 31556 47460 31566
rect 47628 31556 47684 31566
rect 47404 31554 47572 31556
rect 47404 31502 47406 31554
rect 47458 31502 47572 31554
rect 47404 31500 47572 31502
rect 47404 31490 47460 31500
rect 46844 31054 46846 31106
rect 46898 31054 46900 31106
rect 46844 31042 46900 31054
rect 47516 31332 47572 31500
rect 47628 31462 47684 31500
rect 48188 31332 48244 31726
rect 47516 31276 48244 31332
rect 46284 30994 46340 31006
rect 46284 30942 46286 30994
rect 46338 30942 46340 30994
rect 46284 30884 46340 30942
rect 46620 30994 46676 31006
rect 46620 30942 46622 30994
rect 46674 30942 46676 30994
rect 46284 30818 46340 30828
rect 46396 30882 46452 30894
rect 46396 30830 46398 30882
rect 46450 30830 46452 30882
rect 46396 30772 46452 30830
rect 46396 30706 46452 30716
rect 46620 30772 46676 30942
rect 47516 30996 47572 31276
rect 48300 31220 48356 31836
rect 48860 31836 49028 31892
rect 49196 31890 49252 31892
rect 49196 31838 49198 31890
rect 49250 31838 49252 31890
rect 48076 31164 48356 31220
rect 48748 31778 48804 31790
rect 48748 31726 48750 31778
rect 48802 31726 48804 31778
rect 48748 31220 48804 31726
rect 47628 30996 47684 31006
rect 47516 30994 47684 30996
rect 47516 30942 47630 30994
rect 47682 30942 47684 30994
rect 47516 30940 47684 30942
rect 47628 30930 47684 30940
rect 48076 30994 48132 31164
rect 48748 31106 48804 31164
rect 48748 31054 48750 31106
rect 48802 31054 48804 31106
rect 48748 31042 48804 31054
rect 48076 30942 48078 30994
rect 48130 30942 48132 30994
rect 48076 30930 48132 30942
rect 48860 30996 48916 31836
rect 49196 31826 49252 31838
rect 49084 31780 49140 31790
rect 48972 31724 49084 31780
rect 48972 31218 49028 31724
rect 49084 31686 49140 31724
rect 48972 31166 48974 31218
rect 49026 31166 49028 31218
rect 48972 31154 49028 31166
rect 49308 31218 49364 32844
rect 49532 32788 49588 33180
rect 49756 34018 49812 34030
rect 49756 33966 49758 34018
rect 49810 33966 49812 34018
rect 49644 32788 49700 32798
rect 49532 32786 49700 32788
rect 49532 32734 49646 32786
rect 49698 32734 49700 32786
rect 49532 32732 49700 32734
rect 49644 32722 49700 32732
rect 49756 32674 49812 33966
rect 49868 33346 49924 34076
rect 49868 33294 49870 33346
rect 49922 33294 49924 33346
rect 49868 33282 49924 33294
rect 49756 32622 49758 32674
rect 49810 32622 49812 32674
rect 49756 32610 49812 32622
rect 49644 32338 49700 32350
rect 49644 32286 49646 32338
rect 49698 32286 49700 32338
rect 49644 31668 49700 32286
rect 49980 31948 50036 34300
rect 50316 34244 50372 36990
rect 50540 36708 50596 36718
rect 50540 36484 50596 36652
rect 50428 36482 50596 36484
rect 50428 36430 50542 36482
rect 50594 36430 50596 36482
rect 50428 36428 50596 36430
rect 50428 35810 50484 36428
rect 50540 36418 50596 36428
rect 51212 36484 51268 39340
rect 51324 38834 51380 40238
rect 51884 40180 51940 41692
rect 52668 41524 52724 41534
rect 51996 40964 52052 40974
rect 51996 40870 52052 40908
rect 51772 40124 51940 40180
rect 51996 40516 52052 40526
rect 51548 39620 51604 39630
rect 51772 39620 51828 40124
rect 51548 39618 51828 39620
rect 51548 39566 51550 39618
rect 51602 39566 51828 39618
rect 51548 39564 51828 39566
rect 51548 39554 51604 39564
rect 51884 39508 51940 39518
rect 51884 39414 51940 39452
rect 51996 39506 52052 40460
rect 52220 40516 52276 40526
rect 52220 39618 52276 40460
rect 52220 39566 52222 39618
rect 52274 39566 52276 39618
rect 52220 39554 52276 39566
rect 52668 39618 52724 41468
rect 52668 39566 52670 39618
rect 52722 39566 52724 39618
rect 52668 39554 52724 39566
rect 51996 39454 51998 39506
rect 52050 39454 52052 39506
rect 51996 39060 52052 39454
rect 52332 39508 52388 39518
rect 51996 38994 52052 39004
rect 52220 39172 52276 39182
rect 51324 38782 51326 38834
rect 51378 38782 51380 38834
rect 51324 38770 51380 38782
rect 51884 38722 51940 38734
rect 51884 38670 51886 38722
rect 51938 38670 51940 38722
rect 51884 38612 51940 38670
rect 52220 38668 52276 39116
rect 51884 38546 51940 38556
rect 51996 38612 52276 38668
rect 51996 38050 52052 38612
rect 51996 37998 51998 38050
rect 52050 37998 52052 38050
rect 51996 37986 52052 37998
rect 51884 37828 51940 37838
rect 51884 37826 52276 37828
rect 51884 37774 51886 37826
rect 51938 37774 52276 37826
rect 51884 37772 52276 37774
rect 51884 37762 51940 37772
rect 51548 37268 51604 37278
rect 51436 36484 51492 36494
rect 51212 36482 51436 36484
rect 51212 36430 51214 36482
rect 51266 36430 51436 36482
rect 51212 36428 51436 36430
rect 51212 36418 51268 36428
rect 50556 36092 50820 36102
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50556 36026 50820 36036
rect 50428 35758 50430 35810
rect 50482 35758 50484 35810
rect 50428 35746 50484 35758
rect 51436 35700 51492 36428
rect 51548 36484 51604 37212
rect 52220 37154 52276 37772
rect 52220 37102 52222 37154
rect 52274 37102 52276 37154
rect 52220 37044 52276 37102
rect 52220 36978 52276 36988
rect 51548 36482 51828 36484
rect 51548 36430 51550 36482
rect 51602 36430 51828 36482
rect 51548 36428 51828 36430
rect 51548 36418 51604 36428
rect 51772 35810 51828 36428
rect 52332 36036 52388 39452
rect 52444 39060 52500 39070
rect 52444 38966 52500 39004
rect 52780 39058 52836 41692
rect 52892 41682 52948 41692
rect 53004 40628 53060 42478
rect 54124 41188 54180 42700
rect 54348 42084 54404 42094
rect 54348 41990 54404 42028
rect 54236 41970 54292 41982
rect 54236 41918 54238 41970
rect 54290 41918 54292 41970
rect 54236 41860 54292 41918
rect 54236 41794 54292 41804
rect 54236 41188 54292 41198
rect 54124 41186 54292 41188
rect 54124 41134 54238 41186
rect 54290 41134 54292 41186
rect 54124 41132 54292 41134
rect 53004 40562 53060 40572
rect 53116 41074 53172 41086
rect 53116 41022 53118 41074
rect 53170 41022 53172 41074
rect 53004 39508 53060 39518
rect 53004 39414 53060 39452
rect 53116 39172 53172 41022
rect 54124 40628 54180 40638
rect 53228 40516 53284 40526
rect 53228 40402 53284 40460
rect 53228 40350 53230 40402
rect 53282 40350 53284 40402
rect 53228 40338 53284 40350
rect 53340 40404 53396 40414
rect 53340 40290 53396 40348
rect 54012 40404 54068 40414
rect 54012 40310 54068 40348
rect 53340 40238 53342 40290
rect 53394 40238 53396 40290
rect 53340 40226 53396 40238
rect 53676 40290 53732 40302
rect 53676 40238 53678 40290
rect 53730 40238 53732 40290
rect 52780 39006 52782 39058
rect 52834 39006 52836 39058
rect 52780 38994 52836 39006
rect 53004 39116 53116 39172
rect 52668 37266 52724 37278
rect 52668 37214 52670 37266
rect 52722 37214 52724 37266
rect 52668 36706 52724 37214
rect 52668 36654 52670 36706
rect 52722 36654 52724 36706
rect 52668 36642 52724 36654
rect 53004 36708 53060 39116
rect 53116 39106 53172 39116
rect 53452 39620 53508 39630
rect 53116 38948 53172 38958
rect 53116 38946 53396 38948
rect 53116 38894 53118 38946
rect 53170 38894 53396 38946
rect 53116 38892 53396 38894
rect 53116 38882 53172 38892
rect 53004 36614 53060 36652
rect 53228 36484 53284 36494
rect 53228 36390 53284 36428
rect 51772 35758 51774 35810
rect 51826 35758 51828 35810
rect 51772 35746 51828 35758
rect 52108 35980 52388 36036
rect 51548 35700 51604 35710
rect 52108 35700 52164 35980
rect 51436 35698 51604 35700
rect 51436 35646 51550 35698
rect 51602 35646 51604 35698
rect 51436 35644 51604 35646
rect 51548 35634 51604 35644
rect 51884 35644 52164 35700
rect 52332 35812 52388 35822
rect 51884 34916 51940 35644
rect 51884 34822 51940 34860
rect 51996 35476 52052 35486
rect 51996 34802 52052 35420
rect 51996 34750 51998 34802
rect 52050 34750 52052 34802
rect 51996 34738 52052 34750
rect 52108 35028 52164 35038
rect 50556 34524 50820 34534
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50556 34458 50820 34468
rect 50316 34130 50372 34188
rect 51324 34244 51380 34254
rect 50316 34078 50318 34130
rect 50370 34078 50372 34130
rect 50316 34066 50372 34078
rect 50652 34132 50708 34142
rect 50652 34038 50708 34076
rect 51324 33458 51380 34188
rect 51996 34244 52052 34282
rect 51996 34178 52052 34188
rect 51324 33406 51326 33458
rect 51378 33406 51380 33458
rect 51324 33394 51380 33406
rect 51548 33684 51604 33694
rect 50764 33236 50820 33246
rect 50764 33142 50820 33180
rect 50556 32956 50820 32966
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50556 32890 50820 32900
rect 51548 32674 51604 33628
rect 51660 33124 51716 33134
rect 51660 32786 51716 33068
rect 51660 32734 51662 32786
rect 51714 32734 51716 32786
rect 51660 32722 51716 32734
rect 52108 32788 52164 34972
rect 52220 34916 52276 34926
rect 52332 34916 52388 35756
rect 53116 35476 53172 35486
rect 52220 34914 52388 34916
rect 52220 34862 52222 34914
rect 52274 34862 52388 34914
rect 52220 34860 52388 34862
rect 52444 35474 53172 35476
rect 52444 35422 53118 35474
rect 53170 35422 53172 35474
rect 52444 35420 53172 35422
rect 52220 34850 52276 34860
rect 52444 34132 52500 35420
rect 53116 35410 53172 35420
rect 53340 35252 53396 38892
rect 53452 38836 53508 39564
rect 53564 39060 53620 39070
rect 53564 38966 53620 39004
rect 53452 38834 53620 38836
rect 53452 38782 53454 38834
rect 53506 38782 53620 38834
rect 53452 38780 53620 38782
rect 53452 38770 53508 38780
rect 53228 35196 53396 35252
rect 53452 38612 53508 38622
rect 52668 35028 52724 35038
rect 52668 34934 52724 34972
rect 52780 34916 52836 34926
rect 52780 34802 52836 34860
rect 53004 34804 53060 34814
rect 52780 34750 52782 34802
rect 52834 34750 52836 34802
rect 52780 34738 52836 34750
rect 52892 34802 53060 34804
rect 52892 34750 53006 34802
rect 53058 34750 53060 34802
rect 52892 34748 53060 34750
rect 52780 34354 52836 34366
rect 52780 34302 52782 34354
rect 52834 34302 52836 34354
rect 52444 34038 52500 34076
rect 52668 34244 52724 34254
rect 52332 33236 52388 33246
rect 52220 32788 52276 32798
rect 52108 32786 52276 32788
rect 52108 32734 52222 32786
rect 52274 32734 52276 32786
rect 52108 32732 52276 32734
rect 52220 32722 52276 32732
rect 51548 32622 51550 32674
rect 51602 32622 51604 32674
rect 51548 32610 51604 32622
rect 51884 32564 51940 32574
rect 52108 32564 52164 32574
rect 52332 32564 52388 33180
rect 52668 32676 52724 34188
rect 52556 32674 52724 32676
rect 52556 32622 52670 32674
rect 52722 32622 52724 32674
rect 52556 32620 52724 32622
rect 52780 32676 52836 34302
rect 52892 33684 52948 34748
rect 53004 34738 53060 34748
rect 53116 34692 53172 34702
rect 53004 34132 53060 34142
rect 53116 34132 53172 34636
rect 53228 34468 53284 35196
rect 53452 35140 53508 38556
rect 53340 35084 53508 35140
rect 53340 34580 53396 35084
rect 53452 34916 53508 34926
rect 53452 34822 53508 34860
rect 53340 34524 53508 34580
rect 53228 34412 53396 34468
rect 53340 34244 53396 34412
rect 53340 34150 53396 34188
rect 53452 34354 53508 34524
rect 53452 34302 53454 34354
rect 53506 34302 53508 34354
rect 53004 34130 53172 34132
rect 53004 34078 53006 34130
rect 53058 34078 53172 34130
rect 53004 34076 53172 34078
rect 53004 34066 53060 34076
rect 53452 33908 53508 34302
rect 53116 33852 53508 33908
rect 53004 33684 53060 33694
rect 52892 33628 53004 33684
rect 53004 33618 53060 33628
rect 53116 33236 53172 33852
rect 53004 33234 53172 33236
rect 53004 33182 53118 33234
rect 53170 33182 53172 33234
rect 53004 33180 53172 33182
rect 52780 32620 52948 32676
rect 51884 32562 52052 32564
rect 51884 32510 51886 32562
rect 51938 32510 52052 32562
rect 51884 32508 52052 32510
rect 51884 32498 51940 32508
rect 49868 31892 50036 31948
rect 51548 31892 51604 31902
rect 49532 31666 49700 31668
rect 49532 31614 49646 31666
rect 49698 31614 49700 31666
rect 49532 31612 49700 31614
rect 49532 31444 49588 31612
rect 49644 31602 49700 31612
rect 49756 31780 49812 31790
rect 49308 31166 49310 31218
rect 49362 31166 49364 31218
rect 49308 31154 49364 31166
rect 49420 31388 49588 31444
rect 49756 31444 49812 31724
rect 49196 31106 49252 31118
rect 49196 31054 49198 31106
rect 49250 31054 49252 31106
rect 49196 30996 49252 31054
rect 49420 30996 49476 31388
rect 49756 31378 49812 31388
rect 49532 31220 49588 31230
rect 49532 31106 49588 31164
rect 49532 31054 49534 31106
rect 49586 31054 49588 31106
rect 49532 31042 49588 31054
rect 49868 31108 49924 31892
rect 51548 31798 51604 31836
rect 51996 31892 52052 32508
rect 52164 32508 52388 32564
rect 52444 32562 52500 32574
rect 52444 32510 52446 32562
rect 52498 32510 52500 32562
rect 52108 32470 52164 32508
rect 52332 32004 52388 32014
rect 51996 31826 52052 31836
rect 52108 31948 52332 32004
rect 52108 31890 52164 31948
rect 52332 31938 52388 31948
rect 52108 31838 52110 31890
rect 52162 31838 52164 31890
rect 52108 31826 52164 31838
rect 51884 31778 51940 31790
rect 51884 31726 51886 31778
rect 51938 31726 51940 31778
rect 48860 30940 49028 30996
rect 49196 30940 49476 30996
rect 46620 30706 46676 30716
rect 47180 30884 47236 30894
rect 45724 30380 46228 30436
rect 45612 30322 45668 30334
rect 45612 30270 45614 30322
rect 45666 30270 45668 30322
rect 45612 29876 45668 30270
rect 45724 30210 45780 30380
rect 45724 30158 45726 30210
rect 45778 30158 45780 30210
rect 45724 30146 45780 30158
rect 45612 29810 45668 29820
rect 45836 29652 45892 29662
rect 45836 29558 45892 29596
rect 46060 29650 46116 30380
rect 46284 30212 46340 30222
rect 46284 30118 46340 30156
rect 47180 30210 47236 30828
rect 47180 30158 47182 30210
rect 47234 30158 47236 30210
rect 47180 30146 47236 30158
rect 47740 30772 47796 30782
rect 47740 30210 47796 30716
rect 47740 30158 47742 30210
rect 47794 30158 47796 30210
rect 47740 30146 47796 30158
rect 48972 30660 49028 30940
rect 48972 30210 49028 30604
rect 48972 30158 48974 30210
rect 49026 30158 49028 30210
rect 48972 30146 49028 30158
rect 47068 30098 47124 30110
rect 47068 30046 47070 30098
rect 47122 30046 47124 30098
rect 46396 29988 46452 29998
rect 46396 29894 46452 29932
rect 46620 29986 46676 29998
rect 46620 29934 46622 29986
rect 46674 29934 46676 29986
rect 46060 29598 46062 29650
rect 46114 29598 46116 29650
rect 46060 29586 46116 29598
rect 46172 29876 46228 29886
rect 46172 29538 46228 29820
rect 46172 29486 46174 29538
rect 46226 29486 46228 29538
rect 46172 29474 46228 29486
rect 46620 29540 46676 29934
rect 47068 29876 47124 30046
rect 49868 30098 49924 31052
rect 50204 31556 50260 31566
rect 50204 30994 50260 31500
rect 50556 31388 50820 31398
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50556 31322 50820 31332
rect 51100 31108 51156 31118
rect 51100 31014 51156 31052
rect 51884 31108 51940 31726
rect 52444 31220 52500 32510
rect 52556 31668 52612 32620
rect 52668 32610 52724 32620
rect 52780 32450 52836 32462
rect 52780 32398 52782 32450
rect 52834 32398 52836 32450
rect 52780 32004 52836 32398
rect 52780 31938 52836 31948
rect 52892 31780 52948 32620
rect 53004 32674 53060 33180
rect 53116 33170 53172 33180
rect 53564 33236 53620 38780
rect 53676 37380 53732 40238
rect 54124 39618 54180 40572
rect 54236 40402 54292 41132
rect 54236 40350 54238 40402
rect 54290 40350 54292 40402
rect 54236 40338 54292 40350
rect 54124 39566 54126 39618
rect 54178 39566 54180 39618
rect 54124 39554 54180 39566
rect 54460 38948 54516 42924
rect 54572 39732 54628 43148
rect 54684 42756 54740 43262
rect 55356 43316 55412 43326
rect 55356 43222 55412 43260
rect 54684 42690 54740 42700
rect 55244 42754 55300 42766
rect 55244 42702 55246 42754
rect 55298 42702 55300 42754
rect 54908 42196 54964 42206
rect 54908 41858 54964 42140
rect 54908 41806 54910 41858
rect 54962 41806 54964 41858
rect 54908 41794 54964 41806
rect 55244 41186 55300 42702
rect 55692 42754 55748 43652
rect 57148 43316 57204 43326
rect 57148 42866 57204 43260
rect 57148 42814 57150 42866
rect 57202 42814 57204 42866
rect 57148 42802 57204 42814
rect 55692 42702 55694 42754
rect 55746 42702 55748 42754
rect 55692 42196 55748 42702
rect 56700 42756 56756 42766
rect 56700 42662 56756 42700
rect 55692 42130 55748 42140
rect 55244 41134 55246 41186
rect 55298 41134 55300 41186
rect 54684 40964 54740 40974
rect 54684 40402 54740 40908
rect 55244 40964 55300 41134
rect 55244 40898 55300 40908
rect 55468 41074 55524 41086
rect 55468 41022 55470 41074
rect 55522 41022 55524 41074
rect 54684 40350 54686 40402
rect 54738 40350 54740 40402
rect 54684 40338 54740 40350
rect 55132 40628 55188 40638
rect 54572 39676 55076 39732
rect 54572 39618 54628 39676
rect 54572 39566 54574 39618
rect 54626 39566 54628 39618
rect 54572 39554 54628 39566
rect 54236 38946 54516 38948
rect 54236 38894 54462 38946
rect 54514 38894 54516 38946
rect 54236 38892 54516 38894
rect 53788 38834 53844 38846
rect 53788 38782 53790 38834
rect 53842 38782 53844 38834
rect 53788 38050 53844 38782
rect 54236 38668 54292 38892
rect 54460 38882 54516 38892
rect 54796 39506 54852 39518
rect 54796 39454 54798 39506
rect 54850 39454 54852 39506
rect 54796 38834 54852 39454
rect 55020 39508 55076 39676
rect 55132 39730 55188 40572
rect 55468 40516 55524 41022
rect 55468 40450 55524 40460
rect 55132 39678 55134 39730
rect 55186 39678 55188 39730
rect 55132 39666 55188 39678
rect 55356 39618 55412 39630
rect 55356 39566 55358 39618
rect 55410 39566 55412 39618
rect 55356 39508 55412 39566
rect 55020 39452 55412 39508
rect 55692 39396 55748 39406
rect 54796 38782 54798 38834
rect 54850 38782 54852 38834
rect 54684 38722 54740 38734
rect 54684 38670 54686 38722
rect 54738 38670 54740 38722
rect 54236 38612 54516 38668
rect 53788 37998 53790 38050
rect 53842 37998 53844 38050
rect 53788 37986 53844 37998
rect 54460 38050 54516 38612
rect 54460 37998 54462 38050
rect 54514 37998 54516 38050
rect 53676 37324 54292 37380
rect 54236 37268 54292 37324
rect 53900 37156 53956 37166
rect 53900 37154 54068 37156
rect 53900 37102 53902 37154
rect 53954 37102 54068 37154
rect 53900 37100 54068 37102
rect 53900 37090 53956 37100
rect 53900 34916 53956 34926
rect 53900 34822 53956 34860
rect 53676 34692 53732 34702
rect 54012 34692 54068 37100
rect 54124 37044 54180 37054
rect 54124 36594 54180 36988
rect 54124 36542 54126 36594
rect 54178 36542 54180 36594
rect 54124 36530 54180 36542
rect 54236 36482 54292 37212
rect 54460 37266 54516 37998
rect 54460 37214 54462 37266
rect 54514 37214 54516 37266
rect 54460 37202 54516 37214
rect 54572 37044 54628 37054
rect 54236 36430 54238 36482
rect 54290 36430 54292 36482
rect 53676 34598 53732 34636
rect 53788 34636 54068 34692
rect 54124 36370 54180 36382
rect 54124 36318 54126 36370
rect 54178 36318 54180 36370
rect 53676 34130 53732 34142
rect 53676 34078 53678 34130
rect 53730 34078 53732 34130
rect 53676 33348 53732 34078
rect 53676 33282 53732 33292
rect 53788 33346 53844 34636
rect 54124 33684 54180 36318
rect 54236 34692 54292 36430
rect 54460 36484 54516 36494
rect 54460 35700 54516 36428
rect 54348 35698 54516 35700
rect 54348 35646 54462 35698
rect 54514 35646 54516 35698
rect 54348 35644 54516 35646
rect 54348 35138 54404 35644
rect 54460 35634 54516 35644
rect 54348 35086 54350 35138
rect 54402 35086 54404 35138
rect 54348 35074 54404 35086
rect 54572 35138 54628 36988
rect 54684 35812 54740 38670
rect 54796 37268 54852 38782
rect 55468 39394 55748 39396
rect 55468 39342 55694 39394
rect 55746 39342 55748 39394
rect 55468 39340 55748 39342
rect 55468 38834 55524 39340
rect 55692 39330 55748 39340
rect 55468 38782 55470 38834
rect 55522 38782 55524 38834
rect 55468 38770 55524 38782
rect 55580 38274 55636 38286
rect 55580 38222 55582 38274
rect 55634 38222 55636 38274
rect 55132 38050 55188 38062
rect 55132 37998 55134 38050
rect 55186 37998 55188 38050
rect 55132 37268 55188 37998
rect 55468 37378 55524 37390
rect 55468 37326 55470 37378
rect 55522 37326 55524 37378
rect 54796 37266 55188 37268
rect 54796 37214 54798 37266
rect 54850 37214 55188 37266
rect 54796 37212 55188 37214
rect 55244 37266 55300 37278
rect 55244 37214 55246 37266
rect 55298 37214 55300 37266
rect 54796 37202 54852 37212
rect 55244 37044 55300 37214
rect 55468 37268 55524 37326
rect 55468 37202 55524 37212
rect 55244 36978 55300 36988
rect 55356 37154 55412 37166
rect 55356 37102 55358 37154
rect 55410 37102 55412 37154
rect 55356 36820 55412 37102
rect 55580 37044 55636 38222
rect 57820 37380 57876 37390
rect 57820 37286 57876 37324
rect 58156 37266 58212 37278
rect 58156 37214 58158 37266
rect 58210 37214 58212 37266
rect 55132 36764 55412 36820
rect 55468 36988 55636 37044
rect 56028 37154 56084 37166
rect 56028 37102 56030 37154
rect 56082 37102 56084 37154
rect 54684 35756 54964 35812
rect 54572 35086 54574 35138
rect 54626 35086 54628 35138
rect 54572 35074 54628 35086
rect 54796 34914 54852 34926
rect 54796 34862 54798 34914
rect 54850 34862 54852 34914
rect 54796 34692 54852 34862
rect 54236 34636 54852 34692
rect 54124 33618 54180 33628
rect 54908 33460 54964 35756
rect 55132 35700 55188 36764
rect 55468 36708 55524 36988
rect 55244 36652 55524 36708
rect 55244 36484 55300 36652
rect 55244 36390 55300 36428
rect 55580 36484 55636 36494
rect 56028 36484 56084 37102
rect 57596 37154 57652 37166
rect 57596 37102 57598 37154
rect 57650 37102 57652 37154
rect 57596 37044 57652 37102
rect 57596 36978 57652 36988
rect 58156 37044 58212 37214
rect 58156 36978 58212 36988
rect 55580 36482 56084 36484
rect 55580 36430 55582 36482
rect 55634 36430 56084 36482
rect 55580 36428 56084 36430
rect 57932 36594 57988 36606
rect 57932 36542 57934 36594
rect 57986 36542 57988 36594
rect 55468 35812 55524 35822
rect 55468 35718 55524 35756
rect 55244 35700 55300 35710
rect 55132 35698 55300 35700
rect 55132 35646 55246 35698
rect 55298 35646 55300 35698
rect 55132 35644 55300 35646
rect 55244 35634 55300 35644
rect 55580 35588 55636 36428
rect 57820 35924 57876 35934
rect 57820 35810 57876 35868
rect 57820 35758 57822 35810
rect 57874 35758 57876 35810
rect 57820 35746 57876 35758
rect 57932 35812 57988 36542
rect 57932 35746 57988 35756
rect 58156 35698 58212 35710
rect 58156 35646 58158 35698
rect 58210 35646 58212 35698
rect 55580 35522 55636 35532
rect 57596 35588 57652 35598
rect 58156 35588 58212 35646
rect 57596 35586 58212 35588
rect 57596 35534 57598 35586
rect 57650 35534 58212 35586
rect 57596 35532 58212 35534
rect 57596 35522 57652 35532
rect 58156 35028 58212 35532
rect 58156 34962 58212 34972
rect 54684 33458 54964 33460
rect 54684 33406 54910 33458
rect 54962 33406 54964 33458
rect 54684 33404 54964 33406
rect 54572 33348 54628 33358
rect 53788 33294 53790 33346
rect 53842 33294 53844 33346
rect 53788 33282 53844 33294
rect 54460 33292 54572 33348
rect 53564 33142 53620 33180
rect 54124 33234 54180 33246
rect 54124 33182 54126 33234
rect 54178 33182 54180 33234
rect 53228 33124 53284 33134
rect 53228 33030 53284 33068
rect 53004 32622 53006 32674
rect 53058 32622 53060 32674
rect 53004 32610 53060 32622
rect 53228 32676 53284 32686
rect 53228 32582 53284 32620
rect 53452 32564 53508 32574
rect 52892 31724 53060 31780
rect 52556 31602 52612 31612
rect 52892 31556 52948 31566
rect 52892 31462 52948 31500
rect 52444 31154 52500 31164
rect 51884 31042 51940 31052
rect 50204 30942 50206 30994
rect 50258 30942 50260 30994
rect 50204 30930 50260 30942
rect 50988 30996 51044 31006
rect 49980 30212 50036 30222
rect 50316 30212 50372 30222
rect 49980 30210 50372 30212
rect 49980 30158 49982 30210
rect 50034 30158 50318 30210
rect 50370 30158 50372 30210
rect 49980 30156 50372 30158
rect 49980 30146 50036 30156
rect 50316 30146 50372 30156
rect 50988 30210 51044 30940
rect 51660 30996 51716 31006
rect 51660 30882 51716 30940
rect 51660 30830 51662 30882
rect 51714 30830 51716 30882
rect 51660 30818 51716 30830
rect 52668 30994 52724 31006
rect 52668 30942 52670 30994
rect 52722 30942 52724 30994
rect 52556 30772 52612 30782
rect 52556 30678 52612 30716
rect 51212 30324 51268 30334
rect 51212 30230 51268 30268
rect 52668 30324 52724 30942
rect 53004 30996 53060 31724
rect 53452 31778 53508 32508
rect 54124 32564 54180 33182
rect 54124 32498 54180 32508
rect 54460 32562 54516 33292
rect 54572 33254 54628 33292
rect 54460 32510 54462 32562
rect 54514 32510 54516 32562
rect 54460 32498 54516 32510
rect 54684 32676 54740 33404
rect 54908 33394 54964 33404
rect 57148 33684 57204 33694
rect 55580 33346 55636 33358
rect 55580 33294 55582 33346
rect 55634 33294 55636 33346
rect 55580 32788 55636 33294
rect 55580 32722 55636 32732
rect 56700 32786 56756 32798
rect 56700 32734 56702 32786
rect 56754 32734 56756 32786
rect 54684 32562 54740 32620
rect 54684 32510 54686 32562
rect 54738 32510 54740 32562
rect 54684 32498 54740 32510
rect 54908 32564 54964 32574
rect 56588 32564 56644 32574
rect 54908 32562 55076 32564
rect 54908 32510 54910 32562
rect 54962 32510 55076 32562
rect 54908 32508 55076 32510
rect 54908 32498 54964 32508
rect 53452 31726 53454 31778
rect 53506 31726 53508 31778
rect 53452 31714 53508 31726
rect 54124 31892 54180 31902
rect 54124 31778 54180 31836
rect 54684 31892 54740 31902
rect 54740 31836 54852 31892
rect 54684 31826 54740 31836
rect 54124 31726 54126 31778
rect 54178 31726 54180 31778
rect 54124 31714 54180 31726
rect 54348 31666 54404 31678
rect 54348 31614 54350 31666
rect 54402 31614 54404 31666
rect 53676 31220 53732 31230
rect 54348 31220 54404 31614
rect 53732 31164 53844 31220
rect 53676 31154 53732 31164
rect 53004 30902 53060 30940
rect 53788 30994 53844 31164
rect 54236 31164 54348 31220
rect 53788 30942 53790 30994
rect 53842 30942 53844 30994
rect 53788 30930 53844 30942
rect 54124 30996 54180 31006
rect 54124 30902 54180 30940
rect 52668 30230 52724 30268
rect 53340 30772 53396 30782
rect 50988 30158 50990 30210
rect 51042 30158 51044 30210
rect 50988 30146 51044 30158
rect 53340 30210 53396 30716
rect 53340 30158 53342 30210
rect 53394 30158 53396 30210
rect 53340 30146 53396 30158
rect 49868 30046 49870 30098
rect 49922 30046 49924 30098
rect 49868 30034 49924 30046
rect 54236 30098 54292 31164
rect 54348 31154 54404 31164
rect 54796 31218 54852 31836
rect 54796 31166 54798 31218
rect 54850 31166 54852 31218
rect 54348 30994 54404 31006
rect 54348 30942 54350 30994
rect 54402 30942 54404 30994
rect 54348 30884 54404 30942
rect 54684 30884 54740 30894
rect 54348 30882 54740 30884
rect 54348 30830 54686 30882
rect 54738 30830 54740 30882
rect 54348 30828 54740 30830
rect 54684 30818 54740 30828
rect 54796 30322 54852 31166
rect 55020 30772 55076 32508
rect 56588 32470 56644 32508
rect 55580 31780 55636 31790
rect 55580 31686 55636 31724
rect 56700 30996 56756 32734
rect 57148 32562 57204 33628
rect 57820 33458 57876 33470
rect 57820 33406 57822 33458
rect 57874 33406 57876 33458
rect 57260 33124 57316 33134
rect 57260 32674 57316 33068
rect 57260 32622 57262 32674
rect 57314 32622 57316 32674
rect 57260 32610 57316 32622
rect 57148 32510 57150 32562
rect 57202 32510 57204 32562
rect 57148 32498 57204 32510
rect 56700 30930 56756 30940
rect 57820 30996 57876 33406
rect 57932 32340 57988 32350
rect 57932 31890 57988 32284
rect 57932 31838 57934 31890
rect 57986 31838 57988 31890
rect 57932 31826 57988 31838
rect 57820 30930 57876 30940
rect 57932 31668 57988 31678
rect 55020 30678 55076 30716
rect 57932 30434 57988 31612
rect 57932 30382 57934 30434
rect 57986 30382 57988 30434
rect 57932 30370 57988 30382
rect 54796 30270 54798 30322
rect 54850 30270 54852 30322
rect 54796 30258 54852 30270
rect 54236 30046 54238 30098
rect 54290 30046 54292 30098
rect 54236 30034 54292 30046
rect 55580 30210 55636 30222
rect 55580 30158 55582 30210
rect 55634 30158 55636 30210
rect 48972 29988 49028 29998
rect 48972 29894 49028 29932
rect 47068 29810 47124 29820
rect 50556 29820 50820 29830
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50556 29754 50820 29764
rect 55580 29764 55636 30158
rect 55580 29698 55636 29708
rect 46620 29474 46676 29484
rect 45500 29374 45502 29426
rect 45554 29374 45556 29426
rect 45500 29362 45556 29374
rect 49756 28868 49812 28878
rect 49756 28754 49812 28812
rect 49756 28702 49758 28754
rect 49810 28702 49812 28754
rect 49756 28690 49812 28702
rect 57932 28754 57988 28766
rect 57932 28702 57934 28754
rect 57986 28702 57988 28754
rect 50316 28642 50372 28654
rect 50316 28590 50318 28642
rect 50370 28590 50372 28642
rect 44492 27918 44494 27970
rect 44546 27918 44548 27970
rect 44492 27906 44548 27918
rect 48748 28196 48804 28206
rect 48748 27970 48804 28140
rect 48748 27918 48750 27970
rect 48802 27918 48804 27970
rect 48748 27906 48804 27918
rect 45164 27860 45220 27870
rect 45164 27858 45332 27860
rect 45164 27806 45166 27858
rect 45218 27806 45332 27858
rect 45164 27804 45332 27806
rect 45164 27794 45220 27804
rect 43820 27694 43822 27746
rect 43874 27694 43876 27746
rect 43820 27682 43876 27694
rect 43260 27570 43316 27580
rect 43148 27188 43204 27198
rect 42812 26852 42868 26862
rect 42476 26516 42532 26526
rect 41916 26514 42532 26516
rect 41916 26462 42478 26514
rect 42530 26462 42532 26514
rect 41916 26460 42532 26462
rect 41916 26402 41972 26460
rect 42476 26450 42532 26460
rect 41916 26350 41918 26402
rect 41970 26350 41972 26402
rect 41916 26338 41972 26350
rect 42812 26402 42868 26796
rect 43148 26516 43204 27132
rect 43148 26450 43204 26460
rect 45276 26964 45332 27804
rect 46284 27858 46340 27870
rect 46284 27806 46286 27858
rect 46338 27806 46340 27858
rect 45388 27748 45444 27758
rect 45388 27746 45556 27748
rect 45388 27694 45390 27746
rect 45442 27694 45556 27746
rect 45388 27692 45556 27694
rect 45388 27682 45444 27692
rect 42812 26350 42814 26402
rect 42866 26350 42868 26402
rect 42812 26338 42868 26350
rect 41020 26126 41022 26178
rect 41074 26126 41076 26178
rect 39900 25778 39956 25788
rect 39452 25554 39508 25564
rect 38332 25442 38388 25452
rect 40236 25508 40292 25518
rect 40684 25508 40740 25518
rect 40236 25414 40292 25452
rect 40460 25452 40684 25508
rect 39004 25396 39060 25406
rect 39004 25282 39060 25340
rect 39004 25230 39006 25282
rect 39058 25230 39060 25282
rect 39004 24836 39060 25230
rect 39452 25284 39508 25294
rect 39452 25190 39508 25228
rect 39900 25284 39956 25294
rect 39900 25190 39956 25228
rect 39228 24836 39284 24846
rect 39900 24836 39956 24846
rect 39004 24780 39228 24836
rect 39228 24610 39284 24780
rect 39228 24558 39230 24610
rect 39282 24558 39284 24610
rect 39228 24546 39284 24558
rect 39452 24834 39956 24836
rect 39452 24782 39902 24834
rect 39954 24782 39956 24834
rect 39452 24780 39956 24782
rect 37772 24108 38276 24164
rect 37100 23826 37268 23828
rect 37100 23774 37102 23826
rect 37154 23774 37268 23826
rect 37100 23772 37268 23774
rect 37660 23940 37716 23950
rect 37660 23826 37716 23884
rect 37772 23938 37828 24108
rect 38220 24050 38276 24108
rect 38220 23998 38222 24050
rect 38274 23998 38276 24050
rect 38220 23986 38276 23998
rect 37772 23886 37774 23938
rect 37826 23886 37828 23938
rect 37772 23874 37828 23886
rect 38108 23940 38164 23950
rect 37660 23774 37662 23826
rect 37714 23774 37716 23826
rect 37100 23762 37156 23772
rect 37660 23762 37716 23774
rect 37436 23716 37492 23726
rect 37436 23622 37492 23660
rect 37100 23156 37156 23166
rect 36540 22372 36596 22382
rect 36540 22278 36596 22316
rect 36316 22258 36484 22260
rect 36316 22206 36318 22258
rect 36370 22206 36484 22258
rect 36316 22204 36484 22206
rect 36316 22194 36372 22204
rect 35084 22146 35140 22158
rect 35084 22094 35086 22146
rect 35138 22094 35140 22146
rect 34860 21812 34916 21822
rect 35084 21812 35140 22094
rect 34860 21810 35140 21812
rect 34860 21758 34862 21810
rect 34914 21758 35140 21810
rect 34860 21756 35140 21758
rect 34860 21746 34916 21756
rect 35644 21698 35700 21710
rect 35644 21646 35646 21698
rect 35698 21646 35700 21698
rect 35084 21586 35140 21598
rect 35084 21534 35086 21586
rect 35138 21534 35140 21586
rect 34972 21474 35028 21486
rect 34972 21422 34974 21474
rect 35026 21422 35028 21474
rect 34972 20132 35028 21422
rect 35084 20916 35140 21534
rect 35532 21588 35588 21598
rect 35644 21588 35700 21646
rect 35532 21586 35700 21588
rect 35532 21534 35534 21586
rect 35586 21534 35700 21586
rect 35532 21532 35700 21534
rect 35868 21698 35924 21710
rect 35868 21646 35870 21698
rect 35922 21646 35924 21698
rect 35532 21522 35588 21532
rect 35868 21476 35924 21646
rect 35980 21700 36036 21710
rect 36428 21700 36484 22204
rect 36988 22258 37044 22270
rect 36988 22206 36990 22258
rect 37042 22206 37044 22258
rect 36988 22148 37044 22206
rect 36988 22082 37044 22092
rect 37100 21924 37156 23100
rect 38108 23042 38164 23884
rect 39340 23828 39396 23838
rect 39340 23734 39396 23772
rect 38556 23492 38612 23502
rect 38556 23378 38612 23436
rect 38556 23326 38558 23378
rect 38610 23326 38612 23378
rect 38556 23314 38612 23326
rect 38108 22990 38110 23042
rect 38162 22990 38164 23042
rect 38108 22978 38164 22990
rect 38668 23156 38724 23166
rect 37884 22482 37940 22494
rect 37884 22430 37886 22482
rect 37938 22430 37940 22482
rect 37436 22372 37492 22382
rect 37436 22278 37492 22316
rect 36988 21868 37156 21924
rect 36036 21644 36148 21700
rect 36428 21644 36596 21700
rect 35980 21606 36036 21644
rect 35868 21410 35924 21420
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 35084 20850 35140 20860
rect 35756 20914 35812 20926
rect 35756 20862 35758 20914
rect 35810 20862 35812 20914
rect 35644 20692 35700 20702
rect 35196 20132 35252 20142
rect 34972 20130 35252 20132
rect 34972 20078 35198 20130
rect 35250 20078 35252 20130
rect 34972 20076 35252 20078
rect 35196 20066 35252 20076
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 35644 18788 35700 20636
rect 35756 20468 35812 20862
rect 36092 20802 36148 21644
rect 36204 21588 36260 21598
rect 36204 21026 36260 21532
rect 36428 21476 36484 21486
rect 36428 21382 36484 21420
rect 36204 20974 36206 21026
rect 36258 20974 36260 21026
rect 36204 20962 36260 20974
rect 36092 20750 36094 20802
rect 36146 20750 36148 20802
rect 36092 20738 36148 20750
rect 36204 20580 36260 20590
rect 36204 20578 36372 20580
rect 36204 20526 36206 20578
rect 36258 20526 36372 20578
rect 36204 20524 36372 20526
rect 36204 20468 36260 20524
rect 35756 20412 36260 20468
rect 36204 19572 36260 19582
rect 36092 19516 36204 19572
rect 35420 18732 35924 18788
rect 35420 18674 35476 18732
rect 35420 18622 35422 18674
rect 35474 18622 35476 18674
rect 35420 18610 35476 18622
rect 34972 18564 35028 18574
rect 34860 17892 34916 17902
rect 34748 17890 34916 17892
rect 34748 17838 34862 17890
rect 34914 17838 34916 17890
rect 34748 17836 34916 17838
rect 34860 17826 34916 17836
rect 34524 17614 34526 17666
rect 34578 17614 34580 17666
rect 34524 17602 34580 17614
rect 34972 17106 35028 18508
rect 35084 18562 35140 18574
rect 35084 18510 35086 18562
rect 35138 18510 35140 18562
rect 35084 18452 35140 18510
rect 35084 17668 35140 18396
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 35308 17668 35364 17678
rect 35532 17668 35588 18732
rect 35868 18674 35924 18732
rect 35868 18622 35870 18674
rect 35922 18622 35924 18674
rect 35868 18610 35924 18622
rect 35980 18450 36036 18462
rect 35980 18398 35982 18450
rect 36034 18398 36036 18450
rect 35980 18340 36036 18398
rect 35980 18274 36036 18284
rect 35868 18228 35924 18238
rect 35868 18134 35924 18172
rect 35084 17666 35364 17668
rect 35084 17614 35310 17666
rect 35362 17614 35364 17666
rect 35084 17612 35364 17614
rect 35308 17602 35364 17612
rect 35420 17612 35588 17668
rect 35644 17668 35700 17678
rect 34972 17054 34974 17106
rect 35026 17054 35028 17106
rect 34524 16884 34580 16894
rect 34524 16882 34916 16884
rect 34524 16830 34526 16882
rect 34578 16830 34916 16882
rect 34524 16828 34916 16830
rect 34524 16818 34580 16828
rect 34636 16660 34692 16670
rect 34636 16658 34804 16660
rect 34636 16606 34638 16658
rect 34690 16606 34804 16658
rect 34636 16604 34804 16606
rect 34636 16594 34692 16604
rect 33404 15988 33460 15998
rect 33404 15894 33460 15932
rect 33292 15874 33348 15886
rect 34076 15876 34132 15886
rect 33292 15822 33294 15874
rect 33346 15822 33348 15874
rect 33068 15316 33124 15326
rect 33292 15316 33348 15822
rect 33124 15260 33348 15316
rect 33628 15874 34132 15876
rect 33628 15822 34078 15874
rect 34130 15822 34132 15874
rect 33628 15820 34132 15822
rect 33068 14754 33124 15260
rect 33628 15148 33684 15820
rect 34076 15810 34132 15820
rect 34188 15428 34244 15438
rect 33852 15372 34188 15428
rect 33740 15316 33796 15326
rect 33740 15222 33796 15260
rect 33068 14702 33070 14754
rect 33122 14702 33124 14754
rect 33068 14690 33124 14702
rect 33516 15092 33684 15148
rect 32396 14530 32452 14542
rect 32396 14478 32398 14530
rect 32450 14478 32452 14530
rect 32396 13746 32452 14478
rect 33516 14418 33572 15092
rect 33516 14366 33518 14418
rect 33570 14366 33572 14418
rect 32732 14308 32788 14318
rect 32732 14214 32788 14252
rect 32956 14308 33012 14318
rect 33516 14308 33572 14366
rect 32956 14306 33572 14308
rect 32956 14254 32958 14306
rect 33010 14254 33572 14306
rect 32956 14252 33572 14254
rect 32956 14242 33012 14252
rect 32508 13972 32564 13982
rect 32508 13878 32564 13916
rect 32396 13694 32398 13746
rect 32450 13694 32452 13746
rect 32396 11394 32452 13694
rect 33180 13636 33236 13646
rect 33180 13074 33236 13580
rect 33516 13300 33572 14252
rect 33628 14530 33684 14542
rect 33628 14478 33630 14530
rect 33682 14478 33684 14530
rect 33628 14308 33684 14478
rect 33628 13524 33684 14252
rect 33852 14306 33908 15372
rect 34188 15362 34244 15372
rect 33852 14254 33854 14306
rect 33906 14254 33908 14306
rect 33852 13746 33908 14254
rect 33852 13694 33854 13746
rect 33906 13694 33908 13746
rect 33852 13682 33908 13694
rect 34076 15202 34132 15214
rect 34076 15150 34078 15202
rect 34130 15150 34132 15202
rect 34076 13636 34132 15150
rect 34300 15204 34356 16044
rect 34412 16436 34468 16446
rect 34412 15986 34468 16380
rect 34412 15934 34414 15986
rect 34466 15934 34468 15986
rect 34412 15922 34468 15934
rect 34636 15988 34692 15998
rect 34636 15538 34692 15932
rect 34748 15652 34804 16604
rect 34860 16212 34916 16828
rect 34972 16772 35028 17054
rect 35308 17108 35364 17118
rect 35420 17108 35476 17612
rect 35644 17574 35700 17612
rect 35980 17668 36036 17678
rect 36092 17668 36148 19516
rect 36204 19506 36260 19516
rect 35980 17666 36260 17668
rect 35980 17614 35982 17666
rect 36034 17614 36260 17666
rect 35980 17612 36260 17614
rect 35980 17602 36036 17612
rect 35308 17106 35476 17108
rect 35308 17054 35310 17106
rect 35362 17054 35476 17106
rect 35308 17052 35476 17054
rect 35532 17442 35588 17454
rect 35532 17390 35534 17442
rect 35586 17390 35588 17442
rect 35532 17108 35588 17390
rect 35756 17444 35812 17454
rect 35756 17350 35812 17388
rect 35308 17042 35364 17052
rect 35532 17042 35588 17052
rect 35756 16884 35812 16894
rect 35756 16882 36036 16884
rect 35756 16830 35758 16882
rect 35810 16830 36036 16882
rect 35756 16828 36036 16830
rect 35756 16818 35812 16828
rect 34972 16436 35028 16716
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 34972 16370 35028 16380
rect 35308 16324 35364 16334
rect 34860 16156 35252 16212
rect 34972 15988 35028 15998
rect 34972 15986 35140 15988
rect 34972 15934 34974 15986
rect 35026 15934 35140 15986
rect 34972 15932 35140 15934
rect 34972 15922 35028 15932
rect 35084 15876 35140 15932
rect 35084 15810 35140 15820
rect 34860 15652 34916 15662
rect 34748 15596 34860 15652
rect 34860 15586 34916 15596
rect 34636 15486 34638 15538
rect 34690 15486 34692 15538
rect 34636 15474 34692 15486
rect 34860 15428 34916 15438
rect 34860 15334 34916 15372
rect 34972 15314 35028 15326
rect 34972 15262 34974 15314
rect 35026 15262 35028 15314
rect 34412 15204 34468 15214
rect 34300 15202 34468 15204
rect 34300 15150 34414 15202
rect 34466 15150 34468 15202
rect 34300 15148 34468 15150
rect 34412 15138 34468 15148
rect 34860 15092 34916 15102
rect 34524 14532 34580 14542
rect 34524 14438 34580 14476
rect 34748 14530 34804 14542
rect 34748 14478 34750 14530
rect 34802 14478 34804 14530
rect 34076 13570 34132 13580
rect 34188 13860 34244 13870
rect 33628 13458 33684 13468
rect 33516 13244 33684 13300
rect 33180 13022 33182 13074
rect 33234 13022 33236 13074
rect 33180 13010 33236 13022
rect 33180 11506 33236 11518
rect 33180 11454 33182 11506
rect 33234 11454 33236 11506
rect 32396 11342 32398 11394
rect 32450 11342 32452 11394
rect 32396 11330 32452 11342
rect 32956 11394 33012 11406
rect 32956 11342 32958 11394
rect 33010 11342 33012 11394
rect 32508 10724 32564 10734
rect 32508 10630 32564 10668
rect 32284 10108 32452 10164
rect 32284 9938 32340 9950
rect 32284 9886 32286 9938
rect 32338 9886 32340 9938
rect 32284 9828 32340 9886
rect 32284 9762 32340 9772
rect 31164 9426 31220 9436
rect 32060 9602 32116 9614
rect 32060 9550 32062 9602
rect 32114 9550 32116 9602
rect 31052 9380 31108 9390
rect 31052 8370 31108 9324
rect 32060 9380 32116 9550
rect 32060 9314 32116 9324
rect 32172 9268 32228 9660
rect 32284 9604 32340 9614
rect 32284 9510 32340 9548
rect 32396 9492 32452 10108
rect 32956 10052 33012 11342
rect 33180 10612 33236 11454
rect 33516 10612 33572 10622
rect 33180 10610 33572 10612
rect 33180 10558 33518 10610
rect 33570 10558 33572 10610
rect 33180 10556 33572 10558
rect 32956 9938 33012 9996
rect 32956 9886 32958 9938
rect 33010 9886 33012 9938
rect 32956 9874 33012 9886
rect 33068 10500 33124 10510
rect 32620 9826 32676 9838
rect 32620 9774 32622 9826
rect 32674 9774 32676 9826
rect 32396 9436 32564 9492
rect 32172 9202 32228 9212
rect 31164 9156 31220 9166
rect 31164 9154 31780 9156
rect 31164 9102 31166 9154
rect 31218 9102 31780 9154
rect 31164 9100 31780 9102
rect 31164 9090 31220 9100
rect 31052 8318 31054 8370
rect 31106 8318 31108 8370
rect 31052 8306 31108 8318
rect 31164 8930 31220 8942
rect 31164 8878 31166 8930
rect 31218 8878 31220 8930
rect 31164 8146 31220 8878
rect 31388 8820 31444 8830
rect 31388 8726 31444 8764
rect 31164 8094 31166 8146
rect 31218 8094 31220 8146
rect 31164 8082 31220 8094
rect 31388 8260 31444 8270
rect 30492 6580 30548 6590
rect 30492 6486 30548 6524
rect 30940 6132 30996 6636
rect 31388 7588 31444 8204
rect 31388 6690 31444 7532
rect 31724 7476 31780 9100
rect 31836 9154 31892 9166
rect 31836 9102 31838 9154
rect 31890 9102 31892 9154
rect 31836 8372 31892 9102
rect 32172 9044 32228 9054
rect 32172 9042 32340 9044
rect 32172 8990 32174 9042
rect 32226 8990 32340 9042
rect 32172 8988 32340 8990
rect 32172 8978 32228 8988
rect 32284 8820 32340 8988
rect 31892 8316 32004 8372
rect 31836 8306 31892 8316
rect 31948 7476 32004 8316
rect 31724 7474 31892 7476
rect 31724 7422 31726 7474
rect 31778 7422 31892 7474
rect 31724 7420 31892 7422
rect 31724 7410 31780 7420
rect 31836 6692 31892 7420
rect 31948 7382 32004 7420
rect 31388 6638 31390 6690
rect 31442 6638 31444 6690
rect 31388 6626 31444 6638
rect 31500 6690 31892 6692
rect 31500 6638 31838 6690
rect 31890 6638 31892 6690
rect 31500 6636 31892 6638
rect 31052 6466 31108 6478
rect 31500 6468 31556 6636
rect 31836 6626 31892 6636
rect 32172 7250 32228 7262
rect 32172 7198 32174 7250
rect 32226 7198 32228 7250
rect 31052 6414 31054 6466
rect 31106 6414 31108 6466
rect 31052 6356 31108 6414
rect 31052 6290 31108 6300
rect 31164 6412 31556 6468
rect 30940 6076 31108 6132
rect 29484 5854 29486 5906
rect 29538 5854 29540 5906
rect 29484 5842 29540 5854
rect 30044 5906 30100 5918
rect 30044 5854 30046 5906
rect 30098 5854 30100 5906
rect 29260 5794 29316 5806
rect 29260 5742 29262 5794
rect 29314 5742 29316 5794
rect 29260 5124 29316 5742
rect 30044 5460 30100 5854
rect 30044 5394 30100 5404
rect 30492 5906 30548 5918
rect 30492 5854 30494 5906
rect 30546 5854 30548 5906
rect 29260 4788 29316 5068
rect 29708 5124 29764 5134
rect 29708 5030 29764 5068
rect 30044 5124 30100 5134
rect 30044 5010 30100 5068
rect 30044 4958 30046 5010
rect 30098 4958 30100 5010
rect 30044 4946 30100 4958
rect 30492 5012 30548 5854
rect 30940 5908 30996 5918
rect 30940 5814 30996 5852
rect 30940 5572 30996 5582
rect 30940 5234 30996 5516
rect 30940 5182 30942 5234
rect 30994 5182 30996 5234
rect 30940 5170 30996 5182
rect 30492 4946 30548 4956
rect 29260 4722 29316 4732
rect 29372 4898 29428 4910
rect 29372 4846 29374 4898
rect 29426 4846 29428 4898
rect 29372 4564 29428 4846
rect 30380 4900 30436 4910
rect 30380 4806 30436 4844
rect 28812 4508 29428 4564
rect 28812 4338 28868 4508
rect 28812 4286 28814 4338
rect 28866 4286 28868 4338
rect 28812 4274 28868 4286
rect 29484 4116 29540 4126
rect 29484 4022 29540 4060
rect 28700 3390 28702 3442
rect 28754 3390 28756 3442
rect 28700 3378 28756 3390
rect 29260 3666 29316 3678
rect 29260 3614 29262 3666
rect 29314 3614 29316 3666
rect 29260 3388 29316 3614
rect 28252 2044 28532 2100
rect 28924 3332 29316 3388
rect 30268 3668 30324 3678
rect 28252 800 28308 2044
rect 28924 800 28980 3332
rect 30268 800 30324 3612
rect 31052 3556 31108 6076
rect 31164 5346 31220 6412
rect 32060 6356 32116 6366
rect 31164 5294 31166 5346
rect 31218 5294 31220 5346
rect 31164 5282 31220 5294
rect 31388 5906 31444 5918
rect 31388 5854 31390 5906
rect 31442 5854 31444 5906
rect 31388 5236 31444 5854
rect 31836 5794 31892 5806
rect 31836 5742 31838 5794
rect 31890 5742 31892 5794
rect 31836 5684 31892 5742
rect 31836 5618 31892 5628
rect 32060 5460 32116 6300
rect 32172 5796 32228 7198
rect 32284 6244 32340 8764
rect 32396 6692 32452 6702
rect 32396 6598 32452 6636
rect 32284 6188 32452 6244
rect 32172 5730 32228 5740
rect 31836 5404 32116 5460
rect 32172 5460 32228 5470
rect 31500 5236 31556 5246
rect 31388 5180 31500 5236
rect 31500 4340 31556 5180
rect 31612 5124 31668 5134
rect 31612 5030 31668 5068
rect 31724 5010 31780 5022
rect 31724 4958 31726 5010
rect 31778 4958 31780 5010
rect 31724 4900 31780 4958
rect 31836 4900 31892 5404
rect 31948 5236 32004 5246
rect 31948 5122 32004 5180
rect 31948 5070 31950 5122
rect 32002 5070 32004 5122
rect 31948 5058 32004 5070
rect 32060 5124 32116 5134
rect 31836 4844 32004 4900
rect 31724 4450 31780 4844
rect 31724 4398 31726 4450
rect 31778 4398 31780 4450
rect 31724 4386 31780 4398
rect 31948 4450 32004 4844
rect 31948 4398 31950 4450
rect 32002 4398 32004 4450
rect 31948 4386 32004 4398
rect 31612 4340 31668 4350
rect 31500 4338 31668 4340
rect 31500 4286 31614 4338
rect 31666 4286 31668 4338
rect 31500 4284 31668 4286
rect 32060 4340 32116 5068
rect 32172 5122 32228 5404
rect 32172 5070 32174 5122
rect 32226 5070 32228 5122
rect 32172 4564 32228 5070
rect 32172 4498 32228 4508
rect 32284 5236 32340 5246
rect 32172 4340 32228 4350
rect 32060 4338 32228 4340
rect 32060 4286 32174 4338
rect 32226 4286 32228 4338
rect 32060 4284 32228 4286
rect 31612 4274 31668 4284
rect 31164 3556 31220 3566
rect 31052 3554 31220 3556
rect 31052 3502 31166 3554
rect 31218 3502 31220 3554
rect 31052 3500 31220 3502
rect 31164 3490 31220 3500
rect 31612 3556 31668 3566
rect 30940 3444 30996 3454
rect 30940 800 30996 3388
rect 31612 800 31668 3500
rect 32172 3220 32228 4284
rect 32172 3154 32228 3164
rect 32284 800 32340 5180
rect 32396 4564 32452 6188
rect 32508 5122 32564 9436
rect 32620 9380 32676 9774
rect 32732 9826 32788 9838
rect 32732 9774 32734 9826
rect 32786 9774 32788 9826
rect 32732 9716 32788 9774
rect 32732 9650 32788 9660
rect 33068 9826 33124 10444
rect 33068 9774 33070 9826
rect 33122 9774 33124 9826
rect 32620 9314 32676 9324
rect 33068 9156 33124 9774
rect 33404 9940 33460 9950
rect 33404 9826 33460 9884
rect 33404 9774 33406 9826
rect 33458 9774 33460 9826
rect 33404 9762 33460 9774
rect 32620 9100 33124 9156
rect 33180 9154 33236 9166
rect 33180 9102 33182 9154
rect 33234 9102 33236 9154
rect 32620 7698 32676 9100
rect 33068 8820 33124 8830
rect 32844 8818 33124 8820
rect 32844 8766 33070 8818
rect 33122 8766 33124 8818
rect 32844 8764 33124 8766
rect 32844 8146 32900 8764
rect 33068 8754 33124 8764
rect 32844 8094 32846 8146
rect 32898 8094 32900 8146
rect 32844 8082 32900 8094
rect 32620 7646 32622 7698
rect 32674 7646 32676 7698
rect 32620 7634 32676 7646
rect 33068 7588 33124 7598
rect 33068 7494 33124 7532
rect 33180 7252 33236 9102
rect 33404 8818 33460 8830
rect 33404 8766 33406 8818
rect 33458 8766 33460 8818
rect 33404 8148 33460 8766
rect 33516 8370 33572 10556
rect 33628 8708 33684 13244
rect 34188 12962 34244 13804
rect 34748 13860 34804 14478
rect 34748 13794 34804 13804
rect 34188 12910 34190 12962
rect 34242 12910 34244 12962
rect 34188 12898 34244 12910
rect 33852 11844 33908 11854
rect 33628 8642 33684 8652
rect 33740 9604 33796 9614
rect 33740 9042 33796 9548
rect 33740 8990 33742 9042
rect 33794 8990 33796 9042
rect 33740 8484 33796 8990
rect 33740 8418 33796 8428
rect 33516 8318 33518 8370
rect 33570 8318 33572 8370
rect 33516 8306 33572 8318
rect 33740 8260 33796 8270
rect 33740 8148 33796 8204
rect 33404 8092 33796 8148
rect 33292 7476 33348 7486
rect 33292 7382 33348 7420
rect 33740 7474 33796 8092
rect 33740 7422 33742 7474
rect 33794 7422 33796 7474
rect 33740 7410 33796 7422
rect 33516 7252 33572 7262
rect 33180 7196 33516 7252
rect 33516 7158 33572 7196
rect 32732 6690 32788 6702
rect 32732 6638 32734 6690
rect 32786 6638 32788 6690
rect 32732 6580 32788 6638
rect 32732 6514 32788 6524
rect 33628 6580 33684 6590
rect 33628 6578 33796 6580
rect 33628 6526 33630 6578
rect 33682 6526 33796 6578
rect 33628 6524 33796 6526
rect 33628 6514 33684 6524
rect 33516 6132 33572 6142
rect 33068 5906 33124 5918
rect 33068 5854 33070 5906
rect 33122 5854 33124 5906
rect 32620 5796 32676 5806
rect 32620 5794 32788 5796
rect 32620 5742 32622 5794
rect 32674 5742 32788 5794
rect 32620 5740 32788 5742
rect 32620 5730 32676 5740
rect 32508 5070 32510 5122
rect 32562 5070 32564 5122
rect 32508 5058 32564 5070
rect 32620 4564 32676 4574
rect 32396 4562 32676 4564
rect 32396 4510 32622 4562
rect 32674 4510 32676 4562
rect 32396 4508 32676 4510
rect 32620 4498 32676 4508
rect 32396 3668 32452 3678
rect 32396 3574 32452 3612
rect 32620 3556 32676 3566
rect 32732 3556 32788 5740
rect 33068 5348 33124 5854
rect 33516 5794 33572 6076
rect 33740 5908 33796 6524
rect 33852 6468 33908 11788
rect 34076 11506 34132 11518
rect 34076 11454 34078 11506
rect 34130 11454 34132 11506
rect 34076 10724 34132 11454
rect 34860 11506 34916 15036
rect 34972 13972 35028 15262
rect 35196 15148 35252 16156
rect 35308 15986 35364 16268
rect 35532 16100 35588 16110
rect 35532 16006 35588 16044
rect 35868 15988 35924 15998
rect 35308 15934 35310 15986
rect 35362 15934 35364 15986
rect 35308 15922 35364 15934
rect 35756 15932 35868 15988
rect 35756 15876 35812 15932
rect 35868 15894 35924 15932
rect 35644 15540 35700 15550
rect 35756 15540 35812 15820
rect 35980 15652 36036 16828
rect 36204 16882 36260 17612
rect 36204 16830 36206 16882
rect 36258 16830 36260 16882
rect 36204 16818 36260 16830
rect 36092 16772 36148 16782
rect 36092 15986 36148 16716
rect 36204 16100 36260 16110
rect 36204 16006 36260 16044
rect 36092 15934 36094 15986
rect 36146 15934 36148 15986
rect 36092 15922 36148 15934
rect 35980 15596 36148 15652
rect 35644 15538 35812 15540
rect 35644 15486 35646 15538
rect 35698 15486 35812 15538
rect 35644 15484 35812 15486
rect 35644 15474 35700 15484
rect 35084 15092 35252 15148
rect 35980 15314 36036 15326
rect 35980 15262 35982 15314
rect 36034 15262 36036 15314
rect 35980 15092 36036 15262
rect 35084 14756 35140 15092
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35084 14700 35252 14756
rect 35196 14420 35252 14700
rect 35644 14532 35700 14542
rect 35196 14354 35252 14364
rect 35420 14418 35476 14430
rect 35420 14366 35422 14418
rect 35474 14366 35476 14418
rect 34972 13746 35028 13916
rect 34972 13694 34974 13746
rect 35026 13694 35028 13746
rect 34972 13682 35028 13694
rect 35084 14306 35140 14318
rect 35084 14254 35086 14306
rect 35138 14254 35140 14306
rect 35084 13748 35140 14254
rect 35420 13860 35476 14366
rect 35532 14308 35588 14318
rect 35532 14214 35588 14252
rect 35644 14306 35700 14476
rect 35980 14420 36036 15036
rect 36092 14644 36148 15596
rect 36316 15148 36372 20524
rect 36540 18452 36596 21644
rect 36988 19346 37044 21868
rect 37884 21812 37940 22430
rect 37324 21476 37380 21486
rect 37100 20578 37156 20590
rect 37100 20526 37102 20578
rect 37154 20526 37156 20578
rect 37100 20132 37156 20526
rect 37100 20066 37156 20076
rect 37324 19906 37380 21420
rect 37772 20132 37828 20142
rect 37772 20038 37828 20076
rect 37324 19854 37326 19906
rect 37378 19854 37380 19906
rect 37324 19460 37380 19854
rect 37324 19394 37380 19404
rect 36988 19294 36990 19346
rect 37042 19294 37044 19346
rect 36988 19282 37044 19294
rect 37436 19348 37492 19358
rect 37884 19348 37940 21756
rect 38668 21810 38724 23100
rect 39340 21924 39396 21934
rect 38668 21758 38670 21810
rect 38722 21758 38724 21810
rect 38556 21586 38612 21598
rect 38556 21534 38558 21586
rect 38610 21534 38612 21586
rect 38332 21476 38388 21486
rect 38556 21476 38612 21534
rect 38332 21474 38612 21476
rect 38332 21422 38334 21474
rect 38386 21422 38612 21474
rect 38332 21420 38612 21422
rect 38332 21410 38388 21420
rect 38556 21364 38612 21420
rect 38556 21298 38612 21308
rect 38668 19572 38724 21758
rect 39004 21812 39060 21822
rect 38892 21586 38948 21598
rect 38892 21534 38894 21586
rect 38946 21534 38948 21586
rect 38892 20804 38948 21534
rect 39004 21586 39060 21756
rect 39340 21810 39396 21868
rect 39340 21758 39342 21810
rect 39394 21758 39396 21810
rect 39340 21746 39396 21758
rect 39452 21812 39508 24780
rect 39900 24770 39956 24780
rect 40012 24722 40068 24734
rect 40012 24670 40014 24722
rect 40066 24670 40068 24722
rect 39900 24498 39956 24510
rect 39900 24446 39902 24498
rect 39954 24446 39956 24498
rect 39788 24050 39844 24062
rect 39788 23998 39790 24050
rect 39842 23998 39844 24050
rect 39788 23268 39844 23998
rect 39900 23940 39956 24446
rect 40012 24276 40068 24670
rect 40012 24210 40068 24220
rect 39900 23938 40292 23940
rect 39900 23886 39902 23938
rect 39954 23886 40292 23938
rect 39900 23884 40292 23886
rect 39900 23874 39956 23884
rect 40236 23378 40292 23884
rect 40236 23326 40238 23378
rect 40290 23326 40292 23378
rect 40236 23314 40292 23326
rect 40460 23378 40516 25452
rect 40684 25414 40740 25452
rect 41020 25284 41076 26126
rect 41580 26290 41636 26302
rect 41580 26238 41582 26290
rect 41634 26238 41636 26290
rect 41468 26068 41524 26078
rect 41580 26068 41636 26238
rect 41468 26066 41636 26068
rect 41468 26014 41470 26066
rect 41522 26014 41636 26066
rect 41468 26012 41636 26014
rect 42588 26292 42644 26302
rect 41468 26002 41524 26012
rect 41020 25218 41076 25228
rect 41132 25508 41188 25518
rect 41580 25508 41636 25518
rect 41132 25506 41524 25508
rect 41132 25454 41134 25506
rect 41186 25454 41524 25506
rect 41132 25452 41524 25454
rect 41132 25060 41188 25452
rect 40908 25004 41188 25060
rect 40908 23940 40964 25004
rect 41020 24834 41076 24846
rect 41020 24782 41022 24834
rect 41074 24782 41076 24834
rect 41020 24164 41076 24782
rect 41132 24724 41188 24734
rect 41468 24724 41524 25452
rect 41580 25414 41636 25452
rect 41692 25282 41748 25294
rect 41692 25230 41694 25282
rect 41746 25230 41748 25282
rect 41692 24834 41748 25230
rect 41692 24782 41694 24834
rect 41746 24782 41748 24834
rect 41692 24770 41748 24782
rect 42140 25282 42196 25294
rect 42140 25230 42142 25282
rect 42194 25230 42196 25282
rect 41580 24724 41636 24734
rect 41468 24722 41636 24724
rect 41468 24670 41582 24722
rect 41634 24670 41636 24722
rect 41468 24668 41636 24670
rect 41132 24630 41188 24668
rect 41580 24658 41636 24668
rect 41244 24498 41300 24510
rect 41244 24446 41246 24498
rect 41298 24446 41300 24498
rect 41244 24276 41300 24446
rect 42140 24276 42196 25230
rect 42588 24946 42644 26236
rect 43260 26292 43316 26302
rect 43260 26198 43316 26236
rect 44492 26292 44548 26302
rect 44492 26198 44548 26236
rect 45164 26290 45220 26302
rect 45164 26238 45166 26290
rect 45218 26238 45220 26290
rect 43708 26180 43764 26190
rect 44380 26180 44436 26190
rect 43764 26124 43876 26180
rect 43708 26086 43764 26124
rect 42588 24894 42590 24946
rect 42642 24894 42644 24946
rect 42588 24882 42644 24894
rect 43820 24834 43876 26124
rect 44380 26086 44436 26124
rect 44828 25508 44884 25518
rect 44828 25506 45108 25508
rect 44828 25454 44830 25506
rect 44882 25454 45108 25506
rect 44828 25452 45108 25454
rect 44828 25442 44884 25452
rect 43820 24782 43822 24834
rect 43874 24782 43876 24834
rect 43820 24770 43876 24782
rect 44940 25282 44996 25294
rect 44940 25230 44942 25282
rect 44994 25230 44996 25282
rect 42476 24724 42532 24734
rect 42476 24630 42532 24668
rect 44268 24724 44324 24734
rect 44940 24724 44996 25230
rect 44268 24722 44996 24724
rect 44268 24670 44270 24722
rect 44322 24670 44996 24722
rect 44268 24668 44996 24670
rect 44156 24610 44212 24622
rect 44156 24558 44158 24610
rect 44210 24558 44212 24610
rect 41244 24220 41636 24276
rect 41020 24108 41524 24164
rect 41020 23940 41076 23950
rect 40908 23938 41076 23940
rect 40908 23886 41022 23938
rect 41074 23886 41076 23938
rect 40908 23884 41076 23886
rect 41020 23874 41076 23884
rect 41468 23938 41524 24108
rect 41468 23886 41470 23938
rect 41522 23886 41524 23938
rect 40460 23326 40462 23378
rect 40514 23326 40516 23378
rect 40460 23314 40516 23326
rect 41020 23380 41076 23390
rect 41020 23286 41076 23324
rect 41468 23378 41524 23886
rect 41580 23940 41636 24220
rect 41916 23940 41972 23950
rect 41580 23938 41972 23940
rect 41580 23886 41918 23938
rect 41970 23886 41972 23938
rect 41580 23884 41972 23886
rect 41468 23326 41470 23378
rect 41522 23326 41524 23378
rect 41468 23314 41524 23326
rect 40124 23268 40180 23278
rect 39564 23266 40180 23268
rect 39564 23214 40126 23266
rect 40178 23214 40180 23266
rect 39564 23212 40180 23214
rect 39564 22482 39620 23212
rect 40124 23202 40180 23212
rect 40908 23156 40964 23166
rect 40908 23062 40964 23100
rect 41244 23156 41300 23166
rect 41580 23156 41636 23166
rect 41244 23154 41636 23156
rect 41244 23102 41246 23154
rect 41298 23102 41582 23154
rect 41634 23102 41636 23154
rect 41244 23100 41636 23102
rect 41244 23090 41300 23100
rect 41580 23090 41636 23100
rect 40236 23044 40292 23054
rect 39564 22430 39566 22482
rect 39618 22430 39620 22482
rect 39564 22418 39620 22430
rect 40124 22988 40236 23044
rect 40012 22370 40068 22382
rect 40012 22318 40014 22370
rect 40066 22318 40068 22370
rect 40012 22148 40068 22318
rect 40012 21924 40068 22092
rect 39788 21868 40068 21924
rect 40124 21924 40180 22988
rect 40236 22978 40292 22988
rect 41132 22484 41188 22494
rect 41916 22484 41972 23884
rect 42140 23380 42196 24220
rect 44044 24276 44100 24286
rect 42140 23286 42196 23324
rect 43036 23828 43092 23838
rect 43036 23154 43092 23772
rect 43932 23828 43988 23838
rect 43932 23734 43988 23772
rect 44044 23826 44100 24220
rect 44156 24052 44212 24558
rect 44156 23986 44212 23996
rect 44268 23938 44324 24668
rect 44940 24276 44996 24286
rect 44940 24050 44996 24220
rect 44940 23998 44942 24050
rect 44994 23998 44996 24050
rect 44940 23986 44996 23998
rect 45052 24052 45108 25452
rect 45164 25506 45220 26238
rect 45276 26178 45332 26908
rect 45276 26126 45278 26178
rect 45330 26126 45332 26178
rect 45276 26114 45332 26126
rect 45500 27074 45556 27692
rect 45948 27634 46004 27646
rect 45948 27582 45950 27634
rect 46002 27582 46004 27634
rect 45948 27300 46004 27582
rect 45948 27234 46004 27244
rect 45500 27022 45502 27074
rect 45554 27022 45556 27074
rect 45500 25730 45556 27022
rect 45612 26964 45668 27002
rect 45612 26898 45668 26908
rect 45948 26404 46004 26414
rect 45500 25678 45502 25730
rect 45554 25678 45556 25730
rect 45500 25666 45556 25678
rect 45836 26402 46004 26404
rect 45836 26350 45950 26402
rect 46002 26350 46004 26402
rect 45836 26348 46004 26350
rect 45164 25454 45166 25506
rect 45218 25454 45220 25506
rect 45164 25442 45220 25454
rect 45612 25508 45668 25518
rect 45836 25508 45892 26348
rect 45948 26338 46004 26348
rect 46060 26290 46116 26302
rect 46060 26238 46062 26290
rect 46114 26238 46116 26290
rect 45668 25452 45892 25508
rect 45948 26066 46004 26078
rect 45948 26014 45950 26066
rect 46002 26014 46004 26066
rect 45948 25506 46004 26014
rect 46060 25844 46116 26238
rect 46284 26068 46340 27806
rect 47964 27860 48020 27870
rect 47964 27858 48132 27860
rect 47964 27806 47966 27858
rect 48018 27806 48132 27858
rect 47964 27804 48132 27806
rect 47964 27794 48020 27804
rect 47628 27746 47684 27758
rect 47628 27694 47630 27746
rect 47682 27694 47684 27746
rect 46508 27076 46564 27086
rect 46508 26850 46564 27020
rect 46620 27074 46676 27086
rect 46620 27022 46622 27074
rect 46674 27022 46676 27074
rect 46620 26908 46676 27022
rect 47404 27074 47460 27086
rect 47404 27022 47406 27074
rect 47458 27022 47460 27074
rect 46620 26852 47012 26908
rect 46508 26798 46510 26850
rect 46562 26798 46564 26850
rect 46508 26786 46564 26798
rect 46284 26002 46340 26012
rect 46060 25788 46452 25844
rect 45948 25454 45950 25506
rect 46002 25454 46004 25506
rect 45388 24948 45444 24958
rect 45388 24722 45444 24892
rect 45612 24946 45668 25452
rect 45948 25442 46004 25454
rect 46284 25618 46340 25630
rect 46284 25566 46286 25618
rect 46338 25566 46340 25618
rect 46284 25396 46340 25566
rect 46396 25508 46452 25788
rect 46956 25618 47012 26852
rect 47404 26292 47460 27022
rect 47628 26852 47684 27694
rect 47964 27188 48020 27198
rect 47628 26786 47684 26796
rect 47740 27186 48020 27188
rect 47740 27134 47966 27186
rect 48018 27134 48020 27186
rect 47740 27132 48020 27134
rect 47740 26628 47796 27132
rect 47964 27122 48020 27132
rect 48076 27076 48132 27804
rect 49196 27858 49252 27870
rect 50316 27860 50372 28590
rect 50652 28644 50708 28654
rect 51100 28644 51156 28654
rect 50652 28642 51044 28644
rect 50652 28590 50654 28642
rect 50706 28590 51044 28642
rect 50652 28588 51044 28590
rect 50652 28578 50708 28588
rect 50556 28252 50820 28262
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50556 28186 50820 28196
rect 49196 27806 49198 27858
rect 49250 27806 49252 27858
rect 48076 26982 48132 27020
rect 49084 27746 49140 27758
rect 49084 27694 49086 27746
rect 49138 27694 49140 27746
rect 49084 27074 49140 27694
rect 49084 27022 49086 27074
rect 49138 27022 49140 27074
rect 48748 26964 48804 27002
rect 48748 26898 48804 26908
rect 47516 26572 47796 26628
rect 47852 26852 47908 26862
rect 47516 26514 47572 26572
rect 47516 26462 47518 26514
rect 47570 26462 47572 26514
rect 47516 26450 47572 26462
rect 47740 26292 47796 26302
rect 47852 26292 47908 26796
rect 47404 26236 47572 26292
rect 46956 25566 46958 25618
rect 47010 25566 47012 25618
rect 46956 25554 47012 25566
rect 47404 26068 47460 26078
rect 47404 25620 47460 26012
rect 47404 25554 47460 25564
rect 46732 25508 46788 25518
rect 46396 25506 46788 25508
rect 46396 25454 46734 25506
rect 46786 25454 46788 25506
rect 46396 25452 46788 25454
rect 46284 25330 46340 25340
rect 45612 24894 45614 24946
rect 45666 24894 45668 24946
rect 45612 24882 45668 24894
rect 46060 24948 46116 24958
rect 46060 24854 46116 24892
rect 45388 24670 45390 24722
rect 45442 24670 45444 24722
rect 45388 24276 45444 24670
rect 45388 24210 45444 24220
rect 45052 23986 45108 23996
rect 45836 24052 45892 24062
rect 45836 23958 45892 23996
rect 44268 23886 44270 23938
rect 44322 23886 44324 23938
rect 44268 23874 44324 23886
rect 46284 23938 46340 23950
rect 46284 23886 46286 23938
rect 46338 23886 46340 23938
rect 44044 23774 44046 23826
rect 44098 23774 44100 23826
rect 44044 23762 44100 23774
rect 45276 23604 45332 23614
rect 44044 23378 44100 23390
rect 44044 23326 44046 23378
rect 44098 23326 44100 23378
rect 43036 23102 43038 23154
rect 43090 23102 43092 23154
rect 42812 23044 42868 23054
rect 42812 22950 42868 22988
rect 42028 22484 42084 22494
rect 41132 22482 41860 22484
rect 41132 22430 41134 22482
rect 41186 22430 41860 22482
rect 41132 22428 41860 22430
rect 41916 22482 42084 22484
rect 41916 22430 42030 22482
rect 42082 22430 42084 22482
rect 41916 22428 42084 22430
rect 41132 22418 41188 22428
rect 40460 22370 40516 22382
rect 40460 22318 40462 22370
rect 40514 22318 40516 22370
rect 40460 22260 40516 22318
rect 40460 22194 40516 22204
rect 40908 22370 40964 22382
rect 40908 22318 40910 22370
rect 40962 22318 40964 22370
rect 40908 22148 40964 22318
rect 41244 22260 41300 22270
rect 41300 22204 41412 22260
rect 41244 22166 41300 22204
rect 40908 22082 40964 22092
rect 39564 21812 39620 21822
rect 39452 21810 39620 21812
rect 39452 21758 39566 21810
rect 39618 21758 39620 21810
rect 39452 21756 39620 21758
rect 39004 21534 39006 21586
rect 39058 21534 39060 21586
rect 39004 21522 39060 21534
rect 39564 20916 39620 21756
rect 39676 21812 39732 21822
rect 39788 21812 39844 21868
rect 39676 21810 39844 21812
rect 39676 21758 39678 21810
rect 39730 21758 39844 21810
rect 39676 21756 39844 21758
rect 39676 21746 39732 21756
rect 39900 21700 39956 21710
rect 40124 21700 40180 21868
rect 39900 21698 40180 21700
rect 39900 21646 39902 21698
rect 39954 21646 40180 21698
rect 39900 21644 40180 21646
rect 40348 21756 41076 21812
rect 39900 21634 39956 21644
rect 40236 21586 40292 21598
rect 40236 21534 40238 21586
rect 40290 21534 40292 21586
rect 40236 21364 40292 21534
rect 40236 21298 40292 21308
rect 39564 20850 39620 20860
rect 38892 20748 39508 20804
rect 39452 20692 39508 20748
rect 40012 20802 40068 20814
rect 40012 20750 40014 20802
rect 40066 20750 40068 20802
rect 39452 20690 39844 20692
rect 39452 20638 39454 20690
rect 39506 20638 39844 20690
rect 39452 20636 39844 20638
rect 39452 20626 39508 20636
rect 39788 20130 39844 20636
rect 39788 20078 39790 20130
rect 39842 20078 39844 20130
rect 39788 20066 39844 20078
rect 40012 20020 40068 20750
rect 40348 20242 40404 21756
rect 41020 21698 41076 21756
rect 41020 21646 41022 21698
rect 41074 21646 41076 21698
rect 41020 21634 41076 21646
rect 40348 20190 40350 20242
rect 40402 20190 40404 20242
rect 40348 20178 40404 20190
rect 40908 21586 40964 21598
rect 40908 21534 40910 21586
rect 40962 21534 40964 21586
rect 40124 20132 40180 20142
rect 40124 20130 40292 20132
rect 40124 20078 40126 20130
rect 40178 20078 40292 20130
rect 40124 20076 40292 20078
rect 40124 20066 40180 20076
rect 40012 19954 40068 19964
rect 40236 20018 40292 20076
rect 40908 20130 40964 21534
rect 41356 20914 41412 22204
rect 41804 21586 41860 22428
rect 42028 22418 42084 22428
rect 42588 22372 42644 22382
rect 42588 22278 42644 22316
rect 41916 21812 41972 21822
rect 41916 21718 41972 21756
rect 41804 21534 41806 21586
rect 41858 21534 41860 21586
rect 41804 21522 41860 21534
rect 42476 21474 42532 21486
rect 42476 21422 42478 21474
rect 42530 21422 42532 21474
rect 42476 21364 42532 21422
rect 42476 21298 42532 21308
rect 41356 20862 41358 20914
rect 41410 20862 41412 20914
rect 41356 20850 41412 20862
rect 40908 20078 40910 20130
rect 40962 20078 40964 20130
rect 40908 20066 40964 20078
rect 41132 20690 41188 20702
rect 41132 20638 41134 20690
rect 41186 20638 41188 20690
rect 40236 19966 40238 20018
rect 40290 19966 40292 20018
rect 40236 19954 40292 19966
rect 40796 20020 40852 20030
rect 38668 19506 38724 19516
rect 39900 19572 39956 19582
rect 39004 19460 39060 19470
rect 38332 19348 38388 19358
rect 37436 19346 37604 19348
rect 37436 19294 37438 19346
rect 37490 19294 37604 19346
rect 37436 19292 37604 19294
rect 37884 19346 38388 19348
rect 37884 19294 38334 19346
rect 38386 19294 38388 19346
rect 37884 19292 38388 19294
rect 37436 19282 37492 19292
rect 37324 19236 37380 19246
rect 37212 18788 37268 18798
rect 37212 18674 37268 18732
rect 37212 18622 37214 18674
rect 37266 18622 37268 18674
rect 37212 18610 37268 18622
rect 36988 18564 37044 18574
rect 36988 18470 37044 18508
rect 36540 18386 36596 18396
rect 36428 18340 36484 18350
rect 36428 16324 36484 18284
rect 37324 18338 37380 19180
rect 37324 18286 37326 18338
rect 37378 18286 37380 18338
rect 37324 18274 37380 18286
rect 37436 18450 37492 18462
rect 37436 18398 37438 18450
rect 37490 18398 37492 18450
rect 37436 17554 37492 18398
rect 37548 17892 37604 19292
rect 38332 19282 38388 19292
rect 37660 19236 37716 19246
rect 38780 19236 38836 19246
rect 37660 19234 37828 19236
rect 37660 19182 37662 19234
rect 37714 19182 37828 19234
rect 37660 19180 37828 19182
rect 37660 19170 37716 19180
rect 37772 18340 37828 19180
rect 38780 19142 38836 19180
rect 37884 18564 37940 18574
rect 37884 18470 37940 18508
rect 38892 18564 38948 18574
rect 38332 18452 38388 18462
rect 38332 18358 38388 18396
rect 38892 18450 38948 18508
rect 38892 18398 38894 18450
rect 38946 18398 38948 18450
rect 38892 18386 38948 18398
rect 37884 18340 37940 18350
rect 37772 18284 37884 18340
rect 37884 18246 37940 18284
rect 38556 18340 38612 18350
rect 37548 17798 37604 17836
rect 38556 17666 38612 18284
rect 38556 17614 38558 17666
rect 38610 17614 38612 17666
rect 38556 17602 38612 17614
rect 38780 17668 38836 17678
rect 38780 17574 38836 17612
rect 37436 17502 37438 17554
rect 37490 17502 37492 17554
rect 36540 17442 36596 17454
rect 36540 17390 36542 17442
rect 36594 17390 36596 17442
rect 36540 17108 36596 17390
rect 37100 17444 37156 17454
rect 37100 17350 37156 17388
rect 37436 17220 37492 17502
rect 38332 17556 38388 17566
rect 38108 17444 38164 17454
rect 37436 17164 37828 17220
rect 36540 17042 36596 17052
rect 37548 16994 37604 17006
rect 37548 16942 37550 16994
rect 37602 16942 37604 16994
rect 36764 16884 36820 16894
rect 36820 16828 36932 16884
rect 36764 16790 36820 16828
rect 36428 16258 36484 16268
rect 36876 15540 36932 16828
rect 37324 16660 37380 16670
rect 37212 16658 37380 16660
rect 37212 16606 37326 16658
rect 37378 16606 37380 16658
rect 37212 16604 37380 16606
rect 37100 16100 37156 16110
rect 37212 16100 37268 16604
rect 37324 16594 37380 16604
rect 37100 16098 37268 16100
rect 37100 16046 37102 16098
rect 37154 16046 37268 16098
rect 37100 16044 37268 16046
rect 37324 16100 37380 16110
rect 37548 16100 37604 16942
rect 37380 16044 37604 16100
rect 37660 16658 37716 16670
rect 37660 16606 37662 16658
rect 37714 16606 37716 16658
rect 36876 15484 37044 15540
rect 36876 15314 36932 15326
rect 36876 15262 36878 15314
rect 36930 15262 36932 15314
rect 36540 15202 36596 15214
rect 36540 15150 36542 15202
rect 36594 15150 36596 15202
rect 36316 15092 36484 15148
rect 36092 14588 36372 14644
rect 36204 14420 36260 14430
rect 35980 14418 36260 14420
rect 35980 14366 36206 14418
rect 36258 14366 36260 14418
rect 35980 14364 36260 14366
rect 35644 14254 35646 14306
rect 35698 14254 35700 14306
rect 35644 13972 35700 14254
rect 35420 13794 35476 13804
rect 35532 13916 35700 13972
rect 36204 13972 36260 14364
rect 35084 13682 35140 13692
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35532 13188 35588 13916
rect 36204 13906 36260 13916
rect 36316 14306 36372 14588
rect 36316 14254 36318 14306
rect 36370 14254 36372 14306
rect 35644 13746 35700 13758
rect 35644 13694 35646 13746
rect 35698 13694 35700 13746
rect 35644 13636 35700 13694
rect 35644 13570 35700 13580
rect 35084 13132 35588 13188
rect 35084 12962 35140 13132
rect 35084 12910 35086 12962
rect 35138 12910 35140 12962
rect 35084 11620 35140 12910
rect 35308 12852 35364 12862
rect 35308 12758 35364 12796
rect 36316 12740 36372 14254
rect 36428 14084 36484 15092
rect 36540 14532 36596 15150
rect 36540 14466 36596 14476
rect 36876 14644 36932 15262
rect 36988 15092 37044 15484
rect 36988 15026 37044 15036
rect 36764 14420 36820 14430
rect 36540 14308 36596 14318
rect 36764 14308 36820 14364
rect 36540 14306 36820 14308
rect 36540 14254 36542 14306
rect 36594 14254 36820 14306
rect 36540 14252 36820 14254
rect 36540 14242 36596 14252
rect 36428 14028 36820 14084
rect 36652 13748 36708 13758
rect 36204 12684 36372 12740
rect 36428 13746 36708 13748
rect 36428 13694 36654 13746
rect 36706 13694 36708 13746
rect 36428 13692 36708 13694
rect 36428 12852 36484 13692
rect 36652 13682 36708 13692
rect 36764 13524 36820 14028
rect 36876 13634 36932 14588
rect 36988 14644 37044 14654
rect 37100 14644 37156 16044
rect 37324 16006 37380 16044
rect 37660 15876 37716 16606
rect 37772 16212 37828 17164
rect 37996 16212 38052 16222
rect 37772 16210 38052 16212
rect 37772 16158 37998 16210
rect 38050 16158 38052 16210
rect 37772 16156 38052 16158
rect 37996 16146 38052 16156
rect 37660 15810 37716 15820
rect 37660 15652 37716 15662
rect 37324 15316 37380 15326
rect 37324 15222 37380 15260
rect 37660 15314 37716 15596
rect 37660 15262 37662 15314
rect 37714 15262 37716 15314
rect 37660 15250 37716 15262
rect 37772 15426 37828 15438
rect 37772 15374 37774 15426
rect 37826 15374 37828 15426
rect 37772 15316 37828 15374
rect 37772 15250 37828 15260
rect 38108 14756 38164 17388
rect 38332 17106 38388 17500
rect 38332 17054 38334 17106
rect 38386 17054 38388 17106
rect 38332 17042 38388 17054
rect 38780 17444 38836 17454
rect 38668 16658 38724 16670
rect 38668 16606 38670 16658
rect 38722 16606 38724 16658
rect 38668 16100 38724 16606
rect 38780 16210 38836 17388
rect 38780 16158 38782 16210
rect 38834 16158 38836 16210
rect 38780 16146 38836 16158
rect 38892 16770 38948 16782
rect 38892 16718 38894 16770
rect 38946 16718 38948 16770
rect 38668 16034 38724 16044
rect 38892 15540 38948 16718
rect 38892 15474 38948 15484
rect 39004 15148 39060 19404
rect 39228 19234 39284 19246
rect 39228 19182 39230 19234
rect 39282 19182 39284 19234
rect 39116 18788 39172 18798
rect 39116 18674 39172 18732
rect 39116 18622 39118 18674
rect 39170 18622 39172 18674
rect 39116 18610 39172 18622
rect 39228 17668 39284 19182
rect 39676 19010 39732 19022
rect 39676 18958 39678 19010
rect 39730 18958 39732 19010
rect 39676 18564 39732 18958
rect 39676 18498 39732 18508
rect 39900 18562 39956 19516
rect 40572 19348 40628 19358
rect 40236 19292 40572 19348
rect 40012 19012 40068 19022
rect 40236 19012 40292 19292
rect 40572 19254 40628 19292
rect 40012 19010 40292 19012
rect 40012 18958 40014 19010
rect 40066 18958 40292 19010
rect 40012 18956 40292 18958
rect 40012 18946 40068 18956
rect 39900 18510 39902 18562
rect 39954 18510 39956 18562
rect 39900 18498 39956 18510
rect 40236 18450 40292 18956
rect 40236 18398 40238 18450
rect 40290 18398 40292 18450
rect 40236 18386 40292 18398
rect 40348 18340 40404 18350
rect 40348 18246 40404 18284
rect 40796 17778 40852 19964
rect 41132 19908 41188 20638
rect 42476 20130 42532 20142
rect 42476 20078 42478 20130
rect 42530 20078 42532 20130
rect 41356 20020 41412 20030
rect 41356 19926 41412 19964
rect 42364 20018 42420 20030
rect 42364 19966 42366 20018
rect 42418 19966 42420 20018
rect 41132 19842 41188 19852
rect 41692 19908 41748 19918
rect 41692 19814 41748 19852
rect 42364 19908 42420 19966
rect 42364 19842 42420 19852
rect 42476 20020 42532 20078
rect 42476 19684 42532 19964
rect 42252 19628 42532 19684
rect 42588 20132 42980 20188
rect 41020 19348 41076 19358
rect 41020 19254 41076 19292
rect 42028 19236 42084 19246
rect 42252 19236 42308 19628
rect 42364 19460 42420 19470
rect 42588 19460 42644 20132
rect 42924 20130 42980 20132
rect 42924 20078 42926 20130
rect 42978 20078 42980 20130
rect 42700 20020 42756 20030
rect 42700 19926 42756 19964
rect 42924 19908 42980 20078
rect 42924 19842 42980 19852
rect 43036 19796 43092 23102
rect 43708 23154 43764 23166
rect 43708 23102 43710 23154
rect 43762 23102 43764 23154
rect 43372 22930 43428 22942
rect 43372 22878 43374 22930
rect 43426 22878 43428 22930
rect 43372 22372 43428 22878
rect 43596 22372 43652 22382
rect 43708 22372 43764 23102
rect 43932 23156 43988 23166
rect 43932 23062 43988 23100
rect 43372 22370 43764 22372
rect 43372 22318 43598 22370
rect 43650 22318 43764 22370
rect 43372 22316 43764 22318
rect 43372 21924 43428 21934
rect 43372 20802 43428 21868
rect 43596 21364 43652 22316
rect 43932 22258 43988 22270
rect 43932 22206 43934 22258
rect 43986 22206 43988 22258
rect 43932 21924 43988 22206
rect 43708 21868 43988 21924
rect 43708 21812 43764 21868
rect 44044 21812 44100 23326
rect 44268 23154 44324 23166
rect 44268 23102 44270 23154
rect 44322 23102 44324 23154
rect 44268 22484 44324 23102
rect 44268 21924 44324 22428
rect 44604 22820 44660 22830
rect 44268 21858 44324 21868
rect 44492 21924 44548 21934
rect 43708 21586 43764 21756
rect 43708 21534 43710 21586
rect 43762 21534 43764 21586
rect 43708 21522 43764 21534
rect 43932 21756 44100 21812
rect 43932 21474 43988 21756
rect 44380 21588 44436 21598
rect 43932 21422 43934 21474
rect 43986 21422 43988 21474
rect 43932 21410 43988 21422
rect 44044 21586 44436 21588
rect 44044 21534 44382 21586
rect 44434 21534 44436 21586
rect 44044 21532 44436 21534
rect 43596 21308 43876 21364
rect 43372 20750 43374 20802
rect 43426 20750 43428 20802
rect 43148 20020 43204 20030
rect 43148 19926 43204 19964
rect 43260 19908 43316 19918
rect 43372 19908 43428 20750
rect 43708 20804 43764 20814
rect 43708 20710 43764 20748
rect 43820 20692 43876 21308
rect 44044 21026 44100 21532
rect 44380 21522 44436 21532
rect 44044 20974 44046 21026
rect 44098 20974 44100 21026
rect 44044 20962 44100 20974
rect 43932 20692 43988 20702
rect 43820 20690 43988 20692
rect 43820 20638 43934 20690
rect 43986 20638 43988 20690
rect 43820 20636 43988 20638
rect 43932 20626 43988 20636
rect 43820 20132 43876 20142
rect 43820 20038 43876 20076
rect 43260 19906 43428 19908
rect 43260 19854 43262 19906
rect 43314 19854 43428 19906
rect 43260 19852 43428 19854
rect 43484 20018 43540 20030
rect 43484 19966 43486 20018
rect 43538 19966 43540 20018
rect 43260 19842 43316 19852
rect 43484 19796 43540 19966
rect 43596 20020 43652 20030
rect 43596 19926 43652 19964
rect 43932 20018 43988 20030
rect 43932 19966 43934 20018
rect 43986 19966 43988 20018
rect 43932 19908 43988 19966
rect 43932 19842 43988 19852
rect 44156 20018 44212 20030
rect 44156 19966 44158 20018
rect 44210 19966 44212 20018
rect 43036 19740 43204 19796
rect 42364 19458 42644 19460
rect 42364 19406 42366 19458
rect 42418 19406 42644 19458
rect 42364 19404 42644 19406
rect 42812 19460 42868 19470
rect 42364 19394 42420 19404
rect 42812 19366 42868 19404
rect 42588 19236 42644 19246
rect 43036 19236 43092 19740
rect 43148 19572 43204 19740
rect 43484 19730 43540 19740
rect 44156 19796 44212 19966
rect 43596 19684 43652 19694
rect 43148 19516 43540 19572
rect 42252 19234 42644 19236
rect 42252 19182 42590 19234
rect 42642 19182 42644 19234
rect 42252 19180 42644 19182
rect 42028 19142 42084 19180
rect 42588 19170 42644 19180
rect 42700 19180 43092 19236
rect 43484 19234 43540 19516
rect 43484 19182 43486 19234
rect 43538 19182 43540 19234
rect 41804 19124 41860 19134
rect 41804 19030 41860 19068
rect 42252 19012 42308 19022
rect 42700 19012 42756 19180
rect 43484 19170 43540 19182
rect 42252 19010 42756 19012
rect 42252 18958 42254 19010
rect 42306 18958 42756 19010
rect 42252 18956 42756 18958
rect 43148 19012 43204 19022
rect 42252 18946 42308 18956
rect 42364 18674 42420 18956
rect 43148 18918 43204 18956
rect 42364 18622 42366 18674
rect 42418 18622 42420 18674
rect 42364 18610 42420 18622
rect 41132 18450 41188 18462
rect 41132 18398 41134 18450
rect 41186 18398 41188 18450
rect 41132 17780 41188 18398
rect 41916 18452 41972 18462
rect 40796 17726 40798 17778
rect 40850 17726 40852 17778
rect 40796 17714 40852 17726
rect 40908 17724 41188 17780
rect 41356 18340 41412 18350
rect 39228 17444 39284 17612
rect 40348 17668 40404 17678
rect 40348 17574 40404 17612
rect 39228 17378 39284 17388
rect 39564 16996 39620 17006
rect 39452 15876 39508 15886
rect 39452 15314 39508 15820
rect 39452 15262 39454 15314
rect 39506 15262 39508 15314
rect 39452 15250 39508 15262
rect 39564 15148 39620 16940
rect 39788 16884 39844 16894
rect 39788 16790 39844 16828
rect 40460 16884 40516 16894
rect 40460 16790 40516 16828
rect 39900 16772 39956 16782
rect 39900 16678 39956 16716
rect 39004 15092 39172 15148
rect 38108 14690 38164 14700
rect 36988 14642 37156 14644
rect 36988 14590 36990 14642
rect 37042 14590 37156 14642
rect 36988 14588 37156 14590
rect 38332 14644 38388 14654
rect 36988 14578 37044 14588
rect 37212 14532 37268 14542
rect 37212 14418 37268 14476
rect 37212 14366 37214 14418
rect 37266 14366 37268 14418
rect 36876 13582 36878 13634
rect 36930 13582 36932 13634
rect 36876 13570 36932 13582
rect 37100 13972 37156 13982
rect 36204 12290 36260 12684
rect 36428 12628 36484 12796
rect 36204 12238 36206 12290
rect 36258 12238 36260 12290
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 36204 11620 36260 12238
rect 36316 12572 36484 12628
rect 36652 13468 36820 13524
rect 36316 12066 36372 12572
rect 36316 12014 36318 12066
rect 36370 12014 36372 12066
rect 36316 12002 36372 12014
rect 36428 12180 36484 12190
rect 36316 11620 36372 11630
rect 35084 11564 35364 11620
rect 36204 11564 36316 11620
rect 34860 11454 34862 11506
rect 34914 11454 34916 11506
rect 34860 11442 34916 11454
rect 34076 10610 34132 10668
rect 34412 11394 34468 11406
rect 34412 11342 34414 11394
rect 34466 11342 34468 11394
rect 34076 10558 34078 10610
rect 34130 10558 34132 10610
rect 34076 10546 34132 10558
rect 34300 10612 34356 10622
rect 34412 10612 34468 11342
rect 35308 10836 35364 11564
rect 36316 11554 36372 11564
rect 36204 11396 36260 11406
rect 36428 11396 36484 12124
rect 36204 11394 36484 11396
rect 36204 11342 36206 11394
rect 36258 11342 36484 11394
rect 36204 11340 36484 11342
rect 36204 11330 36260 11340
rect 36540 11284 36596 11294
rect 36540 11190 36596 11228
rect 36316 11172 36372 11182
rect 36316 11078 36372 11116
rect 35420 10836 35476 10846
rect 35308 10780 35420 10836
rect 35420 10770 35476 10780
rect 35084 10612 35140 10622
rect 34412 10610 35140 10612
rect 34412 10558 35086 10610
rect 35138 10558 35140 10610
rect 34412 10556 35140 10558
rect 34300 9940 34356 10556
rect 34860 9940 34916 10556
rect 35084 10546 35140 10556
rect 36428 10612 36484 10622
rect 36428 10518 36484 10556
rect 36540 10498 36596 10510
rect 36540 10446 36542 10498
rect 36594 10446 36596 10498
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 34300 9884 34468 9940
rect 33964 9380 34020 9390
rect 33964 9044 34020 9324
rect 34300 9268 34356 9278
rect 34412 9268 34468 9884
rect 34860 9846 34916 9884
rect 35420 10052 35476 10062
rect 34748 9826 34804 9838
rect 34748 9774 34750 9826
rect 34802 9774 34804 9826
rect 34300 9266 34468 9268
rect 34300 9214 34302 9266
rect 34354 9214 34468 9266
rect 34300 9212 34468 9214
rect 34524 9714 34580 9726
rect 34524 9662 34526 9714
rect 34578 9662 34580 9714
rect 34300 9202 34356 9212
rect 34188 9044 34244 9054
rect 33964 9042 34188 9044
rect 33964 8990 33966 9042
rect 34018 8990 34188 9042
rect 33964 8988 34188 8990
rect 33964 8978 34020 8988
rect 34076 8258 34132 8270
rect 34076 8206 34078 8258
rect 34130 8206 34132 8258
rect 34076 7476 34132 8206
rect 34188 7698 34244 8988
rect 34524 8708 34580 9662
rect 34748 9716 34804 9774
rect 35084 9828 35140 9838
rect 35084 9734 35140 9772
rect 35420 9826 35476 9996
rect 35420 9774 35422 9826
rect 35474 9774 35476 9826
rect 35420 9762 35476 9774
rect 35644 9828 35700 9838
rect 34748 9650 34804 9660
rect 35420 9604 35476 9614
rect 35420 9510 35476 9548
rect 35196 9268 35252 9278
rect 35196 9174 35252 9212
rect 35308 9154 35364 9166
rect 35308 9102 35310 9154
rect 35362 9102 35364 9154
rect 35308 8820 35364 9102
rect 35644 9042 35700 9772
rect 35756 9716 35812 9726
rect 35756 9714 36148 9716
rect 35756 9662 35758 9714
rect 35810 9662 36148 9714
rect 35756 9660 36148 9662
rect 35756 9650 35812 9660
rect 36092 9266 36148 9660
rect 36092 9214 36094 9266
rect 36146 9214 36148 9266
rect 36092 9202 36148 9214
rect 36540 9268 36596 10446
rect 36540 9154 36596 9212
rect 36540 9102 36542 9154
rect 36594 9102 36596 9154
rect 36540 9090 36596 9102
rect 35644 8990 35646 9042
rect 35698 8990 35700 9042
rect 35644 8978 35700 8990
rect 35868 9044 35924 9054
rect 35868 8950 35924 8988
rect 36204 9042 36260 9054
rect 36204 8990 36206 9042
rect 36258 8990 36260 9042
rect 34524 8642 34580 8652
rect 35084 8764 35364 8820
rect 34412 8484 34468 8494
rect 34412 8390 34468 8428
rect 34188 7646 34190 7698
rect 34242 7646 34244 7698
rect 34188 7634 34244 7646
rect 34300 8258 34356 8270
rect 34300 8206 34302 8258
rect 34354 8206 34356 8258
rect 34300 7588 34356 8206
rect 34860 8036 34916 8046
rect 34860 7698 34916 7980
rect 34860 7646 34862 7698
rect 34914 7646 34916 7698
rect 34860 7634 34916 7646
rect 34300 7522 34356 7532
rect 34076 7410 34132 7420
rect 34636 7474 34692 7486
rect 34636 7422 34638 7474
rect 34690 7422 34692 7474
rect 34636 7252 34692 7422
rect 34636 7186 34692 7196
rect 33852 6402 33908 6412
rect 34300 6692 34356 6702
rect 34188 6020 34244 6030
rect 34188 5926 34244 5964
rect 34076 5908 34132 5918
rect 33796 5906 34132 5908
rect 33796 5854 34078 5906
rect 34130 5854 34132 5906
rect 33796 5852 34132 5854
rect 33740 5814 33796 5852
rect 33516 5742 33518 5794
rect 33570 5742 33572 5794
rect 33516 5730 33572 5742
rect 33068 5282 33124 5292
rect 33516 5236 33572 5246
rect 33516 5142 33572 5180
rect 32676 3500 32788 3556
rect 32956 4788 33012 4798
rect 32620 3490 32676 3500
rect 32956 800 33012 4732
rect 33964 4450 34020 5852
rect 34076 5842 34132 5852
rect 34300 5572 34356 6636
rect 35084 6692 35140 8764
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 36204 8484 36260 8990
rect 36204 8418 36260 8428
rect 36428 8372 36484 8382
rect 36428 8278 36484 8316
rect 35532 8258 35588 8270
rect 35532 8206 35534 8258
rect 35586 8206 35588 8258
rect 35532 8036 35588 8206
rect 35756 8260 35812 8270
rect 35756 8166 35812 8204
rect 36092 8148 36148 8158
rect 35532 7970 35588 7980
rect 35980 8146 36148 8148
rect 35980 8094 36094 8146
rect 36146 8094 36148 8146
rect 35980 8092 36148 8094
rect 35644 7476 35700 7486
rect 35868 7476 35924 7486
rect 35532 7474 35700 7476
rect 35532 7422 35646 7474
rect 35698 7422 35700 7474
rect 35532 7420 35700 7422
rect 35308 7252 35364 7290
rect 35308 7186 35364 7196
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35084 6626 35140 6636
rect 34524 6578 34580 6590
rect 34524 6526 34526 6578
rect 34578 6526 34580 6578
rect 34412 5908 34468 5918
rect 34412 5814 34468 5852
rect 34300 4788 34356 5516
rect 34524 5684 34580 6526
rect 34524 4900 34580 5628
rect 34524 4834 34580 4844
rect 34636 6468 34692 6478
rect 34412 4788 34468 4798
rect 34300 4732 34412 4788
rect 33964 4398 33966 4450
rect 34018 4398 34020 4450
rect 33964 4340 34020 4398
rect 33964 4274 34020 4284
rect 34412 4338 34468 4732
rect 34412 4286 34414 4338
rect 34466 4286 34468 4338
rect 34412 4274 34468 4286
rect 33628 4116 33684 4126
rect 33628 800 33684 4060
rect 34636 3554 34692 6412
rect 34972 6018 35028 6030
rect 34972 5966 34974 6018
rect 35026 5966 35028 6018
rect 34860 4452 34916 4462
rect 34860 4358 34916 4396
rect 34972 4226 35028 5966
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 34972 4174 34974 4226
rect 35026 4174 35028 4226
rect 34972 4162 35028 4174
rect 35084 5012 35140 5022
rect 34636 3502 34638 3554
rect 34690 3502 34692 3554
rect 34636 3490 34692 3502
rect 34972 3780 35028 3790
rect 34300 2548 34356 2558
rect 34300 800 34356 2492
rect 34972 800 35028 3724
rect 35084 3442 35140 4956
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 35308 3556 35364 3566
rect 35308 3462 35364 3500
rect 35084 3390 35086 3442
rect 35138 3390 35140 3442
rect 35084 3378 35140 3390
rect 35532 3220 35588 7420
rect 35644 7410 35700 7420
rect 35756 7474 35924 7476
rect 35756 7422 35870 7474
rect 35922 7422 35924 7474
rect 35756 7420 35924 7422
rect 35644 6580 35700 6590
rect 35644 5124 35700 6524
rect 35756 5348 35812 7420
rect 35868 7410 35924 7420
rect 35868 6804 35924 6814
rect 35980 6804 36036 8092
rect 36092 8082 36148 8092
rect 36316 8036 36372 8046
rect 36372 7980 36484 8036
rect 36316 7942 36372 7980
rect 35924 6748 36036 6804
rect 36204 7474 36260 7486
rect 36204 7422 36206 7474
rect 36258 7422 36260 7474
rect 35868 6130 35924 6748
rect 35868 6078 35870 6130
rect 35922 6078 35924 6130
rect 35868 6066 35924 6078
rect 36092 6578 36148 6590
rect 36092 6526 36094 6578
rect 36146 6526 36148 6578
rect 36092 5906 36148 6526
rect 36204 6356 36260 7422
rect 36204 6290 36260 6300
rect 36316 7474 36372 7486
rect 36316 7422 36318 7474
rect 36370 7422 36372 7474
rect 36092 5854 36094 5906
rect 36146 5854 36148 5906
rect 36092 5842 36148 5854
rect 36316 6132 36372 7422
rect 36428 7476 36484 7980
rect 36428 7410 36484 7420
rect 36540 7252 36596 7262
rect 36428 6468 36484 6478
rect 36428 6374 36484 6412
rect 35756 5282 35812 5292
rect 35868 5796 35924 5806
rect 35868 5234 35924 5740
rect 35868 5182 35870 5234
rect 35922 5182 35924 5234
rect 35868 5170 35924 5182
rect 35756 5124 35812 5134
rect 35644 5068 35756 5124
rect 35756 5030 35812 5068
rect 35980 4900 36036 4910
rect 35532 3154 35588 3164
rect 35644 3668 35700 3678
rect 35644 800 35700 3612
rect 35980 3332 36036 4844
rect 36204 4900 36260 4910
rect 36204 4806 36260 4844
rect 36316 4564 36372 6076
rect 36540 5906 36596 7196
rect 36540 5854 36542 5906
rect 36594 5854 36596 5906
rect 36540 5842 36596 5854
rect 36652 5684 36708 13468
rect 36764 13300 36820 13310
rect 36764 12290 36820 13244
rect 37100 12738 37156 13916
rect 37212 13524 37268 14366
rect 38332 14530 38388 14588
rect 38332 14478 38334 14530
rect 38386 14478 38388 14530
rect 37772 14308 37828 14318
rect 37548 13748 37604 13758
rect 37548 13654 37604 13692
rect 37772 13746 37828 14252
rect 37772 13694 37774 13746
rect 37826 13694 37828 13746
rect 37772 13682 37828 13694
rect 38332 13748 38388 14478
rect 38668 14420 38724 14430
rect 38668 14326 38724 14364
rect 37212 13458 37268 13468
rect 38220 13524 38276 13534
rect 38220 12962 38276 13468
rect 38220 12910 38222 12962
rect 38274 12910 38276 12962
rect 38220 12898 38276 12910
rect 38332 12850 38388 13692
rect 38332 12798 38334 12850
rect 38386 12798 38388 12850
rect 38332 12786 38388 12798
rect 38444 13860 38500 13870
rect 37100 12686 37102 12738
rect 37154 12686 37156 12738
rect 37100 12628 37156 12686
rect 37100 12562 37156 12572
rect 38108 12740 38164 12750
rect 37660 12516 37716 12526
rect 37660 12402 37716 12460
rect 37660 12350 37662 12402
rect 37714 12350 37716 12402
rect 37660 12338 37716 12350
rect 36764 12238 36766 12290
rect 36818 12238 36820 12290
rect 36764 12068 36820 12238
rect 37100 12180 37156 12190
rect 37548 12180 37604 12190
rect 37156 12178 37604 12180
rect 37156 12126 37550 12178
rect 37602 12126 37604 12178
rect 37156 12124 37604 12126
rect 37100 12086 37156 12124
rect 36764 12002 36820 12012
rect 37548 11844 37604 12124
rect 37548 11778 37604 11788
rect 37884 12178 37940 12190
rect 38108 12180 38164 12684
rect 38444 12628 38500 13804
rect 38556 12852 38612 12862
rect 38556 12758 38612 12796
rect 38780 12740 38836 12750
rect 38780 12646 38836 12684
rect 37884 12126 37886 12178
rect 37938 12126 37940 12178
rect 36540 5628 36708 5684
rect 36764 11620 36820 11630
rect 36428 5236 36484 5246
rect 36428 5122 36484 5180
rect 36428 5070 36430 5122
rect 36482 5070 36484 5122
rect 36428 5058 36484 5070
rect 36316 4338 36372 4508
rect 36316 4286 36318 4338
rect 36370 4286 36372 4338
rect 36316 4274 36372 4286
rect 35980 3266 36036 3276
rect 36316 3892 36372 3902
rect 36316 800 36372 3836
rect 36428 3556 36484 3566
rect 36540 3556 36596 5628
rect 36764 5236 36820 11564
rect 37772 11394 37828 11406
rect 37772 11342 37774 11394
rect 37826 11342 37828 11394
rect 37324 11284 37380 11294
rect 37324 11190 37380 11228
rect 37436 10836 37492 10846
rect 37436 10386 37492 10780
rect 37772 10500 37828 11342
rect 37884 10724 37940 12126
rect 37884 10658 37940 10668
rect 37996 12178 38164 12180
rect 37996 12126 38110 12178
rect 38162 12126 38164 12178
rect 37996 12124 38164 12126
rect 37996 11172 38052 12124
rect 38108 12114 38164 12124
rect 38220 12572 38500 12628
rect 38220 11956 38276 12572
rect 38332 12292 38388 12302
rect 38332 12198 38388 12236
rect 38892 12292 38948 12302
rect 38892 12198 38948 12236
rect 38444 12180 38500 12190
rect 38444 12086 38500 12124
rect 37772 10434 37828 10444
rect 37436 10334 37438 10386
rect 37490 10334 37492 10386
rect 37436 10322 37492 10334
rect 37996 10164 38052 11116
rect 38108 11900 38276 11956
rect 38108 10610 38164 11900
rect 38892 11396 38948 11406
rect 38892 11302 38948 11340
rect 38220 10836 38276 10846
rect 38220 10722 38276 10780
rect 38220 10670 38222 10722
rect 38274 10670 38276 10722
rect 38220 10658 38276 10670
rect 38332 10668 38668 10724
rect 38108 10558 38110 10610
rect 38162 10558 38164 10610
rect 38108 10388 38164 10558
rect 38108 10332 38276 10388
rect 37996 10098 38052 10108
rect 38220 10052 38276 10332
rect 38108 9996 38276 10052
rect 37100 9938 37156 9950
rect 37100 9886 37102 9938
rect 37154 9886 37156 9938
rect 37100 9716 37156 9886
rect 37548 9828 37604 9838
rect 37548 9734 37604 9772
rect 37884 9716 37940 9726
rect 37100 9380 37156 9660
rect 37660 9660 37884 9716
rect 37100 9324 37380 9380
rect 37212 9156 37268 9166
rect 37212 9062 37268 9100
rect 36988 9042 37044 9054
rect 36988 8990 36990 9042
rect 37042 8990 37044 9042
rect 36988 7700 37044 8990
rect 37100 8372 37156 8382
rect 37100 8278 37156 8316
rect 37324 8372 37380 9324
rect 37324 8306 37380 8316
rect 37660 9154 37716 9660
rect 37884 9622 37940 9660
rect 37884 9268 37940 9278
rect 37660 9102 37662 9154
rect 37714 9102 37716 9154
rect 37660 8146 37716 9102
rect 37772 9156 37828 9166
rect 37772 9062 37828 9100
rect 37884 9042 37940 9212
rect 37884 8990 37886 9042
rect 37938 8990 37940 9042
rect 37660 8094 37662 8146
rect 37714 8094 37716 8146
rect 37660 8082 37716 8094
rect 37772 8260 37828 8270
rect 36988 7644 37156 7700
rect 37100 7586 37156 7644
rect 37100 7534 37102 7586
rect 37154 7534 37156 7586
rect 36988 7476 37044 7486
rect 36988 6802 37044 7420
rect 36988 6750 36990 6802
rect 37042 6750 37044 6802
rect 36988 6738 37044 6750
rect 37100 6244 37156 7534
rect 37212 7474 37268 7486
rect 37212 7422 37214 7474
rect 37266 7422 37268 7474
rect 37212 6804 37268 7422
rect 37548 7476 37604 7486
rect 37548 7382 37604 7420
rect 37436 6916 37492 6926
rect 37436 6822 37492 6860
rect 37212 6710 37268 6748
rect 37100 6178 37156 6188
rect 37772 5906 37828 8204
rect 37884 6914 37940 8990
rect 38108 8484 38164 9996
rect 38108 8418 38164 8428
rect 38220 9828 38276 9838
rect 38220 7140 38276 9772
rect 38332 9266 38388 10668
rect 38612 10612 38668 10668
rect 39004 10612 39060 10622
rect 38612 10610 39060 10612
rect 38612 10558 39006 10610
rect 39058 10558 39060 10610
rect 38612 10556 39060 10558
rect 39004 10546 39060 10556
rect 38444 10500 38500 10510
rect 38444 10498 38612 10500
rect 38444 10446 38446 10498
rect 38498 10446 38612 10498
rect 38444 10444 38612 10446
rect 38444 10434 38500 10444
rect 38556 10276 38612 10444
rect 38556 10210 38612 10220
rect 38332 9214 38334 9266
rect 38386 9214 38388 9266
rect 38332 9202 38388 9214
rect 38444 10164 38500 10174
rect 38444 9826 38500 10108
rect 38892 9940 38948 9950
rect 38892 9846 38948 9884
rect 38444 9774 38446 9826
rect 38498 9774 38500 9826
rect 38444 7252 38500 9774
rect 38780 9602 38836 9614
rect 38780 9550 38782 9602
rect 38834 9550 38836 9602
rect 38668 9268 38724 9278
rect 38668 9154 38724 9212
rect 38780 9266 38836 9550
rect 39004 9604 39060 9614
rect 39004 9510 39060 9548
rect 38780 9214 38782 9266
rect 38834 9214 38836 9266
rect 38780 9202 38836 9214
rect 38668 9102 38670 9154
rect 38722 9102 38724 9154
rect 38668 9090 38724 9102
rect 39004 9156 39060 9166
rect 39004 9062 39060 9100
rect 38556 8258 38612 8270
rect 38556 8206 38558 8258
rect 38610 8206 38612 8258
rect 38556 7476 38612 8206
rect 39004 7476 39060 7486
rect 38556 7474 38724 7476
rect 38556 7422 38558 7474
rect 38610 7422 38724 7474
rect 38556 7420 38724 7422
rect 38556 7410 38612 7420
rect 38444 7186 38500 7196
rect 38220 7074 38276 7084
rect 37884 6862 37886 6914
rect 37938 6862 37940 6914
rect 37884 6850 37940 6862
rect 38556 7028 38612 7038
rect 38556 6578 38612 6972
rect 38556 6526 38558 6578
rect 38610 6526 38612 6578
rect 38556 6514 38612 6526
rect 38668 6916 38724 7420
rect 38668 6018 38724 6860
rect 39004 6690 39060 7420
rect 39004 6638 39006 6690
rect 39058 6638 39060 6690
rect 39004 6626 39060 6638
rect 39116 6692 39172 15092
rect 39340 15092 39620 15148
rect 39788 16100 39844 16110
rect 39340 13076 39396 15092
rect 39788 14754 39844 16044
rect 40908 15764 40964 17724
rect 41356 17668 41412 18284
rect 41244 17666 41412 17668
rect 41244 17614 41358 17666
rect 41410 17614 41412 17666
rect 41244 17612 41412 17614
rect 41244 17332 41300 17612
rect 41356 17602 41412 17612
rect 41468 18338 41524 18350
rect 41468 18286 41470 18338
rect 41522 18286 41524 18338
rect 41020 17276 41300 17332
rect 41020 15986 41076 17276
rect 41020 15934 41022 15986
rect 41074 15934 41076 15986
rect 41020 15922 41076 15934
rect 41132 16210 41188 16222
rect 41132 16158 41134 16210
rect 41186 16158 41188 16210
rect 41132 15764 41188 16158
rect 40908 15708 41188 15764
rect 39900 15540 39956 15550
rect 39900 15446 39956 15484
rect 41132 15540 41188 15708
rect 41132 15202 41188 15484
rect 41468 16100 41524 18286
rect 41692 18340 41748 18350
rect 41692 18246 41748 18284
rect 41468 15314 41524 16044
rect 41580 16994 41636 17006
rect 41580 16942 41582 16994
rect 41634 16942 41636 16994
rect 41580 16098 41636 16942
rect 41580 16046 41582 16098
rect 41634 16046 41636 16098
rect 41580 16034 41636 16046
rect 41692 16770 41748 16782
rect 41692 16718 41694 16770
rect 41746 16718 41748 16770
rect 41692 15428 41748 16718
rect 41804 16212 41860 16222
rect 41804 15986 41860 16156
rect 41916 16098 41972 18396
rect 42140 18450 42196 18462
rect 42140 18398 42142 18450
rect 42194 18398 42196 18450
rect 42140 17332 42196 18398
rect 42812 18452 42868 18462
rect 42252 18340 42308 18350
rect 42252 17778 42308 18284
rect 42700 18340 42756 18350
rect 42812 18340 42868 18396
rect 43148 18450 43204 18462
rect 43148 18398 43150 18450
rect 43202 18398 43204 18450
rect 42700 18338 42868 18340
rect 42700 18286 42702 18338
rect 42754 18286 42868 18338
rect 42700 18284 42868 18286
rect 43036 18338 43092 18350
rect 43036 18286 43038 18338
rect 43090 18286 43092 18338
rect 42700 18274 42756 18284
rect 42252 17726 42254 17778
rect 42306 17726 42308 17778
rect 42252 17714 42308 17726
rect 42476 17668 42532 17678
rect 42476 17574 42532 17612
rect 42140 17276 42308 17332
rect 42140 17108 42196 17118
rect 41916 16046 41918 16098
rect 41970 16046 41972 16098
rect 41916 16034 41972 16046
rect 42028 16772 42084 16782
rect 41804 15934 41806 15986
rect 41858 15934 41860 15986
rect 41804 15922 41860 15934
rect 41692 15362 41748 15372
rect 41468 15262 41470 15314
rect 41522 15262 41524 15314
rect 41468 15250 41524 15262
rect 42028 15316 42084 16716
rect 41132 15150 41134 15202
rect 41186 15150 41188 15202
rect 41132 15138 41188 15150
rect 39788 14702 39790 14754
rect 39842 14702 39844 14754
rect 39788 14690 39844 14702
rect 41132 14530 41188 14542
rect 41132 14478 41134 14530
rect 41186 14478 41188 14530
rect 41132 13972 41188 14478
rect 42028 14418 42084 15260
rect 42028 14366 42030 14418
rect 42082 14366 42084 14418
rect 42028 14354 42084 14366
rect 41132 13916 41748 13972
rect 39564 13748 39620 13758
rect 39564 13654 39620 13692
rect 41132 13748 41188 13758
rect 40124 13636 40180 13646
rect 40124 13542 40180 13580
rect 39788 13524 39844 13534
rect 39844 13468 39956 13524
rect 39788 13430 39844 13468
rect 39340 13074 39844 13076
rect 39340 13022 39342 13074
rect 39394 13022 39844 13074
rect 39340 13020 39844 13022
rect 39340 13010 39396 13020
rect 39676 12852 39732 12862
rect 39676 12758 39732 12796
rect 39340 12404 39396 12414
rect 39340 12290 39396 12348
rect 39340 12238 39342 12290
rect 39394 12238 39396 12290
rect 39340 12226 39396 12238
rect 39788 12290 39844 13020
rect 39788 12238 39790 12290
rect 39842 12238 39844 12290
rect 39788 12226 39844 12238
rect 39900 11618 39956 13468
rect 41132 13074 41188 13692
rect 41132 13022 41134 13074
rect 41186 13022 41188 13074
rect 41132 13010 41188 13022
rect 41244 13746 41300 13758
rect 41244 13694 41246 13746
rect 41298 13694 41300 13746
rect 40124 12962 40180 12974
rect 40124 12910 40126 12962
rect 40178 12910 40180 12962
rect 39900 11566 39902 11618
rect 39954 11566 39956 11618
rect 39900 11554 39956 11566
rect 40012 12628 40068 12638
rect 40012 11508 40068 12572
rect 40124 12402 40180 12910
rect 40124 12350 40126 12402
rect 40178 12350 40180 12402
rect 40124 12338 40180 12350
rect 40460 12516 40516 12526
rect 40012 11442 40068 11452
rect 40236 12180 40292 12190
rect 40236 11506 40292 12124
rect 40236 11454 40238 11506
rect 40290 11454 40292 11506
rect 40236 11442 40292 11454
rect 40348 11396 40404 11406
rect 39564 10724 39620 10734
rect 39228 10722 39620 10724
rect 39228 10670 39566 10722
rect 39618 10670 39620 10722
rect 39228 10668 39620 10670
rect 39228 9716 39284 10668
rect 39564 10658 39620 10668
rect 39788 10610 39844 10622
rect 39788 10558 39790 10610
rect 39842 10558 39844 10610
rect 39452 10386 39508 10398
rect 39452 10334 39454 10386
rect 39506 10334 39508 10386
rect 39452 9826 39508 10334
rect 39452 9774 39454 9826
rect 39506 9774 39508 9826
rect 39452 9762 39508 9774
rect 39228 9154 39284 9660
rect 39228 9102 39230 9154
rect 39282 9102 39284 9154
rect 39228 9090 39284 9102
rect 39340 9156 39396 9166
rect 39340 7586 39396 9100
rect 39788 9156 39844 10558
rect 40012 10610 40068 10622
rect 40012 10558 40014 10610
rect 40066 10558 40068 10610
rect 40012 9268 40068 10558
rect 40348 9380 40404 11340
rect 40012 9202 40068 9212
rect 40124 9324 40404 9380
rect 39788 9090 39844 9100
rect 40124 8932 40180 9324
rect 40348 9156 40404 9166
rect 40348 9062 40404 9100
rect 39900 8818 39956 8830
rect 39900 8766 39902 8818
rect 39954 8766 39956 8818
rect 39452 8484 39508 8494
rect 39452 8390 39508 8428
rect 39340 7534 39342 7586
rect 39394 7534 39396 7586
rect 39340 7522 39396 7534
rect 39788 7812 39844 7822
rect 39116 6626 39172 6636
rect 39228 7474 39284 7486
rect 39228 7422 39230 7474
rect 39282 7422 39284 7474
rect 39228 6132 39284 7422
rect 39452 7476 39508 7486
rect 39452 7382 39508 7420
rect 39228 6066 39284 6076
rect 39452 6692 39508 6702
rect 38668 5966 38670 6018
rect 38722 5966 38724 6018
rect 38668 5954 38724 5966
rect 37772 5854 37774 5906
rect 37826 5854 37828 5906
rect 36764 5170 36820 5180
rect 37436 5234 37492 5246
rect 37436 5182 37438 5234
rect 37490 5182 37492 5234
rect 36652 5124 36708 5134
rect 36652 4450 36708 5068
rect 36652 4398 36654 4450
rect 36706 4398 36708 4450
rect 36652 4386 36708 4398
rect 36988 4340 37044 4350
rect 36988 4246 37044 4284
rect 36988 3668 37044 3678
rect 36988 3574 37044 3612
rect 36428 3554 36596 3556
rect 36428 3502 36430 3554
rect 36482 3502 36596 3554
rect 36428 3500 36596 3502
rect 36428 3490 36484 3500
rect 37436 3388 37492 5182
rect 37772 4562 37828 5854
rect 39340 5906 39396 5918
rect 39340 5854 39342 5906
rect 39394 5854 39396 5906
rect 39340 5460 39396 5854
rect 39004 5348 39060 5358
rect 37772 4510 37774 4562
rect 37826 4510 37828 4562
rect 37772 4498 37828 4510
rect 38892 5124 38948 5134
rect 37100 3332 37492 3388
rect 37660 4004 37716 4014
rect 37100 980 37156 3332
rect 36988 924 37156 980
rect 36988 800 37044 924
rect 37660 800 37716 3948
rect 38332 3556 38388 3566
rect 38332 800 38388 3500
rect 38892 3442 38948 5068
rect 39004 4450 39060 5292
rect 39228 5236 39284 5246
rect 39004 4398 39006 4450
rect 39058 4398 39060 4450
rect 39004 3668 39060 4398
rect 39004 3602 39060 3612
rect 39116 4788 39172 4798
rect 39116 3554 39172 4732
rect 39228 4564 39284 5180
rect 39228 4338 39284 4508
rect 39228 4286 39230 4338
rect 39282 4286 39284 4338
rect 39228 4274 39284 4286
rect 39116 3502 39118 3554
rect 39170 3502 39172 3554
rect 39116 3490 39172 3502
rect 39340 3556 39396 5404
rect 39452 5124 39508 6636
rect 39788 6244 39844 7756
rect 39900 7476 39956 8766
rect 40012 8818 40068 8830
rect 40012 8766 40014 8818
rect 40066 8766 40068 8818
rect 40012 8260 40068 8766
rect 40012 8194 40068 8204
rect 40124 8036 40180 8876
rect 39900 7382 39956 7420
rect 40012 7980 40180 8036
rect 40236 8818 40292 8830
rect 40236 8766 40238 8818
rect 40290 8766 40292 8818
rect 40236 8034 40292 8766
rect 40236 7982 40238 8034
rect 40290 7982 40292 8034
rect 40012 6356 40068 7980
rect 40236 7588 40292 7982
rect 40460 8146 40516 12460
rect 41244 11732 41300 13694
rect 41580 13746 41636 13758
rect 41580 13694 41582 13746
rect 41634 13694 41636 13746
rect 41468 13636 41524 13646
rect 41468 13188 41524 13580
rect 41356 13132 41468 13188
rect 41356 12178 41412 13132
rect 41468 13122 41524 13132
rect 41580 12740 41636 13694
rect 41356 12126 41358 12178
rect 41410 12126 41412 12178
rect 41356 12114 41412 12126
rect 41468 12292 41524 12302
rect 41580 12292 41636 12684
rect 41524 12236 41636 12292
rect 41692 12962 41748 13916
rect 41692 12910 41694 12962
rect 41746 12910 41748 12962
rect 41468 12178 41524 12236
rect 41468 12126 41470 12178
rect 41522 12126 41524 12178
rect 41468 12114 41524 12126
rect 41244 11666 41300 11676
rect 40908 11396 40964 11406
rect 40908 11394 41188 11396
rect 40908 11342 40910 11394
rect 40962 11342 41188 11394
rect 40908 11340 41188 11342
rect 40908 11330 40964 11340
rect 40572 10724 40628 10734
rect 40572 9714 40628 10668
rect 41132 9940 41188 11340
rect 41244 10836 41300 10846
rect 41692 10836 41748 12910
rect 41804 13524 41860 13534
rect 41804 12402 41860 13468
rect 41916 13522 41972 13534
rect 41916 13470 41918 13522
rect 41970 13470 41972 13522
rect 41916 12852 41972 13470
rect 41916 12786 41972 12796
rect 41804 12350 41806 12402
rect 41858 12350 41860 12402
rect 41804 12338 41860 12350
rect 41916 12066 41972 12078
rect 41916 12014 41918 12066
rect 41970 12014 41972 12066
rect 41916 11732 41972 12014
rect 41972 11676 42084 11732
rect 41916 11638 41972 11676
rect 41244 10834 41748 10836
rect 41244 10782 41246 10834
rect 41298 10782 41748 10834
rect 41244 10780 41748 10782
rect 41244 10770 41300 10780
rect 41580 10610 41636 10622
rect 41580 10558 41582 10610
rect 41634 10558 41636 10610
rect 40572 9662 40574 9714
rect 40626 9662 40628 9714
rect 40572 9650 40628 9662
rect 40796 9826 40852 9838
rect 40796 9774 40798 9826
rect 40850 9774 40852 9826
rect 40796 9380 40852 9774
rect 40796 9324 41076 9380
rect 40908 9042 40964 9054
rect 40908 8990 40910 9042
rect 40962 8990 40964 9042
rect 40908 8932 40964 8990
rect 41020 9044 41076 9324
rect 41020 8950 41076 8988
rect 41132 9042 41188 9884
rect 41468 10500 41524 10510
rect 41244 9156 41300 9166
rect 41300 9100 41412 9156
rect 41244 9090 41300 9100
rect 41132 8990 41134 9042
rect 41186 8990 41188 9042
rect 41132 8978 41188 8990
rect 41356 9042 41412 9100
rect 41356 8990 41358 9042
rect 41410 8990 41412 9042
rect 41356 8978 41412 8990
rect 40908 8866 40964 8876
rect 41468 8820 41524 10444
rect 41244 8764 41524 8820
rect 41580 9940 41636 10558
rect 41580 9826 41636 9884
rect 41580 9774 41582 9826
rect 41634 9774 41636 9826
rect 40796 8372 40852 8382
rect 40796 8258 40852 8316
rect 40796 8206 40798 8258
rect 40850 8206 40852 8258
rect 40796 8194 40852 8206
rect 41132 8260 41188 8270
rect 40460 8094 40462 8146
rect 40514 8094 40516 8146
rect 40460 7812 40516 8094
rect 40460 7746 40516 7756
rect 41132 7700 41188 8204
rect 41132 7634 41188 7644
rect 40236 7028 40292 7532
rect 40236 6962 40292 6972
rect 40348 7532 40740 7588
rect 40348 6802 40404 7532
rect 40684 7476 40740 7532
rect 41132 7476 41188 7486
rect 40684 7474 41188 7476
rect 40684 7422 41134 7474
rect 41186 7422 41188 7474
rect 40684 7420 41188 7422
rect 41132 7410 41188 7420
rect 41244 7362 41300 8764
rect 41244 7310 41246 7362
rect 41298 7310 41300 7362
rect 41244 7298 41300 7310
rect 41468 7364 41524 7374
rect 40348 6750 40350 6802
rect 40402 6750 40404 6802
rect 40348 6738 40404 6750
rect 40684 7252 40740 7262
rect 40124 6580 40180 6590
rect 40124 6578 40628 6580
rect 40124 6526 40126 6578
rect 40178 6526 40628 6578
rect 40124 6524 40628 6526
rect 40124 6514 40180 6524
rect 40012 6300 40180 6356
rect 39788 6188 40068 6244
rect 39788 6020 39844 6188
rect 40012 6130 40068 6188
rect 40012 6078 40014 6130
rect 40066 6078 40068 6130
rect 40012 6066 40068 6078
rect 39788 5954 39844 5964
rect 39452 5030 39508 5068
rect 39564 5796 39620 5806
rect 39564 3780 39620 5740
rect 40124 5234 40180 6300
rect 40236 5906 40292 5918
rect 40236 5854 40238 5906
rect 40290 5854 40292 5906
rect 40236 5348 40292 5854
rect 40236 5282 40292 5292
rect 40124 5182 40126 5234
rect 40178 5182 40180 5234
rect 40124 5170 40180 5182
rect 40348 5124 40404 5134
rect 40348 4562 40404 5068
rect 40572 5124 40628 6524
rect 40684 6578 40740 7196
rect 40684 6526 40686 6578
rect 40738 6526 40740 6578
rect 40684 6514 40740 6526
rect 41020 6580 41076 6590
rect 41020 6486 41076 6524
rect 41356 6244 41412 6254
rect 40908 6132 40964 6142
rect 40964 6076 41076 6132
rect 40908 6066 40964 6076
rect 40572 5030 40628 5068
rect 41020 6018 41076 6076
rect 41020 5966 41022 6018
rect 41074 5966 41076 6018
rect 40348 4510 40350 4562
rect 40402 4510 40404 4562
rect 40348 4498 40404 4510
rect 40908 4452 40964 4462
rect 40908 4358 40964 4396
rect 40012 3780 40068 3790
rect 39564 3778 40068 3780
rect 39564 3726 40014 3778
rect 40066 3726 40068 3778
rect 39564 3724 40068 3726
rect 40012 3714 40068 3724
rect 40348 3668 40404 3678
rect 40908 3668 40964 3678
rect 41020 3668 41076 5966
rect 41356 5908 41412 6188
rect 41468 6020 41524 7308
rect 41580 6802 41636 9774
rect 42028 9602 42084 11676
rect 42028 9550 42030 9602
rect 42082 9550 42084 9602
rect 42028 9538 42084 9550
rect 41804 9042 41860 9054
rect 41804 8990 41806 9042
rect 41858 8990 41860 9042
rect 41580 6750 41582 6802
rect 41634 6750 41636 6802
rect 41580 6738 41636 6750
rect 41692 8034 41748 8046
rect 41692 7982 41694 8034
rect 41746 7982 41748 8034
rect 41692 6132 41748 7982
rect 41804 8036 41860 8990
rect 42028 9042 42084 9054
rect 42028 8990 42030 9042
rect 42082 8990 42084 9042
rect 42028 8148 42084 8990
rect 42028 8082 42084 8092
rect 41804 7970 41860 7980
rect 42140 7364 42196 17052
rect 42252 16996 42308 17276
rect 42252 16212 42308 16940
rect 43036 16996 43092 18286
rect 43036 16902 43092 16940
rect 42252 16146 42308 16156
rect 43148 15428 43204 18398
rect 43596 17106 43652 19628
rect 43708 19236 43764 19246
rect 43708 19142 43764 19180
rect 43820 19124 43876 19134
rect 43820 18452 43876 19068
rect 44156 18900 44212 19740
rect 44268 19124 44324 19162
rect 44268 19058 44324 19068
rect 44268 18900 44324 18910
rect 44156 18844 44268 18900
rect 44268 18834 44324 18844
rect 44156 18564 44212 18574
rect 44156 18470 44212 18508
rect 44268 18564 44324 18574
rect 44492 18564 44548 21868
rect 44604 21474 44660 22764
rect 45276 22596 45332 23548
rect 45276 22530 45332 22540
rect 45388 23156 45444 23166
rect 45164 22484 45220 22494
rect 45164 22390 45220 22428
rect 44828 22372 44884 22382
rect 44828 22278 44884 22316
rect 45388 22370 45444 23100
rect 46284 22820 46340 23886
rect 46284 22754 46340 22764
rect 46396 23154 46452 23166
rect 46396 23102 46398 23154
rect 46450 23102 46452 23154
rect 46396 23044 46452 23102
rect 46396 22596 46452 22988
rect 45388 22318 45390 22370
rect 45442 22318 45444 22370
rect 45388 21812 45444 22318
rect 46060 22540 46452 22596
rect 45948 22258 46004 22270
rect 45948 22206 45950 22258
rect 46002 22206 46004 22258
rect 45948 21924 46004 22206
rect 46060 22258 46116 22540
rect 46060 22206 46062 22258
rect 46114 22206 46116 22258
rect 46060 22194 46116 22206
rect 46284 22372 46340 22382
rect 45948 21858 46004 21868
rect 45164 21756 45444 21812
rect 44604 21422 44606 21474
rect 44658 21422 44660 21474
rect 44604 21410 44660 21422
rect 45052 21700 45108 21710
rect 45164 21700 45220 21756
rect 45052 21698 45220 21700
rect 45052 21646 45054 21698
rect 45106 21646 45220 21698
rect 45052 21644 45220 21646
rect 46284 21698 46340 22316
rect 46620 21924 46676 25452
rect 46732 25442 46788 25452
rect 47180 25508 47236 25518
rect 47516 25508 47572 26236
rect 47796 26236 47908 26292
rect 47740 26198 47796 26236
rect 47628 25508 47684 25518
rect 47516 25506 47684 25508
rect 47516 25454 47630 25506
rect 47682 25454 47684 25506
rect 47516 25452 47684 25454
rect 47180 25414 47236 25452
rect 47628 25442 47684 25452
rect 47404 25396 47460 25406
rect 47404 25302 47460 25340
rect 47852 25394 47908 26236
rect 49084 26066 49140 27022
rect 49196 26964 49252 27806
rect 49196 26898 49252 26908
rect 49980 27804 50316 27860
rect 49980 26850 50036 27804
rect 50316 27794 50372 27804
rect 50988 27858 51044 28588
rect 51100 28550 51156 28588
rect 51772 28642 51828 28654
rect 51772 28590 51774 28642
rect 51826 28590 51828 28642
rect 51772 28196 51828 28590
rect 51772 28130 51828 28140
rect 51996 28642 52052 28654
rect 51996 28590 51998 28642
rect 52050 28590 52052 28642
rect 50988 27806 50990 27858
rect 51042 27806 51044 27858
rect 49980 26798 49982 26850
rect 50034 26798 50036 26850
rect 49980 26786 50036 26798
rect 50204 27074 50260 27086
rect 50204 27022 50206 27074
rect 50258 27022 50260 27074
rect 50204 26516 50260 27022
rect 50988 27074 51044 27806
rect 51212 27860 51268 27870
rect 51884 27860 51940 27870
rect 51212 27766 51268 27804
rect 51660 27858 51940 27860
rect 51660 27806 51886 27858
rect 51938 27806 51940 27858
rect 51660 27804 51940 27806
rect 51996 27860 52052 28590
rect 55580 28644 55636 28654
rect 55580 28550 55636 28588
rect 57932 28308 57988 28702
rect 57932 28242 57988 28252
rect 52780 28196 52836 28206
rect 52668 28084 52724 28094
rect 52668 27990 52724 28028
rect 52108 27860 52164 27870
rect 51996 27804 52108 27860
rect 50988 27022 50990 27074
rect 51042 27022 51044 27074
rect 50988 27010 51044 27022
rect 50556 26684 50820 26694
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50556 26618 50820 26628
rect 49868 26460 50260 26516
rect 51660 26514 51716 27804
rect 51884 27794 51940 27804
rect 52108 27746 52164 27804
rect 52108 27694 52110 27746
rect 52162 27694 52164 27746
rect 52108 27682 52164 27694
rect 52556 27858 52612 27870
rect 52556 27806 52558 27858
rect 52610 27806 52612 27858
rect 51772 27244 52052 27300
rect 51772 27186 51828 27244
rect 51772 27134 51774 27186
rect 51826 27134 51828 27186
rect 51772 27122 51828 27134
rect 51660 26462 51662 26514
rect 51714 26462 51716 26514
rect 49644 26290 49700 26302
rect 49644 26238 49646 26290
rect 49698 26238 49700 26290
rect 49084 26014 49086 26066
rect 49138 26014 49140 26066
rect 49084 26002 49140 26014
rect 49420 26178 49476 26190
rect 49420 26126 49422 26178
rect 49474 26126 49476 26178
rect 49420 25956 49476 26126
rect 47964 25620 48020 25630
rect 47964 25506 48020 25564
rect 47964 25454 47966 25506
rect 48018 25454 48020 25506
rect 47964 25442 48020 25454
rect 48636 25508 48692 25518
rect 49420 25508 49476 25900
rect 49644 25732 49700 26238
rect 49644 25666 49700 25676
rect 49756 26068 49812 26078
rect 49532 25508 49588 25518
rect 49420 25506 49588 25508
rect 49420 25454 49534 25506
rect 49586 25454 49588 25506
rect 49420 25452 49588 25454
rect 48636 25414 48692 25452
rect 49532 25442 49588 25452
rect 47852 25342 47854 25394
rect 47906 25342 47908 25394
rect 47852 25330 47908 25342
rect 48412 25396 48468 25406
rect 47740 24612 47796 24622
rect 46732 23940 46788 23950
rect 46732 23938 46900 23940
rect 46732 23886 46734 23938
rect 46786 23886 46900 23938
rect 46732 23884 46900 23886
rect 46732 23874 46788 23884
rect 46732 23716 46788 23726
rect 46732 23378 46788 23660
rect 46844 23492 46900 23884
rect 47516 23938 47572 23950
rect 47516 23886 47518 23938
rect 47570 23886 47572 23938
rect 47516 23716 47572 23886
rect 47516 23650 47572 23660
rect 47740 23714 47796 24556
rect 48412 24050 48468 25340
rect 49644 25396 49700 25406
rect 48860 25284 48916 25294
rect 48860 25190 48916 25228
rect 49644 24948 49700 25340
rect 49756 25394 49812 26012
rect 49868 25956 49924 26460
rect 51660 26450 51716 26462
rect 51884 27074 51940 27086
rect 51884 27022 51886 27074
rect 51938 27022 51940 27074
rect 50316 26404 50372 26414
rect 50316 26310 50372 26348
rect 51884 26402 51940 27022
rect 51884 26350 51886 26402
rect 51938 26350 51940 26402
rect 50092 26292 50148 26302
rect 50092 26198 50148 26236
rect 50428 26290 50484 26302
rect 50428 26238 50430 26290
rect 50482 26238 50484 26290
rect 49868 25900 50036 25956
rect 49980 25618 50036 25900
rect 49980 25566 49982 25618
rect 50034 25566 50036 25618
rect 49980 25554 50036 25566
rect 50316 25732 50372 25742
rect 49756 25342 49758 25394
rect 49810 25342 49812 25394
rect 49756 25284 49812 25342
rect 49868 25508 49924 25518
rect 49868 25284 49924 25452
rect 50204 25508 50260 25518
rect 50204 25414 50260 25452
rect 50316 25506 50372 25676
rect 50316 25454 50318 25506
rect 50370 25454 50372 25506
rect 50316 25442 50372 25454
rect 50428 25396 50484 26238
rect 51884 25732 51940 26350
rect 51996 26404 52052 27244
rect 51996 26310 52052 26348
rect 52444 26852 52500 26862
rect 52444 26402 52500 26796
rect 52556 26514 52612 27806
rect 52668 27188 52724 27198
rect 52780 27188 52836 28140
rect 53228 28196 53284 28206
rect 53228 27970 53284 28140
rect 53228 27918 53230 27970
rect 53282 27918 53284 27970
rect 53228 27906 53284 27918
rect 53116 27860 53172 27870
rect 53116 27766 53172 27804
rect 57596 27746 57652 27758
rect 57596 27694 57598 27746
rect 57650 27694 57652 27746
rect 52668 27186 52836 27188
rect 52668 27134 52670 27186
rect 52722 27134 52836 27186
rect 52668 27132 52836 27134
rect 54348 27132 54628 27188
rect 52668 27122 52724 27132
rect 53116 27076 53172 27086
rect 52892 27074 53172 27076
rect 52892 27022 53118 27074
rect 53170 27022 53172 27074
rect 52892 27020 53172 27022
rect 52892 26852 52948 27020
rect 53116 27010 53172 27020
rect 53564 27074 53620 27086
rect 53564 27022 53566 27074
rect 53618 27022 53620 27074
rect 53564 26964 53620 27022
rect 52892 26786 52948 26796
rect 53116 26852 53620 26908
rect 54348 26962 54404 27132
rect 54348 26910 54350 26962
rect 54402 26910 54404 26962
rect 54348 26898 54404 26910
rect 54460 26964 54516 27002
rect 54460 26898 54516 26908
rect 53116 26628 53172 26852
rect 52556 26462 52558 26514
rect 52610 26462 52612 26514
rect 52556 26450 52612 26462
rect 52668 26572 53172 26628
rect 52444 26350 52446 26402
rect 52498 26350 52500 26402
rect 52444 26180 52500 26350
rect 52668 26402 52724 26572
rect 52668 26350 52670 26402
rect 52722 26350 52724 26402
rect 52668 26338 52724 26350
rect 53116 26402 53172 26414
rect 53116 26350 53118 26402
rect 53170 26350 53172 26402
rect 52892 26290 52948 26302
rect 52892 26238 52894 26290
rect 52946 26238 52948 26290
rect 52892 26180 52948 26238
rect 52444 26124 52948 26180
rect 53116 26068 53172 26350
rect 54124 26404 54180 26414
rect 54124 26310 54180 26348
rect 53228 26292 53284 26302
rect 53564 26292 53620 26302
rect 53228 26290 53564 26292
rect 53228 26238 53230 26290
rect 53282 26238 53564 26290
rect 53228 26236 53564 26238
rect 53228 26226 53284 26236
rect 51884 25666 51940 25676
rect 52780 25732 52836 25742
rect 52780 25638 52836 25676
rect 52108 25620 52164 25630
rect 52164 25564 52276 25620
rect 52108 25554 52164 25564
rect 50652 25508 50708 25518
rect 50652 25414 50708 25452
rect 51548 25508 51604 25518
rect 49980 25284 50036 25294
rect 50428 25284 50484 25340
rect 49868 25228 49980 25284
rect 49756 25218 49812 25228
rect 49980 25218 50036 25228
rect 50204 25228 50484 25284
rect 50540 25284 50596 25322
rect 49420 24892 49700 24948
rect 49084 24724 49140 24734
rect 49084 24630 49140 24668
rect 49420 24722 49476 24892
rect 49980 24724 50036 24734
rect 49420 24670 49422 24722
rect 49474 24670 49476 24722
rect 49420 24658 49476 24670
rect 49868 24668 49980 24724
rect 49644 24612 49700 24622
rect 49644 24610 49812 24612
rect 49644 24558 49646 24610
rect 49698 24558 49812 24610
rect 49644 24556 49812 24558
rect 49644 24546 49700 24556
rect 48412 23998 48414 24050
rect 48466 23998 48468 24050
rect 48412 23986 48468 23998
rect 49084 23940 49140 23950
rect 49084 23938 49700 23940
rect 49084 23886 49086 23938
rect 49138 23886 49700 23938
rect 49084 23884 49700 23886
rect 49084 23874 49140 23884
rect 47740 23662 47742 23714
rect 47794 23662 47796 23714
rect 47740 23604 47796 23662
rect 47740 23538 47796 23548
rect 46844 23436 47348 23492
rect 46732 23326 46734 23378
rect 46786 23326 46788 23378
rect 46732 23314 46788 23326
rect 47068 23266 47124 23278
rect 47068 23214 47070 23266
rect 47122 23214 47124 23266
rect 47068 22820 47124 23214
rect 47292 23156 47348 23436
rect 48076 23380 48132 23390
rect 48076 23286 48132 23324
rect 47404 23156 47460 23166
rect 47292 23154 47460 23156
rect 47292 23102 47406 23154
rect 47458 23102 47460 23154
rect 47292 23100 47460 23102
rect 47068 22754 47124 22764
rect 47404 22148 47460 23100
rect 48188 23154 48244 23166
rect 48188 23102 48190 23154
rect 48242 23102 48244 23154
rect 47628 22652 47908 22708
rect 47516 22372 47572 22382
rect 47516 22278 47572 22316
rect 47404 22082 47460 22092
rect 46620 21858 46676 21868
rect 47180 21700 47236 21710
rect 46284 21646 46286 21698
rect 46338 21646 46340 21698
rect 45052 20804 45108 21644
rect 46284 21634 46340 21646
rect 47068 21644 47180 21700
rect 45052 20738 45108 20748
rect 45276 21586 45332 21598
rect 45276 21534 45278 21586
rect 45330 21534 45332 21586
rect 45276 20692 45332 21534
rect 45948 21476 46004 21486
rect 45948 21474 46116 21476
rect 45948 21422 45950 21474
rect 46002 21422 46116 21474
rect 45948 21420 46116 21422
rect 45948 21410 46004 21420
rect 46060 21026 46116 21420
rect 46060 20974 46062 21026
rect 46114 20974 46116 21026
rect 46060 20962 46116 20974
rect 46172 20860 46900 20916
rect 45276 19346 45332 20636
rect 45948 20692 46004 20702
rect 45948 20598 46004 20636
rect 46060 20692 46116 20702
rect 46172 20692 46228 20860
rect 46060 20690 46228 20692
rect 46060 20638 46062 20690
rect 46114 20638 46228 20690
rect 46060 20636 46228 20638
rect 46060 20626 46116 20636
rect 46284 19458 46340 20860
rect 46844 20804 46900 20860
rect 46956 20804 47012 20814
rect 46844 20802 47012 20804
rect 46844 20750 46958 20802
rect 47010 20750 47012 20802
rect 46844 20748 47012 20750
rect 46956 20738 47012 20748
rect 46732 20692 46788 20702
rect 46732 20598 46788 20636
rect 46956 20580 47012 20590
rect 47068 20580 47124 21644
rect 47180 21634 47236 21644
rect 46956 20578 47124 20580
rect 46956 20526 46958 20578
rect 47010 20526 47124 20578
rect 46956 20524 47124 20526
rect 47292 21586 47348 21598
rect 47292 21534 47294 21586
rect 47346 21534 47348 21586
rect 47292 20690 47348 21534
rect 47292 20638 47294 20690
rect 47346 20638 47348 20690
rect 46956 20514 47012 20524
rect 46284 19406 46286 19458
rect 46338 19406 46340 19458
rect 46284 19394 46340 19406
rect 45276 19294 45278 19346
rect 45330 19294 45332 19346
rect 45276 19282 45332 19294
rect 45612 19348 45668 19358
rect 45164 19234 45220 19246
rect 45164 19182 45166 19234
rect 45218 19182 45220 19234
rect 45052 19124 45108 19134
rect 45164 19124 45220 19182
rect 45108 19068 45220 19124
rect 45052 19058 45108 19068
rect 44940 19010 44996 19022
rect 44940 18958 44942 19010
rect 44994 18958 44996 19010
rect 44940 18674 44996 18958
rect 45388 19012 45444 19022
rect 45388 18918 45444 18956
rect 44940 18622 44942 18674
rect 44994 18622 44996 18674
rect 44940 18610 44996 18622
rect 45164 18900 45220 18910
rect 44268 18562 44548 18564
rect 44268 18510 44270 18562
rect 44322 18510 44548 18562
rect 44268 18508 44548 18510
rect 43820 18386 43876 18396
rect 44156 18228 44212 18238
rect 44156 18134 44212 18172
rect 43596 17054 43598 17106
rect 43650 17054 43652 17106
rect 43596 17042 43652 17054
rect 43484 16324 43540 16334
rect 43148 15362 43204 15372
rect 43260 16322 43540 16324
rect 43260 16270 43486 16322
rect 43538 16270 43540 16322
rect 43260 16268 43540 16270
rect 42924 15316 42980 15326
rect 42924 15222 42980 15260
rect 42476 14642 42532 14654
rect 42476 14590 42478 14642
rect 42530 14590 42532 14642
rect 42364 13188 42420 13198
rect 42364 13094 42420 13132
rect 42476 13074 42532 14590
rect 43036 14420 43092 14430
rect 43036 13748 43092 14364
rect 43036 13682 43092 13692
rect 43148 14306 43204 14318
rect 43148 14254 43150 14306
rect 43202 14254 43204 14306
rect 43148 13634 43204 14254
rect 43260 13860 43316 16268
rect 43484 16258 43540 16268
rect 44044 16100 44100 16110
rect 44044 16098 44212 16100
rect 44044 16046 44046 16098
rect 44098 16046 44212 16098
rect 44044 16044 44212 16046
rect 44044 16034 44100 16044
rect 43372 15988 43428 15998
rect 43372 15894 43428 15932
rect 43484 15876 43540 15886
rect 43484 15782 43540 15820
rect 44156 15876 44212 16044
rect 44268 15986 44324 18508
rect 45164 17778 45220 18844
rect 45276 18452 45332 18462
rect 45276 18358 45332 18396
rect 45164 17726 45166 17778
rect 45218 17726 45220 17778
rect 45164 17714 45220 17726
rect 45276 17668 45332 17678
rect 45276 16098 45332 17612
rect 45276 16046 45278 16098
rect 45330 16046 45332 16098
rect 44268 15934 44270 15986
rect 44322 15934 44324 15986
rect 44268 15922 44324 15934
rect 44940 15988 44996 15998
rect 44940 15894 44996 15932
rect 43596 15316 43652 15326
rect 43596 15202 43652 15260
rect 43596 15150 43598 15202
rect 43650 15150 43652 15202
rect 43596 15138 43652 15150
rect 43932 15314 43988 15326
rect 43932 15262 43934 15314
rect 43986 15262 43988 15314
rect 43820 14756 43876 14766
rect 43372 14754 43876 14756
rect 43372 14702 43822 14754
rect 43874 14702 43876 14754
rect 43372 14700 43876 14702
rect 43372 14530 43428 14700
rect 43372 14478 43374 14530
rect 43426 14478 43428 14530
rect 43372 14466 43428 14478
rect 43260 13794 43316 13804
rect 43148 13582 43150 13634
rect 43202 13582 43204 13634
rect 43148 13570 43204 13582
rect 43484 13186 43540 14700
rect 43820 14690 43876 14700
rect 43708 14532 43764 14542
rect 43708 14438 43764 14476
rect 43596 13860 43652 13870
rect 43596 13766 43652 13804
rect 43932 13524 43988 15262
rect 44044 14530 44100 14542
rect 44044 14478 44046 14530
rect 44098 14478 44100 14530
rect 44044 14420 44100 14478
rect 44044 14354 44100 14364
rect 43932 13458 43988 13468
rect 43484 13134 43486 13186
rect 43538 13134 43540 13186
rect 43484 13122 43540 13134
rect 44156 13076 44212 15820
rect 44380 15202 44436 15214
rect 44380 15150 44382 15202
rect 44434 15150 44436 15202
rect 44268 14530 44324 14542
rect 44268 14478 44270 14530
rect 44322 14478 44324 14530
rect 44268 13748 44324 14478
rect 44380 14420 44436 15150
rect 44940 14532 44996 14542
rect 44940 14438 44996 14476
rect 44380 14354 44436 14364
rect 44716 13748 44772 13758
rect 44268 13746 44772 13748
rect 44268 13694 44718 13746
rect 44770 13694 44772 13746
rect 44268 13692 44772 13694
rect 42476 13022 42478 13074
rect 42530 13022 42532 13074
rect 42476 13010 42532 13022
rect 43708 13020 44212 13076
rect 42588 12740 42644 12750
rect 42588 12646 42644 12684
rect 42700 12404 42756 12414
rect 42700 12310 42756 12348
rect 43372 12404 43428 12414
rect 43372 12310 43428 12348
rect 43708 12402 43764 13020
rect 44156 12964 44212 13020
rect 44156 12962 44660 12964
rect 44156 12910 44158 12962
rect 44210 12910 44660 12962
rect 44156 12908 44660 12910
rect 44156 12898 44212 12908
rect 43708 12350 43710 12402
rect 43762 12350 43764 12402
rect 43708 12338 43764 12350
rect 43932 12850 43988 12862
rect 43932 12798 43934 12850
rect 43986 12798 43988 12850
rect 42924 12178 42980 12190
rect 42924 12126 42926 12178
rect 42978 12126 42980 12178
rect 42924 12068 42980 12126
rect 43932 12180 43988 12798
rect 44044 12850 44100 12862
rect 44044 12798 44046 12850
rect 44098 12798 44100 12850
rect 44044 12404 44100 12798
rect 44044 12348 44212 12404
rect 44156 12292 44212 12348
rect 44380 12292 44436 12302
rect 44156 12236 44380 12292
rect 44380 12198 44436 12236
rect 44604 12290 44660 12908
rect 44716 12628 44772 13692
rect 45052 12962 45108 12974
rect 45052 12910 45054 12962
rect 45106 12910 45108 12962
rect 44828 12852 44884 12862
rect 44828 12758 44884 12796
rect 44716 12572 44884 12628
rect 44604 12238 44606 12290
rect 44658 12238 44660 12290
rect 44604 12226 44660 12238
rect 44044 12180 44100 12190
rect 43932 12178 44100 12180
rect 43932 12126 44046 12178
rect 44098 12126 44100 12178
rect 43932 12124 44100 12126
rect 42924 12002 42980 12012
rect 43820 12068 43876 12078
rect 43708 11620 43764 11630
rect 42476 10724 42532 10734
rect 42476 10630 42532 10668
rect 43372 10612 43428 10622
rect 43036 10498 43092 10510
rect 43036 10446 43038 10498
rect 43090 10446 43092 10498
rect 43036 9828 43092 10446
rect 43148 9940 43204 9950
rect 43148 9846 43204 9884
rect 43036 9762 43092 9772
rect 43372 9266 43428 10556
rect 43484 9828 43540 9838
rect 43540 9772 43652 9828
rect 43484 9734 43540 9772
rect 43372 9214 43374 9266
rect 43426 9214 43428 9266
rect 43372 9202 43428 9214
rect 43596 9268 43652 9772
rect 43708 9380 43764 11564
rect 43820 11394 43876 12012
rect 43820 11342 43822 11394
rect 43874 11342 43876 11394
rect 43820 11330 43876 11342
rect 43932 11284 43988 11294
rect 43932 11190 43988 11228
rect 43932 9940 43988 9950
rect 44044 9940 44100 12124
rect 44828 11506 44884 12572
rect 45052 12402 45108 12910
rect 45052 12350 45054 12402
rect 45106 12350 45108 12402
rect 45052 12338 45108 12350
rect 44828 11454 44830 11506
rect 44882 11454 44884 11506
rect 44828 11442 44884 11454
rect 44156 11396 44212 11406
rect 44156 11302 44212 11340
rect 44716 11396 44772 11406
rect 44716 10722 44772 11340
rect 44716 10670 44718 10722
rect 44770 10670 44772 10722
rect 44716 10658 44772 10670
rect 44828 11284 44884 11294
rect 43932 9938 44100 9940
rect 43932 9886 43934 9938
rect 43986 9886 44100 9938
rect 43932 9884 44100 9886
rect 44156 9940 44212 9950
rect 43932 9874 43988 9884
rect 43708 9324 44100 9380
rect 43596 9212 43988 9268
rect 42252 9154 42308 9166
rect 42252 9102 42254 9154
rect 42306 9102 42308 9154
rect 42252 8484 42308 9102
rect 42364 9044 42420 9054
rect 42812 9044 42868 9054
rect 42364 9042 42868 9044
rect 42364 8990 42366 9042
rect 42418 8990 42814 9042
rect 42866 8990 42868 9042
rect 42364 8988 42868 8990
rect 42364 8978 42420 8988
rect 42812 8978 42868 8988
rect 43260 9044 43316 9054
rect 43260 8950 43316 8988
rect 43484 9044 43540 9054
rect 43484 8950 43540 8988
rect 42588 8484 42644 8494
rect 42252 8482 42644 8484
rect 42252 8430 42590 8482
rect 42642 8430 42644 8482
rect 42252 8428 42644 8430
rect 42588 8260 42644 8428
rect 43148 8484 43204 8494
rect 42924 8372 42980 8382
rect 43148 8372 43204 8428
rect 42924 8278 42980 8316
rect 43036 8370 43204 8372
rect 43036 8318 43150 8370
rect 43202 8318 43204 8370
rect 43036 8316 43204 8318
rect 42588 8194 42644 8204
rect 42700 8036 42756 8046
rect 42756 7980 42868 8036
rect 42700 7970 42756 7980
rect 42140 7298 42196 7308
rect 42252 7588 42308 7598
rect 42252 7252 42308 7532
rect 42140 6468 42196 6478
rect 41916 6132 41972 6142
rect 41692 6130 41972 6132
rect 41692 6078 41918 6130
rect 41970 6078 41972 6130
rect 41692 6076 41972 6078
rect 41468 5964 41860 6020
rect 41244 5906 41412 5908
rect 41244 5854 41358 5906
rect 41410 5854 41412 5906
rect 41244 5852 41412 5854
rect 41132 5796 41188 5806
rect 41132 4338 41188 5740
rect 41132 4286 41134 4338
rect 41186 4286 41188 4338
rect 41132 4116 41188 4286
rect 41132 4050 41188 4060
rect 41132 3780 41188 3790
rect 41244 3780 41300 5852
rect 41356 5842 41412 5852
rect 41804 5906 41860 5964
rect 41804 5854 41806 5906
rect 41858 5854 41860 5906
rect 41804 5236 41860 5854
rect 41916 5908 41972 6076
rect 41916 5842 41972 5852
rect 41692 5234 41860 5236
rect 41692 5182 41806 5234
rect 41858 5182 41860 5234
rect 41692 5180 41860 5182
rect 41132 3778 41300 3780
rect 41132 3726 41134 3778
rect 41186 3726 41300 3778
rect 41132 3724 41300 3726
rect 41468 5124 41524 5134
rect 41468 3778 41524 5068
rect 41692 4562 41748 5180
rect 41804 5170 41860 5180
rect 41692 4510 41694 4562
rect 41746 4510 41748 4562
rect 41692 4498 41748 4510
rect 42028 4228 42084 4238
rect 42028 4134 42084 4172
rect 41468 3726 41470 3778
rect 41522 3726 41524 3778
rect 41132 3714 41188 3724
rect 41468 3714 41524 3726
rect 42140 3780 42196 6412
rect 42252 5122 42308 7196
rect 42700 6804 42756 6814
rect 42700 6690 42756 6748
rect 42700 6638 42702 6690
rect 42754 6638 42756 6690
rect 42700 6626 42756 6638
rect 42700 6132 42756 6142
rect 42812 6132 42868 7980
rect 42924 7474 42980 7486
rect 42924 7422 42926 7474
rect 42978 7422 42980 7474
rect 42924 7252 42980 7422
rect 42924 7186 42980 7196
rect 42700 6130 42868 6132
rect 42700 6078 42702 6130
rect 42754 6078 42868 6130
rect 42700 6076 42868 6078
rect 42924 6356 42980 6366
rect 42700 6066 42756 6076
rect 42588 6020 42644 6030
rect 42476 5796 42532 5806
rect 42476 5702 42532 5740
rect 42252 5070 42254 5122
rect 42306 5070 42308 5122
rect 42252 5058 42308 5070
rect 42252 4340 42308 4350
rect 42476 4340 42532 4350
rect 42588 4340 42644 5964
rect 42924 4564 42980 6300
rect 43036 5122 43092 8316
rect 43148 8306 43204 8316
rect 43484 8260 43540 8270
rect 43372 7700 43428 7710
rect 43148 6692 43204 6702
rect 43148 5906 43204 6636
rect 43148 5854 43150 5906
rect 43202 5854 43204 5906
rect 43148 5842 43204 5854
rect 43372 5906 43428 7644
rect 43484 6578 43540 8204
rect 43596 7362 43652 9212
rect 43932 9154 43988 9212
rect 43932 9102 43934 9154
rect 43986 9102 43988 9154
rect 43932 9090 43988 9102
rect 43708 8148 43764 8158
rect 43708 8054 43764 8092
rect 43820 8146 43876 8158
rect 43820 8094 43822 8146
rect 43874 8094 43876 8146
rect 43820 8036 43876 8094
rect 43820 7970 43876 7980
rect 43932 7476 43988 7486
rect 43932 7382 43988 7420
rect 43596 7310 43598 7362
rect 43650 7310 43652 7362
rect 43596 7298 43652 7310
rect 43820 7364 43876 7374
rect 43484 6526 43486 6578
rect 43538 6526 43540 6578
rect 43484 6514 43540 6526
rect 43372 5854 43374 5906
rect 43426 5854 43428 5906
rect 43372 5842 43428 5854
rect 43596 6020 43652 6030
rect 43596 5906 43652 5964
rect 43596 5854 43598 5906
rect 43650 5854 43652 5906
rect 43596 5842 43652 5854
rect 43820 5684 43876 7308
rect 43932 6916 43988 6926
rect 43932 5684 43988 6860
rect 44044 6132 44100 9324
rect 44156 9042 44212 9884
rect 44828 9938 44884 11228
rect 45276 11284 45332 16046
rect 45500 15988 45556 15998
rect 45500 15894 45556 15932
rect 45388 14530 45444 14542
rect 45388 14478 45390 14530
rect 45442 14478 45444 14530
rect 45388 13860 45444 14478
rect 45388 13794 45444 13804
rect 45276 11218 45332 11228
rect 45500 11394 45556 11406
rect 45500 11342 45502 11394
rect 45554 11342 45556 11394
rect 45500 10724 45556 11342
rect 45500 10658 45556 10668
rect 44940 10612 44996 10622
rect 44940 10518 44996 10556
rect 44828 9886 44830 9938
rect 44882 9886 44884 9938
rect 44828 9874 44884 9886
rect 45276 9826 45332 9838
rect 45276 9774 45278 9826
rect 45330 9774 45332 9826
rect 44828 9266 44884 9278
rect 44828 9214 44830 9266
rect 44882 9214 44884 9266
rect 44716 9044 44772 9054
rect 44156 8990 44158 9042
rect 44210 8990 44212 9042
rect 44156 8978 44212 8990
rect 44268 9042 44772 9044
rect 44268 8990 44718 9042
rect 44770 8990 44772 9042
rect 44268 8988 44772 8990
rect 44268 8482 44324 8988
rect 44716 8978 44772 8988
rect 44828 8708 44884 9214
rect 44828 8642 44884 8652
rect 44940 9044 44996 9054
rect 44268 8430 44270 8482
rect 44322 8430 44324 8482
rect 44268 8418 44324 8430
rect 44940 8370 44996 8988
rect 45276 8484 45332 9774
rect 45276 8418 45332 8428
rect 44940 8318 44942 8370
rect 44994 8318 44996 8370
rect 44940 8306 44996 8318
rect 44716 8258 44772 8270
rect 44716 8206 44718 8258
rect 44770 8206 44772 8258
rect 44716 8036 44772 8206
rect 45052 8258 45108 8270
rect 45052 8206 45054 8258
rect 45106 8206 45108 8258
rect 45052 8148 45108 8206
rect 45276 8260 45332 8270
rect 45276 8166 45332 8204
rect 45052 8082 45108 8092
rect 44716 7970 44772 7980
rect 44380 7700 44436 7710
rect 44380 7364 44436 7644
rect 44380 7362 44884 7364
rect 44380 7310 44382 7362
rect 44434 7310 44884 7362
rect 44380 7308 44884 7310
rect 44380 7298 44436 7308
rect 44828 6914 44884 7308
rect 45612 6916 45668 19292
rect 46620 19348 46676 19358
rect 47180 19348 47236 19358
rect 46620 19346 47236 19348
rect 46620 19294 46622 19346
rect 46674 19294 47182 19346
rect 47234 19294 47236 19346
rect 46620 19292 47236 19294
rect 46620 19282 46676 19292
rect 46844 19122 46900 19134
rect 46844 19070 46846 19122
rect 46898 19070 46900 19122
rect 46844 19012 46900 19070
rect 46172 18562 46228 18574
rect 46172 18510 46174 18562
rect 46226 18510 46228 18562
rect 46172 18228 46228 18510
rect 46620 18340 46676 18350
rect 46620 18246 46676 18284
rect 46172 18162 46228 18172
rect 46844 18228 46900 18956
rect 47180 18562 47236 19292
rect 47292 18676 47348 20638
rect 47628 20244 47684 22652
rect 47852 22594 47908 22652
rect 47852 22542 47854 22594
rect 47906 22542 47908 22594
rect 47852 22530 47908 22542
rect 47740 22482 47796 22494
rect 47740 22430 47742 22482
rect 47794 22430 47796 22482
rect 47740 22372 47796 22430
rect 47852 22372 47908 22382
rect 47740 22316 47852 22372
rect 47852 22306 47908 22316
rect 47740 22148 47796 22158
rect 47740 21810 47796 22092
rect 47852 22148 47908 22158
rect 48188 22148 48244 23102
rect 49644 23044 49700 23884
rect 49756 23716 49812 24556
rect 49868 23940 49924 24668
rect 49980 24630 50036 24668
rect 49868 23846 49924 23884
rect 49756 23650 49812 23660
rect 49980 23826 50036 23838
rect 49980 23774 49982 23826
rect 50034 23774 50036 23826
rect 49980 23380 50036 23774
rect 49980 23314 50036 23324
rect 49644 22988 50036 23044
rect 49980 22594 50036 22988
rect 49980 22542 49982 22594
rect 50034 22542 50036 22594
rect 49980 22530 50036 22542
rect 47852 22146 48244 22148
rect 47852 22094 47854 22146
rect 47906 22094 48244 22146
rect 47852 22092 48244 22094
rect 49756 22148 49812 22158
rect 47852 22082 47908 22092
rect 47740 21758 47742 21810
rect 47794 21758 47796 21810
rect 47740 21746 47796 21758
rect 49644 21812 49700 21822
rect 49532 21586 49588 21598
rect 49532 21534 49534 21586
rect 49586 21534 49588 21586
rect 49084 20804 49140 20814
rect 49084 20802 49252 20804
rect 49084 20750 49086 20802
rect 49138 20750 49252 20802
rect 49084 20748 49252 20750
rect 49084 20738 49140 20748
rect 47628 20178 47684 20188
rect 48412 20578 48468 20590
rect 48412 20526 48414 20578
rect 48466 20526 48468 20578
rect 48412 20132 48468 20526
rect 48524 20580 48580 20590
rect 48524 20486 48580 20524
rect 48636 20578 48692 20590
rect 48636 20526 48638 20578
rect 48690 20526 48692 20578
rect 48412 20066 48468 20076
rect 48524 20356 48580 20366
rect 47516 19460 47572 19470
rect 47516 19366 47572 19404
rect 48412 19236 48468 19246
rect 48524 19236 48580 20300
rect 48636 19796 48692 20526
rect 48748 20244 48804 20254
rect 48748 20130 48804 20188
rect 48748 20078 48750 20130
rect 48802 20078 48804 20130
rect 48748 20066 48804 20078
rect 49084 20132 49140 20142
rect 49084 20018 49140 20076
rect 49084 19966 49086 20018
rect 49138 19966 49140 20018
rect 49084 19954 49140 19966
rect 49196 20020 49252 20748
rect 49308 20690 49364 20702
rect 49308 20638 49310 20690
rect 49362 20638 49364 20690
rect 49308 20356 49364 20638
rect 49308 20290 49364 20300
rect 49308 20020 49364 20030
rect 49196 20018 49364 20020
rect 49196 19966 49310 20018
rect 49362 19966 49364 20018
rect 49196 19964 49364 19966
rect 48860 19796 48916 19806
rect 48636 19794 48916 19796
rect 48636 19742 48862 19794
rect 48914 19742 48916 19794
rect 48636 19740 48916 19742
rect 48860 19460 48916 19740
rect 48860 19394 48916 19404
rect 48412 19234 48580 19236
rect 48412 19182 48414 19234
rect 48466 19182 48580 19234
rect 48412 19180 48580 19182
rect 47404 19012 47460 19022
rect 47404 18918 47460 18956
rect 47292 18610 47348 18620
rect 47180 18510 47182 18562
rect 47234 18510 47236 18562
rect 47180 18498 47236 18510
rect 47404 18452 47460 18462
rect 47404 18358 47460 18396
rect 47740 18450 47796 18462
rect 47740 18398 47742 18450
rect 47794 18398 47796 18450
rect 45836 17668 45892 17678
rect 45836 17666 46452 17668
rect 45836 17614 45838 17666
rect 45890 17614 46452 17666
rect 45836 17612 46452 17614
rect 45836 17602 45892 17612
rect 45948 16996 46004 17006
rect 45948 15428 46004 16940
rect 46396 16324 46452 17612
rect 46844 17554 46900 18172
rect 46844 17502 46846 17554
rect 46898 17502 46900 17554
rect 46844 17490 46900 17502
rect 47292 18340 47348 18350
rect 47292 17778 47348 18284
rect 47740 18340 47796 18398
rect 47740 18274 47796 18284
rect 47852 18452 47908 18462
rect 47292 17726 47294 17778
rect 47346 17726 47348 17778
rect 46620 16994 46676 17006
rect 46620 16942 46622 16994
rect 46674 16942 46676 16994
rect 46508 16324 46564 16334
rect 46396 16322 46564 16324
rect 46396 16270 46510 16322
rect 46562 16270 46564 16322
rect 46396 16268 46564 16270
rect 45836 15426 46004 15428
rect 45836 15374 45950 15426
rect 46002 15374 46004 15426
rect 45836 15372 46004 15374
rect 45724 15316 45780 15326
rect 45724 15222 45780 15260
rect 45724 14530 45780 14542
rect 45724 14478 45726 14530
rect 45778 14478 45780 14530
rect 45724 13748 45780 14478
rect 45836 13858 45892 15372
rect 45948 15362 46004 15372
rect 46172 15316 46228 15326
rect 46172 14530 46228 15260
rect 46172 14478 46174 14530
rect 46226 14478 46228 14530
rect 46172 14466 46228 14478
rect 46508 14532 46564 16268
rect 46620 15988 46676 16942
rect 46844 16882 46900 16894
rect 46844 16830 46846 16882
rect 46898 16830 46900 16882
rect 46844 16548 46900 16830
rect 46844 16482 46900 16492
rect 46620 15922 46676 15932
rect 47292 15202 47348 17726
rect 47852 17106 47908 18396
rect 48412 17668 48468 19180
rect 48524 19010 48580 19022
rect 48524 18958 48526 19010
rect 48578 18958 48580 19010
rect 48524 18788 48580 18958
rect 48524 18722 48580 18732
rect 48748 19010 48804 19022
rect 48748 18958 48750 19010
rect 48802 18958 48804 19010
rect 48748 18452 48804 18958
rect 48972 18452 49028 18462
rect 48748 18450 49028 18452
rect 48748 18398 48974 18450
rect 49026 18398 49028 18450
rect 48748 18396 49028 18398
rect 48412 17602 48468 17612
rect 48524 17780 48580 17790
rect 47852 17054 47854 17106
rect 47906 17054 47908 17106
rect 47852 17042 47908 17054
rect 47964 16994 48020 17006
rect 47964 16942 47966 16994
rect 48018 16942 48020 16994
rect 47852 16098 47908 16110
rect 47852 16046 47854 16098
rect 47906 16046 47908 16098
rect 47516 15316 47572 15326
rect 47516 15222 47572 15260
rect 47852 15316 47908 16046
rect 47852 15250 47908 15260
rect 47292 15150 47294 15202
rect 47346 15150 47348 15202
rect 47292 15148 47348 15150
rect 47292 15092 47460 15148
rect 47068 14756 47124 14766
rect 47124 14700 47236 14756
rect 47068 14690 47124 14700
rect 46508 14466 46564 14476
rect 45836 13806 45838 13858
rect 45890 13806 45892 13858
rect 45836 13794 45892 13806
rect 45724 13074 45780 13692
rect 45724 13022 45726 13074
rect 45778 13022 45780 13074
rect 45724 13010 45780 13022
rect 46620 12964 46676 12974
rect 46284 12962 46676 12964
rect 46284 12910 46622 12962
rect 46674 12910 46676 12962
rect 46284 12908 46676 12910
rect 45836 11508 45892 11518
rect 45724 9042 45780 9054
rect 45724 8990 45726 9042
rect 45778 8990 45780 9042
rect 45724 8372 45780 8990
rect 45724 8306 45780 8316
rect 45724 8148 45780 8158
rect 45724 7700 45780 8092
rect 45724 7606 45780 7644
rect 45836 7476 45892 11452
rect 46060 10724 46116 10734
rect 46116 10668 46228 10724
rect 46060 10630 46116 10668
rect 46060 9156 46116 9166
rect 46060 9062 46116 9100
rect 46172 8370 46228 10668
rect 46284 10722 46340 12908
rect 46620 12898 46676 12908
rect 47068 12178 47124 12190
rect 47068 12126 47070 12178
rect 47122 12126 47124 12178
rect 46284 10670 46286 10722
rect 46338 10670 46340 10722
rect 46284 10658 46340 10670
rect 46396 11844 46452 11854
rect 46396 11394 46452 11788
rect 47068 11844 47124 12126
rect 47068 11778 47124 11788
rect 46396 11342 46398 11394
rect 46450 11342 46452 11394
rect 46396 8708 46452 11342
rect 46732 11396 46788 11406
rect 46732 11282 46788 11340
rect 46732 11230 46734 11282
rect 46786 11230 46788 11282
rect 46732 11218 46788 11230
rect 47068 10610 47124 10622
rect 47068 10558 47070 10610
rect 47122 10558 47124 10610
rect 47068 9266 47124 10558
rect 47180 9380 47236 14700
rect 47404 14642 47460 15092
rect 47404 14590 47406 14642
rect 47458 14590 47460 14642
rect 47404 14578 47460 14590
rect 47628 14980 47684 14990
rect 47516 14532 47572 14542
rect 47516 14438 47572 14476
rect 47628 13972 47684 14924
rect 47516 13916 47684 13972
rect 47292 13748 47348 13758
rect 47292 13654 47348 13692
rect 47516 12964 47572 13916
rect 47628 13748 47684 13758
rect 47628 13746 47796 13748
rect 47628 13694 47630 13746
rect 47682 13694 47796 13746
rect 47628 13692 47796 13694
rect 47628 13682 47684 13692
rect 47292 12962 47572 12964
rect 47292 12910 47518 12962
rect 47570 12910 47572 12962
rect 47292 12908 47572 12910
rect 47292 10834 47348 12908
rect 47516 12898 47572 12908
rect 47628 12738 47684 12750
rect 47628 12686 47630 12738
rect 47682 12686 47684 12738
rect 47292 10782 47294 10834
rect 47346 10782 47348 10834
rect 47292 10770 47348 10782
rect 47404 12178 47460 12190
rect 47404 12126 47406 12178
rect 47458 12126 47460 12178
rect 47404 10724 47460 12126
rect 47628 12180 47684 12686
rect 47740 12516 47796 13692
rect 47964 13634 48020 16942
rect 48524 14756 48580 17724
rect 48748 17554 48804 18396
rect 48972 18386 49028 18396
rect 49084 18340 49140 18350
rect 49084 17780 49140 18284
rect 49308 18228 49364 19964
rect 49420 19236 49476 19246
rect 49420 19122 49476 19180
rect 49420 19070 49422 19122
rect 49474 19070 49476 19122
rect 49420 19058 49476 19070
rect 49532 19012 49588 21534
rect 49644 20690 49700 21756
rect 49756 21810 49812 22092
rect 49756 21758 49758 21810
rect 49810 21758 49812 21810
rect 49756 21746 49812 21758
rect 50204 21812 50260 25228
rect 50540 25218 50596 25228
rect 50556 25116 50820 25126
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50556 25050 50820 25060
rect 50316 24722 50372 24734
rect 50316 24670 50318 24722
rect 50370 24670 50372 24722
rect 50316 23828 50372 24670
rect 50652 24722 50708 24734
rect 50652 24670 50654 24722
rect 50706 24670 50708 24722
rect 50316 22820 50372 23772
rect 50428 24610 50484 24622
rect 50428 24558 50430 24610
rect 50482 24558 50484 24610
rect 50428 23380 50484 24558
rect 50652 24164 50708 24670
rect 50652 24108 51380 24164
rect 50988 23940 51044 23950
rect 50988 23826 51044 23884
rect 50988 23774 50990 23826
rect 51042 23774 51044 23826
rect 50988 23762 51044 23774
rect 51212 23828 51268 23838
rect 51324 23828 51380 24108
rect 51436 23828 51492 23838
rect 51324 23826 51492 23828
rect 51324 23774 51438 23826
rect 51490 23774 51492 23826
rect 51324 23772 51492 23774
rect 51212 23734 51268 23772
rect 50876 23714 50932 23726
rect 50876 23662 50878 23714
rect 50930 23662 50932 23714
rect 50556 23548 50820 23558
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50556 23482 50820 23492
rect 50428 23324 50596 23380
rect 50428 23156 50484 23166
rect 50428 23062 50484 23100
rect 50540 23042 50596 23324
rect 50876 23154 50932 23662
rect 50876 23102 50878 23154
rect 50930 23102 50932 23154
rect 50876 23090 50932 23102
rect 50540 22990 50542 23042
rect 50594 22990 50596 23042
rect 50540 22978 50596 22990
rect 51100 22930 51156 22942
rect 51100 22878 51102 22930
rect 51154 22878 51156 22930
rect 50316 22764 50596 22820
rect 50540 22484 50596 22764
rect 50540 22390 50596 22428
rect 50316 22372 50372 22382
rect 50428 22372 50484 22382
rect 50316 22370 50428 22372
rect 50316 22318 50318 22370
rect 50370 22318 50428 22370
rect 50316 22316 50428 22318
rect 50316 22306 50372 22316
rect 50204 21746 50260 21756
rect 50428 20914 50484 22316
rect 51100 22260 51156 22878
rect 51436 22372 51492 23772
rect 51436 22306 51492 22316
rect 51100 22194 51156 22204
rect 51324 22258 51380 22270
rect 51324 22206 51326 22258
rect 51378 22206 51380 22258
rect 50556 21980 50820 21990
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50556 21914 50820 21924
rect 51324 21924 51380 22206
rect 51324 21858 51380 21868
rect 51436 22146 51492 22158
rect 51436 22094 51438 22146
rect 51490 22094 51492 22146
rect 50988 21812 51044 21822
rect 51436 21812 51492 22094
rect 51548 22148 51604 25452
rect 52108 25284 52164 25294
rect 52108 24948 52164 25228
rect 51996 24892 52164 24948
rect 51996 24724 52052 24892
rect 51996 24658 52052 24668
rect 52108 24724 52164 24734
rect 52220 24724 52276 25564
rect 52780 25396 52836 25406
rect 52780 25302 52836 25340
rect 52892 25394 52948 25406
rect 52892 25342 52894 25394
rect 52946 25342 52948 25394
rect 52892 24948 52948 25342
rect 53116 25396 53172 26012
rect 53564 25506 53620 26236
rect 53788 26180 53844 26190
rect 53564 25454 53566 25506
rect 53618 25454 53620 25506
rect 53564 25442 53620 25454
rect 53676 26124 53788 26180
rect 53116 25330 53172 25340
rect 53676 25394 53732 26124
rect 53788 26086 53844 26124
rect 54572 26180 54628 27132
rect 55580 27076 55636 27086
rect 55580 26982 55636 27020
rect 54684 26962 54740 26974
rect 54684 26910 54686 26962
rect 54738 26910 54740 26962
rect 54684 26908 54740 26910
rect 54908 26962 54964 26974
rect 54908 26910 54910 26962
rect 54962 26910 54964 26962
rect 54684 26852 54852 26908
rect 54796 26290 54852 26852
rect 54908 26516 54964 26910
rect 57596 26908 57652 27694
rect 57932 27636 57988 27646
rect 57932 27298 57988 27580
rect 57932 27246 57934 27298
rect 57986 27246 57988 27298
rect 57932 27234 57988 27246
rect 57484 26852 57540 26862
rect 57596 26852 58212 26908
rect 54908 26450 54964 26460
rect 55580 26516 55636 26526
rect 55580 26422 55636 26460
rect 55356 26292 55412 26302
rect 54796 26238 54798 26290
rect 54850 26238 54852 26290
rect 54572 26178 54740 26180
rect 54572 26126 54574 26178
rect 54626 26126 54740 26178
rect 54572 26124 54740 26126
rect 54572 26114 54628 26124
rect 53900 25676 54628 25732
rect 53900 25506 53956 25676
rect 53900 25454 53902 25506
rect 53954 25454 53956 25506
rect 53900 25442 53956 25454
rect 54572 25506 54628 25676
rect 54684 25730 54740 26124
rect 54684 25678 54686 25730
rect 54738 25678 54740 25730
rect 54684 25666 54740 25678
rect 54572 25454 54574 25506
rect 54626 25454 54628 25506
rect 54572 25442 54628 25454
rect 53676 25342 53678 25394
rect 53730 25342 53732 25394
rect 53676 25284 53732 25342
rect 53676 25218 53732 25228
rect 52108 24722 52276 24724
rect 52108 24670 52110 24722
rect 52162 24670 52276 24722
rect 52108 24668 52276 24670
rect 52332 24892 52948 24948
rect 52108 24658 52164 24668
rect 52332 24052 52388 24892
rect 52556 24722 52612 24734
rect 52556 24670 52558 24722
rect 52610 24670 52612 24722
rect 52108 23996 52500 24052
rect 52108 23938 52164 23996
rect 52108 23886 52110 23938
rect 52162 23886 52164 23938
rect 52108 23874 52164 23886
rect 51884 23828 51940 23838
rect 51772 23772 51884 23828
rect 51772 23714 51828 23772
rect 51884 23762 51940 23772
rect 51772 23662 51774 23714
rect 51826 23662 51828 23714
rect 51772 23650 51828 23662
rect 51996 23716 52052 23726
rect 51660 23044 51716 23054
rect 51660 22370 51716 22988
rect 51660 22318 51662 22370
rect 51714 22318 51716 22370
rect 51660 22306 51716 22318
rect 51884 22372 51940 22382
rect 51548 22082 51604 22092
rect 51884 22148 51940 22316
rect 51996 22258 52052 23660
rect 52332 23266 52388 23278
rect 52332 23214 52334 23266
rect 52386 23214 52388 23266
rect 52108 23044 52164 23054
rect 52108 22950 52164 22988
rect 52220 22372 52276 22382
rect 52332 22372 52388 23214
rect 52220 22370 52388 22372
rect 52220 22318 52222 22370
rect 52274 22318 52388 22370
rect 52220 22316 52388 22318
rect 52220 22306 52276 22316
rect 51996 22206 51998 22258
rect 52050 22206 52052 22258
rect 51996 22194 52052 22206
rect 51884 22082 51940 22092
rect 51044 21756 51156 21812
rect 50988 21718 51044 21756
rect 50764 21698 50820 21710
rect 50764 21646 50766 21698
rect 50818 21646 50820 21698
rect 50652 21364 50708 21374
rect 50428 20862 50430 20914
rect 50482 20862 50484 20914
rect 50428 20850 50484 20862
rect 50540 21362 50708 21364
rect 50540 21310 50654 21362
rect 50706 21310 50708 21362
rect 50540 21308 50708 21310
rect 50540 20804 50596 21308
rect 50652 21298 50708 21308
rect 50764 21028 50820 21646
rect 50764 20972 51044 21028
rect 50540 20748 50932 20804
rect 49644 20638 49646 20690
rect 49698 20638 49700 20690
rect 49644 20626 49700 20638
rect 50092 20690 50148 20702
rect 50092 20638 50094 20690
rect 50146 20638 50148 20690
rect 50092 20020 50148 20638
rect 50540 20690 50596 20748
rect 50540 20638 50542 20690
rect 50594 20638 50596 20690
rect 50540 20626 50596 20638
rect 50316 20580 50372 20590
rect 50316 20188 50372 20524
rect 50876 20468 50932 20748
rect 50988 20692 51044 20972
rect 51100 20802 51156 21756
rect 51436 21746 51492 21756
rect 51996 21924 52052 21934
rect 51996 21810 52052 21868
rect 51996 21758 51998 21810
rect 52050 21758 52052 21810
rect 51996 21746 52052 21758
rect 51884 21700 51940 21710
rect 51884 21606 51940 21644
rect 51100 20750 51102 20802
rect 51154 20750 51156 20802
rect 51100 20738 51156 20750
rect 51212 21586 51268 21598
rect 51212 21534 51214 21586
rect 51266 21534 51268 21586
rect 50988 20598 51044 20636
rect 51212 20692 51268 21534
rect 52108 21586 52164 21598
rect 52108 21534 52110 21586
rect 52162 21534 52164 21586
rect 52108 21140 52164 21534
rect 51660 21084 52164 21140
rect 51660 21026 51716 21084
rect 51660 20974 51662 21026
rect 51714 20974 51716 21026
rect 51660 20962 51716 20974
rect 51212 20690 51492 20692
rect 51212 20638 51214 20690
rect 51266 20638 51492 20690
rect 51212 20636 51492 20638
rect 51212 20626 51268 20636
rect 50556 20412 50820 20422
rect 50876 20412 51380 20468
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50556 20346 50820 20356
rect 50316 20132 50932 20188
rect 50092 19954 50148 19964
rect 50876 20018 50932 20132
rect 51324 20130 51380 20412
rect 51324 20078 51326 20130
rect 51378 20078 51380 20130
rect 51324 20066 51380 20078
rect 50876 19966 50878 20018
rect 50930 19966 50932 20018
rect 50876 19954 50932 19966
rect 51100 20020 51156 20030
rect 51100 20018 51268 20020
rect 51100 19966 51102 20018
rect 51154 19966 51268 20018
rect 51100 19964 51268 19966
rect 51100 19954 51156 19964
rect 51212 19908 51268 19964
rect 51212 19842 51268 19852
rect 50428 19346 50484 19358
rect 50428 19294 50430 19346
rect 50482 19294 50484 19346
rect 49532 18946 49588 18956
rect 49644 19234 49700 19246
rect 49644 19182 49646 19234
rect 49698 19182 49700 19234
rect 49644 18788 49700 19182
rect 50428 18900 50484 19294
rect 51212 19348 51268 19358
rect 51436 19348 51492 20636
rect 51212 19346 51492 19348
rect 51212 19294 51214 19346
rect 51266 19294 51492 19346
rect 51212 19292 51492 19294
rect 51548 20020 51604 20030
rect 51212 19282 51268 19292
rect 50764 19236 50820 19246
rect 50764 19234 50932 19236
rect 50764 19182 50766 19234
rect 50818 19182 50932 19234
rect 50764 19180 50932 19182
rect 50764 19170 50820 19180
rect 49644 18564 49700 18732
rect 49644 18498 49700 18508
rect 50316 18844 50484 18900
rect 50556 18844 50820 18854
rect 49308 18162 49364 18172
rect 50316 18450 50372 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50556 18778 50820 18788
rect 50316 18398 50318 18450
rect 50370 18398 50372 18450
rect 49084 17714 49140 17724
rect 48748 17502 48750 17554
rect 48802 17502 48804 17554
rect 48748 17490 48804 17502
rect 50316 17556 50372 18398
rect 50316 17462 50372 17500
rect 50428 18676 50484 18686
rect 50428 17442 50484 18620
rect 50764 18676 50820 18686
rect 50540 18228 50596 18238
rect 50540 18134 50596 18172
rect 50764 17668 50820 18620
rect 50876 18340 50932 19180
rect 50876 18274 50932 18284
rect 50988 18564 51044 18574
rect 50876 17668 50932 17678
rect 50764 17666 50932 17668
rect 50764 17614 50878 17666
rect 50930 17614 50932 17666
rect 50764 17612 50932 17614
rect 50428 17390 50430 17442
rect 50482 17390 50484 17442
rect 50428 17378 50484 17390
rect 50556 17276 50820 17286
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50556 17210 50820 17220
rect 50876 16660 50932 17612
rect 50988 17554 51044 18508
rect 51548 18562 51604 19964
rect 52444 20020 52500 23996
rect 52556 22260 52612 24670
rect 53452 24722 53508 24734
rect 53452 24670 53454 24722
rect 53506 24670 53508 24722
rect 53004 24610 53060 24622
rect 53004 24558 53006 24610
rect 53058 24558 53060 24610
rect 53004 23380 53060 24558
rect 53452 24052 53508 24670
rect 53452 23986 53508 23996
rect 53676 24052 53732 24062
rect 53676 23938 53732 23996
rect 53676 23886 53678 23938
rect 53730 23886 53732 23938
rect 53676 23874 53732 23886
rect 53452 23828 53508 23838
rect 53452 23734 53508 23772
rect 54796 23604 54852 26238
rect 55132 26236 55356 26292
rect 55020 25618 55076 25630
rect 55020 25566 55022 25618
rect 55074 25566 55076 25618
rect 55020 25508 55076 25566
rect 55020 25442 55076 25452
rect 55020 23940 55076 23950
rect 55020 23826 55076 23884
rect 55020 23774 55022 23826
rect 55074 23774 55076 23826
rect 55020 23762 55076 23774
rect 54796 23538 54852 23548
rect 53004 23314 53060 23324
rect 53900 23380 53956 23390
rect 53340 23156 53396 23166
rect 53004 22484 53060 22494
rect 52556 22194 52612 22204
rect 52668 22258 52724 22270
rect 52668 22206 52670 22258
rect 52722 22206 52724 22258
rect 52668 21924 52724 22206
rect 53004 22260 53060 22428
rect 53004 22258 53284 22260
rect 53004 22206 53006 22258
rect 53058 22206 53284 22258
rect 53004 22204 53284 22206
rect 53004 22194 53060 22204
rect 52668 21858 52724 21868
rect 53004 21812 53060 21822
rect 53004 21698 53060 21756
rect 53228 21810 53284 22204
rect 53228 21758 53230 21810
rect 53282 21758 53284 21810
rect 53228 21746 53284 21758
rect 53004 21646 53006 21698
rect 53058 21646 53060 21698
rect 52556 21588 52612 21598
rect 52556 21586 52836 21588
rect 52556 21534 52558 21586
rect 52610 21534 52836 21586
rect 52556 21532 52836 21534
rect 52556 21522 52612 21532
rect 52444 19954 52500 19964
rect 51548 18510 51550 18562
rect 51602 18510 51604 18562
rect 51548 18498 51604 18510
rect 50988 17502 50990 17554
rect 51042 17502 51044 17554
rect 50988 17490 51044 17502
rect 52108 18452 52164 18462
rect 51212 17444 51268 17454
rect 51212 17350 51268 17388
rect 52108 17444 52164 18396
rect 52220 18452 52276 18462
rect 52220 18450 52388 18452
rect 52220 18398 52222 18450
rect 52274 18398 52388 18450
rect 52220 18396 52388 18398
rect 52220 18386 52276 18396
rect 52108 16994 52164 17388
rect 52108 16942 52110 16994
rect 52162 16942 52164 16994
rect 52108 16930 52164 16942
rect 52220 17556 52276 17566
rect 50428 16604 50932 16660
rect 51660 16772 51716 16782
rect 49084 16548 49140 16558
rect 49140 16492 49252 16548
rect 48972 15988 49028 15998
rect 48972 15894 49028 15932
rect 48748 15316 48804 15354
rect 48748 15250 48804 15260
rect 49084 15314 49140 16492
rect 49196 16210 49252 16492
rect 49196 16158 49198 16210
rect 49250 16158 49252 16210
rect 49196 16146 49252 16158
rect 50204 16324 50260 16334
rect 49980 16100 50036 16110
rect 49308 15988 49364 15998
rect 49084 15262 49086 15314
rect 49138 15262 49140 15314
rect 48524 14662 48580 14700
rect 48300 14532 48356 14542
rect 48300 13970 48356 14476
rect 49084 14420 49140 15262
rect 48300 13918 48302 13970
rect 48354 13918 48356 13970
rect 48300 13906 48356 13918
rect 48748 14364 49140 14420
rect 49196 15316 49252 15326
rect 48748 13858 48804 14364
rect 48748 13806 48750 13858
rect 48802 13806 48804 13858
rect 48748 13794 48804 13806
rect 47964 13582 47966 13634
rect 48018 13582 48020 13634
rect 47964 12964 48020 13582
rect 48972 13748 49028 13758
rect 48972 13074 49028 13692
rect 48972 13022 48974 13074
rect 49026 13022 49028 13074
rect 48972 13010 49028 13022
rect 49084 13746 49140 13758
rect 49084 13694 49086 13746
rect 49138 13694 49140 13746
rect 48412 12964 48468 12974
rect 47964 12962 48468 12964
rect 47964 12910 48414 12962
rect 48466 12910 48468 12962
rect 47964 12908 48468 12910
rect 47852 12740 47908 12750
rect 47852 12646 47908 12684
rect 48076 12628 48132 12638
rect 48076 12516 48132 12572
rect 47740 12460 48132 12516
rect 47628 12114 47684 12124
rect 47964 12180 48020 12190
rect 47964 12086 48020 12124
rect 47516 12066 47572 12078
rect 47516 12014 47518 12066
rect 47570 12014 47572 12066
rect 47516 11506 47572 12014
rect 48076 11618 48132 12460
rect 48188 12292 48244 12302
rect 48188 12198 48244 12236
rect 48076 11566 48078 11618
rect 48130 11566 48132 11618
rect 48076 11554 48132 11566
rect 48412 11620 48468 12908
rect 48748 12962 48804 12974
rect 48748 12910 48750 12962
rect 48802 12910 48804 12962
rect 48748 12628 48804 12910
rect 48748 12562 48804 12572
rect 49084 12628 49140 13694
rect 49084 12562 49140 12572
rect 49196 12404 49252 15260
rect 49308 14530 49364 15932
rect 49868 15988 49924 15998
rect 49868 15426 49924 15932
rect 49980 15538 50036 16044
rect 50092 15988 50148 15998
rect 50204 15988 50260 16268
rect 50092 15986 50260 15988
rect 50092 15934 50094 15986
rect 50146 15934 50260 15986
rect 50092 15932 50260 15934
rect 50092 15922 50148 15932
rect 49980 15486 49982 15538
rect 50034 15486 50036 15538
rect 49980 15474 50036 15486
rect 50204 15540 50260 15932
rect 50428 15876 50484 16604
rect 50764 16156 50932 16212
rect 50764 16100 50820 16156
rect 50764 16034 50820 16044
rect 50204 15474 50260 15484
rect 50316 15820 50484 15876
rect 49868 15374 49870 15426
rect 49922 15374 49924 15426
rect 49420 15092 49476 15102
rect 49420 14998 49476 15036
rect 49308 14478 49310 14530
rect 49362 14478 49364 14530
rect 49308 14466 49364 14478
rect 49420 12852 49476 12862
rect 49420 12758 49476 12796
rect 49868 12852 49924 15374
rect 50316 15428 50372 15820
rect 50876 15764 50932 16156
rect 51100 16098 51156 16110
rect 51100 16046 51102 16098
rect 51154 16046 51156 16098
rect 50988 15988 51044 15998
rect 50988 15894 51044 15932
rect 51100 15876 51156 16046
rect 51100 15820 51492 15876
rect 50556 15708 50820 15718
rect 50876 15708 51156 15764
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50556 15642 50820 15652
rect 50540 15540 50596 15550
rect 50540 15446 50596 15484
rect 50428 15428 50484 15438
rect 50316 15426 50484 15428
rect 50316 15374 50430 15426
rect 50482 15374 50484 15426
rect 50316 15372 50484 15374
rect 50204 15314 50260 15326
rect 50204 15262 50206 15314
rect 50258 15262 50260 15314
rect 50204 13634 50260 15262
rect 50428 14980 50484 15372
rect 50764 15316 50820 15326
rect 50764 15314 50932 15316
rect 50764 15262 50766 15314
rect 50818 15262 50932 15314
rect 50764 15260 50932 15262
rect 50764 15250 50820 15260
rect 50428 14914 50484 14924
rect 50764 15092 50820 15102
rect 50764 14642 50820 15036
rect 50764 14590 50766 14642
rect 50818 14590 50820 14642
rect 50764 14578 50820 14590
rect 50428 14532 50484 14542
rect 50428 14438 50484 14476
rect 50556 14140 50820 14150
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50556 14074 50820 14084
rect 50764 13860 50820 13870
rect 50876 13860 50932 15260
rect 50988 15314 51044 15326
rect 50988 15262 50990 15314
rect 51042 15262 51044 15314
rect 50988 14868 51044 15262
rect 50988 14802 51044 14812
rect 50820 13804 50932 13860
rect 50764 13766 50820 13804
rect 50204 13582 50206 13634
rect 50258 13582 50260 13634
rect 50204 13570 50260 13582
rect 50988 12964 51044 12974
rect 50988 12870 51044 12908
rect 49868 12786 49924 12796
rect 51100 12850 51156 15708
rect 51436 13748 51492 15820
rect 51548 15874 51604 15886
rect 51548 15822 51550 15874
rect 51602 15822 51604 15874
rect 51548 14644 51604 15822
rect 51660 15202 51716 16716
rect 51660 15150 51662 15202
rect 51714 15150 51716 15202
rect 51660 15138 51716 15150
rect 52220 15314 52276 17500
rect 52332 17108 52388 18396
rect 52780 17780 52836 21532
rect 52892 20692 52948 20702
rect 52892 20130 52948 20636
rect 52892 20078 52894 20130
rect 52946 20078 52948 20130
rect 52892 20066 52948 20078
rect 53004 19458 53060 21646
rect 53340 21474 53396 23100
rect 53564 23154 53620 23166
rect 53564 23102 53566 23154
rect 53618 23102 53620 23154
rect 53452 22260 53508 22270
rect 53452 22166 53508 22204
rect 53340 21422 53342 21474
rect 53394 21422 53396 21474
rect 53340 21410 53396 21422
rect 53564 21586 53620 23102
rect 53900 22370 53956 23324
rect 55020 23268 55076 23278
rect 54684 23156 54740 23166
rect 55020 23156 55076 23212
rect 54684 23062 54740 23100
rect 54796 23100 55076 23156
rect 53900 22318 53902 22370
rect 53954 22318 53956 22370
rect 53900 22306 53956 22318
rect 54460 22930 54516 22942
rect 54796 22932 54852 23100
rect 55132 23044 55188 26236
rect 55356 26198 55412 26236
rect 55692 26290 55748 26302
rect 55692 26238 55694 26290
rect 55746 26238 55748 26290
rect 55692 26180 55748 26238
rect 55916 26290 55972 26302
rect 56588 26292 56644 26302
rect 55916 26238 55918 26290
rect 55970 26238 55972 26290
rect 55748 26124 55860 26180
rect 55692 26114 55748 26124
rect 55580 25844 55636 25854
rect 55468 25508 55524 25518
rect 55356 24498 55412 24510
rect 55356 24446 55358 24498
rect 55410 24446 55412 24498
rect 55356 24276 55412 24446
rect 55356 24210 55412 24220
rect 55244 23826 55300 23838
rect 55244 23774 55246 23826
rect 55298 23774 55300 23826
rect 55244 23716 55300 23774
rect 55468 23716 55524 25452
rect 55580 25506 55636 25788
rect 55580 25454 55582 25506
rect 55634 25454 55636 25506
rect 55580 25442 55636 25454
rect 55580 24836 55636 24846
rect 55580 24164 55636 24780
rect 55580 23938 55636 24108
rect 55580 23886 55582 23938
rect 55634 23886 55636 23938
rect 55580 23874 55636 23886
rect 55692 23828 55748 23838
rect 55468 23660 55636 23716
rect 55244 23650 55300 23660
rect 55468 23492 55524 23502
rect 54460 22878 54462 22930
rect 54514 22878 54516 22930
rect 54460 22370 54516 22878
rect 54460 22318 54462 22370
rect 54514 22318 54516 22370
rect 54460 22306 54516 22318
rect 54572 22876 54852 22932
rect 54908 22988 55188 23044
rect 55244 23154 55300 23166
rect 55244 23102 55246 23154
rect 55298 23102 55300 23154
rect 54348 22148 54404 22158
rect 54348 22054 54404 22092
rect 54348 21812 54404 21822
rect 54348 21718 54404 21756
rect 53564 21534 53566 21586
rect 53618 21534 53620 21586
rect 53004 19406 53006 19458
rect 53058 19406 53060 19458
rect 53004 19394 53060 19406
rect 53116 20018 53172 20030
rect 53116 19966 53118 20018
rect 53170 19966 53172 20018
rect 53116 19236 53172 19966
rect 53564 19460 53620 21534
rect 54572 21588 54628 22876
rect 54908 22370 54964 22988
rect 55132 22372 55188 22382
rect 54908 22318 54910 22370
rect 54962 22318 54964 22370
rect 54684 21812 54740 21822
rect 54908 21812 54964 22318
rect 54684 21810 54964 21812
rect 54684 21758 54686 21810
rect 54738 21758 54964 21810
rect 54684 21756 54964 21758
rect 55020 22370 55188 22372
rect 55020 22318 55134 22370
rect 55186 22318 55188 22370
rect 55020 22316 55188 22318
rect 54684 21746 54740 21756
rect 54796 21588 54852 21598
rect 54572 21532 54796 21588
rect 54124 20020 54180 20030
rect 53788 19908 53844 19918
rect 53788 19814 53844 19852
rect 54124 19460 54180 19964
rect 54236 20020 54292 20030
rect 54236 20018 54404 20020
rect 54236 19966 54238 20018
rect 54290 19966 54404 20018
rect 54236 19964 54404 19966
rect 54236 19954 54292 19964
rect 54348 19572 54404 19964
rect 54796 19906 54852 21532
rect 54908 21586 54964 21598
rect 54908 21534 54910 21586
rect 54962 21534 54964 21586
rect 54908 20188 54964 21534
rect 55020 20692 55076 22316
rect 55132 22306 55188 22316
rect 55244 22372 55300 23102
rect 55468 23154 55524 23436
rect 55468 23102 55470 23154
rect 55522 23102 55524 23154
rect 55468 22484 55524 23102
rect 55244 22306 55300 22316
rect 55356 22428 55524 22484
rect 55132 22146 55188 22158
rect 55132 22094 55134 22146
rect 55186 22094 55188 22146
rect 55132 21812 55188 22094
rect 55356 22036 55412 22428
rect 55468 22260 55524 22270
rect 55580 22260 55636 23660
rect 55692 22372 55748 23772
rect 55804 23492 55860 26124
rect 55916 25508 55972 26238
rect 55916 25442 55972 25452
rect 56140 26290 56644 26292
rect 56140 26238 56590 26290
rect 56642 26238 56644 26290
rect 56140 26236 56644 26238
rect 55804 23426 55860 23436
rect 56140 24052 56196 26236
rect 56588 26226 56644 26236
rect 57372 26178 57428 26190
rect 57372 26126 57374 26178
rect 57426 26126 57428 26178
rect 56140 23378 56196 23996
rect 56140 23326 56142 23378
rect 56194 23326 56196 23378
rect 56140 23314 56196 23326
rect 56588 26066 56644 26078
rect 56588 26014 56590 26066
rect 56642 26014 56644 26066
rect 55804 23268 55860 23278
rect 55804 23174 55860 23212
rect 55916 23266 55972 23278
rect 55916 23214 55918 23266
rect 55970 23214 55972 23266
rect 55916 23156 55972 23214
rect 55916 23100 56532 23156
rect 56252 22372 56308 22382
rect 55692 22370 56308 22372
rect 55692 22318 56254 22370
rect 56306 22318 56308 22370
rect 55692 22316 56308 22318
rect 56252 22306 56308 22316
rect 55580 22204 55748 22260
rect 55468 22166 55524 22204
rect 55356 21970 55412 21980
rect 55132 21756 55636 21812
rect 55580 21586 55636 21756
rect 55580 21534 55582 21586
rect 55634 21534 55636 21586
rect 55580 21522 55636 21534
rect 55692 21474 55748 22204
rect 55692 21422 55694 21474
rect 55746 21422 55748 21474
rect 55692 21410 55748 21422
rect 55804 21924 55860 21934
rect 55804 21026 55860 21868
rect 56476 21812 56532 23100
rect 56588 22482 56644 26014
rect 56924 26066 56980 26078
rect 56924 26014 56926 26066
rect 56978 26014 56980 26066
rect 56700 25956 56756 25966
rect 56700 24610 56756 25900
rect 56700 24558 56702 24610
rect 56754 24558 56756 24610
rect 56700 24546 56756 24558
rect 56924 24276 56980 26014
rect 57372 25844 57428 26126
rect 57372 25778 57428 25788
rect 57484 25730 57540 26796
rect 57484 25678 57486 25730
rect 57538 25678 57540 25730
rect 57484 25666 57540 25678
rect 57820 26402 57876 26414
rect 57820 26350 57822 26402
rect 57874 26350 57876 26402
rect 57820 25396 57876 26350
rect 57820 25330 57876 25340
rect 58156 26290 58212 26852
rect 58156 26238 58158 26290
rect 58210 26238 58212 26290
rect 57932 24948 57988 24958
rect 56700 24220 56980 24276
rect 57148 24722 57204 24734
rect 57148 24670 57150 24722
rect 57202 24670 57204 24722
rect 56700 23940 56756 24220
rect 56700 23042 56756 23884
rect 56700 22990 56702 23042
rect 56754 22990 56756 23042
rect 56700 22978 56756 22990
rect 56812 23604 56868 23614
rect 56812 22594 56868 23548
rect 57036 23156 57092 23166
rect 56812 22542 56814 22594
rect 56866 22542 56868 22594
rect 56812 22530 56868 22542
rect 56924 23154 57092 23156
rect 56924 23102 57038 23154
rect 57090 23102 57092 23154
rect 56924 23100 57092 23102
rect 56588 22430 56590 22482
rect 56642 22430 56644 22482
rect 56588 22418 56644 22430
rect 56812 22370 56868 22382
rect 56812 22318 56814 22370
rect 56866 22318 56868 22370
rect 56476 21756 56756 21812
rect 55916 21700 55972 21710
rect 55916 21606 55972 21644
rect 55804 20974 55806 21026
rect 55858 20974 55860 21026
rect 55804 20962 55860 20974
rect 55020 20626 55076 20636
rect 55692 20690 55748 20702
rect 55692 20638 55694 20690
rect 55746 20638 55748 20690
rect 55692 20188 55748 20638
rect 55804 20692 55860 20702
rect 55804 20598 55860 20636
rect 54908 20132 55748 20188
rect 56476 20242 56532 21756
rect 56700 21698 56756 21756
rect 56700 21646 56702 21698
rect 56754 21646 56756 21698
rect 56700 21634 56756 21646
rect 56812 21700 56868 22318
rect 56588 21588 56644 21598
rect 56588 21494 56644 21532
rect 56812 21474 56868 21644
rect 56812 21422 56814 21474
rect 56866 21422 56868 21474
rect 56812 21410 56868 21422
rect 56924 21924 56980 23100
rect 57036 23090 57092 23100
rect 57148 22370 57204 24670
rect 57372 24610 57428 24622
rect 57372 24558 57374 24610
rect 57426 24558 57428 24610
rect 57372 23716 57428 24558
rect 57932 24162 57988 24892
rect 57932 24110 57934 24162
rect 57986 24110 57988 24162
rect 57932 24098 57988 24110
rect 58044 24164 58100 24174
rect 57148 22318 57150 22370
rect 57202 22318 57204 22370
rect 57148 22148 57204 22318
rect 57148 22082 57204 22092
rect 57260 23042 57316 23054
rect 57260 22990 57262 23042
rect 57314 22990 57316 23042
rect 57260 22260 57316 22990
rect 57372 22370 57428 23660
rect 58044 23380 58100 24108
rect 58156 23604 58212 26238
rect 58156 23538 58212 23548
rect 58156 23380 58212 23390
rect 58044 23378 58212 23380
rect 58044 23326 58158 23378
rect 58210 23326 58212 23378
rect 58044 23324 58212 23326
rect 58156 23314 58212 23324
rect 57372 22318 57374 22370
rect 57426 22318 57428 22370
rect 57372 22306 57428 22318
rect 57260 21924 57316 22204
rect 56812 20804 56868 20814
rect 56924 20804 56980 21868
rect 56812 20802 56980 20804
rect 56812 20750 56814 20802
rect 56866 20750 56980 20802
rect 56812 20748 56980 20750
rect 57036 21868 57316 21924
rect 57036 20802 57092 21868
rect 57484 21588 57540 21598
rect 57260 21586 57540 21588
rect 57260 21534 57486 21586
rect 57538 21534 57540 21586
rect 57260 21532 57540 21534
rect 57260 20914 57316 21532
rect 57484 21522 57540 21532
rect 58156 21588 58212 21598
rect 57260 20862 57262 20914
rect 57314 20862 57316 20914
rect 57260 20850 57316 20862
rect 57820 21364 57876 21374
rect 57036 20750 57038 20802
rect 57090 20750 57092 20802
rect 56812 20738 56868 20748
rect 57036 20692 57092 20750
rect 56476 20190 56478 20242
rect 56530 20190 56532 20242
rect 56476 20178 56532 20190
rect 56924 20636 57092 20692
rect 57820 20690 57876 21308
rect 58156 20804 58212 21532
rect 58156 20802 58324 20804
rect 58156 20750 58158 20802
rect 58210 20750 58324 20802
rect 58156 20748 58324 20750
rect 58156 20738 58212 20748
rect 57820 20638 57822 20690
rect 57874 20638 57876 20690
rect 55020 20020 55076 20030
rect 55020 20018 55188 20020
rect 55020 19966 55022 20018
rect 55074 19966 55188 20018
rect 55020 19964 55188 19966
rect 55020 19954 55076 19964
rect 54796 19854 54798 19906
rect 54850 19854 54852 19906
rect 54796 19842 54852 19854
rect 54348 19516 54964 19572
rect 53564 19394 53620 19404
rect 53676 19458 54180 19460
rect 53676 19406 54126 19458
rect 54178 19406 54180 19458
rect 53676 19404 54180 19406
rect 53116 19170 53172 19180
rect 53340 19234 53396 19246
rect 53340 19182 53342 19234
rect 53394 19182 53396 19234
rect 53340 18564 53396 19182
rect 53340 18498 53396 18508
rect 53564 19124 53620 19134
rect 53564 18452 53620 19068
rect 53564 18358 53620 18396
rect 53452 18340 53508 18350
rect 52780 17724 53396 17780
rect 52444 17108 52500 17118
rect 52332 17052 52444 17108
rect 52444 17042 52500 17052
rect 53228 17108 53284 17118
rect 53228 16882 53284 17052
rect 53340 17106 53396 17724
rect 53340 17054 53342 17106
rect 53394 17054 53396 17106
rect 53340 17042 53396 17054
rect 53228 16830 53230 16882
rect 53282 16830 53284 16882
rect 53228 16818 53284 16830
rect 53340 16772 53396 16782
rect 53452 16772 53508 18284
rect 53676 18228 53732 19404
rect 54124 19394 54180 19404
rect 54460 19348 54516 19358
rect 54460 19254 54516 19292
rect 54908 19346 54964 19516
rect 54908 19294 54910 19346
rect 54962 19294 54964 19346
rect 54908 19282 54964 19294
rect 53900 19236 53956 19246
rect 53900 19142 53956 19180
rect 54796 19122 54852 19134
rect 54796 19070 54798 19122
rect 54850 19070 54852 19122
rect 54124 18564 54180 18574
rect 54124 18470 54180 18508
rect 54796 18564 54852 19070
rect 55020 19124 55076 19134
rect 55020 19030 55076 19068
rect 54796 18498 54852 18508
rect 54572 18450 54628 18462
rect 54572 18398 54574 18450
rect 54626 18398 54628 18450
rect 54572 18340 54628 18398
rect 55132 18452 55188 19964
rect 55132 18386 55188 18396
rect 54572 18274 54628 18284
rect 55020 18340 55076 18350
rect 55020 18246 55076 18284
rect 53396 16716 53508 16772
rect 53564 18172 53732 18228
rect 53340 16706 53396 16716
rect 53228 16324 53284 16334
rect 53228 16210 53284 16268
rect 53228 16158 53230 16210
rect 53282 16158 53284 16210
rect 53228 16146 53284 16158
rect 53564 15988 53620 18172
rect 55356 18116 55412 20132
rect 56700 20130 56756 20142
rect 56700 20078 56702 20130
rect 56754 20078 56756 20130
rect 55804 19460 55860 19470
rect 55804 19366 55860 19404
rect 56700 19348 56756 20078
rect 56700 19282 56756 19292
rect 56812 20018 56868 20030
rect 56812 19966 56814 20018
rect 56866 19966 56868 20018
rect 56140 19234 56196 19246
rect 56140 19182 56142 19234
rect 56194 19182 56196 19234
rect 54908 18060 55412 18116
rect 55580 18452 55636 18462
rect 54572 16882 54628 16894
rect 54572 16830 54574 16882
rect 54626 16830 54628 16882
rect 53116 15986 53620 15988
rect 53116 15934 53566 15986
rect 53618 15934 53620 15986
rect 53116 15932 53620 15934
rect 52220 15262 52222 15314
rect 52274 15262 52276 15314
rect 52220 15148 52276 15262
rect 52780 15314 52836 15326
rect 52780 15262 52782 15314
rect 52834 15262 52836 15314
rect 52220 15092 52724 15148
rect 51548 14578 51604 14588
rect 52668 13858 52724 15092
rect 52780 14754 52836 15262
rect 52780 14702 52782 14754
rect 52834 14702 52836 14754
rect 52780 14690 52836 14702
rect 52892 14644 52948 14654
rect 52892 14550 52948 14588
rect 52668 13806 52670 13858
rect 52722 13806 52724 13858
rect 52668 13794 52724 13806
rect 53004 14530 53060 14542
rect 53004 14478 53006 14530
rect 53058 14478 53060 14530
rect 51996 13748 52052 13758
rect 51436 13746 52052 13748
rect 51436 13694 51998 13746
rect 52050 13694 52052 13746
rect 51436 13692 52052 13694
rect 51660 13524 51716 13534
rect 51660 13074 51716 13468
rect 51660 13022 51662 13074
rect 51714 13022 51716 13074
rect 51660 13010 51716 13022
rect 51996 12964 52052 13692
rect 53004 13524 53060 14478
rect 53004 13458 53060 13468
rect 52108 12964 52164 12974
rect 51996 12962 52164 12964
rect 51996 12910 52110 12962
rect 52162 12910 52164 12962
rect 51996 12908 52164 12910
rect 51100 12798 51102 12850
rect 51154 12798 51156 12850
rect 49532 12740 49588 12750
rect 49588 12684 49700 12740
rect 49532 12674 49588 12684
rect 49084 12348 49252 12404
rect 49084 11954 49140 12348
rect 49644 12180 49700 12684
rect 50556 12572 50820 12582
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 51100 12516 51156 12798
rect 50556 12506 50820 12516
rect 50876 12460 51156 12516
rect 50764 12404 50820 12414
rect 50876 12404 50932 12460
rect 50764 12402 50932 12404
rect 50764 12350 50766 12402
rect 50818 12350 50932 12402
rect 50764 12348 50932 12350
rect 51884 12404 51940 12414
rect 50764 12338 50820 12348
rect 51884 12310 51940 12348
rect 51660 12292 51716 12302
rect 51660 12198 51716 12236
rect 52108 12290 52164 12908
rect 53004 12852 53060 12862
rect 53116 12852 53172 15932
rect 53564 15922 53620 15932
rect 53676 16324 53732 16334
rect 53676 15986 53732 16268
rect 54572 16324 54628 16830
rect 54572 16258 54628 16268
rect 54908 16882 54964 18060
rect 55580 17778 55636 18396
rect 55580 17726 55582 17778
rect 55634 17726 55636 17778
rect 55580 17714 55636 17726
rect 55916 18340 55972 18350
rect 55916 17108 55972 18284
rect 56140 17668 56196 19182
rect 56588 18564 56644 18574
rect 56812 18564 56868 19966
rect 56588 18562 56868 18564
rect 56588 18510 56590 18562
rect 56642 18510 56868 18562
rect 56588 18508 56868 18510
rect 56588 18498 56644 18508
rect 56140 17574 56196 17612
rect 54908 16830 54910 16882
rect 54962 16830 54964 16882
rect 53676 15934 53678 15986
rect 53730 15934 53732 15986
rect 53676 15922 53732 15934
rect 53900 15988 53956 15998
rect 54236 15988 54292 15998
rect 53900 15986 54292 15988
rect 53900 15934 53902 15986
rect 53954 15934 54238 15986
rect 54290 15934 54292 15986
rect 53900 15932 54292 15934
rect 53900 15922 53956 15932
rect 54012 15426 54068 15932
rect 54236 15922 54292 15932
rect 54348 15876 54404 15886
rect 54348 15782 54404 15820
rect 54012 15374 54014 15426
rect 54066 15374 54068 15426
rect 54012 15362 54068 15374
rect 53788 15202 53844 15214
rect 53788 15150 53790 15202
rect 53842 15150 53844 15202
rect 53788 15148 53844 15150
rect 54908 15148 54964 16830
rect 55020 16994 55076 17006
rect 55020 16942 55022 16994
rect 55074 16942 55076 16994
rect 55020 16324 55076 16942
rect 55580 16996 55636 17006
rect 55244 16884 55300 16894
rect 55468 16884 55524 16894
rect 55244 16882 55468 16884
rect 55244 16830 55246 16882
rect 55298 16830 55468 16882
rect 55244 16828 55468 16830
rect 55244 16818 55300 16828
rect 55468 16790 55524 16828
rect 55020 16258 55076 16268
rect 55132 16772 55188 16782
rect 55132 16098 55188 16716
rect 55580 16322 55636 16940
rect 55580 16270 55582 16322
rect 55634 16270 55636 16322
rect 55580 16258 55636 16270
rect 55692 16658 55748 16670
rect 55692 16606 55694 16658
rect 55746 16606 55748 16658
rect 55132 16046 55134 16098
rect 55186 16046 55188 16098
rect 55132 16034 55188 16046
rect 55356 16210 55412 16222
rect 55356 16158 55358 16210
rect 55410 16158 55412 16210
rect 55244 15316 55300 15326
rect 53452 15092 53844 15148
rect 54572 15092 54964 15148
rect 55020 15314 55300 15316
rect 55020 15262 55246 15314
rect 55298 15262 55300 15314
rect 55020 15260 55300 15262
rect 53228 14530 53284 14542
rect 53228 14478 53230 14530
rect 53282 14478 53284 14530
rect 53228 13860 53284 14478
rect 53452 13970 53508 15092
rect 53452 13918 53454 13970
rect 53506 13918 53508 13970
rect 53452 13906 53508 13918
rect 54236 14530 54292 14542
rect 54460 14532 54516 14542
rect 54236 14478 54238 14530
rect 54290 14478 54292 14530
rect 53228 13794 53284 13804
rect 53676 13748 53732 13758
rect 53340 13524 53396 13534
rect 53340 13430 53396 13468
rect 53676 13186 53732 13692
rect 54236 13748 54292 14478
rect 54236 13682 54292 13692
rect 54348 14530 54516 14532
rect 54348 14478 54462 14530
rect 54514 14478 54516 14530
rect 54348 14476 54516 14478
rect 54348 13746 54404 14476
rect 54460 14466 54516 14476
rect 54460 14308 54516 14318
rect 54460 13970 54516 14252
rect 54572 14084 54628 15092
rect 54684 14530 54740 14542
rect 54684 14478 54686 14530
rect 54738 14478 54740 14530
rect 54684 14196 54740 14478
rect 55020 14196 55076 15260
rect 55244 15250 55300 15260
rect 55356 15148 55412 16158
rect 55692 16100 55748 16606
rect 55804 16100 55860 16110
rect 55692 16044 55804 16100
rect 55804 16034 55860 16044
rect 55804 15876 55860 15886
rect 55132 15092 55188 15102
rect 55356 15092 55524 15148
rect 55132 14756 55188 15036
rect 55132 14754 55300 14756
rect 55132 14702 55134 14754
rect 55186 14702 55300 14754
rect 55132 14700 55300 14702
rect 55132 14690 55188 14700
rect 55244 14530 55300 14700
rect 55468 14642 55524 15092
rect 55468 14590 55470 14642
rect 55522 14590 55524 14642
rect 55468 14578 55524 14590
rect 55244 14478 55246 14530
rect 55298 14478 55300 14530
rect 55244 14466 55300 14478
rect 55804 14530 55860 15820
rect 55916 15426 55972 17052
rect 56924 17106 56980 20636
rect 57820 20626 57876 20638
rect 58268 20242 58324 20748
rect 58268 20190 58270 20242
rect 58322 20190 58324 20242
rect 58268 20178 58324 20190
rect 57484 19348 57540 19358
rect 56924 17054 56926 17106
rect 56978 17054 56980 17106
rect 56924 17042 56980 17054
rect 57148 19234 57204 19246
rect 57484 19236 57540 19292
rect 57148 19182 57150 19234
rect 57202 19182 57204 19234
rect 57148 18450 57204 19182
rect 57148 18398 57150 18450
rect 57202 18398 57204 18450
rect 57148 17666 57204 18398
rect 57148 17614 57150 17666
rect 57202 17614 57204 17666
rect 57148 16996 57204 17614
rect 57372 19234 57540 19236
rect 57372 19182 57486 19234
rect 57538 19182 57540 19234
rect 57372 19180 57540 19182
rect 57372 17554 57428 19180
rect 57484 19170 57540 19180
rect 57372 17502 57374 17554
rect 57426 17502 57428 17554
rect 57372 17490 57428 17502
rect 57484 18338 57540 18350
rect 57484 18286 57486 18338
rect 57538 18286 57540 18338
rect 57484 17668 57540 18286
rect 57372 16996 57428 17006
rect 57148 16940 57372 16996
rect 57372 16902 57428 16940
rect 56028 16884 56084 16894
rect 56700 16884 56756 16894
rect 56028 16882 56756 16884
rect 56028 16830 56030 16882
rect 56082 16830 56702 16882
rect 56754 16830 56756 16882
rect 56028 16828 56756 16830
rect 56028 16818 56084 16828
rect 56700 16818 56756 16828
rect 56812 16884 56868 16894
rect 57484 16884 57540 17612
rect 57820 16884 57876 16894
rect 57484 16882 57876 16884
rect 57484 16830 57822 16882
rect 57874 16830 57876 16882
rect 57484 16828 57876 16830
rect 55916 15374 55918 15426
rect 55970 15374 55972 15426
rect 55916 15362 55972 15374
rect 56028 16100 56084 16110
rect 55804 14478 55806 14530
rect 55858 14478 55860 14530
rect 55804 14466 55860 14478
rect 56028 14532 56084 16044
rect 56140 16098 56196 16110
rect 56140 16046 56142 16098
rect 56194 16046 56196 16098
rect 56140 15540 56196 16046
rect 56476 16100 56532 16110
rect 56476 16006 56532 16044
rect 56812 16098 56868 16828
rect 57820 16212 57876 16828
rect 57932 16212 57988 16222
rect 57820 16210 57988 16212
rect 57820 16158 57934 16210
rect 57986 16158 57988 16210
rect 57820 16156 57988 16158
rect 57932 16146 57988 16156
rect 56812 16046 56814 16098
rect 56866 16046 56868 16098
rect 56812 16034 56868 16046
rect 56588 15876 56644 15886
rect 56476 15540 56532 15550
rect 56140 15538 56532 15540
rect 56140 15486 56478 15538
rect 56530 15486 56532 15538
rect 56140 15484 56532 15486
rect 56476 15474 56532 15484
rect 56588 15538 56644 15820
rect 56588 15486 56590 15538
rect 56642 15486 56644 15538
rect 56588 15474 56644 15486
rect 56812 15314 56868 15326
rect 56812 15262 56814 15314
rect 56866 15262 56868 15314
rect 56812 15148 56868 15262
rect 56476 15092 56868 15148
rect 57036 15314 57092 15326
rect 57036 15262 57038 15314
rect 57090 15262 57092 15314
rect 57036 15204 57092 15262
rect 57036 15138 57092 15148
rect 56140 14532 56196 14542
rect 56028 14530 56196 14532
rect 56028 14478 56142 14530
rect 56194 14478 56196 14530
rect 56028 14476 56196 14478
rect 56140 14466 56196 14476
rect 55692 14418 55748 14430
rect 55692 14366 55694 14418
rect 55746 14366 55748 14418
rect 55692 14308 55748 14366
rect 56476 14418 56532 15092
rect 56476 14366 56478 14418
rect 56530 14366 56532 14418
rect 56364 14308 56420 14318
rect 55692 14242 55748 14252
rect 55804 14306 56420 14308
rect 55804 14254 56366 14306
rect 56418 14254 56420 14306
rect 55804 14252 56420 14254
rect 54684 14140 55076 14196
rect 54572 14028 54964 14084
rect 54460 13918 54462 13970
rect 54514 13918 54516 13970
rect 54460 13906 54516 13918
rect 54796 13860 54852 13870
rect 54348 13694 54350 13746
rect 54402 13694 54404 13746
rect 54348 13524 54404 13694
rect 54572 13748 54628 13758
rect 54572 13654 54628 13692
rect 54348 13458 54404 13468
rect 54572 13524 54628 13534
rect 53676 13134 53678 13186
rect 53730 13134 53732 13186
rect 53676 13122 53732 13134
rect 54572 12962 54628 13468
rect 54796 12964 54852 13804
rect 54572 12910 54574 12962
rect 54626 12910 54628 12962
rect 53004 12850 53172 12852
rect 53004 12798 53006 12850
rect 53058 12798 53172 12850
rect 53004 12796 53172 12798
rect 53340 12850 53396 12862
rect 53340 12798 53342 12850
rect 53394 12798 53396 12850
rect 53004 12786 53060 12796
rect 52108 12238 52110 12290
rect 52162 12238 52164 12290
rect 52108 12226 52164 12238
rect 52668 12738 52724 12750
rect 52668 12686 52670 12738
rect 52722 12686 52724 12738
rect 49644 12086 49700 12124
rect 50204 12180 50260 12190
rect 50204 12086 50260 12124
rect 50876 12180 50932 12190
rect 49532 12068 49588 12078
rect 49084 11902 49086 11954
rect 49138 11902 49140 11954
rect 49084 11890 49140 11902
rect 49196 12012 49532 12068
rect 48636 11620 48692 11630
rect 48412 11618 48692 11620
rect 48412 11566 48638 11618
rect 48690 11566 48692 11618
rect 48412 11564 48692 11566
rect 48636 11554 48692 11564
rect 47516 11454 47518 11506
rect 47570 11454 47572 11506
rect 47516 11442 47572 11454
rect 47628 11396 47684 11406
rect 47628 11302 47684 11340
rect 47852 10836 47908 10846
rect 47852 10742 47908 10780
rect 47404 10612 47460 10668
rect 49196 10722 49252 12012
rect 49532 11974 49588 12012
rect 50428 12068 50484 12078
rect 50428 11974 50484 12012
rect 49196 10670 49198 10722
rect 49250 10670 49252 10722
rect 49196 10658 49252 10670
rect 49868 11396 49924 11406
rect 49868 10836 49924 11340
rect 47516 10612 47572 10622
rect 47404 10610 47572 10612
rect 47404 10558 47518 10610
rect 47570 10558 47572 10610
rect 47404 10556 47572 10558
rect 47516 10546 47572 10556
rect 47852 10612 47908 10622
rect 47852 10518 47908 10556
rect 48188 10610 48244 10622
rect 48188 10558 48190 10610
rect 48242 10558 48244 10610
rect 47180 9324 47572 9380
rect 47068 9214 47070 9266
rect 47122 9214 47124 9266
rect 46396 8642 46452 8652
rect 46844 9042 46900 9054
rect 46844 8990 46846 9042
rect 46898 8990 46900 9042
rect 46844 8484 46900 8990
rect 46844 8418 46900 8428
rect 46172 8318 46174 8370
rect 46226 8318 46228 8370
rect 46172 8306 46228 8318
rect 47068 7924 47124 9214
rect 47180 9156 47236 9166
rect 47180 9062 47236 9100
rect 47404 8820 47460 8830
rect 47292 8260 47348 8270
rect 46956 7868 47124 7924
rect 47180 8204 47292 8260
rect 44828 6862 44830 6914
rect 44882 6862 44884 6914
rect 44828 6850 44884 6862
rect 45276 6860 45668 6916
rect 45724 7420 45892 7476
rect 46060 7474 46116 7486
rect 46060 7422 46062 7474
rect 46114 7422 46116 7474
rect 44156 6802 44212 6814
rect 44156 6750 44158 6802
rect 44210 6750 44212 6802
rect 44156 6692 44212 6750
rect 44940 6804 44996 6814
rect 44940 6710 44996 6748
rect 44156 6626 44212 6636
rect 45052 6468 45108 6478
rect 44940 6466 45108 6468
rect 44940 6414 45054 6466
rect 45106 6414 45108 6466
rect 44940 6412 45108 6414
rect 44044 6076 44212 6132
rect 44044 5908 44100 5918
rect 44156 5908 44212 6076
rect 44604 6020 44660 6030
rect 44940 6020 44996 6412
rect 45052 6402 45108 6412
rect 45276 6244 45332 6860
rect 44660 5964 44996 6020
rect 45052 6188 45332 6244
rect 45388 6692 45444 6702
rect 44156 5852 44548 5908
rect 44044 5814 44100 5852
rect 44380 5684 44436 5694
rect 43932 5628 44100 5684
rect 43820 5618 43876 5628
rect 43708 5572 43764 5582
rect 43036 5070 43038 5122
rect 43090 5070 43092 5122
rect 43036 4788 43092 5070
rect 43484 5348 43540 5358
rect 43708 5348 43764 5516
rect 43484 5122 43540 5292
rect 43484 5070 43486 5122
rect 43538 5070 43540 5122
rect 43484 5058 43540 5070
rect 43596 5292 43764 5348
rect 43932 5460 43988 5470
rect 43596 5122 43652 5292
rect 43820 5124 43876 5134
rect 43596 5070 43598 5122
rect 43650 5070 43652 5122
rect 43596 5058 43652 5070
rect 43708 5068 43820 5124
rect 43260 4900 43316 4910
rect 43260 4806 43316 4844
rect 43372 4898 43428 4910
rect 43708 4900 43764 5068
rect 43820 5058 43876 5068
rect 43932 5122 43988 5404
rect 43932 5070 43934 5122
rect 43986 5070 43988 5122
rect 43932 5058 43988 5070
rect 43372 4846 43374 4898
rect 43426 4846 43428 4898
rect 43036 4676 43092 4732
rect 43036 4620 43316 4676
rect 42924 4498 42980 4508
rect 42252 4338 42644 4340
rect 42252 4286 42254 4338
rect 42306 4286 42478 4338
rect 42530 4286 42644 4338
rect 42252 4284 42644 4286
rect 42700 4340 42756 4350
rect 43148 4340 43204 4350
rect 42756 4284 43092 4340
rect 42252 4274 42308 4284
rect 42476 4274 42532 4284
rect 42700 4246 42756 4284
rect 40348 3666 41076 3668
rect 40348 3614 40350 3666
rect 40402 3614 40910 3666
rect 40962 3614 41076 3666
rect 40348 3612 41076 3614
rect 41804 3668 41860 3678
rect 40348 3602 40404 3612
rect 40908 3602 40964 3612
rect 41804 3574 41860 3612
rect 39788 3556 39844 3566
rect 39340 3554 39844 3556
rect 39340 3502 39790 3554
rect 39842 3502 39844 3554
rect 39340 3500 39844 3502
rect 42140 3556 42196 3724
rect 42252 3556 42308 3566
rect 42140 3554 42308 3556
rect 42140 3502 42254 3554
rect 42306 3502 42308 3554
rect 42140 3500 42308 3502
rect 39788 3490 39844 3500
rect 42252 3490 42308 3500
rect 38892 3390 38894 3442
rect 38946 3390 38948 3442
rect 38892 3378 38948 3390
rect 39004 3444 39060 3454
rect 39004 800 39060 3388
rect 42700 3442 42756 3454
rect 42700 3390 42702 3442
rect 42754 3390 42756 3442
rect 42700 3220 42756 3390
rect 43036 3442 43092 4284
rect 43148 4246 43204 4284
rect 43260 4338 43316 4620
rect 43260 4286 43262 4338
rect 43314 4286 43316 4338
rect 43260 4274 43316 4286
rect 43372 4228 43428 4846
rect 43372 4162 43428 4172
rect 43484 4844 43764 4900
rect 43820 4900 43876 4910
rect 43484 4338 43540 4844
rect 43484 4286 43486 4338
rect 43538 4286 43540 4338
rect 43036 3390 43038 3442
rect 43090 3390 43092 3442
rect 43036 3378 43092 3390
rect 43148 3668 43204 3678
rect 42700 3154 42756 3164
rect 39676 2660 39732 2670
rect 39676 800 39732 2604
rect 43148 1876 43204 3612
rect 43484 3332 43540 4286
rect 43596 4564 43652 4574
rect 43596 3442 43652 4508
rect 43820 4562 43876 4844
rect 43820 4510 43822 4562
rect 43874 4510 43876 4562
rect 43820 4498 43876 4510
rect 43596 3390 43598 3442
rect 43650 3390 43652 3442
rect 43596 3378 43652 3390
rect 43932 3780 43988 3790
rect 43932 3554 43988 3724
rect 43932 3502 43934 3554
rect 43986 3502 43988 3554
rect 43484 3266 43540 3276
rect 43932 2548 43988 3502
rect 44044 3444 44100 5628
rect 44492 5684 44548 5852
rect 44604 5906 44660 5964
rect 44604 5854 44606 5906
rect 44658 5854 44660 5906
rect 44604 5842 44660 5854
rect 44492 5628 44772 5684
rect 44380 5348 44436 5628
rect 44380 5292 44660 5348
rect 44156 5236 44212 5246
rect 44156 5010 44212 5180
rect 44604 5124 44660 5292
rect 44380 5068 44660 5124
rect 44156 4958 44158 5010
rect 44210 4958 44212 5010
rect 44156 4946 44212 4958
rect 44268 5012 44324 5022
rect 44268 4918 44324 4956
rect 44380 4338 44436 5068
rect 44716 4562 44772 5628
rect 44828 5124 44884 5134
rect 44828 5030 44884 5068
rect 44716 4510 44718 4562
rect 44770 4510 44772 4562
rect 44716 4498 44772 4510
rect 44380 4286 44382 4338
rect 44434 4286 44436 4338
rect 44380 4274 44436 4286
rect 44940 4338 44996 4350
rect 44940 4286 44942 4338
rect 44994 4286 44996 4338
rect 44940 4004 44996 4286
rect 44940 3938 44996 3948
rect 44492 3892 44548 3902
rect 44492 3554 44548 3836
rect 44492 3502 44494 3554
rect 44546 3502 44548 3554
rect 44492 3490 44548 3502
rect 44268 3444 44324 3454
rect 44044 3442 44324 3444
rect 44044 3390 44270 3442
rect 44322 3390 44324 3442
rect 44044 3388 44324 3390
rect 44268 3378 44324 3388
rect 44940 3444 44996 3454
rect 45052 3444 45108 6188
rect 45388 5906 45444 6636
rect 45612 6468 45668 6478
rect 45612 6374 45668 6412
rect 45388 5854 45390 5906
rect 45442 5854 45444 5906
rect 45164 5796 45220 5806
rect 45164 5702 45220 5740
rect 45164 5348 45220 5358
rect 45164 5010 45220 5292
rect 45388 5236 45444 5854
rect 45612 5236 45668 5246
rect 45388 5234 45668 5236
rect 45388 5182 45614 5234
rect 45666 5182 45668 5234
rect 45388 5180 45668 5182
rect 45612 5170 45668 5180
rect 45164 4958 45166 5010
rect 45218 4958 45220 5010
rect 45164 4946 45220 4958
rect 45612 5012 45668 5022
rect 45388 4788 45444 4798
rect 45388 4562 45444 4732
rect 45388 4510 45390 4562
rect 45442 4510 45444 4562
rect 45388 4498 45444 4510
rect 45612 4340 45668 4956
rect 45612 4246 45668 4284
rect 45164 3556 45220 3566
rect 45164 3462 45220 3500
rect 44940 3442 45108 3444
rect 44940 3390 44942 3442
rect 44994 3390 45108 3442
rect 44940 3388 45108 3390
rect 45612 3444 45668 3454
rect 45724 3444 45780 7420
rect 46060 7364 46116 7422
rect 46060 6692 46116 7308
rect 46844 7476 46900 7486
rect 46396 6692 46452 6702
rect 46060 6690 46452 6692
rect 46060 6638 46398 6690
rect 46450 6638 46452 6690
rect 46060 6636 46452 6638
rect 46060 6468 46116 6478
rect 46060 6132 46116 6412
rect 45836 6130 46116 6132
rect 45836 6078 46062 6130
rect 46114 6078 46116 6130
rect 45836 6076 46116 6078
rect 45836 5572 45892 6076
rect 46060 6066 46116 6076
rect 45948 5906 46004 5918
rect 45948 5854 45950 5906
rect 46002 5854 46004 5906
rect 45948 5684 46004 5854
rect 46396 5796 46452 6636
rect 46844 6578 46900 7420
rect 46956 7364 47012 7868
rect 47068 7700 47124 7710
rect 47068 7586 47124 7644
rect 47068 7534 47070 7586
rect 47122 7534 47124 7586
rect 47068 7522 47124 7534
rect 47180 7588 47236 8204
rect 47292 8166 47348 8204
rect 47180 7586 47348 7588
rect 47180 7534 47182 7586
rect 47234 7534 47348 7586
rect 47180 7532 47348 7534
rect 47180 7522 47236 7532
rect 46956 7308 47124 7364
rect 46844 6526 46846 6578
rect 46898 6526 46900 6578
rect 46844 6020 46900 6526
rect 47068 6468 47124 7308
rect 47292 6692 47348 7532
rect 47292 6598 47348 6636
rect 47068 6402 47124 6412
rect 47404 6466 47460 8764
rect 47516 6580 47572 9324
rect 48188 9268 48244 10558
rect 49868 10610 49924 10780
rect 49868 10558 49870 10610
rect 49922 10558 49924 10610
rect 49868 10546 49924 10558
rect 49980 11394 50036 11406
rect 49980 11342 49982 11394
rect 50034 11342 50036 11394
rect 49980 10500 50036 11342
rect 50764 11396 50820 11406
rect 50764 11302 50820 11340
rect 50876 11282 50932 12124
rect 50876 11230 50878 11282
rect 50930 11230 50932 11282
rect 50876 11218 50932 11230
rect 51548 12180 51604 12190
rect 50556 11004 50820 11014
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50556 10938 50820 10948
rect 50092 10500 50148 10510
rect 49980 10498 50148 10500
rect 49980 10446 50094 10498
rect 50146 10446 50148 10498
rect 49980 10444 50148 10446
rect 50092 9828 50148 10444
rect 51212 9940 51268 9950
rect 50092 9762 50148 9772
rect 51100 9884 51212 9940
rect 50556 9436 50820 9446
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50556 9370 50820 9380
rect 48188 9202 48244 9212
rect 48860 9268 48916 9278
rect 48860 9174 48916 9212
rect 49756 9156 49812 9166
rect 49756 9154 49924 9156
rect 49756 9102 49758 9154
rect 49810 9102 49924 9154
rect 49756 9100 49924 9102
rect 49756 9090 49812 9100
rect 48748 9042 48804 9054
rect 48748 8990 48750 9042
rect 48802 8990 48804 9042
rect 48300 8372 48356 8382
rect 48300 8146 48356 8316
rect 48300 8094 48302 8146
rect 48354 8094 48356 8146
rect 48300 8082 48356 8094
rect 48300 7924 48356 7934
rect 47628 7700 47684 7710
rect 47628 7606 47684 7644
rect 48300 7698 48356 7868
rect 48300 7646 48302 7698
rect 48354 7646 48356 7698
rect 48300 7634 48356 7646
rect 48748 7700 48804 8990
rect 49644 8932 49700 8942
rect 48972 8820 49028 8830
rect 48972 8726 49028 8764
rect 49196 8818 49252 8830
rect 49196 8766 49198 8818
rect 49250 8766 49252 8818
rect 49196 8596 49252 8766
rect 49196 8530 49252 8540
rect 49532 8484 49588 8494
rect 48860 8372 48916 8382
rect 49420 8372 49476 8382
rect 48860 8370 49476 8372
rect 48860 8318 48862 8370
rect 48914 8318 49422 8370
rect 49474 8318 49476 8370
rect 48860 8316 49476 8318
rect 48860 7924 48916 8316
rect 49420 8306 49476 8316
rect 49532 8148 49588 8428
rect 49308 8092 49588 8148
rect 48860 7858 48916 7868
rect 48972 8036 49028 8046
rect 48076 7586 48132 7598
rect 48076 7534 48078 7586
rect 48130 7534 48132 7586
rect 47964 7474 48020 7486
rect 47964 7422 47966 7474
rect 48018 7422 48020 7474
rect 47964 7364 48020 7422
rect 48076 7476 48132 7534
rect 48076 7410 48132 7420
rect 48748 7474 48804 7644
rect 48748 7422 48750 7474
rect 48802 7422 48804 7474
rect 48748 7410 48804 7422
rect 48972 7474 49028 7980
rect 48972 7422 48974 7474
rect 49026 7422 49028 7474
rect 48972 7410 49028 7422
rect 49308 7474 49364 8092
rect 49532 7700 49588 7710
rect 49644 7700 49700 8876
rect 49756 8484 49812 8494
rect 49756 8258 49812 8428
rect 49756 8206 49758 8258
rect 49810 8206 49812 8258
rect 49756 8194 49812 8206
rect 49756 8036 49812 8046
rect 49868 8036 49924 9100
rect 50652 9154 50708 9166
rect 50652 9102 50654 9154
rect 50706 9102 50708 9154
rect 49980 9042 50036 9054
rect 49980 8990 49982 9042
rect 50034 8990 50036 9042
rect 49980 8820 50036 8990
rect 49980 8754 50036 8764
rect 50428 8820 50484 8830
rect 50428 8726 50484 8764
rect 49812 7980 49924 8036
rect 49980 8596 50036 8606
rect 49756 7970 49812 7980
rect 49532 7698 49700 7700
rect 49532 7646 49534 7698
rect 49586 7646 49700 7698
rect 49532 7644 49700 7646
rect 49532 7634 49588 7644
rect 49308 7422 49310 7474
rect 49362 7422 49364 7474
rect 49308 7410 49364 7422
rect 49420 7476 49476 7486
rect 49420 7382 49476 7420
rect 49644 7476 49700 7486
rect 49980 7476 50036 8540
rect 50652 8036 50708 9102
rect 50764 8820 50820 8830
rect 50764 8818 51044 8820
rect 50764 8766 50766 8818
rect 50818 8766 51044 8818
rect 50764 8764 51044 8766
rect 50764 8754 50820 8764
rect 50876 8260 50932 8270
rect 50876 8166 50932 8204
rect 50652 7980 50932 8036
rect 50556 7868 50820 7878
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50556 7802 50820 7812
rect 50764 7700 50820 7710
rect 50652 7644 50764 7700
rect 50204 7588 50260 7598
rect 50204 7494 50260 7532
rect 50428 7586 50484 7598
rect 50428 7534 50430 7586
rect 50482 7534 50484 7586
rect 49644 7474 50036 7476
rect 49644 7422 49646 7474
rect 49698 7422 50036 7474
rect 49644 7420 50036 7422
rect 49644 7410 49700 7420
rect 47964 7298 48020 7308
rect 50428 6916 50484 7534
rect 50540 7588 50596 7598
rect 50652 7588 50708 7644
rect 50764 7634 50820 7644
rect 50540 7586 50708 7588
rect 50540 7534 50542 7586
rect 50594 7534 50708 7586
rect 50540 7532 50708 7534
rect 50540 7522 50596 7532
rect 50428 6860 50596 6916
rect 47516 6514 47572 6524
rect 49308 6692 49364 6702
rect 47404 6414 47406 6466
rect 47458 6414 47460 6466
rect 47404 6402 47460 6414
rect 48860 6132 48916 6142
rect 48860 6130 49140 6132
rect 48860 6078 48862 6130
rect 48914 6078 49140 6130
rect 48860 6076 49140 6078
rect 48860 6066 48916 6076
rect 46844 5964 47236 6020
rect 46396 5730 46452 5740
rect 46620 5794 46676 5806
rect 46620 5742 46622 5794
rect 46674 5742 46676 5794
rect 45948 5618 46004 5628
rect 46060 5682 46116 5694
rect 46060 5630 46062 5682
rect 46114 5630 46116 5682
rect 45836 4900 45892 5516
rect 45948 5234 46004 5246
rect 45948 5182 45950 5234
rect 46002 5182 46004 5234
rect 45948 5124 46004 5182
rect 45948 5058 46004 5068
rect 46060 5236 46116 5630
rect 46620 5684 46676 5742
rect 46620 5618 46676 5628
rect 47068 5794 47124 5806
rect 47068 5742 47070 5794
rect 47122 5742 47124 5794
rect 46956 5236 47012 5246
rect 46060 5234 47012 5236
rect 46060 5182 46958 5234
rect 47010 5182 47012 5234
rect 46060 5180 47012 5182
rect 46060 5122 46116 5180
rect 46956 5170 47012 5180
rect 46060 5070 46062 5122
rect 46114 5070 46116 5122
rect 46060 5058 46116 5070
rect 45836 4844 46116 4900
rect 46060 4562 46116 4844
rect 46060 4510 46062 4562
rect 46114 4510 46116 4562
rect 46060 4498 46116 4510
rect 46396 4452 46452 4462
rect 46396 4358 46452 4396
rect 46284 4340 46340 4350
rect 45612 3442 45780 3444
rect 45612 3390 45614 3442
rect 45666 3390 45780 3442
rect 45612 3388 45780 3390
rect 45948 4228 46004 4238
rect 45948 3554 46004 4172
rect 45948 3502 45950 3554
rect 46002 3502 46004 3554
rect 44940 3378 44996 3388
rect 45612 3378 45668 3388
rect 45948 3332 46004 3502
rect 46284 3442 46340 4284
rect 46844 4226 46900 4238
rect 46844 4174 46846 4226
rect 46898 4174 46900 4226
rect 46844 3780 46900 4174
rect 46844 3714 46900 3724
rect 46284 3390 46286 3442
rect 46338 3390 46340 3442
rect 46284 3378 46340 3390
rect 46620 3556 46676 3566
rect 47068 3556 47124 5742
rect 47180 5348 47236 5964
rect 48972 5908 49028 5918
rect 48972 5814 49028 5852
rect 48860 5684 48916 5694
rect 48860 5590 48916 5628
rect 47516 5348 47572 5358
rect 47180 5346 47572 5348
rect 47180 5294 47518 5346
rect 47570 5294 47572 5346
rect 47180 5292 47572 5294
rect 47516 5282 47572 5292
rect 47964 5348 48020 5358
rect 47180 5124 47236 5134
rect 47740 5124 47796 5134
rect 47236 5122 47796 5124
rect 47236 5070 47742 5122
rect 47794 5070 47796 5122
rect 47236 5068 47796 5070
rect 47180 5030 47236 5068
rect 47740 5058 47796 5068
rect 47964 5010 48020 5292
rect 49084 5348 49140 6076
rect 49308 6018 49364 6636
rect 50428 6692 50484 6702
rect 49308 5966 49310 6018
rect 49362 5966 49364 6018
rect 49308 5954 49364 5966
rect 49532 6580 49588 6590
rect 47964 4958 47966 5010
rect 48018 4958 48020 5010
rect 47964 4946 48020 4958
rect 48076 5124 48132 5134
rect 48076 5010 48132 5068
rect 48076 4958 48078 5010
rect 48130 4958 48132 5010
rect 48076 4946 48132 4958
rect 48412 5124 48468 5134
rect 47404 4452 47460 4462
rect 47292 4226 47348 4238
rect 47292 4174 47294 4226
rect 47346 4174 47348 4226
rect 47292 4004 47348 4174
rect 47292 3938 47348 3948
rect 46620 3554 47124 3556
rect 46620 3502 46622 3554
rect 46674 3502 47124 3554
rect 46620 3500 47124 3502
rect 47292 3556 47348 3566
rect 46620 3388 46676 3500
rect 47292 3388 47348 3500
rect 45948 3266 46004 3276
rect 46508 3332 46676 3388
rect 47068 3332 47348 3388
rect 47404 3442 47460 4396
rect 47740 4226 47796 4238
rect 47740 4174 47742 4226
rect 47794 4174 47796 4226
rect 47740 3892 47796 4174
rect 48188 4228 48244 4238
rect 48188 4134 48244 4172
rect 47740 3826 47796 3836
rect 47628 3668 47684 3678
rect 47628 3554 47684 3612
rect 47628 3502 47630 3554
rect 47682 3502 47684 3554
rect 47628 3490 47684 3502
rect 48188 3556 48244 3566
rect 48188 3462 48244 3500
rect 47404 3390 47406 3442
rect 47458 3390 47460 3442
rect 47404 3378 47460 3390
rect 48412 3442 48468 5068
rect 49084 5122 49140 5292
rect 49532 5234 49588 6524
rect 50316 6580 50372 6590
rect 50316 6486 50372 6524
rect 49980 6468 50036 6478
rect 49868 6466 50036 6468
rect 49868 6414 49982 6466
rect 50034 6414 50036 6466
rect 49868 6412 50036 6414
rect 49868 6132 49924 6412
rect 49980 6402 50036 6412
rect 49868 5796 49924 6076
rect 49868 5730 49924 5740
rect 49980 5906 50036 5918
rect 49980 5854 49982 5906
rect 50034 5854 50036 5906
rect 49980 5684 50036 5854
rect 49980 5618 50036 5628
rect 50204 5908 50260 5918
rect 49532 5182 49534 5234
rect 49586 5182 49588 5234
rect 49532 5170 49588 5182
rect 49084 5070 49086 5122
rect 49138 5070 49140 5122
rect 49084 5058 49140 5070
rect 49980 5124 50036 5134
rect 49980 5030 50036 5068
rect 48860 4226 48916 4238
rect 48860 4174 48862 4226
rect 48914 4174 48916 4226
rect 48860 3556 48916 4174
rect 49756 4226 49812 4238
rect 49756 4174 49758 4226
rect 49810 4174 49812 4226
rect 49308 3668 49364 3678
rect 49308 3574 49364 3612
rect 48860 3490 48916 3500
rect 49756 3556 49812 4174
rect 49980 3556 50036 3566
rect 49756 3554 50036 3556
rect 49756 3502 49982 3554
rect 50034 3502 50036 3554
rect 49756 3500 50036 3502
rect 48412 3390 48414 3442
rect 48466 3390 48468 3442
rect 48412 3378 48468 3390
rect 48748 3444 48804 3454
rect 48748 3332 48804 3388
rect 48860 3332 48916 3342
rect 46508 2660 46564 3332
rect 46508 2594 46564 2604
rect 43932 2482 43988 2492
rect 43036 1820 43204 1876
rect 43036 800 43092 1820
rect 47068 800 47124 3332
rect 48748 3330 48916 3332
rect 48748 3278 48862 3330
rect 48914 3278 48916 3330
rect 48748 3276 48916 3278
rect 48860 3266 48916 3276
rect 49756 800 49812 3500
rect 49980 3490 50036 3500
rect 50204 3444 50260 5852
rect 50428 5906 50484 6636
rect 50540 6468 50596 6860
rect 50652 6690 50708 7532
rect 50876 6916 50932 7980
rect 50988 7362 51044 8764
rect 51100 7700 51156 9884
rect 51212 9874 51268 9884
rect 51548 9828 51604 12124
rect 52668 12180 52724 12686
rect 52668 12114 52724 12124
rect 52892 12178 52948 12190
rect 52892 12126 52894 12178
rect 52946 12126 52948 12178
rect 52892 11506 52948 12126
rect 52892 11454 52894 11506
rect 52946 11454 52948 11506
rect 52892 10724 52948 11454
rect 53228 12068 53284 12078
rect 53340 12068 53396 12798
rect 53564 12738 53620 12750
rect 53564 12686 53566 12738
rect 53618 12686 53620 12738
rect 53564 12404 53620 12686
rect 53620 12348 53956 12404
rect 53564 12338 53620 12348
rect 53900 12178 53956 12348
rect 53900 12126 53902 12178
rect 53954 12126 53956 12178
rect 53900 12114 53956 12126
rect 53788 12068 53844 12078
rect 53340 12012 53732 12068
rect 53228 11396 53284 12012
rect 53676 11506 53732 12012
rect 53788 11974 53844 12012
rect 54572 11956 54628 12910
rect 53676 11454 53678 11506
rect 53730 11454 53732 11506
rect 53676 11442 53732 11454
rect 53900 11900 54628 11956
rect 54684 12962 54852 12964
rect 54684 12910 54798 12962
rect 54850 12910 54852 12962
rect 54684 12908 54852 12910
rect 54684 11956 54740 12908
rect 54796 12898 54852 12908
rect 54908 12628 54964 14028
rect 55020 13746 55076 14140
rect 55580 13972 55636 13982
rect 55804 13972 55860 14252
rect 56364 14242 56420 14252
rect 56476 14308 56532 14366
rect 56476 14242 56532 14252
rect 55580 13970 55860 13972
rect 55580 13918 55582 13970
rect 55634 13918 55860 13970
rect 55580 13916 55860 13918
rect 55580 13906 55636 13916
rect 55356 13860 55412 13870
rect 55356 13766 55412 13804
rect 55020 13694 55022 13746
rect 55074 13694 55076 13746
rect 55020 13076 55076 13694
rect 55244 13746 55300 13758
rect 55244 13694 55246 13746
rect 55298 13694 55300 13746
rect 55132 13524 55188 13534
rect 55244 13524 55300 13694
rect 55188 13468 55300 13524
rect 55132 13458 55188 13468
rect 55468 13076 55524 13086
rect 55020 13074 55524 13076
rect 55020 13022 55470 13074
rect 55522 13022 55524 13074
rect 55020 13020 55524 13022
rect 55468 13010 55524 13020
rect 54796 12572 55076 12628
rect 54796 12290 54852 12572
rect 54796 12238 54798 12290
rect 54850 12238 54852 12290
rect 54796 12226 54852 12238
rect 54908 12292 54964 12302
rect 54908 12198 54964 12236
rect 54908 11956 54964 11966
rect 54684 11954 54964 11956
rect 54684 11902 54910 11954
rect 54962 11902 54964 11954
rect 54684 11900 54964 11902
rect 53228 11394 53396 11396
rect 53228 11342 53230 11394
rect 53282 11342 53396 11394
rect 53228 11340 53396 11342
rect 53228 11330 53284 11340
rect 52556 9828 52612 9838
rect 51548 9772 52052 9828
rect 51996 9714 52052 9772
rect 51996 9662 51998 9714
rect 52050 9662 52052 9714
rect 51660 9604 51716 9614
rect 51100 7634 51156 7644
rect 51212 9602 51716 9604
rect 51212 9550 51662 9602
rect 51714 9550 51716 9602
rect 51212 9548 51716 9550
rect 51212 9042 51268 9548
rect 51660 9538 51716 9548
rect 51884 9602 51940 9614
rect 51884 9550 51886 9602
rect 51938 9550 51940 9602
rect 51884 9268 51940 9550
rect 51884 9202 51940 9212
rect 51212 8990 51214 9042
rect 51266 8990 51268 9042
rect 51212 7586 51268 8990
rect 51436 9042 51492 9054
rect 51436 8990 51438 9042
rect 51490 8990 51492 9042
rect 51436 8372 51492 8990
rect 51548 9044 51604 9054
rect 51548 8950 51604 8988
rect 51772 9042 51828 9054
rect 51772 8990 51774 9042
rect 51826 8990 51828 9042
rect 51436 8306 51492 8316
rect 51772 8260 51828 8990
rect 51772 8194 51828 8204
rect 51212 7534 51214 7586
rect 51266 7534 51268 7586
rect 51212 7522 51268 7534
rect 51436 8146 51492 8158
rect 51436 8094 51438 8146
rect 51490 8094 51492 8146
rect 51436 7476 51492 8094
rect 51436 7410 51492 7420
rect 50988 7310 50990 7362
rect 51042 7310 51044 7362
rect 50988 7298 51044 7310
rect 50764 6804 50820 6814
rect 50876 6804 50932 6860
rect 50764 6802 50932 6804
rect 50764 6750 50766 6802
rect 50818 6750 50932 6802
rect 50764 6748 50932 6750
rect 50764 6738 50820 6748
rect 50652 6638 50654 6690
rect 50706 6638 50708 6690
rect 50652 6468 50708 6638
rect 51436 6692 51492 6702
rect 51436 6580 51492 6636
rect 51436 6524 51828 6580
rect 50652 6412 51716 6468
rect 50540 6402 50596 6412
rect 50556 6300 50820 6310
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50556 6234 50820 6244
rect 51660 6130 51716 6412
rect 51660 6078 51662 6130
rect 51714 6078 51716 6130
rect 51660 6066 51716 6078
rect 51772 6132 51828 6524
rect 51884 6132 51940 6142
rect 51772 6130 51940 6132
rect 51772 6078 51886 6130
rect 51938 6078 51940 6130
rect 51772 6076 51940 6078
rect 51884 6066 51940 6076
rect 51996 6020 52052 9662
rect 52108 9156 52164 9194
rect 52108 9090 52164 9100
rect 52556 9042 52612 9772
rect 52892 9266 52948 10668
rect 53228 10836 53284 10846
rect 53228 9940 53284 10780
rect 53340 10834 53396 11340
rect 53340 10782 53342 10834
rect 53394 10782 53396 10834
rect 53340 10770 53396 10782
rect 53900 10834 53956 11900
rect 54908 11890 54964 11900
rect 53900 10782 53902 10834
rect 53954 10782 53956 10834
rect 53900 10770 53956 10782
rect 54012 11282 54068 11294
rect 54012 11230 54014 11282
rect 54066 11230 54068 11282
rect 54012 10836 54068 11230
rect 54124 11170 54180 11182
rect 54124 11118 54126 11170
rect 54178 11118 54180 11170
rect 54124 10836 54180 11118
rect 54236 10836 54292 10846
rect 54124 10834 54292 10836
rect 54124 10782 54238 10834
rect 54290 10782 54292 10834
rect 54124 10780 54292 10782
rect 54012 10770 54068 10780
rect 54236 10770 54292 10780
rect 55020 10834 55076 12572
rect 55020 10782 55022 10834
rect 55074 10782 55076 10834
rect 55020 10770 55076 10782
rect 53788 10724 53844 10734
rect 53788 10630 53844 10668
rect 54012 10610 54068 10622
rect 54012 10558 54014 10610
rect 54066 10558 54068 10610
rect 53452 10388 53508 10398
rect 53452 10294 53508 10332
rect 54012 10388 54068 10558
rect 54012 10052 54068 10332
rect 54684 10610 54740 10622
rect 54684 10558 54686 10610
rect 54738 10558 54740 10610
rect 54460 10052 54516 10062
rect 54012 10050 54516 10052
rect 54012 9998 54462 10050
rect 54514 9998 54516 10050
rect 54012 9996 54516 9998
rect 54460 9986 54516 9996
rect 53452 9940 53508 9950
rect 53228 9938 53508 9940
rect 53228 9886 53454 9938
rect 53506 9886 53508 9938
rect 53228 9884 53508 9886
rect 53452 9874 53508 9884
rect 53676 9940 53732 9950
rect 52892 9214 52894 9266
rect 52946 9214 52948 9266
rect 52892 9202 52948 9214
rect 53116 9828 53172 9838
rect 52556 8990 52558 9042
rect 52610 8990 52612 9042
rect 52556 8708 52612 8990
rect 52892 9044 52948 9054
rect 52892 8950 52948 8988
rect 52556 8642 52612 8652
rect 52556 8372 52612 8382
rect 52556 8278 52612 8316
rect 53004 8260 53060 8270
rect 52780 8258 53060 8260
rect 52780 8206 53006 8258
rect 53058 8206 53060 8258
rect 52780 8204 53060 8206
rect 52444 7588 52500 7598
rect 52444 7476 52500 7532
rect 52780 7476 52836 8204
rect 53004 8148 53060 8204
rect 53004 8082 53060 8092
rect 52444 7474 52836 7476
rect 52444 7422 52446 7474
rect 52498 7422 52836 7474
rect 52444 7420 52836 7422
rect 52444 7410 52500 7420
rect 52780 6914 52836 7420
rect 52780 6862 52782 6914
rect 52834 6862 52836 6914
rect 52780 6850 52836 6862
rect 52892 8036 52948 8046
rect 52892 6914 52948 7980
rect 52892 6862 52894 6914
rect 52946 6862 52948 6914
rect 52892 6850 52948 6862
rect 53004 6916 53060 6926
rect 53116 6916 53172 9772
rect 53676 9826 53732 9884
rect 54684 9940 54740 10558
rect 54684 9874 54740 9884
rect 53676 9774 53678 9826
rect 53730 9774 53732 9826
rect 53676 9762 53732 9774
rect 53900 9826 53956 9838
rect 53900 9774 53902 9826
rect 53954 9774 53956 9826
rect 53228 9714 53284 9726
rect 53228 9662 53230 9714
rect 53282 9662 53284 9714
rect 53228 9268 53284 9662
rect 53228 9202 53284 9212
rect 53900 9268 53956 9774
rect 54124 9828 54180 9838
rect 54124 9734 54180 9772
rect 53900 9202 53956 9212
rect 53340 8708 53396 8718
rect 53228 8258 53284 8270
rect 53228 8206 53230 8258
rect 53282 8206 53284 8258
rect 53228 8036 53284 8206
rect 53228 7970 53284 7980
rect 53340 7698 53396 8652
rect 53340 7646 53342 7698
rect 53394 7646 53396 7698
rect 53340 7634 53396 7646
rect 53452 8372 53508 8382
rect 53452 8258 53508 8316
rect 54012 8372 54068 8382
rect 53452 8206 53454 8258
rect 53506 8206 53508 8258
rect 53228 6916 53284 6926
rect 53116 6914 53284 6916
rect 53116 6862 53230 6914
rect 53282 6862 53284 6914
rect 53116 6860 53284 6862
rect 53004 6804 53060 6860
rect 53228 6850 53284 6860
rect 53452 6916 53508 8206
rect 53900 8260 53956 8270
rect 53900 8166 53956 8204
rect 54012 8258 54068 8316
rect 54012 8206 54014 8258
rect 54066 8206 54068 8258
rect 54012 8194 54068 8206
rect 54236 8148 54292 8158
rect 54236 8054 54292 8092
rect 53788 8036 53844 8046
rect 53788 7942 53844 7980
rect 53452 6850 53508 6860
rect 53004 6748 53172 6804
rect 53116 6690 53172 6748
rect 53116 6638 53118 6690
rect 53170 6638 53172 6690
rect 53116 6626 53172 6638
rect 52220 6132 52276 6142
rect 52108 6020 52164 6030
rect 51996 6018 52164 6020
rect 51996 5966 52110 6018
rect 52162 5966 52164 6018
rect 51996 5964 52164 5966
rect 50428 5854 50430 5906
rect 50482 5854 50484 5906
rect 50428 5842 50484 5854
rect 51324 5908 51380 5918
rect 51324 5814 51380 5852
rect 50316 5684 50372 5694
rect 50316 5010 50372 5628
rect 52108 5684 52164 5964
rect 52220 6018 52276 6076
rect 52668 6132 52724 6142
rect 52668 6038 52724 6076
rect 52220 5966 52222 6018
rect 52274 5966 52276 6018
rect 52220 5954 52276 5966
rect 52108 5618 52164 5628
rect 50316 4958 50318 5010
rect 50370 4958 50372 5010
rect 50316 4946 50372 4958
rect 50556 4732 50820 4742
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50556 4666 50820 4676
rect 50316 3444 50372 3454
rect 50204 3442 50372 3444
rect 50204 3390 50318 3442
rect 50370 3390 50372 3442
rect 50204 3388 50372 3390
rect 50316 3378 50372 3388
rect 50556 3164 50820 3174
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50556 3098 50820 3108
rect 0 0 112 800
rect 672 0 784 800
rect 1344 0 1456 800
rect 2016 0 2128 800
rect 2688 0 2800 800
rect 3360 0 3472 800
rect 4032 0 4144 800
rect 4704 0 4816 800
rect 5376 0 5488 800
rect 6048 0 6160 800
rect 6720 0 6832 800
rect 7392 0 7504 800
rect 8064 0 8176 800
rect 8736 0 8848 800
rect 9408 0 9520 800
rect 10080 0 10192 800
rect 19488 0 19600 800
rect 22176 0 22288 800
rect 24864 0 24976 800
rect 26880 0 26992 800
rect 28224 0 28336 800
rect 28896 0 29008 800
rect 30240 0 30352 800
rect 30912 0 31024 800
rect 31584 0 31696 800
rect 32256 0 32368 800
rect 32928 0 33040 800
rect 33600 0 33712 800
rect 34272 0 34384 800
rect 34944 0 35056 800
rect 35616 0 35728 800
rect 36288 0 36400 800
rect 36960 0 37072 800
rect 37632 0 37744 800
rect 38304 0 38416 800
rect 38976 0 39088 800
rect 39648 0 39760 800
rect 43008 0 43120 800
rect 47040 0 47152 800
rect 49728 0 49840 800
<< via2 >>
rect 19836 56474 19892 56476
rect 19836 56422 19838 56474
rect 19838 56422 19890 56474
rect 19890 56422 19892 56474
rect 19836 56420 19892 56422
rect 19940 56474 19996 56476
rect 19940 56422 19942 56474
rect 19942 56422 19994 56474
rect 19994 56422 19996 56474
rect 19940 56420 19996 56422
rect 20044 56474 20100 56476
rect 20044 56422 20046 56474
rect 20046 56422 20098 56474
rect 20098 56422 20100 56474
rect 20044 56420 20100 56422
rect 4476 55690 4532 55692
rect 4476 55638 4478 55690
rect 4478 55638 4530 55690
rect 4530 55638 4532 55690
rect 4476 55636 4532 55638
rect 4580 55690 4636 55692
rect 4580 55638 4582 55690
rect 4582 55638 4634 55690
rect 4634 55638 4636 55690
rect 4580 55636 4636 55638
rect 4684 55690 4740 55692
rect 4684 55638 4686 55690
rect 4686 55638 4738 55690
rect 4738 55638 4740 55690
rect 4684 55636 4740 55638
rect 19836 54906 19892 54908
rect 19836 54854 19838 54906
rect 19838 54854 19890 54906
rect 19890 54854 19892 54906
rect 19836 54852 19892 54854
rect 19940 54906 19996 54908
rect 19940 54854 19942 54906
rect 19942 54854 19994 54906
rect 19994 54854 19996 54906
rect 19940 54852 19996 54854
rect 20044 54906 20100 54908
rect 20044 54854 20046 54906
rect 20046 54854 20098 54906
rect 20098 54854 20100 54906
rect 20044 54852 20100 54854
rect 4476 54122 4532 54124
rect 4476 54070 4478 54122
rect 4478 54070 4530 54122
rect 4530 54070 4532 54122
rect 4476 54068 4532 54070
rect 4580 54122 4636 54124
rect 4580 54070 4582 54122
rect 4582 54070 4634 54122
rect 4634 54070 4636 54122
rect 4580 54068 4636 54070
rect 4684 54122 4740 54124
rect 4684 54070 4686 54122
rect 4686 54070 4738 54122
rect 4738 54070 4740 54122
rect 4684 54068 4740 54070
rect 4476 52554 4532 52556
rect 4476 52502 4478 52554
rect 4478 52502 4530 52554
rect 4530 52502 4532 52554
rect 4476 52500 4532 52502
rect 4580 52554 4636 52556
rect 4580 52502 4582 52554
rect 4582 52502 4634 52554
rect 4634 52502 4636 52554
rect 4580 52500 4636 52502
rect 4684 52554 4740 52556
rect 4684 52502 4686 52554
rect 4686 52502 4738 52554
rect 4738 52502 4740 52554
rect 4684 52500 4740 52502
rect 1708 50482 1764 50484
rect 1708 50430 1710 50482
rect 1710 50430 1762 50482
rect 1762 50430 1764 50482
rect 1708 50428 1764 50430
rect 4476 50986 4532 50988
rect 4476 50934 4478 50986
rect 4478 50934 4530 50986
rect 4530 50934 4532 50986
rect 4476 50932 4532 50934
rect 4580 50986 4636 50988
rect 4580 50934 4582 50986
rect 4582 50934 4634 50986
rect 4634 50934 4636 50986
rect 4580 50932 4636 50934
rect 4684 50986 4740 50988
rect 4684 50934 4686 50986
rect 4686 50934 4738 50986
rect 4738 50934 4740 50986
rect 4684 50932 4740 50934
rect 5964 50988 6020 51044
rect 2940 50482 2996 50484
rect 2940 50430 2942 50482
rect 2942 50430 2994 50482
rect 2994 50430 2996 50482
rect 2940 50428 2996 50430
rect 1708 49308 1764 49364
rect 1484 48748 1540 48804
rect 1372 44380 1428 44436
rect 1260 39340 1316 39396
rect 1372 34748 1428 34804
rect 1708 48524 1764 48580
rect 2044 50370 2100 50372
rect 2044 50318 2046 50370
rect 2046 50318 2098 50370
rect 2098 50318 2100 50370
rect 2044 50316 2100 50318
rect 2044 48802 2100 48804
rect 2044 48750 2046 48802
rect 2046 48750 2098 48802
rect 2098 48750 2100 48802
rect 2044 48748 2100 48750
rect 2828 49698 2884 49700
rect 2828 49646 2830 49698
rect 2830 49646 2882 49698
rect 2882 49646 2884 49698
rect 2828 49644 2884 49646
rect 2492 49196 2548 49252
rect 2380 49026 2436 49028
rect 2380 48974 2382 49026
rect 2382 48974 2434 49026
rect 2434 48974 2436 49026
rect 2380 48972 2436 48974
rect 2156 48354 2212 48356
rect 2156 48302 2158 48354
rect 2158 48302 2210 48354
rect 2210 48302 2212 48354
rect 2156 48300 2212 48302
rect 1820 46732 1876 46788
rect 2044 47234 2100 47236
rect 2044 47182 2046 47234
rect 2046 47182 2098 47234
rect 2098 47182 2100 47234
rect 2044 47180 2100 47182
rect 2716 48412 2772 48468
rect 2604 48188 2660 48244
rect 2268 46732 2324 46788
rect 2492 47458 2548 47460
rect 2492 47406 2494 47458
rect 2494 47406 2546 47458
rect 2546 47406 2548 47458
rect 2492 47404 2548 47406
rect 1596 44268 1652 44324
rect 1708 44098 1764 44100
rect 1708 44046 1710 44098
rect 1710 44046 1762 44098
rect 1762 44046 1764 44098
rect 1708 44044 1764 44046
rect 1708 41970 1764 41972
rect 1708 41918 1710 41970
rect 1710 41918 1762 41970
rect 1762 41918 1764 41970
rect 1708 41916 1764 41918
rect 2156 45276 2212 45332
rect 1932 44492 1988 44548
rect 2156 44268 2212 44324
rect 2044 43708 2100 43764
rect 2044 42812 2100 42868
rect 1932 42364 1988 42420
rect 1708 41020 1764 41076
rect 1932 40348 1988 40404
rect 1932 39676 1988 39732
rect 1708 38556 1764 38612
rect 2044 39564 2100 39620
rect 2044 39394 2100 39396
rect 2044 39342 2046 39394
rect 2046 39342 2098 39394
rect 2098 39342 2100 39394
rect 2044 39340 2100 39342
rect 3388 49084 3444 49140
rect 3276 49026 3332 49028
rect 3276 48974 3278 49026
rect 3278 48974 3330 49026
rect 3330 48974 3332 49026
rect 3276 48972 3332 48974
rect 3052 48188 3108 48244
rect 3052 47404 3108 47460
rect 3612 48636 3668 48692
rect 4844 50316 4900 50372
rect 3948 49308 4004 49364
rect 3948 49084 4004 49140
rect 4476 49418 4532 49420
rect 4476 49366 4478 49418
rect 4478 49366 4530 49418
rect 4530 49366 4532 49418
rect 4476 49364 4532 49366
rect 4580 49418 4636 49420
rect 4580 49366 4582 49418
rect 4582 49366 4634 49418
rect 4634 49366 4636 49418
rect 4580 49364 4636 49366
rect 4684 49418 4740 49420
rect 4684 49366 4686 49418
rect 4686 49366 4738 49418
rect 4738 49366 4740 49418
rect 4684 49364 4740 49366
rect 5628 50370 5684 50372
rect 5628 50318 5630 50370
rect 5630 50318 5682 50370
rect 5682 50318 5684 50370
rect 5628 50316 5684 50318
rect 4844 49084 4900 49140
rect 4172 48972 4228 49028
rect 4732 48972 4788 49028
rect 3836 48914 3892 48916
rect 3836 48862 3838 48914
rect 3838 48862 3890 48914
rect 3890 48862 3892 48914
rect 3836 48860 3892 48862
rect 3388 48412 3444 48468
rect 3948 48636 4004 48692
rect 3276 48300 3332 48356
rect 3388 48076 3444 48132
rect 3276 47292 3332 47348
rect 3052 47068 3108 47124
rect 3052 46674 3108 46676
rect 3052 46622 3054 46674
rect 3054 46622 3106 46674
rect 3106 46622 3108 46674
rect 3052 46620 3108 46622
rect 3164 45890 3220 45892
rect 3164 45838 3166 45890
rect 3166 45838 3218 45890
rect 3218 45838 3220 45890
rect 3164 45836 3220 45838
rect 2380 44434 2436 44436
rect 2380 44382 2382 44434
rect 2382 44382 2434 44434
rect 2434 44382 2436 44434
rect 2380 44380 2436 44382
rect 2716 44604 2772 44660
rect 3052 44994 3108 44996
rect 3052 44942 3054 44994
rect 3054 44942 3106 44994
rect 3106 44942 3108 44994
rect 3052 44940 3108 44942
rect 2716 44380 2772 44436
rect 3500 45052 3556 45108
rect 3388 44828 3444 44884
rect 2940 44322 2996 44324
rect 2940 44270 2942 44322
rect 2942 44270 2994 44322
rect 2994 44270 2996 44322
rect 2940 44268 2996 44270
rect 2828 44156 2884 44212
rect 3388 44098 3444 44100
rect 3388 44046 3390 44098
rect 3390 44046 3442 44098
rect 3442 44046 3444 44098
rect 3388 44044 3444 44046
rect 2716 43596 2772 43652
rect 4508 48524 4564 48580
rect 6300 48972 6356 49028
rect 4956 48860 5012 48916
rect 6076 48860 6132 48916
rect 7196 50594 7252 50596
rect 7196 50542 7198 50594
rect 7198 50542 7250 50594
rect 7250 50542 7252 50594
rect 7196 50540 7252 50542
rect 6860 49698 6916 49700
rect 6860 49646 6862 49698
rect 6862 49646 6914 49698
rect 6914 49646 6916 49698
rect 6860 49644 6916 49646
rect 6972 49138 7028 49140
rect 6972 49086 6974 49138
rect 6974 49086 7026 49138
rect 7026 49086 7028 49138
rect 6972 49084 7028 49086
rect 6636 48972 6692 49028
rect 4060 48130 4116 48132
rect 4060 48078 4062 48130
rect 4062 48078 4114 48130
rect 4114 48078 4116 48130
rect 4060 48076 4116 48078
rect 4508 48076 4564 48132
rect 3724 47570 3780 47572
rect 3724 47518 3726 47570
rect 3726 47518 3778 47570
rect 3778 47518 3780 47570
rect 3724 47516 3780 47518
rect 4476 47850 4532 47852
rect 4476 47798 4478 47850
rect 4478 47798 4530 47850
rect 4530 47798 4532 47850
rect 4476 47796 4532 47798
rect 4580 47850 4636 47852
rect 4580 47798 4582 47850
rect 4582 47798 4634 47850
rect 4634 47798 4636 47850
rect 4580 47796 4636 47798
rect 4684 47850 4740 47852
rect 4684 47798 4686 47850
rect 4686 47798 4738 47850
rect 4738 47798 4740 47850
rect 4684 47796 4740 47798
rect 4172 47516 4228 47572
rect 3612 43820 3668 43876
rect 2940 43426 2996 43428
rect 2940 43374 2942 43426
rect 2942 43374 2994 43426
rect 2994 43374 2996 43426
rect 2940 43372 2996 43374
rect 2716 42812 2772 42868
rect 2156 38892 2212 38948
rect 2156 38556 2212 38612
rect 1932 37042 1988 37044
rect 1932 36990 1934 37042
rect 1934 36990 1986 37042
rect 1986 36990 1988 37042
rect 1932 36988 1988 36990
rect 1596 36428 1652 36484
rect 1820 36258 1876 36260
rect 1820 36206 1822 36258
rect 1822 36206 1874 36258
rect 1874 36206 1876 36258
rect 1820 36204 1876 36206
rect 2268 37996 2324 38052
rect 3948 46674 4004 46676
rect 3948 46622 3950 46674
rect 3950 46622 4002 46674
rect 4002 46622 4004 46674
rect 3948 46620 4004 46622
rect 5740 48802 5796 48804
rect 5740 48750 5742 48802
rect 5742 48750 5794 48802
rect 5794 48750 5796 48802
rect 5740 48748 5796 48750
rect 6636 48748 6692 48804
rect 5628 48076 5684 48132
rect 5068 47458 5124 47460
rect 5068 47406 5070 47458
rect 5070 47406 5122 47458
rect 5122 47406 5124 47458
rect 5068 47404 5124 47406
rect 5964 48130 6020 48132
rect 5964 48078 5966 48130
rect 5966 48078 6018 48130
rect 6018 48078 6020 48130
rect 5964 48076 6020 48078
rect 6300 47346 6356 47348
rect 6300 47294 6302 47346
rect 6302 47294 6354 47346
rect 6354 47294 6356 47346
rect 6300 47292 6356 47294
rect 5404 47068 5460 47124
rect 3724 45836 3780 45892
rect 3052 43314 3108 43316
rect 3052 43262 3054 43314
rect 3054 43262 3106 43314
rect 3106 43262 3108 43314
rect 3052 43260 3108 43262
rect 2716 38892 2772 38948
rect 2380 37548 2436 37604
rect 2380 37324 2436 37380
rect 2156 36540 2212 36596
rect 2156 36092 2212 36148
rect 2268 36316 2324 36372
rect 1708 35868 1764 35924
rect 1708 35308 1764 35364
rect 1484 34412 1540 34468
rect 1708 34076 1764 34132
rect 1708 33122 1764 33124
rect 1708 33070 1710 33122
rect 1710 33070 1762 33122
rect 1762 33070 1764 33122
rect 1708 33068 1764 33070
rect 1932 35196 1988 35252
rect 2044 35084 2100 35140
rect 2044 33964 2100 34020
rect 1932 33906 1988 33908
rect 1932 33854 1934 33906
rect 1934 33854 1986 33906
rect 1986 33854 1988 33906
rect 1932 33852 1988 33854
rect 2268 35308 2324 35364
rect 1820 32956 1876 33012
rect 2604 38444 2660 38500
rect 2716 37996 2772 38052
rect 2716 37548 2772 37604
rect 2828 36988 2884 37044
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 4172 46002 4228 46004
rect 4172 45950 4174 46002
rect 4174 45950 4226 46002
rect 4226 45950 4228 46002
rect 4172 45948 4228 45950
rect 4620 45612 4676 45668
rect 4732 45276 4788 45332
rect 3948 44828 4004 44884
rect 5068 45052 5124 45108
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 4620 44322 4676 44324
rect 4620 44270 4622 44322
rect 4622 44270 4674 44322
rect 4674 44270 4676 44322
rect 4620 44268 4676 44270
rect 4620 43650 4676 43652
rect 4620 43598 4622 43650
rect 4622 43598 4674 43650
rect 4674 43598 4676 43650
rect 4620 43596 4676 43598
rect 4060 43538 4116 43540
rect 4060 43486 4062 43538
rect 4062 43486 4114 43538
rect 4114 43486 4116 43538
rect 4060 43484 4116 43486
rect 4844 43484 4900 43540
rect 5068 44380 5124 44436
rect 3836 41692 3892 41748
rect 3948 43372 4004 43428
rect 8316 51490 8372 51492
rect 8316 51438 8318 51490
rect 8318 51438 8370 51490
rect 8370 51438 8372 51490
rect 8316 51436 8372 51438
rect 7644 49868 7700 49924
rect 7756 49644 7812 49700
rect 8204 49868 8260 49924
rect 10108 50988 10164 51044
rect 8764 50706 8820 50708
rect 8764 50654 8766 50706
rect 8766 50654 8818 50706
rect 8818 50654 8820 50706
rect 8764 50652 8820 50654
rect 9212 50594 9268 50596
rect 9212 50542 9214 50594
rect 9214 50542 9266 50594
rect 9266 50542 9268 50594
rect 9212 50540 9268 50542
rect 8316 48860 8372 48916
rect 5628 46060 5684 46116
rect 6300 46060 6356 46116
rect 6412 45778 6468 45780
rect 6412 45726 6414 45778
rect 6414 45726 6466 45778
rect 6466 45726 6468 45778
rect 6412 45724 6468 45726
rect 6860 46674 6916 46676
rect 6860 46622 6862 46674
rect 6862 46622 6914 46674
rect 6914 46622 6916 46674
rect 6860 46620 6916 46622
rect 5852 45052 5908 45108
rect 5628 44940 5684 44996
rect 5964 44828 6020 44884
rect 6412 45276 6468 45332
rect 6300 44210 6356 44212
rect 6300 44158 6302 44210
rect 6302 44158 6354 44210
rect 6354 44158 6356 44210
rect 6300 44156 6356 44158
rect 5852 44098 5908 44100
rect 5852 44046 5854 44098
rect 5854 44046 5906 44098
rect 5906 44046 5908 44098
rect 5852 44044 5908 44046
rect 7196 45106 7252 45108
rect 7196 45054 7198 45106
rect 7198 45054 7250 45106
rect 7250 45054 7252 45106
rect 7196 45052 7252 45054
rect 6412 44044 6468 44100
rect 4284 43260 4340 43316
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 5516 43148 5572 43204
rect 4684 43092 4740 43094
rect 5740 43596 5796 43652
rect 5852 43426 5908 43428
rect 5852 43374 5854 43426
rect 5854 43374 5906 43426
rect 5906 43374 5908 43426
rect 5852 43372 5908 43374
rect 4620 42812 4676 42868
rect 3612 40348 3668 40404
rect 3724 41020 3780 41076
rect 3388 38332 3444 38388
rect 4620 41858 4676 41860
rect 4620 41806 4622 41858
rect 4622 41806 4674 41858
rect 4674 41806 4676 41858
rect 4620 41804 4676 41806
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 4284 41356 4340 41412
rect 4732 41020 4788 41076
rect 4284 40796 4340 40852
rect 4172 40684 4228 40740
rect 3948 40124 4004 40180
rect 4060 40348 4116 40404
rect 3724 37660 3780 37716
rect 3724 37324 3780 37380
rect 2716 36316 2772 36372
rect 2940 36204 2996 36260
rect 2492 36092 2548 36148
rect 2716 36092 2772 36148
rect 2604 35922 2660 35924
rect 2604 35870 2606 35922
rect 2606 35870 2658 35922
rect 2658 35870 2660 35922
rect 2604 35868 2660 35870
rect 2604 35308 2660 35364
rect 2604 35084 2660 35140
rect 3836 36092 3892 36148
rect 4956 40962 5012 40964
rect 4956 40910 4958 40962
rect 4958 40910 5010 40962
rect 5010 40910 5012 40962
rect 4956 40908 5012 40910
rect 5404 41970 5460 41972
rect 5404 41918 5406 41970
rect 5406 41918 5458 41970
rect 5458 41918 5460 41970
rect 5404 41916 5460 41918
rect 4620 40290 4676 40292
rect 4620 40238 4622 40290
rect 4622 40238 4674 40290
rect 4674 40238 4676 40290
rect 4620 40236 4676 40238
rect 4284 40124 4340 40180
rect 4732 40124 4788 40180
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 5068 40460 5124 40516
rect 4620 38834 4676 38836
rect 4620 38782 4622 38834
rect 4622 38782 4674 38834
rect 4674 38782 4676 38834
rect 4620 38780 4676 38782
rect 5180 38780 5236 38836
rect 3276 35420 3332 35476
rect 3500 35196 3556 35252
rect 1260 31724 1316 31780
rect 2492 33068 2548 33124
rect 2716 33292 2772 33348
rect 2492 32674 2548 32676
rect 2492 32622 2494 32674
rect 2494 32622 2546 32674
rect 2546 32622 2548 32674
rect 2492 32620 2548 32622
rect 2380 31836 2436 31892
rect 3276 32786 3332 32788
rect 3276 32734 3278 32786
rect 3278 32734 3330 32786
rect 3330 32734 3332 32786
rect 3276 32732 3332 32734
rect 2716 31276 2772 31332
rect 1932 30940 1988 30996
rect 3052 31500 3108 31556
rect 4060 38444 4116 38500
rect 4172 38220 4228 38276
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 4956 38444 5012 38500
rect 4284 37996 4340 38052
rect 4732 38050 4788 38052
rect 4732 37998 4734 38050
rect 4734 37998 4786 38050
rect 4786 37998 4788 38050
rect 4732 37996 4788 37998
rect 4844 37548 4900 37604
rect 4732 37378 4788 37380
rect 4732 37326 4734 37378
rect 4734 37326 4786 37378
rect 4786 37326 4788 37378
rect 4732 37324 4788 37326
rect 4396 36988 4452 37044
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4844 36876 4900 36932
rect 4684 36820 4740 36822
rect 4620 36370 4676 36372
rect 4620 36318 4622 36370
rect 4622 36318 4674 36370
rect 4674 36318 4676 36370
rect 4620 36316 4676 36318
rect 4284 36092 4340 36148
rect 3836 34972 3892 35028
rect 4060 35196 4116 35252
rect 3724 34188 3780 34244
rect 3500 33852 3556 33908
rect 4396 35474 4452 35476
rect 4396 35422 4398 35474
rect 4398 35422 4450 35474
rect 4450 35422 4452 35474
rect 4396 35420 4452 35422
rect 4284 35308 4340 35364
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4508 34972 4564 35028
rect 4060 34636 4116 34692
rect 5516 39004 5572 39060
rect 6300 41916 6356 41972
rect 6188 41804 6244 41860
rect 6188 41244 6244 41300
rect 6300 40514 6356 40516
rect 6300 40462 6302 40514
rect 6302 40462 6354 40514
rect 6354 40462 6356 40514
rect 6300 40460 6356 40462
rect 6076 40348 6132 40404
rect 6636 44828 6692 44884
rect 6860 44322 6916 44324
rect 6860 44270 6862 44322
rect 6862 44270 6914 44322
rect 6914 44270 6916 44322
rect 6860 44268 6916 44270
rect 7196 44044 7252 44100
rect 7532 48076 7588 48132
rect 7532 47516 7588 47572
rect 9212 48860 9268 48916
rect 8988 48188 9044 48244
rect 9100 48300 9156 48356
rect 7644 46620 7700 46676
rect 7980 47570 8036 47572
rect 7980 47518 7982 47570
rect 7982 47518 8034 47570
rect 8034 47518 8036 47570
rect 7980 47516 8036 47518
rect 8316 47570 8372 47572
rect 8316 47518 8318 47570
rect 8318 47518 8370 47570
rect 8370 47518 8372 47570
rect 8316 47516 8372 47518
rect 8876 47292 8932 47348
rect 8540 46060 8596 46116
rect 8652 45724 8708 45780
rect 7644 44434 7700 44436
rect 7644 44382 7646 44434
rect 7646 44382 7698 44434
rect 7698 44382 7700 44434
rect 7644 44380 7700 44382
rect 7532 44268 7588 44324
rect 6748 43484 6804 43540
rect 6636 41916 6692 41972
rect 6860 42028 6916 42084
rect 6636 40572 6692 40628
rect 6748 41132 6804 41188
rect 5852 40012 5908 40068
rect 5964 39564 6020 39620
rect 5404 38220 5460 38276
rect 5740 38108 5796 38164
rect 5740 37548 5796 37604
rect 5740 37266 5796 37268
rect 5740 37214 5742 37266
rect 5742 37214 5794 37266
rect 5794 37214 5796 37266
rect 5740 37212 5796 37214
rect 5516 36988 5572 37044
rect 5292 35922 5348 35924
rect 5292 35870 5294 35922
rect 5294 35870 5346 35922
rect 5346 35870 5348 35922
rect 5292 35868 5348 35870
rect 6860 40684 6916 40740
rect 6076 38668 6132 38724
rect 6748 37996 6804 38052
rect 6300 37100 6356 37156
rect 6524 36876 6580 36932
rect 6636 36652 6692 36708
rect 6860 37100 6916 37156
rect 5964 35868 6020 35924
rect 5404 35756 5460 35812
rect 5628 35698 5684 35700
rect 5628 35646 5630 35698
rect 5630 35646 5682 35698
rect 5682 35646 5684 35698
rect 5628 35644 5684 35646
rect 4956 35532 5012 35588
rect 4956 34300 5012 34356
rect 6076 35308 6132 35364
rect 6524 36204 6580 36260
rect 8428 44156 8484 44212
rect 7308 43484 7364 43540
rect 8092 43260 8148 43316
rect 8316 41916 8372 41972
rect 8652 41692 8708 41748
rect 8092 41580 8148 41636
rect 7196 41298 7252 41300
rect 7196 41246 7198 41298
rect 7198 41246 7250 41298
rect 7250 41246 7252 41298
rect 7196 41244 7252 41246
rect 7196 40626 7252 40628
rect 7196 40574 7198 40626
rect 7198 40574 7250 40626
rect 7250 40574 7252 40626
rect 7196 40572 7252 40574
rect 7420 41186 7476 41188
rect 7420 41134 7422 41186
rect 7422 41134 7474 41186
rect 7474 41134 7476 41186
rect 7420 41132 7476 41134
rect 7420 40626 7476 40628
rect 7420 40574 7422 40626
rect 7422 40574 7474 40626
rect 7474 40574 7476 40626
rect 7420 40572 7476 40574
rect 7532 40402 7588 40404
rect 7532 40350 7534 40402
rect 7534 40350 7586 40402
rect 7586 40350 7588 40402
rect 7532 40348 7588 40350
rect 8540 41074 8596 41076
rect 8540 41022 8542 41074
rect 8542 41022 8594 41074
rect 8594 41022 8596 41074
rect 8540 41020 8596 41022
rect 8988 45164 9044 45220
rect 9884 48354 9940 48356
rect 9884 48302 9886 48354
rect 9886 48302 9938 48354
rect 9938 48302 9940 48354
rect 9884 48300 9940 48302
rect 12460 52892 12516 52948
rect 11004 52386 11060 52388
rect 11004 52334 11006 52386
rect 11006 52334 11058 52386
rect 11058 52334 11060 52386
rect 11004 52332 11060 52334
rect 11116 52108 11172 52164
rect 10332 51436 10388 51492
rect 10780 51378 10836 51380
rect 10780 51326 10782 51378
rect 10782 51326 10834 51378
rect 10834 51326 10836 51378
rect 10780 51324 10836 51326
rect 12460 52332 12516 52388
rect 11788 52162 11844 52164
rect 11788 52110 11790 52162
rect 11790 52110 11842 52162
rect 11842 52110 11844 52162
rect 11788 52108 11844 52110
rect 12348 52162 12404 52164
rect 12348 52110 12350 52162
rect 12350 52110 12402 52162
rect 12402 52110 12404 52162
rect 12348 52108 12404 52110
rect 12236 52050 12292 52052
rect 12236 51998 12238 52050
rect 12238 51998 12290 52050
rect 12290 51998 12292 52050
rect 12236 51996 12292 51998
rect 11228 51324 11284 51380
rect 11676 49868 11732 49924
rect 10556 48802 10612 48804
rect 10556 48750 10558 48802
rect 10558 48750 10610 48802
rect 10610 48750 10612 48802
rect 10556 48748 10612 48750
rect 9772 47516 9828 47572
rect 9548 47346 9604 47348
rect 9548 47294 9550 47346
rect 9550 47294 9602 47346
rect 9602 47294 9604 47346
rect 9548 47292 9604 47294
rect 9212 47180 9268 47236
rect 10332 47292 10388 47348
rect 9660 46060 9716 46116
rect 9772 45666 9828 45668
rect 9772 45614 9774 45666
rect 9774 45614 9826 45666
rect 9826 45614 9828 45666
rect 9772 45612 9828 45614
rect 9772 45330 9828 45332
rect 9772 45278 9774 45330
rect 9774 45278 9826 45330
rect 9826 45278 9828 45330
rect 9772 45276 9828 45278
rect 9212 45052 9268 45108
rect 9660 44994 9716 44996
rect 9660 44942 9662 44994
rect 9662 44942 9714 44994
rect 9714 44942 9716 44994
rect 9660 44940 9716 44942
rect 9996 44882 10052 44884
rect 9996 44830 9998 44882
rect 9998 44830 10050 44882
rect 10050 44830 10052 44882
rect 9996 44828 10052 44830
rect 10220 46620 10276 46676
rect 9548 44322 9604 44324
rect 9548 44270 9550 44322
rect 9550 44270 9602 44322
rect 9602 44270 9604 44322
rect 9548 44268 9604 44270
rect 10444 45388 10500 45444
rect 9436 44210 9492 44212
rect 9436 44158 9438 44210
rect 9438 44158 9490 44210
rect 9490 44158 9492 44210
rect 9436 44156 9492 44158
rect 8988 41356 9044 41412
rect 8316 40402 8372 40404
rect 8316 40350 8318 40402
rect 8318 40350 8370 40402
rect 8370 40350 8372 40402
rect 8316 40348 8372 40350
rect 8092 39506 8148 39508
rect 8092 39454 8094 39506
rect 8094 39454 8146 39506
rect 8146 39454 8148 39506
rect 8092 39452 8148 39454
rect 8316 38946 8372 38948
rect 8316 38894 8318 38946
rect 8318 38894 8370 38946
rect 8370 38894 8372 38946
rect 8316 38892 8372 38894
rect 6972 36092 7028 36148
rect 7196 35868 7252 35924
rect 6524 35532 6580 35588
rect 6860 35420 6916 35476
rect 5068 34860 5124 34916
rect 3836 33852 3892 33908
rect 3948 34076 4004 34132
rect 3724 33516 3780 33572
rect 3612 31612 3668 31668
rect 3500 31500 3556 31556
rect 3276 30882 3332 30884
rect 3276 30830 3278 30882
rect 3278 30830 3330 30882
rect 3330 30830 3332 30882
rect 3276 30828 3332 30830
rect 2268 30604 2324 30660
rect 1708 30268 1764 30324
rect 1596 28812 1652 28868
rect 1260 28140 1316 28196
rect 1484 22764 1540 22820
rect 1484 22316 1540 22372
rect 1484 18396 1540 18452
rect 1372 18172 1428 18228
rect 1932 29202 1988 29204
rect 1932 29150 1934 29202
rect 1934 29150 1986 29202
rect 1986 29150 1988 29202
rect 1932 29148 1988 29150
rect 3388 30604 3444 30660
rect 2492 29596 2548 29652
rect 2828 29708 2884 29764
rect 2716 29372 2772 29428
rect 1932 28252 1988 28308
rect 2044 28588 2100 28644
rect 2716 28642 2772 28644
rect 2716 28590 2718 28642
rect 2718 28590 2770 28642
rect 2770 28590 2772 28642
rect 2716 28588 2772 28590
rect 2940 28364 2996 28420
rect 1820 27858 1876 27860
rect 1820 27806 1822 27858
rect 1822 27806 1874 27858
rect 1874 27806 1876 27858
rect 1820 27804 1876 27806
rect 2380 27580 2436 27636
rect 1708 27074 1764 27076
rect 1708 27022 1710 27074
rect 1710 27022 1762 27074
rect 1762 27022 1764 27074
rect 1708 27020 1764 27022
rect 2044 27132 2100 27188
rect 3388 28588 3444 28644
rect 3052 28252 3108 28308
rect 3724 31052 3780 31108
rect 4732 34130 4788 34132
rect 4732 34078 4734 34130
rect 4734 34078 4786 34130
rect 4786 34078 4788 34130
rect 4732 34076 4788 34078
rect 4284 33852 4340 33908
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 6972 34860 7028 34916
rect 5852 34636 5908 34692
rect 5292 33516 5348 33572
rect 4060 31836 4116 31892
rect 4956 32732 5012 32788
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4732 31948 4788 32004
rect 4284 31612 4340 31668
rect 4620 31778 4676 31780
rect 4620 31726 4622 31778
rect 4622 31726 4674 31778
rect 4674 31726 4676 31778
rect 4620 31724 4676 31726
rect 4172 31388 4228 31444
rect 3948 30604 4004 30660
rect 4956 31836 5012 31892
rect 4956 31164 5012 31220
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 5404 33964 5460 34020
rect 6300 34748 6356 34804
rect 6188 34690 6244 34692
rect 6188 34638 6190 34690
rect 6190 34638 6242 34690
rect 6242 34638 6244 34690
rect 6188 34636 6244 34638
rect 7644 37884 7700 37940
rect 7420 36652 7476 36708
rect 7868 37266 7924 37268
rect 7868 37214 7870 37266
rect 7870 37214 7922 37266
rect 7922 37214 7924 37266
rect 7868 37212 7924 37214
rect 9100 40796 9156 40852
rect 11564 48412 11620 48468
rect 12572 52220 12628 52276
rect 13468 52946 13524 52948
rect 13468 52894 13470 52946
rect 13470 52894 13522 52946
rect 13522 52894 13524 52946
rect 13468 52892 13524 52894
rect 12796 51996 12852 52052
rect 13244 52220 13300 52276
rect 12348 51324 12404 51380
rect 12460 51154 12516 51156
rect 12460 51102 12462 51154
rect 12462 51102 12514 51154
rect 12514 51102 12516 51154
rect 12460 51100 12516 51102
rect 13692 51100 13748 51156
rect 12012 50652 12068 50708
rect 13916 50540 13972 50596
rect 19836 53338 19892 53340
rect 19836 53286 19838 53338
rect 19838 53286 19890 53338
rect 19890 53286 19892 53338
rect 19836 53284 19892 53286
rect 19940 53338 19996 53340
rect 19940 53286 19942 53338
rect 19942 53286 19994 53338
rect 19994 53286 19996 53338
rect 19940 53284 19996 53286
rect 20044 53338 20100 53340
rect 20044 53286 20046 53338
rect 20046 53286 20098 53338
rect 20098 53286 20100 53338
rect 20044 53284 20100 53286
rect 14924 53004 14980 53060
rect 15596 53058 15652 53060
rect 15596 53006 15598 53058
rect 15598 53006 15650 53058
rect 15650 53006 15652 53058
rect 15596 53004 15652 53006
rect 16156 53058 16212 53060
rect 16156 53006 16158 53058
rect 16158 53006 16210 53058
rect 16210 53006 16212 53058
rect 16156 53004 16212 53006
rect 14588 52274 14644 52276
rect 14588 52222 14590 52274
rect 14590 52222 14642 52274
rect 14642 52222 14644 52274
rect 14588 52220 14644 52222
rect 15260 52220 15316 52276
rect 15148 52162 15204 52164
rect 15148 52110 15150 52162
rect 15150 52110 15202 52162
rect 15202 52110 15204 52162
rect 15148 52108 15204 52110
rect 14476 51378 14532 51380
rect 14476 51326 14478 51378
rect 14478 51326 14530 51378
rect 14530 51326 14532 51378
rect 14476 51324 14532 51326
rect 14140 50092 14196 50148
rect 13580 49922 13636 49924
rect 13580 49870 13582 49922
rect 13582 49870 13634 49922
rect 13634 49870 13636 49922
rect 13580 49868 13636 49870
rect 14028 49868 14084 49924
rect 11788 48636 11844 48692
rect 12908 49698 12964 49700
rect 12908 49646 12910 49698
rect 12910 49646 12962 49698
rect 12962 49646 12964 49698
rect 12908 49644 12964 49646
rect 12348 48748 12404 48804
rect 11900 48412 11956 48468
rect 11900 48188 11956 48244
rect 11228 46620 11284 46676
rect 12796 48242 12852 48244
rect 12796 48190 12798 48242
rect 12798 48190 12850 48242
rect 12850 48190 12852 48242
rect 12796 48188 12852 48190
rect 13692 48636 13748 48692
rect 11116 45276 11172 45332
rect 11340 45612 11396 45668
rect 11900 45612 11956 45668
rect 12124 46674 12180 46676
rect 12124 46622 12126 46674
rect 12126 46622 12178 46674
rect 12178 46622 12180 46674
rect 12124 46620 12180 46622
rect 13916 48300 13972 48356
rect 13916 47740 13972 47796
rect 15484 51436 15540 51492
rect 16604 52274 16660 52276
rect 16604 52222 16606 52274
rect 16606 52222 16658 52274
rect 16658 52222 16660 52274
rect 16604 52220 16660 52222
rect 16380 52108 16436 52164
rect 17276 52332 17332 52388
rect 19628 52946 19684 52948
rect 19628 52894 19630 52946
rect 19630 52894 19682 52946
rect 19682 52894 19684 52946
rect 19628 52892 19684 52894
rect 20636 52946 20692 52948
rect 20636 52894 20638 52946
rect 20638 52894 20690 52946
rect 20690 52894 20692 52946
rect 20636 52892 20692 52894
rect 18396 52834 18452 52836
rect 18396 52782 18398 52834
rect 18398 52782 18450 52834
rect 18450 52782 18452 52834
rect 18396 52780 18452 52782
rect 19180 52834 19236 52836
rect 19180 52782 19182 52834
rect 19182 52782 19234 52834
rect 19234 52782 19236 52834
rect 19180 52780 19236 52782
rect 20076 52444 20132 52500
rect 18060 52332 18116 52388
rect 17948 52220 18004 52276
rect 18620 52220 18676 52276
rect 19740 52220 19796 52276
rect 15484 50988 15540 51044
rect 15708 50428 15764 50484
rect 14140 47628 14196 47684
rect 14700 50092 14756 50148
rect 14700 49084 14756 49140
rect 15148 49644 15204 49700
rect 15372 49084 15428 49140
rect 14700 48914 14756 48916
rect 14700 48862 14702 48914
rect 14702 48862 14754 48914
rect 14754 48862 14756 48914
rect 14700 48860 14756 48862
rect 14588 47570 14644 47572
rect 14588 47518 14590 47570
rect 14590 47518 14642 47570
rect 14642 47518 14644 47570
rect 14588 47516 14644 47518
rect 14700 47346 14756 47348
rect 14700 47294 14702 47346
rect 14702 47294 14754 47346
rect 14754 47294 14756 47346
rect 14700 47292 14756 47294
rect 15036 47180 15092 47236
rect 12796 45724 12852 45780
rect 12012 45276 12068 45332
rect 11340 44828 11396 44884
rect 9324 41580 9380 41636
rect 9772 42530 9828 42532
rect 9772 42478 9774 42530
rect 9774 42478 9826 42530
rect 9826 42478 9828 42530
rect 9772 42476 9828 42478
rect 9660 41580 9716 41636
rect 10108 42530 10164 42532
rect 10108 42478 10110 42530
rect 10110 42478 10162 42530
rect 10162 42478 10164 42530
rect 10108 42476 10164 42478
rect 12348 45164 12404 45220
rect 12124 44994 12180 44996
rect 12124 44942 12126 44994
rect 12126 44942 12178 44994
rect 12178 44942 12180 44994
rect 12124 44940 12180 44942
rect 11340 43426 11396 43428
rect 11340 43374 11342 43426
rect 11342 43374 11394 43426
rect 11394 43374 11396 43426
rect 11340 43372 11396 43374
rect 11228 43148 11284 43204
rect 10444 42028 10500 42084
rect 9884 40908 9940 40964
rect 9324 40684 9380 40740
rect 9212 40572 9268 40628
rect 9100 40514 9156 40516
rect 9100 40462 9102 40514
rect 9102 40462 9154 40514
rect 9154 40462 9156 40514
rect 9100 40460 9156 40462
rect 8988 40124 9044 40180
rect 9100 39618 9156 39620
rect 9100 39566 9102 39618
rect 9102 39566 9154 39618
rect 9154 39566 9156 39618
rect 9100 39564 9156 39566
rect 9436 39004 9492 39060
rect 10668 41970 10724 41972
rect 10668 41918 10670 41970
rect 10670 41918 10722 41970
rect 10722 41918 10724 41970
rect 10668 41916 10724 41918
rect 10892 41692 10948 41748
rect 10108 41186 10164 41188
rect 10108 41134 10110 41186
rect 10110 41134 10162 41186
rect 10162 41134 10164 41186
rect 10108 41132 10164 41134
rect 10668 40460 10724 40516
rect 10892 40348 10948 40404
rect 11116 41020 11172 41076
rect 9996 39340 10052 39396
rect 10108 38892 10164 38948
rect 8988 38444 9044 38500
rect 9772 38444 9828 38500
rect 9212 37938 9268 37940
rect 9212 37886 9214 37938
rect 9214 37886 9266 37938
rect 9266 37886 9268 37938
rect 9212 37884 9268 37886
rect 9548 37884 9604 37940
rect 9884 37826 9940 37828
rect 9884 37774 9886 37826
rect 9886 37774 9938 37826
rect 9938 37774 9940 37826
rect 9884 37772 9940 37774
rect 9884 37324 9940 37380
rect 8316 36988 8372 37044
rect 8204 36258 8260 36260
rect 8204 36206 8206 36258
rect 8206 36206 8258 36258
rect 8258 36206 8260 36258
rect 8204 36204 8260 36206
rect 7756 36092 7812 36148
rect 7756 35644 7812 35700
rect 7308 35084 7364 35140
rect 7196 34300 7252 34356
rect 7756 34802 7812 34804
rect 7756 34750 7758 34802
rect 7758 34750 7810 34802
rect 7810 34750 7812 34802
rect 7756 34748 7812 34750
rect 8652 35868 8708 35924
rect 8764 37100 8820 37156
rect 8652 35698 8708 35700
rect 8652 35646 8654 35698
rect 8654 35646 8706 35698
rect 8706 35646 8708 35698
rect 8652 35644 8708 35646
rect 7980 35474 8036 35476
rect 7980 35422 7982 35474
rect 7982 35422 8034 35474
rect 8034 35422 8036 35474
rect 7980 35420 8036 35422
rect 7980 35084 8036 35140
rect 6076 33516 6132 33572
rect 6188 33404 6244 33460
rect 5852 33180 5908 33236
rect 5516 32786 5572 32788
rect 5516 32734 5518 32786
rect 5518 32734 5570 32786
rect 5570 32734 5572 32786
rect 5516 32732 5572 32734
rect 5292 32620 5348 32676
rect 5964 33346 6020 33348
rect 5964 33294 5966 33346
rect 5966 33294 6018 33346
rect 6018 33294 6020 33346
rect 5964 33292 6020 33294
rect 7644 34300 7700 34356
rect 6748 33292 6804 33348
rect 6188 32956 6244 33012
rect 6188 32284 6244 32340
rect 5628 31890 5684 31892
rect 5628 31838 5630 31890
rect 5630 31838 5682 31890
rect 5682 31838 5684 31890
rect 5628 31836 5684 31838
rect 7644 33292 7700 33348
rect 7756 33234 7812 33236
rect 7756 33182 7758 33234
rect 7758 33182 7810 33234
rect 7810 33182 7812 33234
rect 7756 33180 7812 33182
rect 7308 32956 7364 33012
rect 7420 32732 7476 32788
rect 7868 32732 7924 32788
rect 7644 32620 7700 32676
rect 6860 31836 6916 31892
rect 6524 31724 6580 31780
rect 7868 31948 7924 32004
rect 8876 36988 8932 37044
rect 8652 34636 8708 34692
rect 8428 34130 8484 34132
rect 8428 34078 8430 34130
rect 8430 34078 8482 34130
rect 8482 34078 8484 34130
rect 8428 34076 8484 34078
rect 8988 36428 9044 36484
rect 9548 35644 9604 35700
rect 8988 35474 9044 35476
rect 8988 35422 8990 35474
rect 8990 35422 9042 35474
rect 9042 35422 9044 35474
rect 8988 35420 9044 35422
rect 9660 35308 9716 35364
rect 9772 35420 9828 35476
rect 8428 33458 8484 33460
rect 8428 33406 8430 33458
rect 8430 33406 8482 33458
rect 8482 33406 8484 33458
rect 8428 33404 8484 33406
rect 9212 34748 9268 34804
rect 10556 39394 10612 39396
rect 10556 39342 10558 39394
rect 10558 39342 10610 39394
rect 10610 39342 10612 39394
rect 10556 39340 10612 39342
rect 10444 37772 10500 37828
rect 12348 44322 12404 44324
rect 12348 44270 12350 44322
rect 12350 44270 12402 44322
rect 12402 44270 12404 44322
rect 12348 44268 12404 44270
rect 12572 45218 12628 45220
rect 12572 45166 12574 45218
rect 12574 45166 12626 45218
rect 12626 45166 12628 45218
rect 12572 45164 12628 45166
rect 13804 45724 13860 45780
rect 13580 45612 13636 45668
rect 13468 44268 13524 44324
rect 13916 45276 13972 45332
rect 14140 45164 14196 45220
rect 14028 43762 14084 43764
rect 14028 43710 14030 43762
rect 14030 43710 14082 43762
rect 14082 43710 14084 43762
rect 14028 43708 14084 43710
rect 14364 45276 14420 45332
rect 12908 43372 12964 43428
rect 14028 43372 14084 43428
rect 11564 41804 11620 41860
rect 11564 41186 11620 41188
rect 11564 41134 11566 41186
rect 11566 41134 11618 41186
rect 11618 41134 11620 41186
rect 11564 41132 11620 41134
rect 12684 42530 12740 42532
rect 12684 42478 12686 42530
rect 12686 42478 12738 42530
rect 12738 42478 12740 42530
rect 12684 42476 12740 42478
rect 13804 42476 13860 42532
rect 11900 41132 11956 41188
rect 12012 41804 12068 41860
rect 11788 40460 11844 40516
rect 12236 41074 12292 41076
rect 12236 41022 12238 41074
rect 12238 41022 12290 41074
rect 12290 41022 12292 41074
rect 12236 41020 12292 41022
rect 12460 41132 12516 41188
rect 12796 41970 12852 41972
rect 12796 41918 12798 41970
rect 12798 41918 12850 41970
rect 12850 41918 12852 41970
rect 12796 41916 12852 41918
rect 13356 41916 13412 41972
rect 13916 42028 13972 42084
rect 14252 41804 14308 41860
rect 14364 42028 14420 42084
rect 13356 40572 13412 40628
rect 12460 40348 12516 40404
rect 13244 40402 13300 40404
rect 13244 40350 13246 40402
rect 13246 40350 13298 40402
rect 13298 40350 13300 40402
rect 13244 40348 13300 40350
rect 13244 40124 13300 40180
rect 11340 39618 11396 39620
rect 11340 39566 11342 39618
rect 11342 39566 11394 39618
rect 11394 39566 11396 39618
rect 11340 39564 11396 39566
rect 11452 39452 11508 39508
rect 12908 39452 12964 39508
rect 11228 38946 11284 38948
rect 11228 38894 11230 38946
rect 11230 38894 11282 38946
rect 11282 38894 11284 38946
rect 11228 38892 11284 38894
rect 12124 39058 12180 39060
rect 12124 39006 12126 39058
rect 12126 39006 12178 39058
rect 12178 39006 12180 39058
rect 12124 39004 12180 39006
rect 11788 38892 11844 38948
rect 10780 37772 10836 37828
rect 11228 37436 11284 37492
rect 10220 36482 10276 36484
rect 10220 36430 10222 36482
rect 10222 36430 10274 36482
rect 10274 36430 10276 36482
rect 10220 36428 10276 36430
rect 11116 36428 11172 36484
rect 10668 35980 10724 36036
rect 10892 35922 10948 35924
rect 10892 35870 10894 35922
rect 10894 35870 10946 35922
rect 10946 35870 10948 35922
rect 10892 35868 10948 35870
rect 10332 34860 10388 34916
rect 10108 34690 10164 34692
rect 10108 34638 10110 34690
rect 10110 34638 10162 34690
rect 10162 34638 10164 34690
rect 10108 34636 10164 34638
rect 9996 34242 10052 34244
rect 9996 34190 9998 34242
rect 9998 34190 10050 34242
rect 10050 34190 10052 34242
rect 9996 34188 10052 34190
rect 9212 33964 9268 34020
rect 9884 34076 9940 34132
rect 9100 33404 9156 33460
rect 9324 33852 9380 33908
rect 9324 33516 9380 33572
rect 9548 33292 9604 33348
rect 8092 32956 8148 33012
rect 8540 32562 8596 32564
rect 8540 32510 8542 32562
rect 8542 32510 8594 32562
rect 8594 32510 8596 32562
rect 8540 32508 8596 32510
rect 6524 31554 6580 31556
rect 6524 31502 6526 31554
rect 6526 31502 6578 31554
rect 6578 31502 6580 31554
rect 6524 31500 6580 31502
rect 5852 31164 5908 31220
rect 4284 29932 4340 29988
rect 4284 29484 4340 29540
rect 6636 31164 6692 31220
rect 6076 31052 6132 31108
rect 6412 31052 6468 31108
rect 5404 30882 5460 30884
rect 5404 30830 5406 30882
rect 5406 30830 5458 30882
rect 5458 30830 5460 30882
rect 5404 30828 5460 30830
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 6524 30994 6580 30996
rect 6524 30942 6526 30994
rect 6526 30942 6578 30994
rect 6578 30942 6580 30994
rect 6524 30940 6580 30942
rect 6524 29820 6580 29876
rect 6748 31106 6804 31108
rect 6748 31054 6750 31106
rect 6750 31054 6802 31106
rect 6802 31054 6804 31106
rect 6748 31052 6804 31054
rect 7308 31554 7364 31556
rect 7308 31502 7310 31554
rect 7310 31502 7362 31554
rect 7362 31502 7364 31554
rect 7308 31500 7364 31502
rect 7084 31388 7140 31444
rect 9660 32786 9716 32788
rect 9660 32734 9662 32786
rect 9662 32734 9714 32786
rect 9714 32734 9716 32786
rect 9660 32732 9716 32734
rect 8876 32284 8932 32340
rect 8652 31890 8708 31892
rect 8652 31838 8654 31890
rect 8654 31838 8706 31890
rect 8706 31838 8708 31890
rect 8652 31836 8708 31838
rect 8540 31778 8596 31780
rect 8540 31726 8542 31778
rect 8542 31726 8594 31778
rect 8594 31726 8596 31778
rect 8540 31724 8596 31726
rect 7084 31052 7140 31108
rect 7532 30940 7588 30996
rect 6860 29372 6916 29428
rect 7420 29820 7476 29876
rect 7532 29372 7588 29428
rect 7868 30994 7924 30996
rect 7868 30942 7870 30994
rect 7870 30942 7922 30994
rect 7922 30942 7924 30994
rect 7868 30940 7924 30942
rect 8204 30156 8260 30212
rect 8092 30098 8148 30100
rect 8092 30046 8094 30098
rect 8094 30046 8146 30098
rect 8146 30046 8148 30098
rect 8092 30044 8148 30046
rect 8876 31052 8932 31108
rect 9436 31164 9492 31220
rect 9996 33458 10052 33460
rect 9996 33406 9998 33458
rect 9998 33406 10050 33458
rect 10050 33406 10052 33458
rect 9996 33404 10052 33406
rect 8988 30210 9044 30212
rect 8988 30158 8990 30210
rect 8990 30158 9042 30210
rect 9042 30158 9044 30210
rect 8988 30156 9044 30158
rect 8316 29820 8372 29876
rect 7756 29708 7812 29764
rect 10556 34914 10612 34916
rect 10556 34862 10558 34914
rect 10558 34862 10610 34914
rect 10610 34862 10612 34914
rect 10556 34860 10612 34862
rect 10668 34802 10724 34804
rect 10668 34750 10670 34802
rect 10670 34750 10722 34802
rect 10722 34750 10724 34802
rect 10668 34748 10724 34750
rect 10556 34188 10612 34244
rect 11340 34972 11396 35028
rect 12796 37826 12852 37828
rect 12796 37774 12798 37826
rect 12798 37774 12850 37826
rect 12850 37774 12852 37826
rect 12796 37772 12852 37774
rect 12012 37436 12068 37492
rect 13020 37996 13076 38052
rect 12908 36594 12964 36596
rect 12908 36542 12910 36594
rect 12910 36542 12962 36594
rect 12962 36542 12964 36594
rect 12908 36540 12964 36542
rect 11676 36482 11732 36484
rect 11676 36430 11678 36482
rect 11678 36430 11730 36482
rect 11730 36430 11732 36482
rect 11676 36428 11732 36430
rect 12348 36482 12404 36484
rect 12348 36430 12350 36482
rect 12350 36430 12402 36482
rect 12402 36430 12404 36482
rect 12348 36428 12404 36430
rect 11788 36258 11844 36260
rect 11788 36206 11790 36258
rect 11790 36206 11842 36258
rect 11842 36206 11844 36258
rect 11788 36204 11844 36206
rect 11452 34860 11508 34916
rect 11340 34130 11396 34132
rect 11340 34078 11342 34130
rect 11342 34078 11394 34130
rect 11394 34078 11396 34130
rect 11340 34076 11396 34078
rect 10668 33404 10724 33460
rect 11564 34018 11620 34020
rect 11564 33966 11566 34018
rect 11566 33966 11618 34018
rect 11618 33966 11620 34018
rect 11564 33964 11620 33966
rect 11788 33404 11844 33460
rect 10108 32674 10164 32676
rect 10108 32622 10110 32674
rect 10110 32622 10162 32674
rect 10162 32622 10164 32674
rect 10108 32620 10164 32622
rect 11676 32620 11732 32676
rect 10220 32562 10276 32564
rect 10220 32510 10222 32562
rect 10222 32510 10274 32562
rect 10274 32510 10276 32562
rect 10220 32508 10276 32510
rect 10332 31836 10388 31892
rect 10108 31778 10164 31780
rect 10108 31726 10110 31778
rect 10110 31726 10162 31778
rect 10162 31726 10164 31778
rect 10108 31724 10164 31726
rect 12012 31890 12068 31892
rect 12012 31838 12014 31890
rect 12014 31838 12066 31890
rect 12066 31838 12068 31890
rect 12012 31836 12068 31838
rect 10220 31554 10276 31556
rect 10220 31502 10222 31554
rect 10222 31502 10274 31554
rect 10274 31502 10276 31554
rect 10220 31500 10276 31502
rect 11452 31164 11508 31220
rect 10220 31106 10276 31108
rect 10220 31054 10222 31106
rect 10222 31054 10274 31106
rect 10274 31054 10276 31106
rect 10220 31052 10276 31054
rect 10108 30210 10164 30212
rect 10108 30158 10110 30210
rect 10110 30158 10162 30210
rect 10162 30158 10164 30210
rect 10108 30156 10164 30158
rect 11788 30994 11844 30996
rect 11788 30942 11790 30994
rect 11790 30942 11842 30994
rect 11842 30942 11844 30994
rect 11788 30940 11844 30942
rect 12348 35868 12404 35924
rect 12684 35644 12740 35700
rect 12908 35698 12964 35700
rect 12908 35646 12910 35698
rect 12910 35646 12962 35698
rect 12962 35646 12964 35698
rect 12908 35644 12964 35646
rect 12796 34748 12852 34804
rect 13020 34748 13076 34804
rect 12796 33458 12852 33460
rect 12796 33406 12798 33458
rect 12798 33406 12850 33458
rect 12850 33406 12852 33458
rect 12796 33404 12852 33406
rect 12460 31106 12516 31108
rect 12460 31054 12462 31106
rect 12462 31054 12514 31106
rect 12514 31054 12516 31106
rect 12460 31052 12516 31054
rect 14028 40460 14084 40516
rect 13804 39004 13860 39060
rect 13356 37660 13412 37716
rect 13468 38556 13524 38612
rect 13916 38332 13972 38388
rect 13580 38162 13636 38164
rect 13580 38110 13582 38162
rect 13582 38110 13634 38162
rect 13634 38110 13636 38162
rect 13580 38108 13636 38110
rect 14028 38108 14084 38164
rect 14140 38780 14196 38836
rect 14252 38332 14308 38388
rect 13916 37436 13972 37492
rect 14028 37378 14084 37380
rect 14028 37326 14030 37378
rect 14030 37326 14082 37378
rect 14082 37326 14084 37378
rect 14028 37324 14084 37326
rect 13804 36540 13860 36596
rect 13692 35756 13748 35812
rect 13804 35698 13860 35700
rect 13804 35646 13806 35698
rect 13806 35646 13858 35698
rect 13858 35646 13860 35698
rect 13804 35644 13860 35646
rect 14364 37884 14420 37940
rect 14588 40514 14644 40516
rect 14588 40462 14590 40514
rect 14590 40462 14642 40514
rect 14642 40462 14644 40514
rect 14588 40460 14644 40462
rect 14588 37436 14644 37492
rect 14476 36540 14532 36596
rect 14812 45948 14868 46004
rect 16828 50594 16884 50596
rect 16828 50542 16830 50594
rect 16830 50542 16882 50594
rect 16882 50542 16884 50594
rect 16828 50540 16884 50542
rect 15932 48412 15988 48468
rect 16380 49026 16436 49028
rect 16380 48974 16382 49026
rect 16382 48974 16434 49026
rect 16434 48974 16436 49026
rect 16380 48972 16436 48974
rect 17052 48914 17108 48916
rect 17052 48862 17054 48914
rect 17054 48862 17106 48914
rect 17106 48862 17108 48914
rect 17052 48860 17108 48862
rect 15932 47516 15988 47572
rect 16380 47740 16436 47796
rect 16380 47516 16436 47572
rect 15596 47180 15652 47236
rect 20188 52162 20244 52164
rect 20188 52110 20190 52162
rect 20190 52110 20242 52162
rect 20242 52110 20244 52162
rect 20188 52108 20244 52110
rect 18508 50482 18564 50484
rect 18508 50430 18510 50482
rect 18510 50430 18562 50482
rect 18562 50430 18564 50482
rect 18508 50428 18564 50430
rect 20748 52834 20804 52836
rect 20748 52782 20750 52834
rect 20750 52782 20802 52834
rect 20802 52782 20804 52834
rect 20748 52780 20804 52782
rect 21308 52780 21364 52836
rect 21308 52444 21364 52500
rect 21196 51996 21252 52052
rect 19836 51770 19892 51772
rect 19836 51718 19838 51770
rect 19838 51718 19890 51770
rect 19890 51718 19892 51770
rect 19836 51716 19892 51718
rect 19940 51770 19996 51772
rect 19940 51718 19942 51770
rect 19942 51718 19994 51770
rect 19994 51718 19996 51770
rect 19940 51716 19996 51718
rect 20044 51770 20100 51772
rect 20044 51718 20046 51770
rect 20046 51718 20098 51770
rect 20098 51718 20100 51770
rect 20044 51716 20100 51718
rect 20076 51436 20132 51492
rect 20300 50540 20356 50596
rect 20636 51602 20692 51604
rect 20636 51550 20638 51602
rect 20638 51550 20690 51602
rect 20690 51550 20692 51602
rect 20636 51548 20692 51550
rect 21532 53058 21588 53060
rect 21532 53006 21534 53058
rect 21534 53006 21586 53058
rect 21586 53006 21588 53058
rect 21532 53004 21588 53006
rect 21644 51996 21700 52052
rect 21532 51938 21588 51940
rect 21532 51886 21534 51938
rect 21534 51886 21586 51938
rect 21586 51886 21588 51938
rect 21532 51884 21588 51886
rect 21532 51660 21588 51716
rect 20860 51490 20916 51492
rect 20860 51438 20862 51490
rect 20862 51438 20914 51490
rect 20914 51438 20916 51490
rect 20860 51436 20916 51438
rect 21644 51602 21700 51604
rect 21644 51550 21646 51602
rect 21646 51550 21698 51602
rect 21698 51550 21700 51602
rect 21644 51548 21700 51550
rect 19292 49756 19348 49812
rect 19836 50202 19892 50204
rect 19836 50150 19838 50202
rect 19838 50150 19890 50202
rect 19890 50150 19892 50202
rect 19836 50148 19892 50150
rect 19940 50202 19996 50204
rect 19940 50150 19942 50202
rect 19942 50150 19994 50202
rect 19994 50150 19996 50202
rect 19940 50148 19996 50150
rect 20044 50202 20100 50204
rect 20044 50150 20046 50202
rect 20046 50150 20098 50202
rect 20098 50150 20100 50202
rect 20044 50148 20100 50150
rect 20188 49922 20244 49924
rect 20188 49870 20190 49922
rect 20190 49870 20242 49922
rect 20242 49870 20244 49922
rect 20188 49868 20244 49870
rect 19404 49084 19460 49140
rect 17388 48412 17444 48468
rect 17724 47628 17780 47684
rect 17276 47458 17332 47460
rect 17276 47406 17278 47458
rect 17278 47406 17330 47458
rect 17330 47406 17332 47458
rect 17276 47404 17332 47406
rect 16716 46732 16772 46788
rect 17500 47292 17556 47348
rect 16604 46620 16660 46676
rect 15484 45948 15540 46004
rect 15932 45724 15988 45780
rect 15932 45388 15988 45444
rect 14924 43484 14980 43540
rect 15820 45164 15876 45220
rect 16380 45330 16436 45332
rect 16380 45278 16382 45330
rect 16382 45278 16434 45330
rect 16434 45278 16436 45330
rect 16380 45276 16436 45278
rect 16716 45724 16772 45780
rect 15484 42028 15540 42084
rect 15708 43372 15764 43428
rect 15372 41970 15428 41972
rect 15372 41918 15374 41970
rect 15374 41918 15426 41970
rect 15426 41918 15428 41970
rect 15372 41916 15428 41918
rect 14924 38892 14980 38948
rect 15372 38834 15428 38836
rect 15372 38782 15374 38834
rect 15374 38782 15426 38834
rect 15426 38782 15428 38834
rect 15372 38780 15428 38782
rect 14812 38556 14868 38612
rect 15036 37884 15092 37940
rect 15372 37548 15428 37604
rect 17948 47292 18004 47348
rect 18732 48748 18788 48804
rect 19516 48914 19572 48916
rect 19516 48862 19518 48914
rect 19518 48862 19570 48914
rect 19570 48862 19572 48914
rect 19516 48860 19572 48862
rect 19404 48748 19460 48804
rect 20524 49810 20580 49812
rect 20524 49758 20526 49810
rect 20526 49758 20578 49810
rect 20578 49758 20580 49810
rect 20524 49756 20580 49758
rect 20188 48860 20244 48916
rect 21196 50652 21252 50708
rect 21980 52220 22036 52276
rect 21980 52050 22036 52052
rect 21980 51998 21982 52050
rect 21982 51998 22034 52050
rect 22034 51998 22036 52050
rect 21980 51996 22036 51998
rect 21868 51772 21924 51828
rect 22316 52556 22372 52612
rect 23884 53618 23940 53620
rect 23884 53566 23886 53618
rect 23886 53566 23938 53618
rect 23938 53566 23940 53618
rect 23884 53564 23940 53566
rect 22652 53004 22708 53060
rect 23660 53004 23716 53060
rect 23436 52780 23492 52836
rect 22540 51884 22596 51940
rect 23100 51884 23156 51940
rect 21532 49868 21588 49924
rect 20524 48802 20580 48804
rect 20524 48750 20526 48802
rect 20526 48750 20578 48802
rect 20578 48750 20580 48802
rect 20524 48748 20580 48750
rect 19836 48634 19892 48636
rect 19836 48582 19838 48634
rect 19838 48582 19890 48634
rect 19890 48582 19892 48634
rect 19836 48580 19892 48582
rect 19940 48634 19996 48636
rect 19940 48582 19942 48634
rect 19942 48582 19994 48634
rect 19994 48582 19996 48634
rect 19940 48580 19996 48582
rect 20044 48634 20100 48636
rect 20044 48582 20046 48634
rect 20046 48582 20098 48634
rect 20098 48582 20100 48634
rect 20044 48580 20100 48582
rect 19292 48412 19348 48468
rect 19852 48466 19908 48468
rect 19852 48414 19854 48466
rect 19854 48414 19906 48466
rect 19906 48414 19908 48466
rect 19852 48412 19908 48414
rect 18508 47516 18564 47572
rect 18620 47346 18676 47348
rect 18620 47294 18622 47346
rect 18622 47294 18674 47346
rect 18674 47294 18676 47346
rect 18620 47292 18676 47294
rect 19292 47292 19348 47348
rect 17724 46674 17780 46676
rect 17724 46622 17726 46674
rect 17726 46622 17778 46674
rect 17778 46622 17780 46674
rect 17724 46620 17780 46622
rect 17612 45164 17668 45220
rect 17724 45276 17780 45332
rect 16604 44828 16660 44884
rect 17836 44492 17892 44548
rect 16828 43932 16884 43988
rect 16380 42588 16436 42644
rect 16492 42140 16548 42196
rect 17388 43260 17444 43316
rect 16716 42140 16772 42196
rect 16716 41298 16772 41300
rect 16716 41246 16718 41298
rect 16718 41246 16770 41298
rect 16770 41246 16772 41298
rect 16716 41244 16772 41246
rect 16044 40236 16100 40292
rect 16604 41020 16660 41076
rect 16156 40402 16212 40404
rect 16156 40350 16158 40402
rect 16158 40350 16210 40402
rect 16210 40350 16212 40402
rect 16156 40348 16212 40350
rect 16156 39564 16212 39620
rect 16268 39452 16324 39508
rect 17724 43426 17780 43428
rect 17724 43374 17726 43426
rect 17726 43374 17778 43426
rect 17778 43374 17780 43426
rect 17724 43372 17780 43374
rect 19068 47180 19124 47236
rect 18732 45778 18788 45780
rect 18732 45726 18734 45778
rect 18734 45726 18786 45778
rect 18786 45726 18788 45778
rect 18732 45724 18788 45726
rect 19628 48242 19684 48244
rect 19628 48190 19630 48242
rect 19630 48190 19682 48242
rect 19682 48190 19684 48242
rect 19628 48188 19684 48190
rect 20860 48412 20916 48468
rect 20972 48748 21028 48804
rect 19404 46786 19460 46788
rect 19404 46734 19406 46786
rect 19406 46734 19458 46786
rect 19458 46734 19460 46786
rect 19404 46732 19460 46734
rect 19964 48188 20020 48244
rect 19852 47346 19908 47348
rect 19852 47294 19854 47346
rect 19854 47294 19906 47346
rect 19906 47294 19908 47346
rect 19852 47292 19908 47294
rect 20300 47346 20356 47348
rect 20300 47294 20302 47346
rect 20302 47294 20354 47346
rect 20354 47294 20356 47346
rect 20300 47292 20356 47294
rect 19740 47180 19796 47236
rect 19836 47066 19892 47068
rect 19836 47014 19838 47066
rect 19838 47014 19890 47066
rect 19890 47014 19892 47066
rect 19836 47012 19892 47014
rect 19940 47066 19996 47068
rect 19940 47014 19942 47066
rect 19942 47014 19994 47066
rect 19994 47014 19996 47066
rect 19940 47012 19996 47014
rect 20044 47066 20100 47068
rect 20044 47014 20046 47066
rect 20046 47014 20098 47066
rect 20098 47014 20100 47066
rect 20044 47012 20100 47014
rect 20300 46844 20356 46900
rect 19628 46786 19684 46788
rect 19628 46734 19630 46786
rect 19630 46734 19682 46786
rect 19682 46734 19684 46786
rect 19628 46732 19684 46734
rect 20748 46786 20804 46788
rect 20748 46734 20750 46786
rect 20750 46734 20802 46786
rect 20802 46734 20804 46786
rect 20748 46732 20804 46734
rect 20188 46620 20244 46676
rect 19068 45666 19124 45668
rect 19068 45614 19070 45666
rect 19070 45614 19122 45666
rect 19122 45614 19124 45666
rect 19068 45612 19124 45614
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 18956 45164 19012 45220
rect 19404 44492 19460 44548
rect 19292 44044 19348 44100
rect 18620 43426 18676 43428
rect 18620 43374 18622 43426
rect 18622 43374 18674 43426
rect 18674 43374 18676 43426
rect 18620 43372 18676 43374
rect 17612 42476 17668 42532
rect 17500 41244 17556 41300
rect 17612 41020 17668 41076
rect 18060 42588 18116 42644
rect 20524 46674 20580 46676
rect 20524 46622 20526 46674
rect 20526 46622 20578 46674
rect 20578 46622 20580 46674
rect 20524 46620 20580 46622
rect 20860 46674 20916 46676
rect 20860 46622 20862 46674
rect 20862 46622 20914 46674
rect 20914 46622 20916 46674
rect 20860 46620 20916 46622
rect 22652 50594 22708 50596
rect 22652 50542 22654 50594
rect 22654 50542 22706 50594
rect 22706 50542 22708 50594
rect 22652 50540 22708 50542
rect 21868 48972 21924 49028
rect 21980 49084 22036 49140
rect 21420 48748 21476 48804
rect 21196 48466 21252 48468
rect 21196 48414 21198 48466
rect 21198 48414 21250 48466
rect 21250 48414 21252 48466
rect 21196 48412 21252 48414
rect 21196 47458 21252 47460
rect 21196 47406 21198 47458
rect 21198 47406 21250 47458
rect 21250 47406 21252 47458
rect 21196 47404 21252 47406
rect 21532 47292 21588 47348
rect 21980 47180 22036 47236
rect 20524 45388 20580 45444
rect 19516 43596 19572 43652
rect 19404 43426 19460 43428
rect 19404 43374 19406 43426
rect 19406 43374 19458 43426
rect 19458 43374 19460 43426
rect 19404 43372 19460 43374
rect 19964 44322 20020 44324
rect 19964 44270 19966 44322
rect 19966 44270 20018 44322
rect 20018 44270 20020 44322
rect 19964 44268 20020 44270
rect 20412 44492 20468 44548
rect 19852 44044 19908 44100
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 20076 43650 20132 43652
rect 20076 43598 20078 43650
rect 20078 43598 20130 43650
rect 20130 43598 20132 43650
rect 20076 43596 20132 43598
rect 19740 43426 19796 43428
rect 19740 43374 19742 43426
rect 19742 43374 19794 43426
rect 19794 43374 19796 43426
rect 19740 43372 19796 43374
rect 20412 43372 20468 43428
rect 19180 42642 19236 42644
rect 19180 42590 19182 42642
rect 19182 42590 19234 42642
rect 19234 42590 19236 42642
rect 19180 42588 19236 42590
rect 18956 42476 19012 42532
rect 17948 41186 18004 41188
rect 17948 41134 17950 41186
rect 17950 41134 18002 41186
rect 18002 41134 18004 41186
rect 17948 41132 18004 41134
rect 17836 40908 17892 40964
rect 18732 41186 18788 41188
rect 18732 41134 18734 41186
rect 18734 41134 18786 41186
rect 18786 41134 18788 41186
rect 18732 41132 18788 41134
rect 18844 41074 18900 41076
rect 18844 41022 18846 41074
rect 18846 41022 18898 41074
rect 18898 41022 18900 41074
rect 18844 41020 18900 41022
rect 19292 41074 19348 41076
rect 19292 41022 19294 41074
rect 19294 41022 19346 41074
rect 19346 41022 19348 41074
rect 19292 41020 19348 41022
rect 17388 40124 17444 40180
rect 17724 40236 17780 40292
rect 16828 39618 16884 39620
rect 16828 39566 16830 39618
rect 16830 39566 16882 39618
rect 16882 39566 16884 39618
rect 16828 39564 16884 39566
rect 17500 39618 17556 39620
rect 17500 39566 17502 39618
rect 17502 39566 17554 39618
rect 17554 39566 17556 39618
rect 17500 39564 17556 39566
rect 15932 38946 15988 38948
rect 15932 38894 15934 38946
rect 15934 38894 15986 38946
rect 15986 38894 15988 38946
rect 15932 38892 15988 38894
rect 15596 37772 15652 37828
rect 15932 37436 15988 37492
rect 15596 37266 15652 37268
rect 15596 37214 15598 37266
rect 15598 37214 15650 37266
rect 15650 37214 15652 37266
rect 15596 37212 15652 37214
rect 17388 39058 17444 39060
rect 17388 39006 17390 39058
rect 17390 39006 17442 39058
rect 17442 39006 17444 39058
rect 17388 39004 17444 39006
rect 16380 38946 16436 38948
rect 16380 38894 16382 38946
rect 16382 38894 16434 38946
rect 16434 38894 16436 38946
rect 16380 38892 16436 38894
rect 19068 40908 19124 40964
rect 19068 40572 19124 40628
rect 18284 40460 18340 40516
rect 18172 39676 18228 39732
rect 17836 39506 17892 39508
rect 17836 39454 17838 39506
rect 17838 39454 17890 39506
rect 17890 39454 17892 39506
rect 17836 39452 17892 39454
rect 18508 39564 18564 39620
rect 20524 42642 20580 42644
rect 20524 42590 20526 42642
rect 20526 42590 20578 42642
rect 20578 42590 20580 42642
rect 20524 42588 20580 42590
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 20748 42476 20804 42532
rect 19964 41074 20020 41076
rect 19964 41022 19966 41074
rect 19966 41022 20018 41074
rect 20018 41022 20020 41074
rect 19964 41020 20020 41022
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 21308 44322 21364 44324
rect 21308 44270 21310 44322
rect 21310 44270 21362 44322
rect 21362 44270 21364 44322
rect 21308 44268 21364 44270
rect 24332 53506 24388 53508
rect 24332 53454 24334 53506
rect 24334 53454 24386 53506
rect 24386 53454 24388 53506
rect 24332 53452 24388 53454
rect 23996 52780 24052 52836
rect 23884 52556 23940 52612
rect 22204 48636 22260 48692
rect 24556 52780 24612 52836
rect 27580 55916 27636 55972
rect 27468 55356 27524 55412
rect 25228 53564 25284 53620
rect 25676 53452 25732 53508
rect 24668 52386 24724 52388
rect 24668 52334 24670 52386
rect 24670 52334 24722 52386
rect 24722 52334 24724 52386
rect 24668 52332 24724 52334
rect 24556 52108 24612 52164
rect 22652 49868 22708 49924
rect 22988 49084 23044 49140
rect 22876 49026 22932 49028
rect 22876 48974 22878 49026
rect 22878 48974 22930 49026
rect 22930 48974 22932 49026
rect 22876 48972 22932 48974
rect 24556 50428 24612 50484
rect 22652 48466 22708 48468
rect 22652 48414 22654 48466
rect 22654 48414 22706 48466
rect 22706 48414 22708 48466
rect 22652 48412 22708 48414
rect 22204 46674 22260 46676
rect 22204 46622 22206 46674
rect 22206 46622 22258 46674
rect 22258 46622 22260 46674
rect 22204 46620 22260 46622
rect 22540 46844 22596 46900
rect 22652 47180 22708 47236
rect 22428 46508 22484 46564
rect 21532 45388 21588 45444
rect 22316 45612 22372 45668
rect 21868 45276 21924 45332
rect 23324 46620 23380 46676
rect 23660 46562 23716 46564
rect 23660 46510 23662 46562
rect 23662 46510 23714 46562
rect 23714 46510 23716 46562
rect 23660 46508 23716 46510
rect 23436 46396 23492 46452
rect 21420 42700 21476 42756
rect 22540 43596 22596 43652
rect 22988 43036 23044 43092
rect 21308 42642 21364 42644
rect 21308 42590 21310 42642
rect 21310 42590 21362 42642
rect 21362 42590 21364 42642
rect 21308 42588 21364 42590
rect 21308 40684 21364 40740
rect 19852 40572 19908 40628
rect 19292 40514 19348 40516
rect 19292 40462 19294 40514
rect 19294 40462 19346 40514
rect 19346 40462 19348 40514
rect 19292 40460 19348 40462
rect 18844 40402 18900 40404
rect 18844 40350 18846 40402
rect 18846 40350 18898 40402
rect 18898 40350 18900 40402
rect 18844 40348 18900 40350
rect 19740 40402 19796 40404
rect 19740 40350 19742 40402
rect 19742 40350 19794 40402
rect 19794 40350 19796 40402
rect 19740 40348 19796 40350
rect 20524 40626 20580 40628
rect 20524 40574 20526 40626
rect 20526 40574 20578 40626
rect 20578 40574 20580 40626
rect 20524 40572 20580 40574
rect 20412 40514 20468 40516
rect 20412 40462 20414 40514
rect 20414 40462 20466 40514
rect 20466 40462 20468 40514
rect 20412 40460 20468 40462
rect 20188 40402 20244 40404
rect 20188 40350 20190 40402
rect 20190 40350 20242 40402
rect 20242 40350 20244 40402
rect 20188 40348 20244 40350
rect 22092 42700 22148 42756
rect 21644 42530 21700 42532
rect 21644 42478 21646 42530
rect 21646 42478 21698 42530
rect 21698 42478 21700 42530
rect 21644 42476 21700 42478
rect 22652 42364 22708 42420
rect 21644 41916 21700 41972
rect 21756 41468 21812 41524
rect 21756 40572 21812 40628
rect 22204 41970 22260 41972
rect 22204 41918 22206 41970
rect 22206 41918 22258 41970
rect 22258 41918 22260 41970
rect 22204 41916 22260 41918
rect 22540 41468 22596 41524
rect 22092 40962 22148 40964
rect 22092 40910 22094 40962
rect 22094 40910 22146 40962
rect 22146 40910 22148 40962
rect 22092 40908 22148 40910
rect 20524 40124 20580 40180
rect 20412 39900 20468 39956
rect 18956 39340 19012 39396
rect 19180 39618 19236 39620
rect 19180 39566 19182 39618
rect 19182 39566 19234 39618
rect 19234 39566 19236 39618
rect 19180 39564 19236 39566
rect 17724 38946 17780 38948
rect 17724 38894 17726 38946
rect 17726 38894 17778 38946
rect 17778 38894 17780 38946
rect 17724 38892 17780 38894
rect 18060 39004 18116 39060
rect 17052 38668 17108 38724
rect 16268 37324 16324 37380
rect 16940 38332 16996 38388
rect 15708 37100 15764 37156
rect 14700 36652 14756 36708
rect 15148 36540 15204 36596
rect 15260 36316 15316 36372
rect 14476 35810 14532 35812
rect 14476 35758 14478 35810
rect 14478 35758 14530 35810
rect 14530 35758 14532 35810
rect 14476 35756 14532 35758
rect 13580 35026 13636 35028
rect 13580 34974 13582 35026
rect 13582 34974 13634 35026
rect 13634 34974 13636 35026
rect 13580 34972 13636 34974
rect 14140 34860 14196 34916
rect 13916 34802 13972 34804
rect 13916 34750 13918 34802
rect 13918 34750 13970 34802
rect 13970 34750 13972 34802
rect 13916 34748 13972 34750
rect 13916 34188 13972 34244
rect 13468 32562 13524 32564
rect 13468 32510 13470 32562
rect 13470 32510 13522 32562
rect 13522 32510 13524 32562
rect 13468 32508 13524 32510
rect 15036 34972 15092 35028
rect 15148 34914 15204 34916
rect 15148 34862 15150 34914
rect 15150 34862 15202 34914
rect 15202 34862 15204 34914
rect 15148 34860 15204 34862
rect 14476 34300 14532 34356
rect 15484 35756 15540 35812
rect 15372 35698 15428 35700
rect 15372 35646 15374 35698
rect 15374 35646 15426 35698
rect 15426 35646 15428 35698
rect 15372 35644 15428 35646
rect 14476 33458 14532 33460
rect 14476 33406 14478 33458
rect 14478 33406 14530 33458
rect 14530 33406 14532 33458
rect 14476 33404 14532 33406
rect 13916 31948 13972 32004
rect 13692 31890 13748 31892
rect 13692 31838 13694 31890
rect 13694 31838 13746 31890
rect 13746 31838 13748 31890
rect 13692 31836 13748 31838
rect 13244 30882 13300 30884
rect 13244 30830 13246 30882
rect 13246 30830 13298 30882
rect 13298 30830 13300 30882
rect 13244 30828 13300 30830
rect 12460 30322 12516 30324
rect 12460 30270 12462 30322
rect 12462 30270 12514 30322
rect 12514 30270 12516 30322
rect 12460 30268 12516 30270
rect 14252 31778 14308 31780
rect 14252 31726 14254 31778
rect 14254 31726 14306 31778
rect 14306 31726 14308 31778
rect 14252 31724 14308 31726
rect 15820 36540 15876 36596
rect 16156 36370 16212 36372
rect 16156 36318 16158 36370
rect 16158 36318 16210 36370
rect 16210 36318 16212 36370
rect 16156 36316 16212 36318
rect 16156 35026 16212 35028
rect 16156 34974 16158 35026
rect 16158 34974 16210 35026
rect 16210 34974 16212 35026
rect 16156 34972 16212 34974
rect 16044 34914 16100 34916
rect 16044 34862 16046 34914
rect 16046 34862 16098 34914
rect 16098 34862 16100 34914
rect 16044 34860 16100 34862
rect 16380 34748 16436 34804
rect 15596 34354 15652 34356
rect 15596 34302 15598 34354
rect 15598 34302 15650 34354
rect 15650 34302 15652 34354
rect 15596 34300 15652 34302
rect 17388 38162 17444 38164
rect 17388 38110 17390 38162
rect 17390 38110 17442 38162
rect 17442 38110 17444 38162
rect 17388 38108 17444 38110
rect 17948 37772 18004 37828
rect 17388 37660 17444 37716
rect 17164 36652 17220 36708
rect 17500 37154 17556 37156
rect 17500 37102 17502 37154
rect 17502 37102 17554 37154
rect 17554 37102 17556 37154
rect 17500 37100 17556 37102
rect 19404 39452 19460 39508
rect 19516 38892 19572 38948
rect 18284 37996 18340 38052
rect 18060 36652 18116 36708
rect 18172 37548 18228 37604
rect 18620 37548 18676 37604
rect 18508 36706 18564 36708
rect 18508 36654 18510 36706
rect 18510 36654 18562 36706
rect 18562 36654 18564 36706
rect 18508 36652 18564 36654
rect 18956 37826 19012 37828
rect 18956 37774 18958 37826
rect 18958 37774 19010 37826
rect 19010 37774 19012 37826
rect 18956 37772 19012 37774
rect 20188 39506 20244 39508
rect 20188 39454 20190 39506
rect 20190 39454 20242 39506
rect 20242 39454 20244 39506
rect 20188 39452 20244 39454
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 19964 38834 20020 38836
rect 19964 38782 19966 38834
rect 19966 38782 20018 38834
rect 20018 38782 20020 38834
rect 19964 38780 20020 38782
rect 20636 40012 20692 40068
rect 21308 39394 21364 39396
rect 21308 39342 21310 39394
rect 21310 39342 21362 39394
rect 21362 39342 21364 39394
rect 21308 39340 21364 39342
rect 21532 39564 21588 39620
rect 21644 39506 21700 39508
rect 21644 39454 21646 39506
rect 21646 39454 21698 39506
rect 21698 39454 21700 39506
rect 21644 39452 21700 39454
rect 20636 38892 20692 38948
rect 21420 38892 21476 38948
rect 21308 38722 21364 38724
rect 21308 38670 21310 38722
rect 21310 38670 21362 38722
rect 21362 38670 21364 38722
rect 21308 38668 21364 38670
rect 19740 38050 19796 38052
rect 19740 37998 19742 38050
rect 19742 37998 19794 38050
rect 19794 37998 19796 38050
rect 19740 37996 19796 37998
rect 19628 37548 19684 37604
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 20188 37324 20244 37380
rect 19068 37266 19124 37268
rect 19068 37214 19070 37266
rect 19070 37214 19122 37266
rect 19122 37214 19124 37266
rect 19068 37212 19124 37214
rect 18732 37100 18788 37156
rect 18956 36988 19012 37044
rect 20076 37042 20132 37044
rect 20076 36990 20078 37042
rect 20078 36990 20130 37042
rect 20130 36990 20132 37042
rect 20076 36988 20132 36990
rect 18732 36594 18788 36596
rect 18732 36542 18734 36594
rect 18734 36542 18786 36594
rect 18786 36542 18788 36594
rect 18732 36540 18788 36542
rect 17612 36204 17668 36260
rect 17388 35810 17444 35812
rect 17388 35758 17390 35810
rect 17390 35758 17442 35810
rect 17442 35758 17444 35810
rect 17388 35756 17444 35758
rect 17164 35644 17220 35700
rect 19964 36594 20020 36596
rect 19964 36542 19966 36594
rect 19966 36542 20018 36594
rect 20018 36542 20020 36594
rect 19964 36540 20020 36542
rect 18844 35756 18900 35812
rect 17948 35698 18004 35700
rect 17948 35646 17950 35698
rect 17950 35646 18002 35698
rect 18002 35646 18004 35698
rect 17948 35644 18004 35646
rect 17836 35586 17892 35588
rect 17836 35534 17838 35586
rect 17838 35534 17890 35586
rect 17890 35534 17892 35586
rect 17836 35532 17892 35534
rect 17164 34860 17220 34916
rect 17500 34914 17556 34916
rect 17500 34862 17502 34914
rect 17502 34862 17554 34914
rect 17554 34862 17556 34914
rect 17500 34860 17556 34862
rect 16940 34300 16996 34356
rect 17276 34412 17332 34468
rect 15708 34242 15764 34244
rect 15708 34190 15710 34242
rect 15710 34190 15762 34242
rect 15762 34190 15764 34242
rect 15708 34188 15764 34190
rect 14924 32620 14980 32676
rect 15260 31948 15316 32004
rect 14588 31836 14644 31892
rect 16380 31890 16436 31892
rect 16380 31838 16382 31890
rect 16382 31838 16434 31890
rect 16434 31838 16436 31890
rect 16380 31836 16436 31838
rect 16156 31778 16212 31780
rect 16156 31726 16158 31778
rect 16158 31726 16210 31778
rect 16210 31726 16212 31778
rect 16156 31724 16212 31726
rect 16604 31778 16660 31780
rect 16604 31726 16606 31778
rect 16606 31726 16658 31778
rect 16658 31726 16660 31778
rect 16604 31724 16660 31726
rect 14812 31612 14868 31668
rect 16604 30994 16660 30996
rect 16604 30942 16606 30994
rect 16606 30942 16658 30994
rect 16658 30942 16660 30994
rect 16604 30940 16660 30942
rect 15260 30828 15316 30884
rect 15260 30380 15316 30436
rect 13916 30268 13972 30324
rect 14700 30268 14756 30324
rect 11452 30210 11508 30212
rect 11452 30158 11454 30210
rect 11454 30158 11506 30210
rect 11506 30158 11508 30210
rect 11452 30156 11508 30158
rect 14476 30210 14532 30212
rect 14476 30158 14478 30210
rect 14478 30158 14530 30210
rect 14530 30158 14532 30210
rect 14476 30156 14532 30158
rect 10668 30044 10724 30100
rect 16604 30716 16660 30772
rect 16044 30434 16100 30436
rect 16044 30382 16046 30434
rect 16046 30382 16098 30434
rect 16098 30382 16100 30434
rect 16044 30380 16100 30382
rect 15372 30268 15428 30324
rect 15708 30210 15764 30212
rect 15708 30158 15710 30210
rect 15710 30158 15762 30210
rect 15762 30158 15764 30210
rect 15708 30156 15764 30158
rect 9660 29708 9716 29764
rect 13468 29932 13524 29988
rect 6636 29202 6692 29204
rect 6636 29150 6638 29202
rect 6638 29150 6690 29202
rect 6690 29150 6692 29202
rect 6636 29148 6692 29150
rect 8428 29426 8484 29428
rect 8428 29374 8430 29426
rect 8430 29374 8482 29426
rect 8482 29374 8484 29426
rect 8428 29372 8484 29374
rect 7868 29148 7924 29204
rect 14364 29426 14420 29428
rect 14364 29374 14366 29426
rect 14366 29374 14418 29426
rect 14418 29374 14420 29426
rect 14364 29372 14420 29374
rect 13468 29260 13524 29316
rect 8540 29148 8596 29204
rect 9996 29148 10052 29204
rect 6636 28588 6692 28644
rect 3612 27804 3668 27860
rect 6636 27804 6692 27860
rect 3164 27580 3220 27636
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 2492 26796 2548 26852
rect 2044 26514 2100 26516
rect 2044 26462 2046 26514
rect 2046 26462 2098 26514
rect 2098 26462 2100 26514
rect 2044 26460 2100 26462
rect 1820 26348 1876 26404
rect 3612 27074 3668 27076
rect 3612 27022 3614 27074
rect 3614 27022 3666 27074
rect 3666 27022 3668 27074
rect 3612 27020 3668 27022
rect 5068 27020 5124 27076
rect 3164 26796 3220 26852
rect 3388 26684 3444 26740
rect 2716 26572 2772 26628
rect 4732 26402 4788 26404
rect 4732 26350 4734 26402
rect 4734 26350 4786 26402
rect 4786 26350 4788 26402
rect 4732 26348 4788 26350
rect 2492 26236 2548 26292
rect 3052 26124 3108 26180
rect 3836 26178 3892 26180
rect 3836 26126 3838 26178
rect 3838 26126 3890 26178
rect 3890 26126 3892 26178
rect 3836 26124 3892 26126
rect 4284 26178 4340 26180
rect 4284 26126 4286 26178
rect 4286 26126 4338 26178
rect 4338 26126 4340 26178
rect 4284 26124 4340 26126
rect 2380 26012 2436 26068
rect 1932 24892 1988 24948
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 4844 25676 4900 25732
rect 4284 25506 4340 25508
rect 4284 25454 4286 25506
rect 4286 25454 4338 25506
rect 4338 25454 4340 25506
rect 4284 25452 4340 25454
rect 4620 25340 4676 25396
rect 2380 24220 2436 24276
rect 2380 24050 2436 24052
rect 2380 23998 2382 24050
rect 2382 23998 2434 24050
rect 2434 23998 2436 24050
rect 2380 23996 2436 23998
rect 2156 23772 2212 23828
rect 1932 23548 1988 23604
rect 1708 22876 1764 22932
rect 1708 20802 1764 20804
rect 1708 20750 1710 20802
rect 1710 20750 1762 20802
rect 1762 20750 1764 20802
rect 1708 20748 1764 20750
rect 1708 20188 1764 20244
rect 1932 21532 1988 21588
rect 2044 21308 2100 21364
rect 2268 23154 2324 23156
rect 2268 23102 2270 23154
rect 2270 23102 2322 23154
rect 2322 23102 2324 23154
rect 2268 23100 2324 23102
rect 2268 22764 2324 22820
rect 2604 23996 2660 24052
rect 2716 23884 2772 23940
rect 2940 23826 2996 23828
rect 2940 23774 2942 23826
rect 2942 23774 2994 23826
rect 2994 23774 2996 23826
rect 2940 23772 2996 23774
rect 2828 23660 2884 23716
rect 2828 23042 2884 23044
rect 2828 22990 2830 23042
rect 2830 22990 2882 23042
rect 2882 22990 2884 23042
rect 2828 22988 2884 22990
rect 2716 22258 2772 22260
rect 2716 22206 2718 22258
rect 2718 22206 2770 22258
rect 2770 22206 2772 22258
rect 2716 22204 2772 22206
rect 2604 21980 2660 22036
rect 2716 21586 2772 21588
rect 2716 21534 2718 21586
rect 2718 21534 2770 21586
rect 2770 21534 2772 21586
rect 2716 21532 2772 21534
rect 3164 23100 3220 23156
rect 4956 25452 5012 25508
rect 5404 25452 5460 25508
rect 5740 25788 5796 25844
rect 5180 25340 5236 25396
rect 5628 25394 5684 25396
rect 5628 25342 5630 25394
rect 5630 25342 5682 25394
rect 5682 25342 5684 25394
rect 5628 25340 5684 25342
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 3388 23938 3444 23940
rect 3388 23886 3390 23938
rect 3390 23886 3442 23938
rect 3442 23886 3444 23938
rect 3388 23884 3444 23886
rect 4620 23772 4676 23828
rect 4060 23714 4116 23716
rect 4060 23662 4062 23714
rect 4062 23662 4114 23714
rect 4114 23662 4116 23714
rect 4060 23660 4116 23662
rect 3612 23100 3668 23156
rect 3276 21868 3332 21924
rect 3500 22092 3556 22148
rect 2380 20748 2436 20804
rect 2492 20076 2548 20132
rect 1820 18172 1876 18228
rect 1820 17500 1876 17556
rect 1708 17052 1764 17108
rect 1820 17276 1876 17332
rect 2044 17554 2100 17556
rect 2044 17502 2046 17554
rect 2046 17502 2098 17554
rect 2098 17502 2100 17554
rect 2044 17500 2100 17502
rect 2604 20018 2660 20020
rect 2604 19966 2606 20018
rect 2606 19966 2658 20018
rect 2658 19966 2660 20018
rect 2604 19964 2660 19966
rect 2828 20578 2884 20580
rect 2828 20526 2830 20578
rect 2830 20526 2882 20578
rect 2882 20526 2884 20578
rect 2828 20524 2884 20526
rect 2716 19852 2772 19908
rect 2716 19404 2772 19460
rect 2380 19122 2436 19124
rect 2380 19070 2382 19122
rect 2382 19070 2434 19122
rect 2434 19070 2436 19122
rect 2380 19068 2436 19070
rect 2716 18396 2772 18452
rect 2492 18284 2548 18340
rect 2380 17164 2436 17220
rect 1932 16940 1988 16996
rect 2044 16604 2100 16660
rect 2940 18844 2996 18900
rect 2604 18060 2660 18116
rect 2940 17724 2996 17780
rect 3276 21196 3332 21252
rect 3276 19852 3332 19908
rect 3276 18620 3332 18676
rect 3388 20524 3444 20580
rect 3612 21980 3668 22036
rect 3724 22204 3780 22260
rect 3612 21532 3668 21588
rect 3612 20636 3668 20692
rect 4844 23154 4900 23156
rect 4844 23102 4846 23154
rect 4846 23102 4898 23154
rect 4898 23102 4900 23154
rect 4844 23100 4900 23102
rect 4172 22988 4228 23044
rect 4172 21756 4228 21812
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 5404 25228 5460 25284
rect 5852 25676 5908 25732
rect 6636 25788 6692 25844
rect 5964 25340 6020 25396
rect 6300 25452 6356 25508
rect 5740 24444 5796 24500
rect 5180 23714 5236 23716
rect 5180 23662 5182 23714
rect 5182 23662 5234 23714
rect 5234 23662 5236 23714
rect 5180 23660 5236 23662
rect 5068 21756 5124 21812
rect 6076 24444 6132 24500
rect 6076 23660 6132 23716
rect 6188 23884 6244 23940
rect 6076 22652 6132 22708
rect 5628 21586 5684 21588
rect 5628 21534 5630 21586
rect 5630 21534 5682 21586
rect 5682 21534 5684 21586
rect 5628 21532 5684 21534
rect 5180 20972 5236 21028
rect 3836 20690 3892 20692
rect 3836 20638 3838 20690
rect 3838 20638 3890 20690
rect 3890 20638 3892 20690
rect 3836 20636 3892 20638
rect 4956 20636 5012 20692
rect 3724 20018 3780 20020
rect 3724 19966 3726 20018
rect 3726 19966 3778 20018
rect 3778 19966 3780 20018
rect 3724 19964 3780 19966
rect 3836 20300 3892 20356
rect 3500 19068 3556 19124
rect 3612 19234 3668 19236
rect 3612 19182 3614 19234
rect 3614 19182 3666 19234
rect 3666 19182 3668 19234
rect 3612 19180 3668 19182
rect 4508 20578 4564 20580
rect 4508 20526 4510 20578
rect 4510 20526 4562 20578
rect 4562 20526 4564 20578
rect 4508 20524 4564 20526
rect 4732 20578 4788 20580
rect 4732 20526 4734 20578
rect 4734 20526 4786 20578
rect 4786 20526 4788 20578
rect 4732 20524 4788 20526
rect 4844 20412 4900 20468
rect 5964 20300 6020 20356
rect 5852 20188 5908 20244
rect 5516 20076 5572 20132
rect 5068 20018 5124 20020
rect 5068 19966 5070 20018
rect 5070 19966 5122 20018
rect 5122 19966 5124 20018
rect 5068 19964 5124 19966
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 4172 19180 4228 19236
rect 4956 19180 5012 19236
rect 3724 18674 3780 18676
rect 3724 18622 3726 18674
rect 3726 18622 3778 18674
rect 3778 18622 3780 18674
rect 3724 18620 3780 18622
rect 3388 17836 3444 17892
rect 3836 18284 3892 18340
rect 3388 17612 3444 17668
rect 2940 16940 2996 16996
rect 3164 16828 3220 16884
rect 3164 16156 3220 16212
rect 2940 15932 2996 15988
rect 1708 15708 1764 15764
rect 1708 15148 1764 15204
rect 2268 15708 2324 15764
rect 1932 15090 1988 15092
rect 1932 15038 1934 15090
rect 1934 15038 1986 15090
rect 1986 15038 1988 15090
rect 1932 15036 1988 15038
rect 2044 14700 2100 14756
rect 1820 13916 1876 13972
rect 2828 15874 2884 15876
rect 2828 15822 2830 15874
rect 2830 15822 2882 15874
rect 2882 15822 2884 15874
rect 2828 15820 2884 15822
rect 2492 15036 2548 15092
rect 2604 15372 2660 15428
rect 2604 14588 2660 14644
rect 2828 14476 2884 14532
rect 2044 13692 2100 13748
rect 1708 12850 1764 12852
rect 1708 12798 1710 12850
rect 1710 12798 1762 12850
rect 1762 12798 1764 12850
rect 1708 12796 1764 12798
rect 2380 13468 2436 13524
rect 3052 15148 3108 15204
rect 3500 16828 3556 16884
rect 3612 17500 3668 17556
rect 4060 18674 4116 18676
rect 4060 18622 4062 18674
rect 4062 18622 4114 18674
rect 4114 18622 4116 18674
rect 4060 18620 4116 18622
rect 5292 19180 5348 19236
rect 5180 18844 5236 18900
rect 5068 18508 5124 18564
rect 4508 18284 4564 18340
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 4396 17836 4452 17892
rect 4172 17442 4228 17444
rect 4172 17390 4174 17442
rect 4174 17390 4226 17442
rect 4226 17390 4228 17442
rect 4172 17388 4228 17390
rect 4508 17554 4564 17556
rect 4508 17502 4510 17554
rect 4510 17502 4562 17554
rect 4562 17502 4564 17554
rect 4508 17500 4564 17502
rect 4844 17554 4900 17556
rect 4844 17502 4846 17554
rect 4846 17502 4898 17554
rect 4898 17502 4900 17554
rect 4844 17500 4900 17502
rect 3836 16828 3892 16884
rect 3948 15986 4004 15988
rect 3948 15934 3950 15986
rect 3950 15934 4002 15986
rect 4002 15934 4004 15986
rect 3948 15932 4004 15934
rect 3612 15820 3668 15876
rect 7532 25506 7588 25508
rect 7532 25454 7534 25506
rect 7534 25454 7586 25506
rect 7586 25454 7588 25506
rect 7532 25452 7588 25454
rect 7644 25394 7700 25396
rect 7644 25342 7646 25394
rect 7646 25342 7698 25394
rect 7698 25342 7700 25394
rect 7644 25340 7700 25342
rect 7532 24892 7588 24948
rect 8204 26290 8260 26292
rect 8204 26238 8206 26290
rect 8206 26238 8258 26290
rect 8258 26238 8260 26290
rect 8204 26236 8260 26238
rect 9660 26908 9716 26964
rect 9100 25900 9156 25956
rect 9324 26348 9380 26404
rect 7868 25506 7924 25508
rect 7868 25454 7870 25506
rect 7870 25454 7922 25506
rect 7922 25454 7924 25506
rect 7868 25452 7924 25454
rect 8876 25506 8932 25508
rect 8876 25454 8878 25506
rect 8878 25454 8930 25506
rect 8930 25454 8932 25506
rect 8876 25452 8932 25454
rect 8428 25394 8484 25396
rect 8428 25342 8430 25394
rect 8430 25342 8482 25394
rect 8482 25342 8484 25394
rect 8428 25340 8484 25342
rect 8092 25228 8148 25284
rect 6972 23996 7028 24052
rect 6860 23938 6916 23940
rect 6860 23886 6862 23938
rect 6862 23886 6914 23938
rect 6914 23886 6916 23938
rect 6860 23884 6916 23886
rect 6972 23714 7028 23716
rect 6972 23662 6974 23714
rect 6974 23662 7026 23714
rect 7026 23662 7028 23714
rect 6972 23660 7028 23662
rect 7196 23714 7252 23716
rect 7196 23662 7198 23714
rect 7198 23662 7250 23714
rect 7250 23662 7252 23714
rect 7196 23660 7252 23662
rect 9548 25228 9604 25284
rect 9436 25116 9492 25172
rect 8092 24892 8148 24948
rect 9100 24722 9156 24724
rect 9100 24670 9102 24722
rect 9102 24670 9154 24722
rect 9154 24670 9156 24722
rect 9100 24668 9156 24670
rect 8316 24444 8372 24500
rect 8204 23938 8260 23940
rect 8204 23886 8206 23938
rect 8206 23886 8258 23938
rect 8258 23886 8260 23938
rect 8204 23884 8260 23886
rect 8092 23660 8148 23716
rect 6636 22876 6692 22932
rect 7308 23548 7364 23604
rect 7756 23548 7812 23604
rect 6860 23266 6916 23268
rect 6860 23214 6862 23266
rect 6862 23214 6914 23266
rect 6914 23214 6916 23266
rect 6860 23212 6916 23214
rect 7084 23154 7140 23156
rect 7084 23102 7086 23154
rect 7086 23102 7138 23154
rect 7138 23102 7140 23154
rect 7084 23100 7140 23102
rect 6524 21532 6580 21588
rect 6188 20802 6244 20804
rect 6188 20750 6190 20802
rect 6190 20750 6242 20802
rect 6242 20750 6244 20802
rect 6188 20748 6244 20750
rect 6412 20972 6468 21028
rect 6300 20076 6356 20132
rect 8876 23826 8932 23828
rect 8876 23774 8878 23826
rect 8878 23774 8930 23826
rect 8930 23774 8932 23826
rect 8876 23772 8932 23774
rect 8540 23548 8596 23604
rect 7084 22316 7140 22372
rect 7196 21532 7252 21588
rect 7196 21026 7252 21028
rect 7196 20974 7198 21026
rect 7198 20974 7250 21026
rect 7250 20974 7252 21026
rect 7196 20972 7252 20974
rect 6972 20802 7028 20804
rect 6972 20750 6974 20802
rect 6974 20750 7026 20802
rect 7026 20750 7028 20802
rect 6972 20748 7028 20750
rect 6860 20188 6916 20244
rect 7420 20300 7476 20356
rect 7196 20130 7252 20132
rect 7196 20078 7198 20130
rect 7198 20078 7250 20130
rect 7250 20078 7252 20130
rect 7196 20076 7252 20078
rect 6076 19404 6132 19460
rect 6300 19852 6356 19908
rect 5964 19292 6020 19348
rect 5740 19122 5796 19124
rect 5740 19070 5742 19122
rect 5742 19070 5794 19122
rect 5794 19070 5796 19122
rect 5740 19068 5796 19070
rect 5516 18508 5572 18564
rect 5852 18620 5908 18676
rect 5852 18450 5908 18452
rect 5852 18398 5854 18450
rect 5854 18398 5906 18450
rect 5906 18398 5908 18450
rect 5852 18396 5908 18398
rect 5740 17778 5796 17780
rect 5740 17726 5742 17778
rect 5742 17726 5794 17778
rect 5794 17726 5796 17778
rect 5740 17724 5796 17726
rect 5180 17612 5236 17668
rect 4508 16940 4564 16996
rect 4620 16770 4676 16772
rect 4620 16718 4622 16770
rect 4622 16718 4674 16770
rect 4674 16718 4676 16770
rect 4620 16716 4676 16718
rect 4172 16156 4228 16212
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 4508 16098 4564 16100
rect 4508 16046 4510 16098
rect 4510 16046 4562 16098
rect 4562 16046 4564 16098
rect 4508 16044 4564 16046
rect 4732 15986 4788 15988
rect 4732 15934 4734 15986
rect 4734 15934 4786 15986
rect 4786 15934 4788 15986
rect 4732 15932 4788 15934
rect 4060 15708 4116 15764
rect 4284 15820 4340 15876
rect 3836 15036 3892 15092
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 3612 13970 3668 13972
rect 3612 13918 3614 13970
rect 3614 13918 3666 13970
rect 3666 13918 3668 13970
rect 3612 13916 3668 13918
rect 4060 13634 4116 13636
rect 4060 13582 4062 13634
rect 4062 13582 4114 13634
rect 4114 13582 4116 13634
rect 4060 13580 4116 13582
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 5292 16994 5348 16996
rect 5292 16942 5294 16994
rect 5294 16942 5346 16994
rect 5346 16942 5348 16994
rect 5292 16940 5348 16942
rect 4956 15538 5012 15540
rect 4956 15486 4958 15538
rect 4958 15486 5010 15538
rect 5010 15486 5012 15538
rect 4956 15484 5012 15486
rect 4956 14642 5012 14644
rect 4956 14590 4958 14642
rect 4958 14590 5010 14642
rect 5010 14590 5012 14642
rect 4956 14588 5012 14590
rect 4844 12908 4900 12964
rect 3612 12850 3668 12852
rect 3612 12798 3614 12850
rect 3614 12798 3666 12850
rect 3666 12798 3668 12850
rect 3612 12796 3668 12798
rect 2492 12178 2548 12180
rect 2492 12126 2494 12178
rect 2494 12126 2546 12178
rect 2546 12126 2548 12178
rect 2492 12124 2548 12126
rect 1708 11452 1764 11508
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 2940 11452 2996 11508
rect 1260 11228 1316 11284
rect 2044 11282 2100 11284
rect 2044 11230 2046 11282
rect 2046 11230 2098 11282
rect 2098 11230 2100 11282
rect 2044 11228 2100 11230
rect 1708 10780 1764 10836
rect 2044 10892 2100 10948
rect 2492 10780 2548 10836
rect 5628 16716 5684 16772
rect 5628 16098 5684 16100
rect 5628 16046 5630 16098
rect 5630 16046 5682 16098
rect 5682 16046 5684 16098
rect 5628 16044 5684 16046
rect 6076 19234 6132 19236
rect 6076 19182 6078 19234
rect 6078 19182 6130 19234
rect 6130 19182 6132 19234
rect 6076 19180 6132 19182
rect 7532 19852 7588 19908
rect 6860 19234 6916 19236
rect 6860 19182 6862 19234
rect 6862 19182 6914 19234
rect 6914 19182 6916 19234
rect 6860 19180 6916 19182
rect 8204 23154 8260 23156
rect 8204 23102 8206 23154
rect 8206 23102 8258 23154
rect 8258 23102 8260 23154
rect 8204 23100 8260 23102
rect 8652 23154 8708 23156
rect 8652 23102 8654 23154
rect 8654 23102 8706 23154
rect 8706 23102 8708 23154
rect 8652 23100 8708 23102
rect 8764 22930 8820 22932
rect 8764 22878 8766 22930
rect 8766 22878 8818 22930
rect 8818 22878 8820 22930
rect 8764 22876 8820 22878
rect 7868 20802 7924 20804
rect 7868 20750 7870 20802
rect 7870 20750 7922 20802
rect 7922 20750 7924 20802
rect 7868 20748 7924 20750
rect 8092 20412 8148 20468
rect 8204 20524 8260 20580
rect 8540 20748 8596 20804
rect 6300 18338 6356 18340
rect 6300 18286 6302 18338
rect 6302 18286 6354 18338
rect 6354 18286 6356 18338
rect 6300 18284 6356 18286
rect 6972 17948 7028 18004
rect 6748 17276 6804 17332
rect 6300 17106 6356 17108
rect 6300 17054 6302 17106
rect 6302 17054 6354 17106
rect 6354 17054 6356 17106
rect 6300 17052 6356 17054
rect 7756 18450 7812 18452
rect 7756 18398 7758 18450
rect 7758 18398 7810 18450
rect 7810 18398 7812 18450
rect 7756 18396 7812 18398
rect 7644 17948 7700 18004
rect 7756 17388 7812 17444
rect 6972 16322 7028 16324
rect 6972 16270 6974 16322
rect 6974 16270 7026 16322
rect 7026 16270 7028 16322
rect 6972 16268 7028 16270
rect 5180 15484 5236 15540
rect 5516 15202 5572 15204
rect 5516 15150 5518 15202
rect 5518 15150 5570 15202
rect 5570 15150 5572 15202
rect 5516 15148 5572 15150
rect 5180 12178 5236 12180
rect 5180 12126 5182 12178
rect 5182 12126 5234 12178
rect 5234 12126 5236 12178
rect 5180 12124 5236 12126
rect 5964 15820 6020 15876
rect 6636 16098 6692 16100
rect 6636 16046 6638 16098
rect 6638 16046 6690 16098
rect 6690 16046 6692 16098
rect 6636 16044 6692 16046
rect 5964 15484 6020 15540
rect 6076 14812 6132 14868
rect 6524 15820 6580 15876
rect 6636 15148 6692 15204
rect 7420 16156 7476 16212
rect 7196 15874 7252 15876
rect 7196 15822 7198 15874
rect 7198 15822 7250 15874
rect 7250 15822 7252 15874
rect 7196 15820 7252 15822
rect 7980 16098 8036 16100
rect 7980 16046 7982 16098
rect 7982 16046 8034 16098
rect 8034 16046 8036 16098
rect 7980 16044 8036 16046
rect 8764 20578 8820 20580
rect 8764 20526 8766 20578
rect 8766 20526 8818 20578
rect 8818 20526 8820 20578
rect 8764 20524 8820 20526
rect 8988 22594 9044 22596
rect 8988 22542 8990 22594
rect 8990 22542 9042 22594
rect 9042 22542 9044 22594
rect 8988 22540 9044 22542
rect 14588 28700 14644 28756
rect 15148 29484 15204 29540
rect 16940 31724 16996 31780
rect 17052 31276 17108 31332
rect 16828 29484 16884 29540
rect 15596 29426 15652 29428
rect 15596 29374 15598 29426
rect 15598 29374 15650 29426
rect 15650 29374 15652 29426
rect 15596 29372 15652 29374
rect 15932 29314 15988 29316
rect 15932 29262 15934 29314
rect 15934 29262 15986 29314
rect 15986 29262 15988 29314
rect 15932 29260 15988 29262
rect 15148 28924 15204 28980
rect 15596 28754 15652 28756
rect 15596 28702 15598 28754
rect 15598 28702 15650 28754
rect 15650 28702 15652 28754
rect 15596 28700 15652 28702
rect 16268 28588 16324 28644
rect 17052 28642 17108 28644
rect 17052 28590 17054 28642
rect 17054 28590 17106 28642
rect 17106 28590 17108 28642
rect 17052 28588 17108 28590
rect 17724 35138 17780 35140
rect 17724 35086 17726 35138
rect 17726 35086 17778 35138
rect 17778 35086 17780 35138
rect 17724 35084 17780 35086
rect 19180 35810 19236 35812
rect 19180 35758 19182 35810
rect 19182 35758 19234 35810
rect 19234 35758 19236 35810
rect 19180 35756 19236 35758
rect 20748 37212 20804 37268
rect 20188 36316 20244 36372
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 21532 38834 21588 38836
rect 21532 38782 21534 38834
rect 21534 38782 21586 38834
rect 21586 38782 21588 38834
rect 21532 38780 21588 38782
rect 22428 38834 22484 38836
rect 22428 38782 22430 38834
rect 22430 38782 22482 38834
rect 22482 38782 22484 38834
rect 22428 38780 22484 38782
rect 22204 38722 22260 38724
rect 22204 38670 22206 38722
rect 22206 38670 22258 38722
rect 22258 38670 22260 38722
rect 22204 38668 22260 38670
rect 21196 37324 21252 37380
rect 21532 37266 21588 37268
rect 21532 37214 21534 37266
rect 21534 37214 21586 37266
rect 21586 37214 21588 37266
rect 21532 37212 21588 37214
rect 22764 38610 22820 38612
rect 22764 38558 22766 38610
rect 22766 38558 22818 38610
rect 22818 38558 22820 38610
rect 22764 38556 22820 38558
rect 23100 41970 23156 41972
rect 23100 41918 23102 41970
rect 23102 41918 23154 41970
rect 23154 41918 23156 41970
rect 23100 41916 23156 41918
rect 23324 41468 23380 41524
rect 24332 45276 24388 45332
rect 23884 42700 23940 42756
rect 24220 43596 24276 43652
rect 23772 40908 23828 40964
rect 23324 38556 23380 38612
rect 22876 36988 22932 37044
rect 21644 36258 21700 36260
rect 21644 36206 21646 36258
rect 21646 36206 21698 36258
rect 21698 36206 21700 36258
rect 21644 36204 21700 36206
rect 19068 35138 19124 35140
rect 19068 35086 19070 35138
rect 19070 35086 19122 35138
rect 19122 35086 19124 35138
rect 19068 35084 19124 35086
rect 19292 34972 19348 35028
rect 20188 35026 20244 35028
rect 20188 34974 20190 35026
rect 20190 34974 20242 35026
rect 20242 34974 20244 35026
rect 20188 34972 20244 34974
rect 20412 34972 20468 35028
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19740 34242 19796 34244
rect 19740 34190 19742 34242
rect 19742 34190 19794 34242
rect 19794 34190 19796 34242
rect 19740 34188 19796 34190
rect 17612 34018 17668 34020
rect 17612 33966 17614 34018
rect 17614 33966 17666 34018
rect 17666 33966 17668 34018
rect 17612 33964 17668 33966
rect 19180 33964 19236 34020
rect 17724 33404 17780 33460
rect 17388 32956 17444 33012
rect 19852 33964 19908 34020
rect 19516 33628 19572 33684
rect 20076 33404 20132 33460
rect 20412 34130 20468 34132
rect 20412 34078 20414 34130
rect 20414 34078 20466 34130
rect 20466 34078 20468 34130
rect 20412 34076 20468 34078
rect 17836 33068 17892 33124
rect 18732 33068 18788 33124
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 19180 32732 19236 32788
rect 17500 31836 17556 31892
rect 17388 31388 17444 31444
rect 17724 31052 17780 31108
rect 19180 31724 19236 31780
rect 18172 31666 18228 31668
rect 18172 31614 18174 31666
rect 18174 31614 18226 31666
rect 18226 31614 18228 31666
rect 18172 31612 18228 31614
rect 18732 31666 18788 31668
rect 18732 31614 18734 31666
rect 18734 31614 18786 31666
rect 18786 31614 18788 31666
rect 18732 31612 18788 31614
rect 17948 31276 18004 31332
rect 17948 31052 18004 31108
rect 17836 30716 17892 30772
rect 17388 30380 17444 30436
rect 17948 29484 18004 29540
rect 17388 28924 17444 28980
rect 20636 33180 20692 33236
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 20860 34242 20916 34244
rect 20860 34190 20862 34242
rect 20862 34190 20914 34242
rect 20914 34190 20916 34242
rect 20860 34188 20916 34190
rect 21084 33628 21140 33684
rect 20860 33180 20916 33236
rect 21868 35026 21924 35028
rect 21868 34974 21870 35026
rect 21870 34974 21922 35026
rect 21922 34974 21924 35026
rect 21868 34972 21924 34974
rect 21420 34076 21476 34132
rect 21756 34300 21812 34356
rect 21532 33516 21588 33572
rect 21420 33404 21476 33460
rect 20748 31388 20804 31444
rect 20188 30994 20244 30996
rect 20188 30942 20190 30994
rect 20190 30942 20242 30994
rect 20242 30942 20244 30994
rect 20188 30940 20244 30942
rect 20636 31164 20692 31220
rect 18284 30044 18340 30100
rect 20076 30828 20132 30884
rect 19404 30434 19460 30436
rect 19404 30382 19406 30434
rect 19406 30382 19458 30434
rect 19458 30382 19460 30434
rect 19404 30380 19460 30382
rect 19068 30098 19124 30100
rect 19068 30046 19070 30098
rect 19070 30046 19122 30098
rect 19122 30046 19124 30098
rect 19068 30044 19124 30046
rect 20748 30716 20804 30772
rect 21756 33346 21812 33348
rect 21756 33294 21758 33346
rect 21758 33294 21810 33346
rect 21810 33294 21812 33346
rect 21756 33292 21812 33294
rect 21756 32450 21812 32452
rect 21756 32398 21758 32450
rect 21758 32398 21810 32450
rect 21810 32398 21812 32450
rect 21756 32396 21812 32398
rect 23100 36876 23156 36932
rect 23100 36258 23156 36260
rect 23100 36206 23102 36258
rect 23102 36206 23154 36258
rect 23154 36206 23156 36258
rect 23100 36204 23156 36206
rect 22988 35756 23044 35812
rect 22988 33292 23044 33348
rect 23100 33740 23156 33796
rect 22876 33180 22932 33236
rect 22204 31890 22260 31892
rect 22204 31838 22206 31890
rect 22206 31838 22258 31890
rect 22258 31838 22260 31890
rect 22204 31836 22260 31838
rect 22764 32396 22820 32452
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 20076 29650 20132 29652
rect 20076 29598 20078 29650
rect 20078 29598 20130 29650
rect 20130 29598 20132 29650
rect 20076 29596 20132 29598
rect 20860 30156 20916 30212
rect 22988 31724 23044 31780
rect 24780 51490 24836 51492
rect 24780 51438 24782 51490
rect 24782 51438 24834 51490
rect 24834 51438 24836 51490
rect 24780 51436 24836 51438
rect 24892 48748 24948 48804
rect 24780 45052 24836 45108
rect 24444 40402 24500 40404
rect 24444 40350 24446 40402
rect 24446 40350 24498 40402
rect 24498 40350 24500 40402
rect 24444 40348 24500 40350
rect 23996 39618 24052 39620
rect 23996 39566 23998 39618
rect 23998 39566 24050 39618
rect 24050 39566 24052 39618
rect 23996 39564 24052 39566
rect 23884 39004 23940 39060
rect 23548 38780 23604 38836
rect 24220 38946 24276 38948
rect 24220 38894 24222 38946
rect 24222 38894 24274 38946
rect 24274 38894 24276 38946
rect 24220 38892 24276 38894
rect 23884 37266 23940 37268
rect 23884 37214 23886 37266
rect 23886 37214 23938 37266
rect 23938 37214 23940 37266
rect 23884 37212 23940 37214
rect 24668 43484 24724 43540
rect 24556 39004 24612 39060
rect 25340 52834 25396 52836
rect 25340 52782 25342 52834
rect 25342 52782 25394 52834
rect 25394 52782 25396 52834
rect 25340 52780 25396 52782
rect 26012 52332 26068 52388
rect 26460 52332 26516 52388
rect 26348 52108 26404 52164
rect 25564 51490 25620 51492
rect 25564 51438 25566 51490
rect 25566 51438 25618 51490
rect 25618 51438 25620 51490
rect 25564 51436 25620 51438
rect 25564 51154 25620 51156
rect 25564 51102 25566 51154
rect 25566 51102 25618 51154
rect 25618 51102 25620 51154
rect 25564 51100 25620 51102
rect 26012 50652 26068 50708
rect 25676 50594 25732 50596
rect 25676 50542 25678 50594
rect 25678 50542 25730 50594
rect 25730 50542 25732 50594
rect 25676 50540 25732 50542
rect 25788 50482 25844 50484
rect 25788 50430 25790 50482
rect 25790 50430 25842 50482
rect 25842 50430 25844 50482
rect 25788 50428 25844 50430
rect 27020 52050 27076 52052
rect 27020 51998 27022 52050
rect 27022 51998 27074 52050
rect 27074 51998 27076 52050
rect 27020 51996 27076 51998
rect 27020 51100 27076 51156
rect 28588 55970 28644 55972
rect 28588 55918 28590 55970
rect 28590 55918 28642 55970
rect 28642 55918 28644 55970
rect 28588 55916 28644 55918
rect 28924 55468 28980 55524
rect 28140 55410 28196 55412
rect 28140 55358 28142 55410
rect 28142 55358 28194 55410
rect 28194 55358 28196 55410
rect 28140 55356 28196 55358
rect 28476 55244 28532 55300
rect 29148 54796 29204 54852
rect 28476 54626 28532 54628
rect 28476 54574 28478 54626
rect 28478 54574 28530 54626
rect 28530 54574 28532 54626
rect 28476 54572 28532 54574
rect 27692 53116 27748 53172
rect 27356 51436 27412 51492
rect 26460 50092 26516 50148
rect 25788 49756 25844 49812
rect 25900 49698 25956 49700
rect 25900 49646 25902 49698
rect 25902 49646 25954 49698
rect 25954 49646 25956 49698
rect 25900 49644 25956 49646
rect 26796 49644 26852 49700
rect 25676 48412 25732 48468
rect 26012 48748 26068 48804
rect 25676 48188 25732 48244
rect 25788 48018 25844 48020
rect 25788 47966 25790 48018
rect 25790 47966 25842 48018
rect 25842 47966 25844 48018
rect 25788 47964 25844 47966
rect 25900 47628 25956 47684
rect 25116 43708 25172 43764
rect 25340 43650 25396 43652
rect 25340 43598 25342 43650
rect 25342 43598 25394 43650
rect 25394 43598 25396 43650
rect 25340 43596 25396 43598
rect 25228 43538 25284 43540
rect 25228 43486 25230 43538
rect 25230 43486 25282 43538
rect 25282 43486 25284 43538
rect 25228 43484 25284 43486
rect 26236 48242 26292 48244
rect 26236 48190 26238 48242
rect 26238 48190 26290 48242
rect 26290 48190 26292 48242
rect 26236 48188 26292 48190
rect 26236 47628 26292 47684
rect 26124 46674 26180 46676
rect 26124 46622 26126 46674
rect 26126 46622 26178 46674
rect 26178 46622 26180 46674
rect 26124 46620 26180 46622
rect 26796 48524 26852 48580
rect 27020 47964 27076 48020
rect 27244 49810 27300 49812
rect 27244 49758 27246 49810
rect 27246 49758 27298 49810
rect 27298 49758 27300 49810
rect 27244 49756 27300 49758
rect 27244 48860 27300 48916
rect 26908 46674 26964 46676
rect 26908 46622 26910 46674
rect 26910 46622 26962 46674
rect 26962 46622 26964 46674
rect 26908 46620 26964 46622
rect 25564 43148 25620 43204
rect 26124 45612 26180 45668
rect 27020 46396 27076 46452
rect 26572 45218 26628 45220
rect 26572 45166 26574 45218
rect 26574 45166 26626 45218
rect 26626 45166 26628 45218
rect 26572 45164 26628 45166
rect 26572 44098 26628 44100
rect 26572 44046 26574 44098
rect 26574 44046 26626 44098
rect 26626 44046 26628 44098
rect 26572 44044 26628 44046
rect 27244 45666 27300 45668
rect 27244 45614 27246 45666
rect 27246 45614 27298 45666
rect 27298 45614 27300 45666
rect 27244 45612 27300 45614
rect 28812 53676 28868 53732
rect 27916 50092 27972 50148
rect 28588 49698 28644 49700
rect 28588 49646 28590 49698
rect 28590 49646 28642 49698
rect 28642 49646 28644 49698
rect 28588 49644 28644 49646
rect 27916 48972 27972 49028
rect 28588 49026 28644 49028
rect 28588 48974 28590 49026
rect 28590 48974 28642 49026
rect 28642 48974 28644 49026
rect 28588 48972 28644 48974
rect 28476 48914 28532 48916
rect 28476 48862 28478 48914
rect 28478 48862 28530 48914
rect 28530 48862 28532 48914
rect 28476 48860 28532 48862
rect 27804 46284 27860 46340
rect 27132 45164 27188 45220
rect 26796 45106 26852 45108
rect 26796 45054 26798 45106
rect 26798 45054 26850 45106
rect 26850 45054 26852 45106
rect 26796 45052 26852 45054
rect 26796 43484 26852 43540
rect 25788 42924 25844 42980
rect 25116 40348 25172 40404
rect 25340 42754 25396 42756
rect 25340 42702 25342 42754
rect 25342 42702 25394 42754
rect 25394 42702 25396 42754
rect 25340 42700 25396 42702
rect 26348 43314 26404 43316
rect 26348 43262 26350 43314
rect 26350 43262 26402 43314
rect 26402 43262 26404 43314
rect 26348 43260 26404 43262
rect 26124 43148 26180 43204
rect 26124 42924 26180 42980
rect 26908 43260 26964 43316
rect 25676 41858 25732 41860
rect 25676 41806 25678 41858
rect 25678 41806 25730 41858
rect 25730 41806 25732 41858
rect 25676 41804 25732 41806
rect 26796 42476 26852 42532
rect 25340 40962 25396 40964
rect 25340 40910 25342 40962
rect 25342 40910 25394 40962
rect 25394 40910 25396 40962
rect 25340 40908 25396 40910
rect 26012 40908 26068 40964
rect 25900 40796 25956 40852
rect 25564 40402 25620 40404
rect 25564 40350 25566 40402
rect 25566 40350 25618 40402
rect 25618 40350 25620 40402
rect 25564 40348 25620 40350
rect 25228 39394 25284 39396
rect 25228 39342 25230 39394
rect 25230 39342 25282 39394
rect 25282 39342 25284 39394
rect 25228 39340 25284 39342
rect 25004 38892 25060 38948
rect 24556 37548 24612 37604
rect 24108 36316 24164 36372
rect 25116 38274 25172 38276
rect 25116 38222 25118 38274
rect 25118 38222 25170 38274
rect 25170 38222 25172 38274
rect 25116 38220 25172 38222
rect 24332 36988 24388 37044
rect 25116 37996 25172 38052
rect 25004 37548 25060 37604
rect 23212 33628 23268 33684
rect 23436 35586 23492 35588
rect 23436 35534 23438 35586
rect 23438 35534 23490 35586
rect 23490 35534 23492 35586
rect 23436 35532 23492 35534
rect 23660 35810 23716 35812
rect 23660 35758 23662 35810
rect 23662 35758 23714 35810
rect 23714 35758 23716 35810
rect 23660 35756 23716 35758
rect 25340 38946 25396 38948
rect 25340 38894 25342 38946
rect 25342 38894 25394 38946
rect 25394 38894 25396 38946
rect 25340 38892 25396 38894
rect 26460 40796 26516 40852
rect 25900 39900 25956 39956
rect 25900 39340 25956 39396
rect 26460 39452 26516 39508
rect 25564 38444 25620 38500
rect 25340 38332 25396 38388
rect 25452 38050 25508 38052
rect 25452 37998 25454 38050
rect 25454 37998 25506 38050
rect 25506 37998 25508 38050
rect 25452 37996 25508 37998
rect 25676 38050 25732 38052
rect 25676 37998 25678 38050
rect 25678 37998 25730 38050
rect 25730 37998 25732 38050
rect 25676 37996 25732 37998
rect 25676 37660 25732 37716
rect 23996 34914 24052 34916
rect 23996 34862 23998 34914
rect 23998 34862 24050 34914
rect 24050 34862 24052 34914
rect 23996 34860 24052 34862
rect 24556 35196 24612 35252
rect 25340 35586 25396 35588
rect 25340 35534 25342 35586
rect 25342 35534 25394 35586
rect 25394 35534 25396 35586
rect 25340 35532 25396 35534
rect 24444 34690 24500 34692
rect 24444 34638 24446 34690
rect 24446 34638 24498 34690
rect 24498 34638 24500 34690
rect 24444 34636 24500 34638
rect 23548 34076 23604 34132
rect 23436 32732 23492 32788
rect 24332 34300 24388 34356
rect 24556 34130 24612 34132
rect 24556 34078 24558 34130
rect 24558 34078 24610 34130
rect 24610 34078 24612 34130
rect 24556 34076 24612 34078
rect 23884 34018 23940 34020
rect 23884 33966 23886 34018
rect 23886 33966 23938 34018
rect 23938 33966 23940 34018
rect 23884 33964 23940 33966
rect 23996 32956 24052 33012
rect 20300 29538 20356 29540
rect 20300 29486 20302 29538
rect 20302 29486 20354 29538
rect 20354 29486 20356 29538
rect 20300 29484 20356 29486
rect 20412 29932 20468 29988
rect 17276 28252 17332 28308
rect 18060 28252 18116 28308
rect 16380 28028 16436 28084
rect 17948 28028 18004 28084
rect 17612 27970 17668 27972
rect 17612 27918 17614 27970
rect 17614 27918 17666 27970
rect 17666 27918 17668 27970
rect 17612 27916 17668 27918
rect 16604 27132 16660 27188
rect 17276 27186 17332 27188
rect 17276 27134 17278 27186
rect 17278 27134 17330 27186
rect 17330 27134 17332 27186
rect 17276 27132 17332 27134
rect 19628 29148 19684 29204
rect 19068 28812 19124 28868
rect 18172 28140 18228 28196
rect 18508 28140 18564 28196
rect 19068 27970 19124 27972
rect 19068 27918 19070 27970
rect 19070 27918 19122 27970
rect 19122 27918 19124 27970
rect 19068 27916 19124 27918
rect 18060 27692 18116 27748
rect 9996 26684 10052 26740
rect 15148 26796 15204 26852
rect 12684 26514 12740 26516
rect 12684 26462 12686 26514
rect 12686 26462 12738 26514
rect 12738 26462 12740 26514
rect 12684 26460 12740 26462
rect 14364 26460 14420 26516
rect 9884 26348 9940 26404
rect 11116 26348 11172 26404
rect 10108 26290 10164 26292
rect 10108 26238 10110 26290
rect 10110 26238 10162 26290
rect 10162 26238 10164 26290
rect 10108 26236 10164 26238
rect 11564 26290 11620 26292
rect 11564 26238 11566 26290
rect 11566 26238 11618 26290
rect 11618 26238 11620 26290
rect 11564 26236 11620 26238
rect 12348 26290 12404 26292
rect 12348 26238 12350 26290
rect 12350 26238 12402 26290
rect 12402 26238 12404 26290
rect 12348 26236 12404 26238
rect 13804 26402 13860 26404
rect 13804 26350 13806 26402
rect 13806 26350 13858 26402
rect 13858 26350 13860 26402
rect 13804 26348 13860 26350
rect 14028 26402 14084 26404
rect 14028 26350 14030 26402
rect 14030 26350 14082 26402
rect 14082 26350 14084 26402
rect 14028 26348 14084 26350
rect 13132 26290 13188 26292
rect 13132 26238 13134 26290
rect 13134 26238 13186 26290
rect 13186 26238 13188 26290
rect 13132 26236 13188 26238
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 20188 27858 20244 27860
rect 20188 27806 20190 27858
rect 20190 27806 20242 27858
rect 20242 27806 20244 27858
rect 20188 27804 20244 27806
rect 19964 27634 20020 27636
rect 19964 27582 19966 27634
rect 19966 27582 20018 27634
rect 20018 27582 20020 27634
rect 19964 27580 20020 27582
rect 20188 27356 20244 27412
rect 18620 26962 18676 26964
rect 18620 26910 18622 26962
rect 18622 26910 18674 26962
rect 18674 26910 18676 26962
rect 18620 26908 18676 26910
rect 11452 25900 11508 25956
rect 12684 25900 12740 25956
rect 9996 25506 10052 25508
rect 9996 25454 9998 25506
rect 9998 25454 10050 25506
rect 10050 25454 10052 25506
rect 9996 25452 10052 25454
rect 9772 25340 9828 25396
rect 9772 24722 9828 24724
rect 9772 24670 9774 24722
rect 9774 24670 9826 24722
rect 9826 24670 9828 24722
rect 9772 24668 9828 24670
rect 10668 25394 10724 25396
rect 10668 25342 10670 25394
rect 10670 25342 10722 25394
rect 10722 25342 10724 25394
rect 10668 25340 10724 25342
rect 11004 25282 11060 25284
rect 11004 25230 11006 25282
rect 11006 25230 11058 25282
rect 11058 25230 11060 25282
rect 11004 25228 11060 25230
rect 10108 23436 10164 23492
rect 10108 22540 10164 22596
rect 10444 23714 10500 23716
rect 10444 23662 10446 23714
rect 10446 23662 10498 23714
rect 10498 23662 10500 23714
rect 10444 23660 10500 23662
rect 10780 24556 10836 24612
rect 11564 25116 11620 25172
rect 10780 24050 10836 24052
rect 10780 23998 10782 24050
rect 10782 23998 10834 24050
rect 10834 23998 10836 24050
rect 10780 23996 10836 23998
rect 11564 23996 11620 24052
rect 11228 23100 11284 23156
rect 11340 23660 11396 23716
rect 11788 23884 11844 23940
rect 11676 23548 11732 23604
rect 11676 23378 11732 23380
rect 11676 23326 11678 23378
rect 11678 23326 11730 23378
rect 11730 23326 11732 23378
rect 11676 23324 11732 23326
rect 10668 22370 10724 22372
rect 10668 22318 10670 22370
rect 10670 22318 10722 22370
rect 10722 22318 10724 22370
rect 10668 22316 10724 22318
rect 10444 21532 10500 21588
rect 9324 20802 9380 20804
rect 9324 20750 9326 20802
rect 9326 20750 9378 20802
rect 9378 20750 9380 20802
rect 9324 20748 9380 20750
rect 8988 20690 9044 20692
rect 8988 20638 8990 20690
rect 8990 20638 9042 20690
rect 9042 20638 9044 20690
rect 8988 20636 9044 20638
rect 8876 20412 8932 20468
rect 9772 20690 9828 20692
rect 9772 20638 9774 20690
rect 9774 20638 9826 20690
rect 9826 20638 9828 20690
rect 9772 20636 9828 20638
rect 9884 20578 9940 20580
rect 9884 20526 9886 20578
rect 9886 20526 9938 20578
rect 9938 20526 9940 20578
rect 9884 20524 9940 20526
rect 8540 19852 8596 19908
rect 9100 19964 9156 20020
rect 8316 19234 8372 19236
rect 8316 19182 8318 19234
rect 8318 19182 8370 19234
rect 8370 19182 8372 19234
rect 8316 19180 8372 19182
rect 8764 19068 8820 19124
rect 8988 19180 9044 19236
rect 9436 17948 9492 18004
rect 8876 16268 8932 16324
rect 8652 16098 8708 16100
rect 8652 16046 8654 16098
rect 8654 16046 8706 16098
rect 8706 16046 8708 16098
rect 8652 16044 8708 16046
rect 6860 15484 6916 15540
rect 7532 15260 7588 15316
rect 7644 15708 7700 15764
rect 6524 14812 6580 14868
rect 6860 14812 6916 14868
rect 7756 15484 7812 15540
rect 7644 14700 7700 14756
rect 7308 14306 7364 14308
rect 7308 14254 7310 14306
rect 7310 14254 7362 14306
rect 7362 14254 7364 14306
rect 7308 14252 7364 14254
rect 9212 15372 9268 15428
rect 8092 14252 8148 14308
rect 8204 14028 8260 14084
rect 8316 13858 8372 13860
rect 8316 13806 8318 13858
rect 8318 13806 8370 13858
rect 8370 13806 8372 13858
rect 8316 13804 8372 13806
rect 5740 12962 5796 12964
rect 5740 12910 5742 12962
rect 5742 12910 5794 12962
rect 5794 12910 5796 12962
rect 5740 12908 5796 12910
rect 6300 13074 6356 13076
rect 6300 13022 6302 13074
rect 6302 13022 6354 13074
rect 6354 13022 6356 13074
rect 6300 13020 6356 13022
rect 6076 12908 6132 12964
rect 7420 13692 7476 13748
rect 6860 13020 6916 13076
rect 6748 12962 6804 12964
rect 6748 12910 6750 12962
rect 6750 12910 6802 12962
rect 6802 12910 6804 12962
rect 6748 12908 6804 12910
rect 6188 12178 6244 12180
rect 6188 12126 6190 12178
rect 6190 12126 6242 12178
rect 6242 12126 6244 12178
rect 6188 12124 6244 12126
rect 5964 12012 6020 12068
rect 5068 11228 5124 11284
rect 5740 11676 5796 11732
rect 6748 12066 6804 12068
rect 6748 12014 6750 12066
rect 6750 12014 6802 12066
rect 6802 12014 6804 12066
rect 6748 12012 6804 12014
rect 8540 15260 8596 15316
rect 8764 15202 8820 15204
rect 8764 15150 8766 15202
rect 8766 15150 8818 15202
rect 8818 15150 8820 15202
rect 8764 15148 8820 15150
rect 8540 13746 8596 13748
rect 8540 13694 8542 13746
rect 8542 13694 8594 13746
rect 8594 13694 8596 13746
rect 8540 13692 8596 13694
rect 8764 13692 8820 13748
rect 6972 12178 7028 12180
rect 6972 12126 6974 12178
rect 6974 12126 7026 12178
rect 7026 12126 7028 12178
rect 6972 12124 7028 12126
rect 6300 11394 6356 11396
rect 6300 11342 6302 11394
rect 6302 11342 6354 11394
rect 6354 11342 6356 11394
rect 6300 11340 6356 11342
rect 5740 11282 5796 11284
rect 5740 11230 5742 11282
rect 5742 11230 5794 11282
rect 5794 11230 5796 11282
rect 5740 11228 5796 11230
rect 6076 10780 6132 10836
rect 4844 10668 4900 10724
rect 6188 10722 6244 10724
rect 6188 10670 6190 10722
rect 6190 10670 6242 10722
rect 6242 10670 6244 10722
rect 6188 10668 6244 10670
rect 1708 10108 1764 10164
rect 2492 10108 2548 10164
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 5628 9266 5684 9268
rect 5628 9214 5630 9266
rect 5630 9214 5682 9266
rect 5682 9214 5684 9266
rect 5628 9212 5684 9214
rect 2044 9154 2100 9156
rect 2044 9102 2046 9154
rect 2046 9102 2098 9154
rect 2098 9102 2100 9154
rect 2044 9100 2100 9102
rect 6860 11506 6916 11508
rect 6860 11454 6862 11506
rect 6862 11454 6914 11506
rect 6914 11454 6916 11506
rect 6860 11452 6916 11454
rect 6972 11340 7028 11396
rect 6300 9212 6356 9268
rect 1708 8764 1764 8820
rect 2492 8764 2548 8820
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 6188 8428 6244 8484
rect 7308 11394 7364 11396
rect 7308 11342 7310 11394
rect 7310 11342 7362 11394
rect 7362 11342 7364 11394
rect 7308 11340 7364 11342
rect 10332 20412 10388 20468
rect 11228 21810 11284 21812
rect 11228 21758 11230 21810
rect 11230 21758 11282 21810
rect 11282 21758 11284 21810
rect 11228 21756 11284 21758
rect 11900 23100 11956 23156
rect 11228 21532 11284 21588
rect 11452 22316 11508 22372
rect 10668 20690 10724 20692
rect 10668 20638 10670 20690
rect 10670 20638 10722 20690
rect 10722 20638 10724 20690
rect 10668 20636 10724 20638
rect 11116 20690 11172 20692
rect 11116 20638 11118 20690
rect 11118 20638 11170 20690
rect 11170 20638 11172 20690
rect 11116 20636 11172 20638
rect 10444 20130 10500 20132
rect 10444 20078 10446 20130
rect 10446 20078 10498 20130
rect 10498 20078 10500 20130
rect 10444 20076 10500 20078
rect 10332 20018 10388 20020
rect 10332 19966 10334 20018
rect 10334 19966 10386 20018
rect 10386 19966 10388 20018
rect 10332 19964 10388 19966
rect 9772 19852 9828 19908
rect 9660 14476 9716 14532
rect 10108 17948 10164 18004
rect 10892 18562 10948 18564
rect 10892 18510 10894 18562
rect 10894 18510 10946 18562
rect 10946 18510 10948 18562
rect 10892 18508 10948 18510
rect 10780 16098 10836 16100
rect 10780 16046 10782 16098
rect 10782 16046 10834 16098
rect 10834 16046 10836 16098
rect 10780 16044 10836 16046
rect 11340 20076 11396 20132
rect 11564 21810 11620 21812
rect 11564 21758 11566 21810
rect 11566 21758 11618 21810
rect 11618 21758 11620 21810
rect 11564 21756 11620 21758
rect 12572 25116 12628 25172
rect 14140 26066 14196 26068
rect 14140 26014 14142 26066
rect 14142 26014 14194 26066
rect 14194 26014 14196 26066
rect 14140 26012 14196 26014
rect 14812 26012 14868 26068
rect 12908 25116 12964 25172
rect 13580 25004 13636 25060
rect 13468 24610 13524 24612
rect 13468 24558 13470 24610
rect 13470 24558 13522 24610
rect 13522 24558 13524 24610
rect 13468 24556 13524 24558
rect 12124 23548 12180 23604
rect 12908 24050 12964 24052
rect 12908 23998 12910 24050
rect 12910 23998 12962 24050
rect 12962 23998 12964 24050
rect 12908 23996 12964 23998
rect 13916 23996 13972 24052
rect 13468 23884 13524 23940
rect 12572 23324 12628 23380
rect 12236 22428 12292 22484
rect 12012 21810 12068 21812
rect 12012 21758 12014 21810
rect 12014 21758 12066 21810
rect 12066 21758 12068 21810
rect 12012 21756 12068 21758
rect 12124 21586 12180 21588
rect 12124 21534 12126 21586
rect 12126 21534 12178 21586
rect 12178 21534 12180 21586
rect 12124 21532 12180 21534
rect 13692 23772 13748 23828
rect 12684 23154 12740 23156
rect 12684 23102 12686 23154
rect 12686 23102 12738 23154
rect 12738 23102 12740 23154
rect 12684 23100 12740 23102
rect 13916 23714 13972 23716
rect 13916 23662 13918 23714
rect 13918 23662 13970 23714
rect 13970 23662 13972 23714
rect 13916 23660 13972 23662
rect 14700 25506 14756 25508
rect 14700 25454 14702 25506
rect 14702 25454 14754 25506
rect 14754 25454 14756 25506
rect 14700 25452 14756 25454
rect 15148 25282 15204 25284
rect 15148 25230 15150 25282
rect 15150 25230 15202 25282
rect 15202 25230 15204 25282
rect 15148 25228 15204 25230
rect 14140 25116 14196 25172
rect 15372 25282 15428 25284
rect 15372 25230 15374 25282
rect 15374 25230 15426 25282
rect 15426 25230 15428 25282
rect 15372 25228 15428 25230
rect 15708 25228 15764 25284
rect 15372 24780 15428 24836
rect 14924 23884 14980 23940
rect 14364 23826 14420 23828
rect 14364 23774 14366 23826
rect 14366 23774 14418 23826
rect 14418 23774 14420 23826
rect 14364 23772 14420 23774
rect 14476 23324 14532 23380
rect 15372 23436 15428 23492
rect 14812 23154 14868 23156
rect 14812 23102 14814 23154
rect 14814 23102 14866 23154
rect 14866 23102 14868 23154
rect 14812 23100 14868 23102
rect 12908 22594 12964 22596
rect 12908 22542 12910 22594
rect 12910 22542 12962 22594
rect 12962 22542 12964 22594
rect 12908 22540 12964 22542
rect 13804 22594 13860 22596
rect 13804 22542 13806 22594
rect 13806 22542 13858 22594
rect 13858 22542 13860 22594
rect 13804 22540 13860 22542
rect 15596 23938 15652 23940
rect 15596 23886 15598 23938
rect 15598 23886 15650 23938
rect 15650 23886 15652 23938
rect 15596 23884 15652 23886
rect 17164 24050 17220 24052
rect 17164 23998 17166 24050
rect 17166 23998 17218 24050
rect 17218 23998 17220 24050
rect 17164 23996 17220 23998
rect 15036 23100 15092 23156
rect 14812 22540 14868 22596
rect 12236 21308 12292 21364
rect 12572 21474 12628 21476
rect 12572 21422 12574 21474
rect 12574 21422 12626 21474
rect 12626 21422 12628 21474
rect 12572 21420 12628 21422
rect 11676 20690 11732 20692
rect 11676 20638 11678 20690
rect 11678 20638 11730 20690
rect 11730 20638 11732 20690
rect 11676 20636 11732 20638
rect 11564 19964 11620 20020
rect 11228 19068 11284 19124
rect 11900 20524 11956 20580
rect 11900 18620 11956 18676
rect 11676 15986 11732 15988
rect 11676 15934 11678 15986
rect 11678 15934 11730 15986
rect 11730 15934 11732 15986
rect 11676 15932 11732 15934
rect 11116 15708 11172 15764
rect 11676 15426 11732 15428
rect 11676 15374 11678 15426
rect 11678 15374 11730 15426
rect 11730 15374 11732 15426
rect 11676 15372 11732 15374
rect 12796 20690 12852 20692
rect 12796 20638 12798 20690
rect 12798 20638 12850 20690
rect 12850 20638 12852 20690
rect 12796 20636 12852 20638
rect 13580 21420 13636 21476
rect 14028 20636 14084 20692
rect 12124 18732 12180 18788
rect 12236 18508 12292 18564
rect 12012 18396 12068 18452
rect 11900 16044 11956 16100
rect 12124 17836 12180 17892
rect 12684 20076 12740 20132
rect 13132 20130 13188 20132
rect 13132 20078 13134 20130
rect 13134 20078 13186 20130
rect 13186 20078 13188 20130
rect 13132 20076 13188 20078
rect 12908 19180 12964 19236
rect 12572 18172 12628 18228
rect 12460 17388 12516 17444
rect 10556 15148 10612 15204
rect 10332 14418 10388 14420
rect 10332 14366 10334 14418
rect 10334 14366 10386 14418
rect 10386 14366 10388 14418
rect 10332 14364 10388 14366
rect 10780 14364 10836 14420
rect 10108 13804 10164 13860
rect 9436 13692 9492 13748
rect 9324 12850 9380 12852
rect 9324 12798 9326 12850
rect 9326 12798 9378 12850
rect 9378 12798 9380 12850
rect 9324 12796 9380 12798
rect 9884 13580 9940 13636
rect 8988 12124 9044 12180
rect 8428 11676 8484 11732
rect 8652 11506 8708 11508
rect 8652 11454 8654 11506
rect 8654 11454 8706 11506
rect 8706 11454 8708 11506
rect 8652 11452 8708 11454
rect 7532 11394 7588 11396
rect 7532 11342 7534 11394
rect 7534 11342 7586 11394
rect 7586 11342 7588 11394
rect 7532 11340 7588 11342
rect 7980 11282 8036 11284
rect 7980 11230 7982 11282
rect 7982 11230 8034 11282
rect 8034 11230 8036 11282
rect 7980 11228 8036 11230
rect 7644 10834 7700 10836
rect 7644 10782 7646 10834
rect 7646 10782 7698 10834
rect 7698 10782 7700 10834
rect 7644 10780 7700 10782
rect 6748 9212 6804 9268
rect 7084 9154 7140 9156
rect 7084 9102 7086 9154
rect 7086 9102 7138 9154
rect 7138 9102 7140 9154
rect 7084 9100 7140 9102
rect 6972 8204 7028 8260
rect 7644 9100 7700 9156
rect 7980 9212 8036 9268
rect 7644 8204 7700 8260
rect 9100 9212 9156 9268
rect 8652 9154 8708 9156
rect 8652 9102 8654 9154
rect 8654 9102 8706 9154
rect 8706 9102 8708 9154
rect 8652 9100 8708 9102
rect 8876 8988 8932 9044
rect 8316 8092 8372 8148
rect 8652 8316 8708 8372
rect 8764 8204 8820 8260
rect 8764 7698 8820 7700
rect 8764 7646 8766 7698
rect 8766 7646 8818 7698
rect 8818 7646 8820 7698
rect 8764 7644 8820 7646
rect 8988 7868 9044 7924
rect 9100 7196 9156 7252
rect 9212 8428 9268 8484
rect 9212 7980 9268 8036
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 9660 12012 9716 12068
rect 9772 11228 9828 11284
rect 9996 12124 10052 12180
rect 10220 12066 10276 12068
rect 10220 12014 10222 12066
rect 10222 12014 10274 12066
rect 10274 12014 10276 12066
rect 10220 12012 10276 12014
rect 14252 20076 14308 20132
rect 13468 19068 13524 19124
rect 14476 19404 14532 19460
rect 13468 18732 13524 18788
rect 13356 18396 13412 18452
rect 14476 19234 14532 19236
rect 14476 19182 14478 19234
rect 14478 19182 14530 19234
rect 14530 19182 14532 19234
rect 14476 19180 14532 19182
rect 15036 19122 15092 19124
rect 15036 19070 15038 19122
rect 15038 19070 15090 19122
rect 15090 19070 15092 19122
rect 15036 19068 15092 19070
rect 15260 19516 15316 19572
rect 15260 19292 15316 19348
rect 13132 17388 13188 17444
rect 13804 18450 13860 18452
rect 13804 18398 13806 18450
rect 13806 18398 13858 18450
rect 13858 18398 13860 18450
rect 13804 18396 13860 18398
rect 14588 18172 14644 18228
rect 15484 19068 15540 19124
rect 15372 18396 15428 18452
rect 15036 18338 15092 18340
rect 15036 18286 15038 18338
rect 15038 18286 15090 18338
rect 15090 18286 15092 18338
rect 15036 18284 15092 18286
rect 15484 18284 15540 18340
rect 13692 17836 13748 17892
rect 15148 18172 15204 18228
rect 14476 17724 14532 17780
rect 12796 16044 12852 16100
rect 12908 15260 12964 15316
rect 13244 16770 13300 16772
rect 13244 16718 13246 16770
rect 13246 16718 13298 16770
rect 13298 16718 13300 16770
rect 13244 16716 13300 16718
rect 14364 17388 14420 17444
rect 14140 16828 14196 16884
rect 13692 16098 13748 16100
rect 13692 16046 13694 16098
rect 13694 16046 13746 16098
rect 13746 16046 13748 16098
rect 13692 16044 13748 16046
rect 14028 15986 14084 15988
rect 14028 15934 14030 15986
rect 14030 15934 14082 15986
rect 14082 15934 14084 15986
rect 14028 15932 14084 15934
rect 13580 15260 13636 15316
rect 11340 12178 11396 12180
rect 11340 12126 11342 12178
rect 11342 12126 11394 12178
rect 11394 12126 11396 12178
rect 11340 12124 11396 12126
rect 12572 12850 12628 12852
rect 12572 12798 12574 12850
rect 12574 12798 12626 12850
rect 12626 12798 12628 12850
rect 12572 12796 12628 12798
rect 10444 11676 10500 11732
rect 10220 11394 10276 11396
rect 10220 11342 10222 11394
rect 10222 11342 10274 11394
rect 10274 11342 10276 11394
rect 10220 11340 10276 11342
rect 10108 10610 10164 10612
rect 10108 10558 10110 10610
rect 10110 10558 10162 10610
rect 10162 10558 10164 10610
rect 10108 10556 10164 10558
rect 11452 11618 11508 11620
rect 11452 11566 11454 11618
rect 11454 11566 11506 11618
rect 11506 11566 11508 11618
rect 11452 11564 11508 11566
rect 11788 11564 11844 11620
rect 11340 11340 11396 11396
rect 10444 10108 10500 10164
rect 10892 10556 10948 10612
rect 12236 11394 12292 11396
rect 12236 11342 12238 11394
rect 12238 11342 12290 11394
rect 12290 11342 12292 11394
rect 12236 11340 12292 11342
rect 11564 10498 11620 10500
rect 11564 10446 11566 10498
rect 11566 10446 11618 10498
rect 11618 10446 11620 10498
rect 11564 10444 11620 10446
rect 12124 10498 12180 10500
rect 12124 10446 12126 10498
rect 12126 10446 12178 10498
rect 12178 10446 12180 10498
rect 12124 10444 12180 10446
rect 10780 9772 10836 9828
rect 15484 17724 15540 17780
rect 15484 17388 15540 17444
rect 15036 16882 15092 16884
rect 15036 16830 15038 16882
rect 15038 16830 15090 16882
rect 15090 16830 15092 16882
rect 15036 16828 15092 16830
rect 15260 16716 15316 16772
rect 15148 15314 15204 15316
rect 15148 15262 15150 15314
rect 15150 15262 15202 15314
rect 15202 15262 15204 15314
rect 15148 15260 15204 15262
rect 14924 14476 14980 14532
rect 16492 23436 16548 23492
rect 16716 23772 16772 23828
rect 15820 22428 15876 22484
rect 15820 21756 15876 21812
rect 16156 21756 16212 21812
rect 16492 20748 16548 20804
rect 15820 20188 15876 20244
rect 15932 20076 15988 20132
rect 15820 19292 15876 19348
rect 15708 18844 15764 18900
rect 16156 19964 16212 20020
rect 19068 26572 19124 26628
rect 18172 26236 18228 26292
rect 17500 22652 17556 22708
rect 18060 24722 18116 24724
rect 18060 24670 18062 24722
rect 18062 24670 18114 24722
rect 18114 24670 18116 24722
rect 18060 24668 18116 24670
rect 17836 24556 17892 24612
rect 17836 23996 17892 24052
rect 18284 25452 18340 25508
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 21084 31500 21140 31556
rect 21308 31388 21364 31444
rect 21196 31276 21252 31332
rect 20860 29538 20916 29540
rect 20860 29486 20862 29538
rect 20862 29486 20914 29538
rect 20914 29486 20916 29538
rect 20860 29484 20916 29486
rect 21308 29148 21364 29204
rect 20748 29036 20804 29092
rect 22316 31218 22372 31220
rect 22316 31166 22318 31218
rect 22318 31166 22370 31218
rect 22370 31166 22372 31218
rect 22316 31164 22372 31166
rect 21756 31052 21812 31108
rect 22988 30994 23044 30996
rect 22988 30942 22990 30994
rect 22990 30942 23042 30994
rect 23042 30942 23044 30994
rect 22988 30940 23044 30942
rect 22204 30882 22260 30884
rect 22204 30830 22206 30882
rect 22206 30830 22258 30882
rect 22258 30830 22260 30882
rect 22204 30828 22260 30830
rect 21644 30156 21700 30212
rect 21532 29596 21588 29652
rect 25004 34076 25060 34132
rect 25116 33964 25172 34020
rect 24668 33628 24724 33684
rect 24220 31948 24276 32004
rect 23660 31500 23716 31556
rect 22204 29538 22260 29540
rect 22204 29486 22206 29538
rect 22206 29486 22258 29538
rect 22258 29486 22260 29538
rect 22204 29484 22260 29486
rect 21420 29036 21476 29092
rect 20524 28364 20580 28420
rect 20524 27804 20580 27860
rect 21196 27692 21252 27748
rect 21308 27580 21364 27636
rect 22092 28028 22148 28084
rect 21644 27916 21700 27972
rect 22204 27970 22260 27972
rect 22204 27918 22206 27970
rect 22206 27918 22258 27970
rect 22258 27918 22260 27970
rect 22204 27916 22260 27918
rect 21756 27804 21812 27860
rect 22092 27804 22148 27860
rect 23324 31388 23380 31444
rect 24444 31388 24500 31444
rect 24556 31106 24612 31108
rect 24556 31054 24558 31106
rect 24558 31054 24610 31106
rect 24610 31054 24612 31106
rect 24556 31052 24612 31054
rect 25228 33180 25284 33236
rect 25452 33628 25508 33684
rect 25452 32956 25508 33012
rect 25340 32620 25396 32676
rect 25116 31948 25172 32004
rect 25228 31836 25284 31892
rect 25900 38274 25956 38276
rect 25900 38222 25902 38274
rect 25902 38222 25954 38274
rect 25954 38222 25956 38274
rect 25900 38220 25956 38222
rect 27244 43650 27300 43652
rect 27244 43598 27246 43650
rect 27246 43598 27298 43650
rect 27298 43598 27300 43650
rect 27244 43596 27300 43598
rect 27132 43538 27188 43540
rect 27132 43486 27134 43538
rect 27134 43486 27186 43538
rect 27186 43486 27188 43538
rect 27132 43484 27188 43486
rect 27132 43260 27188 43316
rect 27580 45218 27636 45220
rect 27580 45166 27582 45218
rect 27582 45166 27634 45218
rect 27634 45166 27636 45218
rect 27580 45164 27636 45166
rect 27468 45106 27524 45108
rect 27468 45054 27470 45106
rect 27470 45054 27522 45106
rect 27522 45054 27524 45106
rect 27468 45052 27524 45054
rect 28252 45612 28308 45668
rect 27244 42866 27300 42868
rect 27244 42814 27246 42866
rect 27246 42814 27298 42866
rect 27298 42814 27300 42866
rect 27244 42812 27300 42814
rect 27132 42476 27188 42532
rect 27804 42642 27860 42644
rect 27804 42590 27806 42642
rect 27806 42590 27858 42642
rect 27858 42590 27860 42642
rect 27804 42588 27860 42590
rect 27132 42194 27188 42196
rect 27132 42142 27134 42194
rect 27134 42142 27186 42194
rect 27186 42142 27188 42194
rect 27132 42140 27188 42142
rect 26684 40908 26740 40964
rect 27244 40684 27300 40740
rect 27132 40514 27188 40516
rect 27132 40462 27134 40514
rect 27134 40462 27186 40514
rect 27186 40462 27188 40514
rect 27132 40460 27188 40462
rect 27132 39506 27188 39508
rect 27132 39454 27134 39506
rect 27134 39454 27186 39506
rect 27186 39454 27188 39506
rect 27132 39452 27188 39454
rect 26796 38220 26852 38276
rect 26124 37996 26180 38052
rect 25676 35532 25732 35588
rect 25788 35196 25844 35252
rect 25564 31724 25620 31780
rect 25676 35084 25732 35140
rect 26572 37660 26628 37716
rect 26796 37378 26852 37380
rect 26796 37326 26798 37378
rect 26798 37326 26850 37378
rect 26850 37326 26852 37378
rect 26796 37324 26852 37326
rect 26348 37212 26404 37268
rect 26236 36988 26292 37044
rect 26124 35756 26180 35812
rect 26012 35084 26068 35140
rect 25676 34636 25732 34692
rect 26236 34748 26292 34804
rect 26012 34354 26068 34356
rect 26012 34302 26014 34354
rect 26014 34302 26066 34354
rect 26066 34302 26068 34354
rect 26012 34300 26068 34302
rect 26572 37212 26628 37268
rect 26684 36988 26740 37044
rect 26572 36764 26628 36820
rect 28028 43538 28084 43540
rect 28028 43486 28030 43538
rect 28030 43486 28082 43538
rect 28082 43486 28084 43538
rect 28028 43484 28084 43486
rect 28252 43538 28308 43540
rect 28252 43486 28254 43538
rect 28254 43486 28306 43538
rect 28306 43486 28308 43538
rect 28252 43484 28308 43486
rect 28812 43650 28868 43652
rect 28812 43598 28814 43650
rect 28814 43598 28866 43650
rect 28866 43598 28868 43650
rect 28812 43596 28868 43598
rect 28924 43484 28980 43540
rect 28028 42924 28084 42980
rect 28476 43260 28532 43316
rect 28700 39788 28756 39844
rect 28140 38162 28196 38164
rect 28140 38110 28142 38162
rect 28142 38110 28194 38162
rect 28194 38110 28196 38162
rect 28140 38108 28196 38110
rect 27916 37884 27972 37940
rect 28364 37436 28420 37492
rect 27356 36428 27412 36484
rect 27916 36428 27972 36484
rect 27244 35532 27300 35588
rect 26908 35420 26964 35476
rect 27244 35308 27300 35364
rect 25676 33068 25732 33124
rect 26684 34636 26740 34692
rect 26012 31778 26068 31780
rect 26012 31726 26014 31778
rect 26014 31726 26066 31778
rect 26066 31726 26068 31778
rect 26012 31724 26068 31726
rect 24780 31388 24836 31444
rect 25452 31276 25508 31332
rect 25228 31164 25284 31220
rect 25340 31106 25396 31108
rect 25340 31054 25342 31106
rect 25342 31054 25394 31106
rect 25394 31054 25396 31106
rect 25340 31052 25396 31054
rect 23324 29484 23380 29540
rect 24220 30156 24276 30212
rect 22652 27580 22708 27636
rect 22988 27580 23044 27636
rect 22876 27244 22932 27300
rect 20412 26348 20468 26404
rect 20524 26684 20580 26740
rect 18732 25506 18788 25508
rect 18732 25454 18734 25506
rect 18734 25454 18786 25506
rect 18786 25454 18788 25506
rect 18732 25452 18788 25454
rect 18508 24610 18564 24612
rect 18508 24558 18510 24610
rect 18510 24558 18562 24610
rect 18562 24558 18564 24610
rect 18508 24556 18564 24558
rect 19404 25788 19460 25844
rect 18956 25228 19012 25284
rect 20188 25282 20244 25284
rect 20188 25230 20190 25282
rect 20190 25230 20242 25282
rect 20242 25230 20244 25282
rect 20188 25228 20244 25230
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 19292 24722 19348 24724
rect 19292 24670 19294 24722
rect 19294 24670 19346 24722
rect 19346 24670 19348 24722
rect 19292 24668 19348 24670
rect 19740 24610 19796 24612
rect 19740 24558 19742 24610
rect 19742 24558 19794 24610
rect 19794 24558 19796 24610
rect 19740 24556 19796 24558
rect 23212 26460 23268 26516
rect 20748 26178 20804 26180
rect 20748 26126 20750 26178
rect 20750 26126 20802 26178
rect 20802 26126 20804 26178
rect 20748 26124 20804 26126
rect 19964 23938 20020 23940
rect 19964 23886 19966 23938
rect 19966 23886 20018 23938
rect 20018 23886 20020 23938
rect 19964 23884 20020 23886
rect 18508 23826 18564 23828
rect 18508 23774 18510 23826
rect 18510 23774 18562 23826
rect 18562 23774 18564 23826
rect 18508 23772 18564 23774
rect 18620 23714 18676 23716
rect 18620 23662 18622 23714
rect 18622 23662 18674 23714
rect 18674 23662 18676 23714
rect 18620 23660 18676 23662
rect 17836 22316 17892 22372
rect 17948 21644 18004 21700
rect 17612 21586 17668 21588
rect 17612 21534 17614 21586
rect 17614 21534 17666 21586
rect 17666 21534 17668 21586
rect 17612 21532 17668 21534
rect 16716 20076 16772 20132
rect 16044 19180 16100 19236
rect 16044 18508 16100 18564
rect 15932 17778 15988 17780
rect 15932 17726 15934 17778
rect 15934 17726 15986 17778
rect 15986 17726 15988 17778
rect 15932 17724 15988 17726
rect 16716 19404 16772 19460
rect 16604 18732 16660 18788
rect 16492 18450 16548 18452
rect 16492 18398 16494 18450
rect 16494 18398 16546 18450
rect 16546 18398 16548 18450
rect 16492 18396 16548 18398
rect 17052 19404 17108 19460
rect 18396 22316 18452 22372
rect 18396 21756 18452 21812
rect 18172 21474 18228 21476
rect 18172 21422 18174 21474
rect 18174 21422 18226 21474
rect 18226 21422 18228 21474
rect 18172 21420 18228 21422
rect 17724 20748 17780 20804
rect 17500 18732 17556 18788
rect 17388 18396 17444 18452
rect 18508 19964 18564 20020
rect 18060 19404 18116 19460
rect 17948 19346 18004 19348
rect 17948 19294 17950 19346
rect 17950 19294 18002 19346
rect 18002 19294 18004 19346
rect 17948 19292 18004 19294
rect 18060 18562 18116 18564
rect 18060 18510 18062 18562
rect 18062 18510 18114 18562
rect 18114 18510 18116 18562
rect 18060 18508 18116 18510
rect 16380 17612 16436 17668
rect 17164 17666 17220 17668
rect 17164 17614 17166 17666
rect 17166 17614 17218 17666
rect 17218 17614 17220 17666
rect 17164 17612 17220 17614
rect 15596 16604 15652 16660
rect 16156 17442 16212 17444
rect 16156 17390 16158 17442
rect 16158 17390 16210 17442
rect 16210 17390 16212 17442
rect 16156 17388 16212 17390
rect 15932 15986 15988 15988
rect 15932 15934 15934 15986
rect 15934 15934 15986 15986
rect 15986 15934 15988 15986
rect 15932 15932 15988 15934
rect 16268 16156 16324 16212
rect 15708 15148 15764 15204
rect 16940 16828 16996 16884
rect 16380 16044 16436 16100
rect 16380 15148 16436 15204
rect 16492 15932 16548 15988
rect 17052 15932 17108 15988
rect 17276 15820 17332 15876
rect 12684 11564 12740 11620
rect 12908 11282 12964 11284
rect 12908 11230 12910 11282
rect 12910 11230 12962 11282
rect 12962 11230 12964 11282
rect 12908 11228 12964 11230
rect 12796 10108 12852 10164
rect 12796 9826 12852 9828
rect 12796 9774 12798 9826
rect 12798 9774 12850 9826
rect 12850 9774 12852 9826
rect 12796 9772 12852 9774
rect 9548 9212 9604 9268
rect 9548 8316 9604 8372
rect 9660 8092 9716 8148
rect 9324 7532 9380 7588
rect 9548 7644 9604 7700
rect 10108 9042 10164 9044
rect 10108 8990 10110 9042
rect 10110 8990 10162 9042
rect 10162 8990 10164 9042
rect 10108 8988 10164 8990
rect 9996 8316 10052 8372
rect 11228 8316 11284 8372
rect 11004 8258 11060 8260
rect 11004 8206 11006 8258
rect 11006 8206 11058 8258
rect 11058 8206 11060 8258
rect 11004 8204 11060 8206
rect 9772 7250 9828 7252
rect 9772 7198 9774 7250
rect 9774 7198 9826 7250
rect 9826 7198 9828 7250
rect 9772 7196 9828 7198
rect 11004 7196 11060 7252
rect 11340 6524 11396 6580
rect 12348 8316 12404 8372
rect 11788 8258 11844 8260
rect 11788 8206 11790 8258
rect 11790 8206 11842 8258
rect 11842 8206 11844 8258
rect 11788 8204 11844 8206
rect 13468 11394 13524 11396
rect 13468 11342 13470 11394
rect 13470 11342 13522 11394
rect 13522 11342 13524 11394
rect 13468 11340 13524 11342
rect 14252 11506 14308 11508
rect 14252 11454 14254 11506
rect 14254 11454 14306 11506
rect 14306 11454 14308 11506
rect 14252 11452 14308 11454
rect 13804 11282 13860 11284
rect 13804 11230 13806 11282
rect 13806 11230 13858 11282
rect 13858 11230 13860 11282
rect 13804 11228 13860 11230
rect 14252 10780 14308 10836
rect 13692 9660 13748 9716
rect 14588 12066 14644 12068
rect 14588 12014 14590 12066
rect 14590 12014 14642 12066
rect 14642 12014 14644 12066
rect 14588 12012 14644 12014
rect 15036 11900 15092 11956
rect 14700 11340 14756 11396
rect 14476 9714 14532 9716
rect 14476 9662 14478 9714
rect 14478 9662 14530 9714
rect 14530 9662 14532 9714
rect 14476 9660 14532 9662
rect 19068 22370 19124 22372
rect 19068 22318 19070 22370
rect 19070 22318 19122 22370
rect 19122 22318 19124 22370
rect 19068 22316 19124 22318
rect 19068 21532 19124 21588
rect 19180 21474 19236 21476
rect 19180 21422 19182 21474
rect 19182 21422 19234 21474
rect 19234 21422 19236 21474
rect 19180 21420 19236 21422
rect 19516 23714 19572 23716
rect 19516 23662 19518 23714
rect 19518 23662 19570 23714
rect 19570 23662 19572 23714
rect 19516 23660 19572 23662
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 22988 25730 23044 25732
rect 22988 25678 22990 25730
rect 22990 25678 23042 25730
rect 23042 25678 23044 25730
rect 22988 25676 23044 25678
rect 23548 28028 23604 28084
rect 23436 27244 23492 27300
rect 23660 27580 23716 27636
rect 23548 27020 23604 27076
rect 23436 26796 23492 26852
rect 23324 26236 23380 26292
rect 24220 27580 24276 27636
rect 23884 26572 23940 26628
rect 23660 26012 23716 26068
rect 23884 25900 23940 25956
rect 24220 26178 24276 26180
rect 24220 26126 24222 26178
rect 24222 26126 24274 26178
rect 24274 26126 24276 26178
rect 24220 26124 24276 26126
rect 24668 30940 24724 30996
rect 24444 30156 24500 30212
rect 25228 29986 25284 29988
rect 25228 29934 25230 29986
rect 25230 29934 25282 29986
rect 25282 29934 25284 29986
rect 25228 29932 25284 29934
rect 25452 29650 25508 29652
rect 25452 29598 25454 29650
rect 25454 29598 25506 29650
rect 25506 29598 25508 29650
rect 25452 29596 25508 29598
rect 25116 29036 25172 29092
rect 24668 28028 24724 28084
rect 24668 27356 24724 27412
rect 25004 27186 25060 27188
rect 25004 27134 25006 27186
rect 25006 27134 25058 27186
rect 25058 27134 25060 27186
rect 25004 27132 25060 27134
rect 24556 27020 24612 27076
rect 25116 26908 25172 26964
rect 24332 26012 24388 26068
rect 24892 26124 24948 26180
rect 24444 25900 24500 25956
rect 23548 25340 23604 25396
rect 23212 25228 23268 25284
rect 20860 23884 20916 23940
rect 20412 22988 20468 23044
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 20300 21644 20356 21700
rect 19404 20802 19460 20804
rect 19404 20750 19406 20802
rect 19406 20750 19458 20802
rect 19458 20750 19460 20802
rect 19404 20748 19460 20750
rect 18956 20018 19012 20020
rect 18956 19966 18958 20018
rect 18958 19966 19010 20018
rect 19010 19966 19012 20018
rect 18956 19964 19012 19966
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 19628 20188 19684 20244
rect 19292 20130 19348 20132
rect 19292 20078 19294 20130
rect 19294 20078 19346 20130
rect 19346 20078 19348 20130
rect 19292 20076 19348 20078
rect 20860 21756 20916 21812
rect 20412 21532 20468 21588
rect 20300 20188 20356 20244
rect 20076 20130 20132 20132
rect 20076 20078 20078 20130
rect 20078 20078 20130 20130
rect 20130 20078 20132 20130
rect 20076 20076 20132 20078
rect 20412 19852 20468 19908
rect 21644 24946 21700 24948
rect 21644 24894 21646 24946
rect 21646 24894 21698 24946
rect 21698 24894 21700 24946
rect 21644 24892 21700 24894
rect 22204 24946 22260 24948
rect 22204 24894 22206 24946
rect 22206 24894 22258 24946
rect 22258 24894 22260 24946
rect 22204 24892 22260 24894
rect 23212 23772 23268 23828
rect 23324 24892 23380 24948
rect 24108 24946 24164 24948
rect 24108 24894 24110 24946
rect 24110 24894 24162 24946
rect 24162 24894 24164 24946
rect 24108 24892 24164 24894
rect 23660 24444 23716 24500
rect 24220 24444 24276 24500
rect 23548 24108 23604 24164
rect 24108 24332 24164 24388
rect 22540 23714 22596 23716
rect 22540 23662 22542 23714
rect 22542 23662 22594 23714
rect 22594 23662 22596 23714
rect 22540 23660 22596 23662
rect 22316 23378 22372 23380
rect 22316 23326 22318 23378
rect 22318 23326 22370 23378
rect 22370 23326 22372 23378
rect 22316 23324 22372 23326
rect 21308 23154 21364 23156
rect 21308 23102 21310 23154
rect 21310 23102 21362 23154
rect 21362 23102 21364 23154
rect 21308 23100 21364 23102
rect 21980 23154 22036 23156
rect 21980 23102 21982 23154
rect 21982 23102 22034 23154
rect 22034 23102 22036 23154
rect 21980 23100 22036 23102
rect 21756 23042 21812 23044
rect 21756 22990 21758 23042
rect 21758 22990 21810 23042
rect 21810 22990 21812 23042
rect 21756 22988 21812 22990
rect 21868 22370 21924 22372
rect 21868 22318 21870 22370
rect 21870 22318 21922 22370
rect 21922 22318 21924 22370
rect 21868 22316 21924 22318
rect 22540 23154 22596 23156
rect 22540 23102 22542 23154
rect 22542 23102 22594 23154
rect 22594 23102 22596 23154
rect 22540 23100 22596 23102
rect 22652 22988 22708 23044
rect 22652 22370 22708 22372
rect 22652 22318 22654 22370
rect 22654 22318 22706 22370
rect 22706 22318 22708 22370
rect 22652 22316 22708 22318
rect 21308 21756 21364 21812
rect 21084 20188 21140 20244
rect 20972 19516 21028 19572
rect 22092 22092 22148 22148
rect 21756 21586 21812 21588
rect 21756 21534 21758 21586
rect 21758 21534 21810 21586
rect 21810 21534 21812 21586
rect 21756 21532 21812 21534
rect 19516 19234 19572 19236
rect 19516 19182 19518 19234
rect 19518 19182 19570 19234
rect 19570 19182 19572 19234
rect 19516 19180 19572 19182
rect 19068 18284 19124 18340
rect 20524 19292 20580 19348
rect 19740 19122 19796 19124
rect 19740 19070 19742 19122
rect 19742 19070 19794 19122
rect 19794 19070 19796 19122
rect 19740 19068 19796 19070
rect 20412 18956 20468 19012
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19628 18396 19684 18452
rect 20300 18284 20356 18340
rect 18956 16210 19012 16212
rect 18956 16158 18958 16210
rect 18958 16158 19010 16210
rect 19010 16158 19012 16210
rect 18956 16156 19012 16158
rect 18844 16098 18900 16100
rect 18844 16046 18846 16098
rect 18846 16046 18898 16098
rect 18898 16046 18900 16098
rect 18844 16044 18900 16046
rect 19180 15932 19236 15988
rect 19404 16044 19460 16100
rect 19292 15260 19348 15316
rect 17948 14754 18004 14756
rect 17948 14702 17950 14754
rect 17950 14702 18002 14754
rect 18002 14702 18004 14754
rect 17948 14700 18004 14702
rect 18844 14700 18900 14756
rect 17724 14530 17780 14532
rect 17724 14478 17726 14530
rect 17726 14478 17778 14530
rect 17778 14478 17780 14530
rect 17724 14476 17780 14478
rect 15372 11506 15428 11508
rect 15372 11454 15374 11506
rect 15374 11454 15426 11506
rect 15426 11454 15428 11506
rect 15372 11452 15428 11454
rect 16492 12290 16548 12292
rect 16492 12238 16494 12290
rect 16494 12238 16546 12290
rect 16546 12238 16548 12290
rect 16492 12236 16548 12238
rect 16604 11340 16660 11396
rect 15036 10780 15092 10836
rect 14924 10722 14980 10724
rect 14924 10670 14926 10722
rect 14926 10670 14978 10722
rect 14978 10670 14980 10722
rect 14924 10668 14980 10670
rect 15148 9772 15204 9828
rect 17388 11340 17444 11396
rect 16604 10668 16660 10724
rect 17052 10556 17108 10612
rect 17836 11954 17892 11956
rect 17836 11902 17838 11954
rect 17838 11902 17890 11954
rect 17890 11902 17892 11954
rect 17836 11900 17892 11902
rect 18060 12850 18116 12852
rect 18060 12798 18062 12850
rect 18062 12798 18114 12850
rect 18114 12798 18116 12850
rect 18060 12796 18116 12798
rect 18060 12236 18116 12292
rect 19292 12850 19348 12852
rect 19292 12798 19294 12850
rect 19294 12798 19346 12850
rect 19346 12798 19348 12850
rect 19292 12796 19348 12798
rect 18956 12290 19012 12292
rect 18956 12238 18958 12290
rect 18958 12238 19010 12290
rect 19010 12238 19012 12290
rect 18956 12236 19012 12238
rect 19404 12684 19460 12740
rect 18508 11900 18564 11956
rect 17948 11228 18004 11284
rect 17836 10610 17892 10612
rect 17836 10558 17838 10610
rect 17838 10558 17890 10610
rect 17890 10558 17892 10610
rect 17836 10556 17892 10558
rect 15372 9826 15428 9828
rect 15372 9774 15374 9826
rect 15374 9774 15426 9826
rect 15426 9774 15428 9826
rect 15372 9772 15428 9774
rect 15148 9154 15204 9156
rect 15148 9102 15150 9154
rect 15150 9102 15202 9154
rect 15202 9102 15204 9154
rect 15148 9100 15204 9102
rect 15260 9212 15316 9268
rect 13020 8316 13076 8372
rect 13580 8258 13636 8260
rect 13580 8206 13582 8258
rect 13582 8206 13634 8258
rect 13634 8206 13636 8258
rect 13580 8204 13636 8206
rect 13804 8316 13860 8372
rect 15484 9660 15540 9716
rect 15820 9714 15876 9716
rect 15820 9662 15822 9714
rect 15822 9662 15874 9714
rect 15874 9662 15876 9714
rect 15820 9660 15876 9662
rect 15820 9266 15876 9268
rect 15820 9214 15822 9266
rect 15822 9214 15874 9266
rect 15874 9214 15876 9266
rect 15820 9212 15876 9214
rect 15484 8146 15540 8148
rect 15484 8094 15486 8146
rect 15486 8094 15538 8146
rect 15538 8094 15540 8146
rect 15484 8092 15540 8094
rect 12684 7980 12740 8036
rect 11900 7868 11956 7924
rect 11788 7586 11844 7588
rect 11788 7534 11790 7586
rect 11790 7534 11842 7586
rect 11842 7534 11844 7586
rect 11788 7532 11844 7534
rect 12348 7586 12404 7588
rect 12348 7534 12350 7586
rect 12350 7534 12402 7586
rect 12402 7534 12404 7586
rect 12348 7532 12404 7534
rect 13020 8034 13076 8036
rect 13020 7982 13022 8034
rect 13022 7982 13074 8034
rect 13074 7982 13076 8034
rect 13020 7980 13076 7982
rect 14140 7980 14196 8036
rect 12796 7868 12852 7924
rect 12684 7532 12740 7588
rect 12236 7250 12292 7252
rect 12236 7198 12238 7250
rect 12238 7198 12290 7250
rect 12290 7198 12292 7250
rect 12236 7196 12292 7198
rect 11676 6802 11732 6804
rect 11676 6750 11678 6802
rect 11678 6750 11730 6802
rect 11730 6750 11732 6802
rect 11676 6748 11732 6750
rect 13132 6748 13188 6804
rect 12460 6690 12516 6692
rect 12460 6638 12462 6690
rect 12462 6638 12514 6690
rect 12514 6638 12516 6690
rect 12460 6636 12516 6638
rect 12348 6578 12404 6580
rect 12348 6526 12350 6578
rect 12350 6526 12402 6578
rect 12402 6526 12404 6578
rect 12348 6524 12404 6526
rect 11788 6412 11844 6468
rect 12572 6466 12628 6468
rect 12572 6414 12574 6466
rect 12574 6414 12626 6466
rect 12626 6414 12628 6466
rect 12572 6412 12628 6414
rect 11564 5964 11620 6020
rect 12348 6018 12404 6020
rect 12348 5966 12350 6018
rect 12350 5966 12402 6018
rect 12402 5966 12404 6018
rect 12348 5964 12404 5966
rect 13580 6802 13636 6804
rect 13580 6750 13582 6802
rect 13582 6750 13634 6802
rect 13634 6750 13636 6802
rect 13580 6748 13636 6750
rect 14924 7868 14980 7924
rect 15372 7698 15428 7700
rect 15372 7646 15374 7698
rect 15374 7646 15426 7698
rect 15426 7646 15428 7698
rect 15372 7644 15428 7646
rect 14252 7362 14308 7364
rect 14252 7310 14254 7362
rect 14254 7310 14306 7362
rect 14306 7310 14308 7362
rect 14252 7308 14308 7310
rect 15148 6412 15204 6468
rect 15932 8876 15988 8932
rect 17052 9826 17108 9828
rect 17052 9774 17054 9826
rect 17054 9774 17106 9826
rect 17106 9774 17108 9826
rect 17052 9772 17108 9774
rect 18284 10556 18340 10612
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 20076 16098 20132 16100
rect 20076 16046 20078 16098
rect 20078 16046 20130 16098
rect 20130 16046 20132 16098
rect 20076 16044 20132 16046
rect 20412 17500 20468 17556
rect 20524 18508 20580 18564
rect 20636 19180 20692 19236
rect 20636 17052 20692 17108
rect 20524 15820 20580 15876
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 20300 15314 20356 15316
rect 20300 15262 20302 15314
rect 20302 15262 20354 15314
rect 20354 15262 20356 15314
rect 20300 15260 20356 15262
rect 20076 14642 20132 14644
rect 20076 14590 20078 14642
rect 20078 14590 20130 14642
rect 20130 14590 20132 14642
rect 20076 14588 20132 14590
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 21420 19068 21476 19124
rect 22876 22316 22932 22372
rect 23436 23324 23492 23380
rect 23772 23042 23828 23044
rect 23772 22990 23774 23042
rect 23774 22990 23826 23042
rect 23826 22990 23828 23042
rect 23772 22988 23828 22990
rect 24444 24892 24500 24948
rect 25116 24892 25172 24948
rect 25788 30268 25844 30324
rect 25340 28140 25396 28196
rect 24444 24050 24500 24052
rect 24444 23998 24446 24050
rect 24446 23998 24498 24050
rect 24498 23998 24500 24050
rect 24444 23996 24500 23998
rect 25676 28700 25732 28756
rect 26012 31388 26068 31444
rect 26012 31052 26068 31108
rect 26012 29538 26068 29540
rect 26012 29486 26014 29538
rect 26014 29486 26066 29538
rect 26066 29486 26068 29538
rect 26012 29484 26068 29486
rect 27132 35196 27188 35252
rect 26908 33852 26964 33908
rect 26572 32956 26628 33012
rect 26684 32844 26740 32900
rect 26572 32060 26628 32116
rect 26572 31052 26628 31108
rect 27020 33740 27076 33796
rect 27020 31500 27076 31556
rect 26348 30156 26404 30212
rect 26796 30828 26852 30884
rect 25788 28924 25844 28980
rect 25564 28082 25620 28084
rect 25564 28030 25566 28082
rect 25566 28030 25618 28082
rect 25618 28030 25620 28082
rect 25564 28028 25620 28030
rect 25788 27916 25844 27972
rect 25676 27858 25732 27860
rect 25676 27806 25678 27858
rect 25678 27806 25730 27858
rect 25730 27806 25732 27858
rect 25676 27804 25732 27806
rect 25676 27356 25732 27412
rect 25676 27074 25732 27076
rect 25676 27022 25678 27074
rect 25678 27022 25730 27074
rect 25730 27022 25732 27074
rect 25676 27020 25732 27022
rect 26012 27468 26068 27524
rect 26572 29426 26628 29428
rect 26572 29374 26574 29426
rect 26574 29374 26626 29426
rect 26626 29374 26628 29426
rect 26572 29372 26628 29374
rect 26460 29314 26516 29316
rect 26460 29262 26462 29314
rect 26462 29262 26514 29314
rect 26514 29262 26516 29314
rect 26460 29260 26516 29262
rect 26348 28588 26404 28644
rect 26796 29538 26852 29540
rect 26796 29486 26798 29538
rect 26798 29486 26850 29538
rect 26850 29486 26852 29538
rect 26796 29484 26852 29486
rect 27244 34748 27300 34804
rect 27356 35084 27412 35140
rect 27244 32956 27300 33012
rect 27468 32732 27524 32788
rect 27692 36204 27748 36260
rect 28140 36204 28196 36260
rect 29708 54796 29764 54852
rect 29148 54626 29204 54628
rect 29148 54574 29150 54626
rect 29150 54574 29202 54626
rect 29202 54574 29204 54626
rect 29148 54572 29204 54574
rect 29932 53506 29988 53508
rect 29932 53454 29934 53506
rect 29934 53454 29986 53506
rect 29986 53454 29988 53506
rect 29932 53452 29988 53454
rect 29148 53170 29204 53172
rect 29148 53118 29150 53170
rect 29150 53118 29202 53170
rect 29202 53118 29204 53170
rect 29148 53116 29204 53118
rect 29708 52834 29764 52836
rect 29708 52782 29710 52834
rect 29710 52782 29762 52834
rect 29762 52782 29764 52834
rect 29708 52780 29764 52782
rect 29708 52220 29764 52276
rect 29932 53004 29988 53060
rect 29932 52162 29988 52164
rect 29932 52110 29934 52162
rect 29934 52110 29986 52162
rect 29986 52110 29988 52162
rect 29932 52108 29988 52110
rect 30604 53900 30660 53956
rect 31612 56252 31668 56308
rect 30268 53452 30324 53508
rect 31276 54348 31332 54404
rect 31164 53618 31220 53620
rect 31164 53566 31166 53618
rect 31166 53566 31218 53618
rect 31218 53566 31220 53618
rect 31164 53564 31220 53566
rect 30268 52220 30324 52276
rect 30156 51996 30212 52052
rect 30492 52780 30548 52836
rect 30604 52444 30660 52500
rect 30492 51996 30548 52052
rect 31164 52444 31220 52500
rect 31052 52108 31108 52164
rect 30380 49980 30436 50036
rect 29708 49756 29764 49812
rect 29372 49308 29428 49364
rect 29820 49196 29876 49252
rect 29932 49644 29988 49700
rect 29596 48860 29652 48916
rect 29372 46284 29428 46340
rect 29148 43596 29204 43652
rect 29148 42588 29204 42644
rect 29260 42924 29316 42980
rect 29148 40460 29204 40516
rect 29260 39788 29316 39844
rect 28812 38108 28868 38164
rect 30380 49810 30436 49812
rect 30380 49758 30382 49810
rect 30382 49758 30434 49810
rect 30434 49758 30436 49810
rect 30380 49756 30436 49758
rect 30604 51212 30660 51268
rect 31052 50594 31108 50596
rect 31052 50542 31054 50594
rect 31054 50542 31106 50594
rect 31106 50542 31108 50594
rect 31052 50540 31108 50542
rect 31164 50428 31220 50484
rect 30828 49980 30884 50036
rect 31612 53676 31668 53732
rect 31724 54572 31780 54628
rect 31612 53058 31668 53060
rect 31612 53006 31614 53058
rect 31614 53006 31666 53058
rect 31666 53006 31668 53058
rect 31612 53004 31668 53006
rect 32284 55356 32340 55412
rect 31836 54402 31892 54404
rect 31836 54350 31838 54402
rect 31838 54350 31890 54402
rect 31890 54350 31892 54402
rect 31836 54348 31892 54350
rect 31388 52780 31444 52836
rect 32060 52220 32116 52276
rect 31724 51884 31780 51940
rect 31612 51490 31668 51492
rect 31612 51438 31614 51490
rect 31614 51438 31666 51490
rect 31666 51438 31668 51490
rect 31612 51436 31668 51438
rect 33180 56306 33236 56308
rect 33180 56254 33182 56306
rect 33182 56254 33234 56306
rect 33234 56254 33236 56306
rect 33180 56252 33236 56254
rect 33516 55410 33572 55412
rect 33516 55358 33518 55410
rect 33518 55358 33570 55410
rect 33570 55358 33572 55410
rect 33516 55356 33572 55358
rect 34300 55916 34356 55972
rect 33740 55356 33796 55412
rect 34972 55244 35028 55300
rect 32956 54684 33012 54740
rect 34188 54738 34244 54740
rect 34188 54686 34190 54738
rect 34190 54686 34242 54738
rect 34242 54686 34244 54738
rect 34188 54684 34244 54686
rect 32396 54626 32452 54628
rect 32396 54574 32398 54626
rect 32398 54574 32450 54626
rect 32450 54574 32452 54626
rect 32396 54572 32452 54574
rect 33180 54514 33236 54516
rect 33180 54462 33182 54514
rect 33182 54462 33234 54514
rect 33234 54462 33236 54514
rect 33180 54460 33236 54462
rect 32620 54348 32676 54404
rect 32396 53900 32452 53956
rect 35196 55690 35252 55692
rect 35196 55638 35198 55690
rect 35198 55638 35250 55690
rect 35250 55638 35252 55690
rect 35196 55636 35252 55638
rect 35300 55690 35356 55692
rect 35300 55638 35302 55690
rect 35302 55638 35354 55690
rect 35354 55638 35356 55690
rect 35300 55636 35356 55638
rect 35404 55690 35460 55692
rect 35404 55638 35406 55690
rect 35406 55638 35458 55690
rect 35458 55638 35460 55690
rect 35404 55636 35460 55638
rect 35532 55356 35588 55412
rect 35196 54122 35252 54124
rect 35196 54070 35198 54122
rect 35198 54070 35250 54122
rect 35250 54070 35252 54122
rect 35196 54068 35252 54070
rect 35300 54122 35356 54124
rect 35300 54070 35302 54122
rect 35302 54070 35354 54122
rect 35354 54070 35356 54122
rect 35300 54068 35356 54070
rect 35404 54122 35460 54124
rect 35404 54070 35406 54122
rect 35406 54070 35458 54122
rect 35458 54070 35460 54122
rect 35404 54068 35460 54070
rect 32396 53618 32452 53620
rect 32396 53566 32398 53618
rect 32398 53566 32450 53618
rect 32450 53566 32452 53618
rect 32396 53564 32452 53566
rect 32844 53004 32900 53060
rect 32396 52892 32452 52948
rect 32172 51884 32228 51940
rect 32396 52108 32452 52164
rect 30156 47964 30212 48020
rect 32508 51490 32564 51492
rect 32508 51438 32510 51490
rect 32510 51438 32562 51490
rect 32562 51438 32564 51490
rect 32508 51436 32564 51438
rect 31500 49644 31556 49700
rect 31052 49026 31108 49028
rect 31052 48974 31054 49026
rect 31054 48974 31106 49026
rect 31106 48974 31108 49026
rect 31052 48972 31108 48974
rect 31164 48914 31220 48916
rect 31164 48862 31166 48914
rect 31166 48862 31218 48914
rect 31218 48862 31220 48914
rect 31164 48860 31220 48862
rect 31164 48076 31220 48132
rect 30604 47516 30660 47572
rect 29484 39004 29540 39060
rect 30156 39842 30212 39844
rect 30156 39790 30158 39842
rect 30158 39790 30210 39842
rect 30210 39790 30212 39842
rect 30156 39788 30212 39790
rect 30940 46786 30996 46788
rect 30940 46734 30942 46786
rect 30942 46734 30994 46786
rect 30994 46734 30996 46786
rect 30940 46732 30996 46734
rect 31052 46060 31108 46116
rect 31500 49308 31556 49364
rect 31388 47570 31444 47572
rect 31388 47518 31390 47570
rect 31390 47518 31442 47570
rect 31442 47518 31444 47570
rect 31388 47516 31444 47518
rect 31724 50428 31780 50484
rect 32172 49980 32228 50036
rect 31724 47628 31780 47684
rect 31276 47180 31332 47236
rect 31388 47068 31444 47124
rect 30604 43148 30660 43204
rect 30604 42642 30660 42644
rect 30604 42590 30606 42642
rect 30606 42590 30658 42642
rect 30658 42590 30660 42642
rect 30604 42588 30660 42590
rect 30716 41916 30772 41972
rect 30828 41132 30884 41188
rect 31388 43148 31444 43204
rect 31612 47180 31668 47236
rect 32172 48972 32228 49028
rect 33180 51548 33236 51604
rect 33404 53058 33460 53060
rect 33404 53006 33406 53058
rect 33406 53006 33458 53058
rect 33458 53006 33460 53058
rect 33404 53004 33460 53006
rect 33068 51324 33124 51380
rect 32844 50652 32900 50708
rect 35420 53900 35476 53956
rect 33852 52946 33908 52948
rect 33852 52894 33854 52946
rect 33854 52894 33906 52946
rect 33906 52894 33908 52946
rect 33852 52892 33908 52894
rect 33740 52332 33796 52388
rect 32956 50482 33012 50484
rect 32956 50430 32958 50482
rect 32958 50430 33010 50482
rect 33010 50430 33012 50482
rect 32956 50428 33012 50430
rect 33964 52162 34020 52164
rect 33964 52110 33966 52162
rect 33966 52110 34018 52162
rect 34018 52110 34020 52162
rect 33964 52108 34020 52110
rect 34636 51772 34692 51828
rect 34076 51436 34132 51492
rect 34524 51266 34580 51268
rect 34524 51214 34526 51266
rect 34526 51214 34578 51266
rect 34578 51214 34580 51266
rect 34524 51212 34580 51214
rect 34412 50764 34468 50820
rect 34188 50540 34244 50596
rect 31948 46732 32004 46788
rect 32844 49138 32900 49140
rect 32844 49086 32846 49138
rect 32846 49086 32898 49138
rect 32898 49086 32900 49138
rect 32844 49084 32900 49086
rect 33180 48914 33236 48916
rect 33180 48862 33182 48914
rect 33182 48862 33234 48914
rect 33234 48862 33236 48914
rect 33180 48860 33236 48862
rect 33292 48748 33348 48804
rect 32396 48354 32452 48356
rect 32396 48302 32398 48354
rect 32398 48302 32450 48354
rect 32450 48302 32452 48354
rect 32396 48300 32452 48302
rect 32844 48188 32900 48244
rect 32284 47628 32340 47684
rect 32060 46956 32116 47012
rect 31836 46562 31892 46564
rect 31836 46510 31838 46562
rect 31838 46510 31890 46562
rect 31890 46510 31892 46562
rect 31836 46508 31892 46510
rect 31948 46114 32004 46116
rect 31948 46062 31950 46114
rect 31950 46062 32002 46114
rect 32002 46062 32004 46114
rect 31948 46060 32004 46062
rect 32284 46620 32340 46676
rect 33068 48130 33124 48132
rect 33068 48078 33070 48130
rect 33070 48078 33122 48130
rect 33122 48078 33124 48130
rect 33068 48076 33124 48078
rect 33292 48018 33348 48020
rect 33292 47966 33294 48018
rect 33294 47966 33346 48018
rect 33346 47966 33348 48018
rect 33292 47964 33348 47966
rect 33516 48748 33572 48804
rect 33516 47964 33572 48020
rect 34300 48748 34356 48804
rect 34636 50540 34692 50596
rect 36316 56252 36372 56308
rect 36988 56140 37044 56196
rect 36204 55970 36260 55972
rect 36204 55918 36206 55970
rect 36206 55918 36258 55970
rect 36258 55918 36260 55970
rect 36204 55916 36260 55918
rect 36092 55356 36148 55412
rect 37212 55410 37268 55412
rect 37212 55358 37214 55410
rect 37214 55358 37266 55410
rect 37266 55358 37268 55410
rect 37212 55356 37268 55358
rect 35756 55132 35812 55188
rect 36428 55186 36484 55188
rect 36428 55134 36430 55186
rect 36430 55134 36482 55186
rect 36482 55134 36484 55186
rect 36428 55132 36484 55134
rect 35980 55074 36036 55076
rect 35980 55022 35982 55074
rect 35982 55022 36034 55074
rect 36034 55022 36036 55074
rect 35980 55020 36036 55022
rect 36764 55020 36820 55076
rect 35644 54348 35700 54404
rect 35308 52780 35364 52836
rect 35196 52554 35252 52556
rect 35196 52502 35198 52554
rect 35198 52502 35250 52554
rect 35250 52502 35252 52554
rect 35196 52500 35252 52502
rect 35300 52554 35356 52556
rect 35300 52502 35302 52554
rect 35302 52502 35354 52554
rect 35354 52502 35356 52554
rect 35300 52500 35356 52502
rect 35404 52554 35460 52556
rect 35404 52502 35406 52554
rect 35406 52502 35458 52554
rect 35458 52502 35460 52554
rect 35404 52500 35460 52502
rect 35532 52332 35588 52388
rect 34860 51378 34916 51380
rect 34860 51326 34862 51378
rect 34862 51326 34914 51378
rect 34914 51326 34916 51378
rect 34860 51324 34916 51326
rect 34860 50428 34916 50484
rect 34748 49980 34804 50036
rect 35196 52220 35252 52276
rect 36092 53004 36148 53060
rect 36204 53900 36260 53956
rect 35980 52332 36036 52388
rect 36764 53788 36820 53844
rect 36876 54124 36932 54180
rect 36316 52780 36372 52836
rect 37436 54012 37492 54068
rect 37100 53564 37156 53620
rect 36988 53058 37044 53060
rect 36988 53006 36990 53058
rect 36990 53006 37042 53058
rect 37042 53006 37044 53058
rect 36988 53004 37044 53006
rect 36428 51884 36484 51940
rect 36540 51996 36596 52052
rect 36316 51772 36372 51828
rect 36316 51548 36372 51604
rect 35532 51490 35588 51492
rect 35532 51438 35534 51490
rect 35534 51438 35586 51490
rect 35586 51438 35588 51490
rect 35532 51436 35588 51438
rect 35196 50986 35252 50988
rect 35196 50934 35198 50986
rect 35198 50934 35250 50986
rect 35250 50934 35252 50986
rect 35196 50932 35252 50934
rect 35300 50986 35356 50988
rect 35300 50934 35302 50986
rect 35302 50934 35354 50986
rect 35354 50934 35356 50986
rect 35300 50932 35356 50934
rect 35404 50986 35460 50988
rect 35404 50934 35406 50986
rect 35406 50934 35458 50986
rect 35458 50934 35460 50986
rect 35404 50932 35460 50934
rect 35420 50764 35476 50820
rect 36428 51436 36484 51492
rect 35756 50540 35812 50596
rect 35532 50428 35588 50484
rect 35196 49418 35252 49420
rect 35196 49366 35198 49418
rect 35198 49366 35250 49418
rect 35250 49366 35252 49418
rect 35196 49364 35252 49366
rect 35300 49418 35356 49420
rect 35300 49366 35302 49418
rect 35302 49366 35354 49418
rect 35354 49366 35356 49418
rect 35300 49364 35356 49366
rect 35404 49418 35460 49420
rect 35404 49366 35406 49418
rect 35406 49366 35458 49418
rect 35458 49366 35460 49418
rect 35404 49364 35460 49366
rect 34524 49138 34580 49140
rect 34524 49086 34526 49138
rect 34526 49086 34578 49138
rect 34578 49086 34580 49138
rect 34524 49084 34580 49086
rect 35196 49026 35252 49028
rect 35196 48974 35198 49026
rect 35198 48974 35250 49026
rect 35250 48974 35252 49026
rect 35196 48972 35252 48974
rect 33740 48242 33796 48244
rect 33740 48190 33742 48242
rect 33742 48190 33794 48242
rect 33794 48190 33796 48242
rect 33740 48188 33796 48190
rect 32732 46732 32788 46788
rect 33068 46674 33124 46676
rect 33068 46622 33070 46674
rect 33070 46622 33122 46674
rect 33122 46622 33124 46674
rect 33068 46620 33124 46622
rect 33292 46956 33348 47012
rect 33516 46620 33572 46676
rect 35420 48636 35476 48692
rect 34860 48242 34916 48244
rect 34860 48190 34862 48242
rect 34862 48190 34914 48242
rect 34914 48190 34916 48242
rect 34860 48188 34916 48190
rect 34636 47516 34692 47572
rect 34860 46508 34916 46564
rect 35644 49868 35700 49924
rect 38556 55916 38612 55972
rect 37660 54572 37716 54628
rect 36876 51548 36932 51604
rect 37436 52108 37492 52164
rect 37324 51884 37380 51940
rect 37548 51884 37604 51940
rect 37436 51490 37492 51492
rect 37436 51438 37438 51490
rect 37438 51438 37490 51490
rect 37490 51438 37492 51490
rect 37436 51436 37492 51438
rect 37324 51324 37380 51380
rect 37996 53004 38052 53060
rect 37884 51884 37940 51940
rect 37772 51378 37828 51380
rect 37772 51326 37774 51378
rect 37774 51326 37826 51378
rect 37826 51326 37828 51378
rect 37772 51324 37828 51326
rect 37772 51100 37828 51156
rect 36204 49868 36260 49924
rect 35980 49420 36036 49476
rect 35756 48636 35812 48692
rect 35868 49196 35924 49252
rect 35644 48300 35700 48356
rect 35196 47850 35252 47852
rect 35196 47798 35198 47850
rect 35198 47798 35250 47850
rect 35250 47798 35252 47850
rect 35196 47796 35252 47798
rect 35300 47850 35356 47852
rect 35300 47798 35302 47850
rect 35302 47798 35354 47850
rect 35354 47798 35356 47850
rect 35300 47796 35356 47798
rect 35404 47850 35460 47852
rect 35404 47798 35406 47850
rect 35406 47798 35458 47850
rect 35458 47798 35460 47850
rect 35404 47796 35460 47798
rect 35084 47068 35140 47124
rect 35532 47068 35588 47124
rect 33740 45106 33796 45108
rect 33740 45054 33742 45106
rect 33742 45054 33794 45106
rect 33794 45054 33796 45106
rect 33740 45052 33796 45054
rect 32060 43708 32116 43764
rect 32284 44380 32340 44436
rect 31724 42588 31780 42644
rect 31836 41970 31892 41972
rect 31836 41918 31838 41970
rect 31838 41918 31890 41970
rect 31890 41918 31892 41970
rect 31836 41916 31892 41918
rect 29596 37436 29652 37492
rect 29820 37938 29876 37940
rect 29820 37886 29822 37938
rect 29822 37886 29874 37938
rect 29874 37886 29876 37938
rect 29820 37884 29876 37886
rect 29484 37100 29540 37156
rect 29372 36428 29428 36484
rect 29148 36258 29204 36260
rect 29148 36206 29150 36258
rect 29150 36206 29202 36258
rect 29202 36206 29204 36258
rect 29148 36204 29204 36206
rect 27916 35308 27972 35364
rect 27916 34748 27972 34804
rect 27804 33458 27860 33460
rect 27804 33406 27806 33458
rect 27806 33406 27858 33458
rect 27858 33406 27860 33458
rect 27804 33404 27860 33406
rect 27692 32002 27748 32004
rect 27692 31950 27694 32002
rect 27694 31950 27746 32002
rect 27746 31950 27748 32002
rect 27692 31948 27748 31950
rect 28252 35532 28308 35588
rect 28140 34690 28196 34692
rect 28140 34638 28142 34690
rect 28142 34638 28194 34690
rect 28194 34638 28196 34690
rect 28140 34636 28196 34638
rect 28028 33068 28084 33124
rect 28364 35308 28420 35364
rect 28476 35084 28532 35140
rect 29372 35586 29428 35588
rect 29372 35534 29374 35586
rect 29374 35534 29426 35586
rect 29426 35534 29428 35586
rect 29372 35532 29428 35534
rect 29484 35420 29540 35476
rect 29596 35644 29652 35700
rect 29260 35084 29316 35140
rect 29372 34802 29428 34804
rect 29372 34750 29374 34802
rect 29374 34750 29426 34802
rect 29426 34750 29428 34802
rect 29372 34748 29428 34750
rect 29036 33404 29092 33460
rect 29932 37826 29988 37828
rect 29932 37774 29934 37826
rect 29934 37774 29986 37826
rect 29986 37774 29988 37826
rect 29932 37772 29988 37774
rect 29708 35084 29764 35140
rect 30268 35756 30324 35812
rect 30156 33404 30212 33460
rect 30156 33234 30212 33236
rect 30156 33182 30158 33234
rect 30158 33182 30210 33234
rect 30210 33182 30212 33234
rect 30156 33180 30212 33182
rect 27916 32172 27972 32228
rect 28028 31890 28084 31892
rect 28028 31838 28030 31890
rect 28030 31838 28082 31890
rect 28082 31838 28084 31890
rect 28028 31836 28084 31838
rect 27356 31666 27412 31668
rect 27356 31614 27358 31666
rect 27358 31614 27410 31666
rect 27410 31614 27412 31666
rect 27356 31612 27412 31614
rect 27244 30994 27300 30996
rect 27244 30942 27246 30994
rect 27246 30942 27298 30994
rect 27298 30942 27300 30994
rect 27244 30940 27300 30942
rect 27468 31164 27524 31220
rect 27356 30380 27412 30436
rect 27692 30156 27748 30212
rect 27580 30098 27636 30100
rect 27580 30046 27582 30098
rect 27582 30046 27634 30098
rect 27634 30046 27636 30098
rect 27580 30044 27636 30046
rect 27132 29484 27188 29540
rect 27020 29260 27076 29316
rect 27132 28476 27188 28532
rect 27468 29932 27524 29988
rect 28028 30044 28084 30100
rect 27692 29484 27748 29540
rect 28476 32732 28532 32788
rect 28252 31612 28308 31668
rect 28364 31724 28420 31780
rect 28476 31836 28532 31892
rect 29036 32172 29092 32228
rect 28588 30156 28644 30212
rect 27804 29820 27860 29876
rect 28028 29426 28084 29428
rect 28028 29374 28030 29426
rect 28030 29374 28082 29426
rect 28082 29374 28084 29426
rect 28028 29372 28084 29374
rect 27580 29260 27636 29316
rect 27692 28812 27748 28868
rect 26348 28364 26404 28420
rect 26796 27746 26852 27748
rect 26796 27694 26798 27746
rect 26798 27694 26850 27746
rect 26850 27694 26852 27746
rect 26796 27692 26852 27694
rect 26796 27468 26852 27524
rect 26572 27186 26628 27188
rect 26572 27134 26574 27186
rect 26574 27134 26626 27186
rect 26626 27134 26628 27186
rect 26572 27132 26628 27134
rect 25564 26514 25620 26516
rect 25564 26462 25566 26514
rect 25566 26462 25618 26514
rect 25618 26462 25620 26514
rect 25564 26460 25620 26462
rect 27356 28028 27412 28084
rect 26460 26514 26516 26516
rect 26460 26462 26462 26514
rect 26462 26462 26514 26514
rect 26514 26462 26516 26514
rect 26460 26460 26516 26462
rect 26684 26514 26740 26516
rect 26684 26462 26686 26514
rect 26686 26462 26738 26514
rect 26738 26462 26740 26514
rect 26684 26460 26740 26462
rect 25452 24332 25508 24388
rect 25116 24050 25172 24052
rect 25116 23998 25118 24050
rect 25118 23998 25170 24050
rect 25170 23998 25172 24050
rect 25116 23996 25172 23998
rect 24332 23884 24388 23940
rect 25452 23938 25508 23940
rect 25452 23886 25454 23938
rect 25454 23886 25506 23938
rect 25506 23886 25508 23938
rect 25452 23884 25508 23886
rect 24444 23324 24500 23380
rect 23660 22482 23716 22484
rect 23660 22430 23662 22482
rect 23662 22430 23714 22482
rect 23714 22430 23716 22482
rect 23660 22428 23716 22430
rect 24220 22428 24276 22484
rect 24668 23042 24724 23044
rect 24668 22990 24670 23042
rect 24670 22990 24722 23042
rect 24722 22990 24724 23042
rect 24668 22988 24724 22990
rect 24556 22540 24612 22596
rect 23212 22204 23268 22260
rect 23100 20972 23156 21028
rect 22876 20130 22932 20132
rect 22876 20078 22878 20130
rect 22878 20078 22930 20130
rect 22930 20078 22932 20130
rect 22876 20076 22932 20078
rect 23660 22146 23716 22148
rect 23660 22094 23662 22146
rect 23662 22094 23714 22146
rect 23714 22094 23716 22146
rect 23660 22092 23716 22094
rect 23548 21980 23604 22036
rect 25564 22370 25620 22372
rect 25564 22318 25566 22370
rect 25566 22318 25618 22370
rect 25618 22318 25620 22370
rect 25564 22316 25620 22318
rect 23548 21586 23604 21588
rect 23548 21534 23550 21586
rect 23550 21534 23602 21586
rect 23602 21534 23604 21586
rect 23548 21532 23604 21534
rect 23324 20578 23380 20580
rect 23324 20526 23326 20578
rect 23326 20526 23378 20578
rect 23378 20526 23380 20578
rect 23324 20524 23380 20526
rect 23548 20860 23604 20916
rect 22764 19628 22820 19684
rect 22204 19180 22260 19236
rect 22876 19234 22932 19236
rect 22876 19182 22878 19234
rect 22878 19182 22930 19234
rect 22930 19182 22932 19234
rect 22876 19180 22932 19182
rect 21756 19068 21812 19124
rect 24332 21644 24388 21700
rect 24556 21532 24612 21588
rect 24780 22092 24836 22148
rect 24444 20972 24500 21028
rect 24668 20076 24724 20132
rect 24444 19964 24500 20020
rect 24556 19852 24612 19908
rect 23436 18956 23492 19012
rect 21084 18396 21140 18452
rect 20748 16940 20804 16996
rect 20972 17500 21028 17556
rect 21756 16994 21812 16996
rect 21756 16942 21758 16994
rect 21758 16942 21810 16994
rect 21810 16942 21812 16994
rect 21756 16940 21812 16942
rect 20972 16828 21028 16884
rect 22204 17666 22260 17668
rect 22204 17614 22206 17666
rect 22206 17614 22258 17666
rect 22258 17614 22260 17666
rect 22204 17612 22260 17614
rect 22204 16828 22260 16884
rect 21644 16098 21700 16100
rect 21644 16046 21646 16098
rect 21646 16046 21698 16098
rect 21698 16046 21700 16098
rect 21644 16044 21700 16046
rect 21308 14588 21364 14644
rect 21420 14306 21476 14308
rect 21420 14254 21422 14306
rect 21422 14254 21474 14306
rect 21474 14254 21476 14306
rect 21420 14252 21476 14254
rect 19628 12908 19684 12964
rect 20636 13580 20692 13636
rect 20076 12850 20132 12852
rect 20076 12798 20078 12850
rect 20078 12798 20130 12850
rect 20130 12798 20132 12850
rect 20076 12796 20132 12798
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 21756 13132 21812 13188
rect 20748 12908 20804 12964
rect 21420 12908 21476 12964
rect 19628 12236 19684 12292
rect 19628 11900 19684 11956
rect 20972 12012 21028 12068
rect 20412 11900 20468 11956
rect 18732 11282 18788 11284
rect 18732 11230 18734 11282
rect 18734 11230 18786 11282
rect 18786 11230 18788 11282
rect 18732 11228 18788 11230
rect 19404 10610 19460 10612
rect 19404 10558 19406 10610
rect 19406 10558 19458 10610
rect 19458 10558 19460 10610
rect 19404 10556 19460 10558
rect 16940 9714 16996 9716
rect 16940 9662 16942 9714
rect 16942 9662 16994 9714
rect 16994 9662 16996 9714
rect 16940 9660 16996 9662
rect 16268 8092 16324 8148
rect 16380 9602 16436 9604
rect 16380 9550 16382 9602
rect 16382 9550 16434 9602
rect 16434 9550 16436 9602
rect 16380 9548 16436 9550
rect 15596 7756 15652 7812
rect 16044 7474 16100 7476
rect 16044 7422 16046 7474
rect 16046 7422 16098 7474
rect 16098 7422 16100 7474
rect 16044 7420 16100 7422
rect 16716 8764 16772 8820
rect 17724 9548 17780 9604
rect 17836 9212 17892 9268
rect 17500 8930 17556 8932
rect 17500 8878 17502 8930
rect 17502 8878 17554 8930
rect 17554 8878 17556 8930
rect 17500 8876 17556 8878
rect 17948 8764 18004 8820
rect 17836 8092 17892 8148
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 20748 11394 20804 11396
rect 20748 11342 20750 11394
rect 20750 11342 20802 11394
rect 20802 11342 20804 11394
rect 20748 11340 20804 11342
rect 19180 9266 19236 9268
rect 19180 9214 19182 9266
rect 19182 9214 19234 9266
rect 19234 9214 19236 9266
rect 19180 9212 19236 9214
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 19516 9266 19572 9268
rect 19516 9214 19518 9266
rect 19518 9214 19570 9266
rect 19570 9214 19572 9266
rect 19516 9212 19572 9214
rect 21756 12796 21812 12852
rect 22092 12684 22148 12740
rect 22876 17666 22932 17668
rect 22876 17614 22878 17666
rect 22878 17614 22930 17666
rect 22930 17614 22932 17666
rect 22876 17612 22932 17614
rect 22764 17052 22820 17108
rect 22428 15820 22484 15876
rect 22764 14924 22820 14980
rect 23660 16044 23716 16100
rect 23324 15986 23380 15988
rect 23324 15934 23326 15986
rect 23326 15934 23378 15986
rect 23378 15934 23380 15986
rect 23324 15932 23380 15934
rect 22540 14252 22596 14308
rect 23100 14924 23156 14980
rect 23548 14642 23604 14644
rect 23548 14590 23550 14642
rect 23550 14590 23602 14642
rect 23602 14590 23604 14642
rect 23548 14588 23604 14590
rect 23324 13746 23380 13748
rect 23324 13694 23326 13746
rect 23326 13694 23378 13746
rect 23378 13694 23380 13746
rect 23324 13692 23380 13694
rect 22876 13634 22932 13636
rect 22876 13582 22878 13634
rect 22878 13582 22930 13634
rect 22930 13582 22932 13634
rect 22876 13580 22932 13582
rect 26572 26178 26628 26180
rect 26572 26126 26574 26178
rect 26574 26126 26626 26178
rect 26626 26126 26628 26178
rect 26572 26124 26628 26126
rect 27020 25618 27076 25620
rect 27020 25566 27022 25618
rect 27022 25566 27074 25618
rect 27074 25566 27076 25618
rect 27020 25564 27076 25566
rect 26460 24946 26516 24948
rect 26460 24894 26462 24946
rect 26462 24894 26514 24946
rect 26514 24894 26516 24946
rect 26460 24892 26516 24894
rect 26908 24892 26964 24948
rect 26236 23324 26292 23380
rect 28700 29650 28756 29652
rect 28700 29598 28702 29650
rect 28702 29598 28754 29650
rect 28754 29598 28756 29650
rect 28700 29596 28756 29598
rect 28476 29260 28532 29316
rect 29148 30044 29204 30100
rect 29148 29820 29204 29876
rect 29708 32844 29764 32900
rect 29820 32786 29876 32788
rect 29820 32734 29822 32786
rect 29822 32734 29874 32786
rect 29874 32734 29876 32786
rect 29820 32732 29876 32734
rect 29372 31778 29428 31780
rect 29372 31726 29374 31778
rect 29374 31726 29426 31778
rect 29426 31726 29428 31778
rect 29372 31724 29428 31726
rect 29820 32396 29876 32452
rect 29596 32172 29652 32228
rect 30156 31948 30212 32004
rect 29820 31836 29876 31892
rect 29484 29932 29540 29988
rect 28140 28028 28196 28084
rect 27580 27468 27636 27524
rect 27692 27692 27748 27748
rect 27580 27074 27636 27076
rect 27580 27022 27582 27074
rect 27582 27022 27634 27074
rect 27634 27022 27636 27074
rect 27580 27020 27636 27022
rect 28476 28418 28532 28420
rect 28476 28366 28478 28418
rect 28478 28366 28530 28418
rect 28530 28366 28532 28418
rect 28476 28364 28532 28366
rect 28364 27804 28420 27860
rect 28924 28364 28980 28420
rect 28700 27916 28756 27972
rect 27804 26850 27860 26852
rect 27804 26798 27806 26850
rect 27806 26798 27858 26850
rect 27858 26798 27860 26850
rect 27804 26796 27860 26798
rect 27468 26290 27524 26292
rect 27468 26238 27470 26290
rect 27470 26238 27522 26290
rect 27522 26238 27524 26290
rect 27468 26236 27524 26238
rect 27468 25618 27524 25620
rect 27468 25566 27470 25618
rect 27470 25566 27522 25618
rect 27522 25566 27524 25618
rect 27468 25564 27524 25566
rect 28140 25452 28196 25508
rect 27692 24892 27748 24948
rect 27468 23378 27524 23380
rect 27468 23326 27470 23378
rect 27470 23326 27522 23378
rect 27522 23326 27524 23378
rect 27468 23324 27524 23326
rect 26348 22204 26404 22260
rect 26012 21644 26068 21700
rect 26348 21586 26404 21588
rect 26348 21534 26350 21586
rect 26350 21534 26402 21586
rect 26402 21534 26404 21586
rect 26348 21532 26404 21534
rect 26012 20914 26068 20916
rect 26012 20862 26014 20914
rect 26014 20862 26066 20914
rect 26066 20862 26068 20914
rect 26012 20860 26068 20862
rect 24780 19852 24836 19908
rect 24780 18844 24836 18900
rect 25564 20130 25620 20132
rect 25564 20078 25566 20130
rect 25566 20078 25618 20130
rect 25618 20078 25620 20130
rect 25564 20076 25620 20078
rect 26684 21644 26740 21700
rect 27132 21586 27188 21588
rect 27132 21534 27134 21586
rect 27134 21534 27186 21586
rect 27186 21534 27188 21586
rect 27132 21532 27188 21534
rect 27356 22204 27412 22260
rect 28028 22594 28084 22596
rect 28028 22542 28030 22594
rect 28030 22542 28082 22594
rect 28082 22542 28084 22594
rect 28028 22540 28084 22542
rect 27916 22428 27972 22484
rect 27468 21586 27524 21588
rect 27468 21534 27470 21586
rect 27470 21534 27522 21586
rect 27522 21534 27524 21586
rect 27468 21532 27524 21534
rect 27692 20914 27748 20916
rect 27692 20862 27694 20914
rect 27694 20862 27746 20914
rect 27746 20862 27748 20914
rect 27692 20860 27748 20862
rect 28028 21362 28084 21364
rect 28028 21310 28030 21362
rect 28030 21310 28082 21362
rect 28082 21310 28084 21362
rect 28028 21308 28084 21310
rect 26572 20076 26628 20132
rect 25228 20018 25284 20020
rect 25228 19966 25230 20018
rect 25230 19966 25282 20018
rect 25282 19966 25284 20018
rect 25228 19964 25284 19966
rect 26124 19852 26180 19908
rect 26012 19234 26068 19236
rect 26012 19182 26014 19234
rect 26014 19182 26066 19234
rect 26066 19182 26068 19234
rect 26012 19180 26068 19182
rect 24556 18674 24612 18676
rect 24556 18622 24558 18674
rect 24558 18622 24610 18674
rect 24610 18622 24612 18674
rect 24556 18620 24612 18622
rect 24444 18562 24500 18564
rect 24444 18510 24446 18562
rect 24446 18510 24498 18562
rect 24498 18510 24500 18562
rect 24444 18508 24500 18510
rect 24780 18450 24836 18452
rect 24780 18398 24782 18450
rect 24782 18398 24834 18450
rect 24834 18398 24836 18450
rect 24780 18396 24836 18398
rect 24332 17612 24388 17668
rect 25452 18844 25508 18900
rect 25004 17612 25060 17668
rect 25228 18620 25284 18676
rect 24444 16940 24500 16996
rect 24220 16098 24276 16100
rect 24220 16046 24222 16098
rect 24222 16046 24274 16098
rect 24274 16046 24276 16098
rect 24220 16044 24276 16046
rect 23884 15874 23940 15876
rect 23884 15822 23886 15874
rect 23886 15822 23938 15874
rect 23938 15822 23940 15874
rect 23884 15820 23940 15822
rect 23884 14588 23940 14644
rect 23436 13580 23492 13636
rect 22540 13468 22596 13524
rect 21868 11676 21924 11732
rect 21532 11394 21588 11396
rect 21532 11342 21534 11394
rect 21534 11342 21586 11394
rect 21586 11342 21588 11394
rect 21532 11340 21588 11342
rect 21532 9212 21588 9268
rect 20076 8428 20132 8484
rect 18284 7980 18340 8036
rect 20524 7980 20580 8036
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 19404 7586 19460 7588
rect 19404 7534 19406 7586
rect 19406 7534 19458 7586
rect 19458 7534 19460 7586
rect 19404 7532 19460 7534
rect 20300 7532 20356 7588
rect 16604 7474 16660 7476
rect 16604 7422 16606 7474
rect 16606 7422 16658 7474
rect 16658 7422 16660 7474
rect 16604 7420 16660 7422
rect 18172 7474 18228 7476
rect 18172 7422 18174 7474
rect 18174 7422 18226 7474
rect 18226 7422 18228 7474
rect 18172 7420 18228 7422
rect 15260 6300 15316 6356
rect 16156 6524 16212 6580
rect 16492 6636 16548 6692
rect 18060 6802 18116 6804
rect 18060 6750 18062 6802
rect 18062 6750 18114 6802
rect 18114 6750 18116 6802
rect 18060 6748 18116 6750
rect 17276 6690 17332 6692
rect 17276 6638 17278 6690
rect 17278 6638 17330 6690
rect 17330 6638 17332 6690
rect 17276 6636 17332 6638
rect 16492 6412 16548 6468
rect 17724 6466 17780 6468
rect 17724 6414 17726 6466
rect 17726 6414 17778 6466
rect 17778 6414 17780 6466
rect 17724 6412 17780 6414
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 19964 7474 20020 7476
rect 19964 7422 19966 7474
rect 19966 7422 20018 7474
rect 20018 7422 20020 7474
rect 19964 7420 20020 7422
rect 18732 6690 18788 6692
rect 18732 6638 18734 6690
rect 18734 6638 18786 6690
rect 18786 6638 18788 6690
rect 18732 6636 18788 6638
rect 18396 5740 18452 5796
rect 19404 6636 19460 6692
rect 20524 6636 20580 6692
rect 20188 6412 20244 6468
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 20748 5852 20804 5908
rect 20524 5516 20580 5572
rect 21756 8204 21812 8260
rect 21868 8428 21924 8484
rect 21644 5906 21700 5908
rect 21644 5854 21646 5906
rect 21646 5854 21698 5906
rect 21698 5854 21700 5906
rect 21644 5852 21700 5854
rect 20860 5740 20916 5796
rect 21868 5516 21924 5572
rect 23884 13468 23940 13524
rect 24108 13746 24164 13748
rect 24108 13694 24110 13746
rect 24110 13694 24162 13746
rect 24162 13694 24164 13746
rect 24108 13692 24164 13694
rect 23996 13132 24052 13188
rect 23100 12684 23156 12740
rect 22988 12012 23044 12068
rect 22092 8988 22148 9044
rect 23324 12290 23380 12292
rect 23324 12238 23326 12290
rect 23326 12238 23378 12290
rect 23378 12238 23380 12290
rect 23324 12236 23380 12238
rect 23100 11900 23156 11956
rect 23996 12066 24052 12068
rect 23996 12014 23998 12066
rect 23998 12014 24050 12066
rect 24050 12014 24052 12066
rect 23996 12012 24052 12014
rect 23436 9884 23492 9940
rect 23660 9772 23716 9828
rect 23996 10050 24052 10052
rect 23996 9998 23998 10050
rect 23998 9998 24050 10050
rect 24050 9998 24052 10050
rect 23996 9996 24052 9998
rect 23660 9042 23716 9044
rect 23660 8990 23662 9042
rect 23662 8990 23714 9042
rect 23714 8990 23716 9042
rect 23660 8988 23716 8990
rect 25116 16098 25172 16100
rect 25116 16046 25118 16098
rect 25118 16046 25170 16098
rect 25170 16046 25172 16098
rect 25116 16044 25172 16046
rect 25340 18396 25396 18452
rect 26572 18674 26628 18676
rect 26572 18622 26574 18674
rect 26574 18622 26626 18674
rect 26626 18622 26628 18674
rect 26572 18620 26628 18622
rect 25788 18284 25844 18340
rect 27020 19010 27076 19012
rect 27020 18958 27022 19010
rect 27022 18958 27074 19010
rect 27074 18958 27076 19010
rect 27020 18956 27076 18958
rect 26796 18396 26852 18452
rect 26908 18284 26964 18340
rect 25788 17666 25844 17668
rect 25788 17614 25790 17666
rect 25790 17614 25842 17666
rect 25842 17614 25844 17666
rect 25788 17612 25844 17614
rect 26012 17836 26068 17892
rect 26796 17836 26852 17892
rect 24668 15202 24724 15204
rect 24668 15150 24670 15202
rect 24670 15150 24722 15202
rect 24722 15150 24724 15202
rect 24668 15148 24724 15150
rect 26012 15708 26068 15764
rect 25452 15484 25508 15540
rect 26012 15484 26068 15540
rect 25564 15260 25620 15316
rect 24668 12684 24724 12740
rect 24332 12178 24388 12180
rect 24332 12126 24334 12178
rect 24334 12126 24386 12178
rect 24386 12126 24388 12178
rect 24332 12124 24388 12126
rect 24332 11900 24388 11956
rect 25452 12178 25508 12180
rect 25452 12126 25454 12178
rect 25454 12126 25506 12178
rect 25506 12126 25508 12178
rect 25452 12124 25508 12126
rect 25340 12012 25396 12068
rect 25900 15148 25956 15204
rect 26572 16828 26628 16884
rect 28252 20130 28308 20132
rect 28252 20078 28254 20130
rect 28254 20078 28306 20130
rect 28306 20078 28308 20130
rect 28252 20076 28308 20078
rect 28028 19234 28084 19236
rect 28028 19182 28030 19234
rect 28030 19182 28082 19234
rect 28082 19182 28084 19234
rect 28028 19180 28084 19182
rect 27356 18396 27412 18452
rect 27468 18284 27524 18340
rect 27356 18172 27412 18228
rect 27244 17948 27300 18004
rect 26908 16828 26964 16884
rect 26348 15596 26404 15652
rect 27244 15314 27300 15316
rect 27244 15262 27246 15314
rect 27246 15262 27298 15314
rect 27298 15262 27300 15314
rect 27244 15260 27300 15262
rect 26460 15148 26516 15204
rect 26572 13858 26628 13860
rect 26572 13806 26574 13858
rect 26574 13806 26626 13858
rect 26626 13806 26628 13858
rect 26572 13804 26628 13806
rect 26124 12850 26180 12852
rect 26124 12798 26126 12850
rect 26126 12798 26178 12850
rect 26178 12798 26180 12850
rect 26124 12796 26180 12798
rect 25900 12236 25956 12292
rect 24108 9884 24164 9940
rect 24332 9660 24388 9716
rect 22876 8370 22932 8372
rect 22876 8318 22878 8370
rect 22878 8318 22930 8370
rect 22930 8318 22932 8370
rect 22876 8316 22932 8318
rect 24220 8988 24276 9044
rect 22428 8258 22484 8260
rect 22428 8206 22430 8258
rect 22430 8206 22482 8258
rect 22482 8206 22484 8258
rect 22428 8204 22484 8206
rect 23436 8204 23492 8260
rect 24444 8204 24500 8260
rect 23548 7420 23604 7476
rect 22204 6802 22260 6804
rect 22204 6750 22206 6802
rect 22206 6750 22258 6802
rect 22258 6750 22260 6802
rect 22204 6748 22260 6750
rect 22092 6690 22148 6692
rect 22092 6638 22094 6690
rect 22094 6638 22146 6690
rect 22146 6638 22148 6690
rect 22092 6636 22148 6638
rect 23996 6802 24052 6804
rect 23996 6750 23998 6802
rect 23998 6750 24050 6802
rect 24050 6750 24052 6802
rect 23996 6748 24052 6750
rect 22540 6690 22596 6692
rect 22540 6638 22542 6690
rect 22542 6638 22594 6690
rect 22594 6638 22596 6690
rect 22540 6636 22596 6638
rect 22428 6524 22484 6580
rect 24108 6690 24164 6692
rect 24108 6638 24110 6690
rect 24110 6638 24162 6690
rect 24162 6638 24164 6690
rect 24108 6636 24164 6638
rect 23660 6578 23716 6580
rect 23660 6526 23662 6578
rect 23662 6526 23714 6578
rect 23714 6526 23716 6578
rect 23660 6524 23716 6526
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 25452 9996 25508 10052
rect 24780 9884 24836 9940
rect 24892 9212 24948 9268
rect 25228 9042 25284 9044
rect 25228 8990 25230 9042
rect 25230 8990 25282 9042
rect 25282 8990 25284 9042
rect 25228 8988 25284 8990
rect 25900 9996 25956 10052
rect 25900 9826 25956 9828
rect 25900 9774 25902 9826
rect 25902 9774 25954 9826
rect 25954 9774 25956 9826
rect 25900 9772 25956 9774
rect 26908 12236 26964 12292
rect 27244 14476 27300 14532
rect 27020 12178 27076 12180
rect 27020 12126 27022 12178
rect 27022 12126 27074 12178
rect 27074 12126 27076 12178
rect 27020 12124 27076 12126
rect 26236 11676 26292 11732
rect 26236 9714 26292 9716
rect 26236 9662 26238 9714
rect 26238 9662 26290 9714
rect 26290 9662 26292 9714
rect 26236 9660 26292 9662
rect 26908 9772 26964 9828
rect 26012 9212 26068 9268
rect 25564 8258 25620 8260
rect 25564 8206 25566 8258
rect 25566 8206 25618 8258
rect 25618 8206 25620 8258
rect 25564 8204 25620 8206
rect 26572 8316 26628 8372
rect 24780 6524 24836 6580
rect 25452 7420 25508 7476
rect 26796 8092 26852 8148
rect 26572 7586 26628 7588
rect 26572 7534 26574 7586
rect 26574 7534 26626 7586
rect 26626 7534 26628 7586
rect 26572 7532 26628 7534
rect 26012 7308 26068 7364
rect 28252 18508 28308 18564
rect 27692 18396 27748 18452
rect 28140 17106 28196 17108
rect 28140 17054 28142 17106
rect 28142 17054 28194 17106
rect 28194 17054 28196 17106
rect 28140 17052 28196 17054
rect 28028 16882 28084 16884
rect 28028 16830 28030 16882
rect 28030 16830 28082 16882
rect 28082 16830 28084 16882
rect 28028 16828 28084 16830
rect 28028 16604 28084 16660
rect 27580 16098 27636 16100
rect 27580 16046 27582 16098
rect 27582 16046 27634 16098
rect 27634 16046 27636 16098
rect 27580 16044 27636 16046
rect 28700 22428 28756 22484
rect 29484 28588 29540 28644
rect 29372 27970 29428 27972
rect 29372 27918 29374 27970
rect 29374 27918 29426 27970
rect 29426 27918 29428 27970
rect 29372 27916 29428 27918
rect 31948 41186 32004 41188
rect 31948 41134 31950 41186
rect 31950 41134 32002 41186
rect 32002 41134 32004 41186
rect 31948 41132 32004 41134
rect 31052 39788 31108 39844
rect 31836 40962 31892 40964
rect 31836 40910 31838 40962
rect 31838 40910 31890 40962
rect 31890 40910 31892 40962
rect 31836 40908 31892 40910
rect 32396 41916 32452 41972
rect 32284 41186 32340 41188
rect 32284 41134 32286 41186
rect 32286 41134 32338 41186
rect 32338 41134 32340 41186
rect 32284 41132 32340 41134
rect 32508 40962 32564 40964
rect 32508 40910 32510 40962
rect 32510 40910 32562 40962
rect 32562 40910 32564 40962
rect 32508 40908 32564 40910
rect 30828 39004 30884 39060
rect 31164 39058 31220 39060
rect 31164 39006 31166 39058
rect 31166 39006 31218 39058
rect 31218 39006 31220 39058
rect 31164 39004 31220 39006
rect 30492 37826 30548 37828
rect 30492 37774 30494 37826
rect 30494 37774 30546 37826
rect 30546 37774 30548 37826
rect 30492 37772 30548 37774
rect 30492 37100 30548 37156
rect 30940 37436 30996 37492
rect 30380 34972 30436 35028
rect 31612 37490 31668 37492
rect 31612 37438 31614 37490
rect 31614 37438 31666 37490
rect 31666 37438 31668 37490
rect 31612 37436 31668 37438
rect 31164 37154 31220 37156
rect 31164 37102 31166 37154
rect 31166 37102 31218 37154
rect 31218 37102 31220 37154
rect 31164 37100 31220 37102
rect 31612 36370 31668 36372
rect 31612 36318 31614 36370
rect 31614 36318 31666 36370
rect 31666 36318 31668 36370
rect 31612 36316 31668 36318
rect 30604 34748 30660 34804
rect 31052 34972 31108 35028
rect 31276 34076 31332 34132
rect 31612 34242 31668 34244
rect 31612 34190 31614 34242
rect 31614 34190 31666 34242
rect 31666 34190 31668 34242
rect 31612 34188 31668 34190
rect 31388 33740 31444 33796
rect 31164 33234 31220 33236
rect 31164 33182 31166 33234
rect 31166 33182 31218 33234
rect 31218 33182 31220 33234
rect 31164 33180 31220 33182
rect 30492 32844 30548 32900
rect 30716 31948 30772 32004
rect 31500 32450 31556 32452
rect 31500 32398 31502 32450
rect 31502 32398 31554 32450
rect 31554 32398 31556 32450
rect 31500 32396 31556 32398
rect 32508 40290 32564 40292
rect 32508 40238 32510 40290
rect 32510 40238 32562 40290
rect 32562 40238 32564 40290
rect 32508 40236 32564 40238
rect 32172 36316 32228 36372
rect 32732 39004 32788 39060
rect 32396 38556 32452 38612
rect 32396 37436 32452 37492
rect 32732 37436 32788 37492
rect 33180 43148 33236 43204
rect 33516 44994 33572 44996
rect 33516 44942 33518 44994
rect 33518 44942 33570 44994
rect 33570 44942 33572 44994
rect 33516 44940 33572 44942
rect 33516 44156 33572 44212
rect 33292 42812 33348 42868
rect 34412 44210 34468 44212
rect 34412 44158 34414 44210
rect 34414 44158 34466 44210
rect 34466 44158 34468 44210
rect 34412 44156 34468 44158
rect 33628 43708 33684 43764
rect 33404 41916 33460 41972
rect 33292 41858 33348 41860
rect 33292 41806 33294 41858
rect 33294 41806 33346 41858
rect 33346 41806 33348 41858
rect 33292 41804 33348 41806
rect 33292 41186 33348 41188
rect 33292 41134 33294 41186
rect 33294 41134 33346 41186
rect 33346 41134 33348 41186
rect 33292 41132 33348 41134
rect 34076 43650 34132 43652
rect 34076 43598 34078 43650
rect 34078 43598 34130 43650
rect 34130 43598 34132 43650
rect 34076 43596 34132 43598
rect 33740 43484 33796 43540
rect 34860 45164 34916 45220
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 35308 46060 35364 46116
rect 35308 45164 35364 45220
rect 34972 45052 35028 45108
rect 35532 44828 35588 44884
rect 36092 49026 36148 49028
rect 36092 48974 36094 49026
rect 36094 48974 36146 49026
rect 36146 48974 36148 49026
rect 36092 48972 36148 48974
rect 36092 48748 36148 48804
rect 35644 44940 35700 44996
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 34972 44434 35028 44436
rect 34972 44382 34974 44434
rect 34974 44382 35026 44434
rect 35026 44382 35028 44434
rect 34972 44380 35028 44382
rect 35532 44380 35588 44436
rect 36876 49868 36932 49924
rect 36764 49420 36820 49476
rect 36988 49026 37044 49028
rect 36988 48974 36990 49026
rect 36990 48974 37042 49026
rect 37042 48974 37044 49026
rect 36988 48972 37044 48974
rect 36764 48860 36820 48916
rect 37548 50764 37604 50820
rect 37772 50540 37828 50596
rect 38780 55020 38836 55076
rect 38556 53452 38612 53508
rect 38780 53058 38836 53060
rect 38780 53006 38782 53058
rect 38782 53006 38834 53058
rect 38834 53006 38836 53058
rect 38780 53004 38836 53006
rect 39228 56082 39284 56084
rect 39228 56030 39230 56082
rect 39230 56030 39282 56082
rect 39282 56030 39284 56082
rect 39228 56028 39284 56030
rect 39228 55244 39284 55300
rect 39452 55132 39508 55188
rect 38892 52892 38948 52948
rect 38444 51938 38500 51940
rect 38444 51886 38446 51938
rect 38446 51886 38498 51938
rect 38498 51886 38500 51938
rect 38444 51884 38500 51886
rect 38668 51772 38724 51828
rect 38332 51436 38388 51492
rect 37324 49644 37380 49700
rect 37212 49420 37268 49476
rect 37100 48524 37156 48580
rect 37100 48242 37156 48244
rect 37100 48190 37102 48242
rect 37102 48190 37154 48242
rect 37154 48190 37156 48242
rect 37100 48188 37156 48190
rect 37660 49420 37716 49476
rect 37772 49868 37828 49924
rect 37436 48802 37492 48804
rect 37436 48750 37438 48802
rect 37438 48750 37490 48802
rect 37490 48750 37492 48802
rect 37436 48748 37492 48750
rect 37548 49084 37604 49140
rect 36988 46674 37044 46676
rect 36988 46622 36990 46674
rect 36990 46622 37042 46674
rect 37042 46622 37044 46674
rect 36988 46620 37044 46622
rect 37772 48860 37828 48916
rect 38108 49868 38164 49924
rect 37996 48914 38052 48916
rect 37996 48862 37998 48914
rect 37998 48862 38050 48914
rect 38050 48862 38052 48914
rect 37996 48860 38052 48862
rect 38332 50540 38388 50596
rect 38332 49644 38388 49700
rect 38332 49026 38388 49028
rect 38332 48974 38334 49026
rect 38334 48974 38386 49026
rect 38386 48974 38388 49026
rect 38332 48972 38388 48974
rect 36316 46060 36372 46116
rect 36092 45612 36148 45668
rect 36204 45388 36260 45444
rect 38108 47458 38164 47460
rect 38108 47406 38110 47458
rect 38110 47406 38162 47458
rect 38162 47406 38164 47458
rect 38108 47404 38164 47406
rect 36428 45778 36484 45780
rect 36428 45726 36430 45778
rect 36430 45726 36482 45778
rect 36482 45726 36484 45778
rect 36428 45724 36484 45726
rect 37100 45666 37156 45668
rect 37100 45614 37102 45666
rect 37102 45614 37154 45666
rect 37154 45614 37156 45666
rect 37100 45612 37156 45614
rect 36764 45276 36820 45332
rect 34748 43260 34804 43316
rect 36204 43708 36260 43764
rect 34524 42866 34580 42868
rect 34524 42814 34526 42866
rect 34526 42814 34578 42866
rect 34578 42814 34580 42866
rect 34524 42812 34580 42814
rect 34748 42812 34804 42868
rect 36092 43596 36148 43652
rect 35980 43260 36036 43316
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 35868 43148 35924 43204
rect 34860 42588 34916 42644
rect 35756 42642 35812 42644
rect 35756 42590 35758 42642
rect 35758 42590 35810 42642
rect 35810 42590 35812 42642
rect 35756 42588 35812 42590
rect 36204 43538 36260 43540
rect 36204 43486 36206 43538
rect 36206 43486 36258 43538
rect 36258 43486 36260 43538
rect 36204 43484 36260 43486
rect 37100 43708 37156 43764
rect 36876 43426 36932 43428
rect 36876 43374 36878 43426
rect 36878 43374 36930 43426
rect 36930 43374 36932 43426
rect 36876 43372 36932 43374
rect 34748 41804 34804 41860
rect 33516 41020 33572 41076
rect 33852 40908 33908 40964
rect 33292 40402 33348 40404
rect 33292 40350 33294 40402
rect 33294 40350 33346 40402
rect 33346 40350 33348 40402
rect 33292 40348 33348 40350
rect 33180 38556 33236 38612
rect 32956 36764 33012 36820
rect 33180 36540 33236 36596
rect 31948 35196 32004 35252
rect 32060 34802 32116 34804
rect 32060 34750 32062 34802
rect 32062 34750 32114 34802
rect 32114 34750 32116 34802
rect 32060 34748 32116 34750
rect 32172 34300 32228 34356
rect 32172 34130 32228 34132
rect 32172 34078 32174 34130
rect 32174 34078 32226 34130
rect 32226 34078 32228 34130
rect 32172 34076 32228 34078
rect 31948 33852 32004 33908
rect 31948 33628 32004 33684
rect 31948 33122 32004 33124
rect 31948 33070 31950 33122
rect 31950 33070 32002 33122
rect 32002 33070 32004 33122
rect 31948 33068 32004 33070
rect 32172 32620 32228 32676
rect 31836 31836 31892 31892
rect 30716 30940 30772 30996
rect 30492 30210 30548 30212
rect 30492 30158 30494 30210
rect 30494 30158 30546 30210
rect 30546 30158 30548 30210
rect 30492 30156 30548 30158
rect 30380 29820 30436 29876
rect 30604 29932 30660 29988
rect 30156 29708 30212 29764
rect 30828 30492 30884 30548
rect 30716 29596 30772 29652
rect 31500 31164 31556 31220
rect 31836 30882 31892 30884
rect 31836 30830 31838 30882
rect 31838 30830 31890 30882
rect 31890 30830 31892 30882
rect 31836 30828 31892 30830
rect 31500 30716 31556 30772
rect 32396 33852 32452 33908
rect 32956 34354 33012 34356
rect 32956 34302 32958 34354
rect 32958 34302 33010 34354
rect 33010 34302 33012 34354
rect 32956 34300 33012 34302
rect 33292 35308 33348 35364
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 34636 41074 34692 41076
rect 34636 41022 34638 41074
rect 34638 41022 34690 41074
rect 34690 41022 34692 41074
rect 34636 41020 34692 41022
rect 34412 40962 34468 40964
rect 34412 40910 34414 40962
rect 34414 40910 34466 40962
rect 34466 40910 34468 40962
rect 34412 40908 34468 40910
rect 34076 40402 34132 40404
rect 34076 40350 34078 40402
rect 34078 40350 34130 40402
rect 34130 40350 34132 40402
rect 34076 40348 34132 40350
rect 34412 40290 34468 40292
rect 34412 40238 34414 40290
rect 34414 40238 34466 40290
rect 34466 40238 34468 40290
rect 34412 40236 34468 40238
rect 35420 40626 35476 40628
rect 35420 40574 35422 40626
rect 35422 40574 35474 40626
rect 35474 40574 35476 40626
rect 35420 40572 35476 40574
rect 35308 40236 35364 40292
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 33964 38668 34020 38724
rect 34748 38668 34804 38724
rect 33516 37490 33572 37492
rect 33516 37438 33518 37490
rect 33518 37438 33570 37490
rect 33570 37438 33572 37490
rect 33516 37436 33572 37438
rect 34300 38108 34356 38164
rect 34524 37436 34580 37492
rect 34188 36764 34244 36820
rect 33852 36594 33908 36596
rect 33852 36542 33854 36594
rect 33854 36542 33906 36594
rect 33906 36542 33908 36594
rect 33852 36540 33908 36542
rect 34412 36594 34468 36596
rect 34412 36542 34414 36594
rect 34414 36542 34466 36594
rect 34466 36542 34468 36594
rect 34412 36540 34468 36542
rect 33292 34690 33348 34692
rect 33292 34638 33294 34690
rect 33294 34638 33346 34690
rect 33346 34638 33348 34690
rect 33292 34636 33348 34638
rect 32620 34130 32676 34132
rect 32620 34078 32622 34130
rect 32622 34078 32674 34130
rect 32674 34078 32676 34130
rect 32620 34076 32676 34078
rect 32508 32620 32564 32676
rect 32732 33122 32788 33124
rect 32732 33070 32734 33122
rect 32734 33070 32786 33122
rect 32786 33070 32788 33122
rect 32732 33068 32788 33070
rect 32396 31052 32452 31108
rect 31500 30492 31556 30548
rect 31612 29932 31668 29988
rect 31276 29820 31332 29876
rect 31052 29596 31108 29652
rect 31164 29708 31220 29764
rect 31948 29650 32004 29652
rect 31948 29598 31950 29650
rect 31950 29598 32002 29650
rect 32002 29598 32004 29650
rect 31948 29596 32004 29598
rect 32284 29650 32340 29652
rect 32284 29598 32286 29650
rect 32286 29598 32338 29650
rect 32338 29598 32340 29650
rect 32284 29596 32340 29598
rect 31164 29484 31220 29540
rect 30380 28588 30436 28644
rect 29260 26908 29316 26964
rect 28588 21420 28644 21476
rect 29708 27074 29764 27076
rect 29708 27022 29710 27074
rect 29710 27022 29762 27074
rect 29762 27022 29764 27074
rect 29708 27020 29764 27022
rect 30380 27244 30436 27300
rect 30044 27020 30100 27076
rect 29708 26402 29764 26404
rect 29708 26350 29710 26402
rect 29710 26350 29762 26402
rect 29762 26350 29764 26402
rect 29708 26348 29764 26350
rect 29484 25900 29540 25956
rect 30604 28812 30660 28868
rect 31164 28754 31220 28756
rect 31164 28702 31166 28754
rect 31166 28702 31218 28754
rect 31218 28702 31220 28754
rect 31164 28700 31220 28702
rect 30828 28642 30884 28644
rect 30828 28590 30830 28642
rect 30830 28590 30882 28642
rect 30882 28590 30884 28642
rect 30828 28588 30884 28590
rect 31612 28642 31668 28644
rect 31612 28590 31614 28642
rect 31614 28590 31666 28642
rect 31666 28590 31668 28642
rect 31612 28588 31668 28590
rect 31724 28364 31780 28420
rect 30828 27074 30884 27076
rect 30828 27022 30830 27074
rect 30830 27022 30882 27074
rect 30882 27022 30884 27074
rect 30828 27020 30884 27022
rect 31388 27020 31444 27076
rect 30604 26684 30660 26740
rect 30492 25004 30548 25060
rect 29260 24892 29316 24948
rect 28588 20076 28644 20132
rect 28588 19180 28644 19236
rect 28364 18172 28420 18228
rect 28476 17948 28532 18004
rect 28364 17500 28420 17556
rect 27356 14140 27412 14196
rect 27580 14924 27636 14980
rect 27244 11228 27300 11284
rect 28812 18956 28868 19012
rect 29372 23324 29428 23380
rect 29260 22482 29316 22484
rect 29260 22430 29262 22482
rect 29262 22430 29314 22482
rect 29314 22430 29316 22482
rect 29260 22428 29316 22430
rect 29148 21474 29204 21476
rect 29148 21422 29150 21474
rect 29150 21422 29202 21474
rect 29202 21422 29204 21474
rect 29148 21420 29204 21422
rect 30380 24834 30436 24836
rect 30380 24782 30382 24834
rect 30382 24782 30434 24834
rect 30434 24782 30436 24834
rect 30380 24780 30436 24782
rect 30940 26402 30996 26404
rect 30940 26350 30942 26402
rect 30942 26350 30994 26402
rect 30994 26350 30996 26402
rect 30940 26348 30996 26350
rect 31164 26402 31220 26404
rect 31164 26350 31166 26402
rect 31166 26350 31218 26402
rect 31218 26350 31220 26402
rect 31164 26348 31220 26350
rect 30716 26290 30772 26292
rect 30716 26238 30718 26290
rect 30718 26238 30770 26290
rect 30770 26238 30772 26290
rect 30716 26236 30772 26238
rect 30828 25340 30884 25396
rect 31276 25452 31332 25508
rect 31164 25228 31220 25284
rect 30156 24220 30212 24276
rect 30268 24108 30324 24164
rect 30492 23938 30548 23940
rect 30492 23886 30494 23938
rect 30494 23886 30546 23938
rect 30546 23886 30548 23938
rect 30492 23884 30548 23886
rect 29708 23324 29764 23380
rect 29484 21756 29540 21812
rect 30492 22092 30548 22148
rect 29260 20524 29316 20580
rect 29372 19404 29428 19460
rect 29708 20578 29764 20580
rect 29708 20526 29710 20578
rect 29710 20526 29762 20578
rect 29762 20526 29764 20578
rect 29708 20524 29764 20526
rect 29708 19628 29764 19684
rect 30380 20076 30436 20132
rect 30044 20018 30100 20020
rect 30044 19966 30046 20018
rect 30046 19966 30098 20018
rect 30098 19966 30100 20018
rect 30044 19964 30100 19966
rect 30492 20018 30548 20020
rect 30492 19966 30494 20018
rect 30494 19966 30546 20018
rect 30546 19966 30548 20018
rect 30492 19964 30548 19966
rect 29820 19516 29876 19572
rect 29148 19234 29204 19236
rect 29148 19182 29150 19234
rect 29150 19182 29202 19234
rect 29202 19182 29204 19234
rect 29148 19180 29204 19182
rect 29260 18956 29316 19012
rect 28812 17724 28868 17780
rect 28700 17106 28756 17108
rect 28700 17054 28702 17106
rect 28702 17054 28754 17106
rect 28754 17054 28756 17106
rect 28700 17052 28756 17054
rect 28924 17106 28980 17108
rect 28924 17054 28926 17106
rect 28926 17054 28978 17106
rect 28978 17054 28980 17106
rect 28924 17052 28980 17054
rect 28476 14924 28532 14980
rect 31276 23826 31332 23828
rect 31276 23774 31278 23826
rect 31278 23774 31330 23826
rect 31330 23774 31332 23826
rect 31276 23772 31332 23774
rect 30828 23378 30884 23380
rect 30828 23326 30830 23378
rect 30830 23326 30882 23378
rect 30882 23326 30884 23378
rect 30828 23324 30884 23326
rect 30716 21980 30772 22036
rect 30828 23100 30884 23156
rect 30940 22988 30996 23044
rect 31724 27356 31780 27412
rect 31612 26348 31668 26404
rect 31500 26290 31556 26292
rect 31500 26238 31502 26290
rect 31502 26238 31554 26290
rect 31554 26238 31556 26290
rect 31500 26236 31556 26238
rect 31836 26290 31892 26292
rect 31836 26238 31838 26290
rect 31838 26238 31890 26290
rect 31890 26238 31892 26290
rect 31836 26236 31892 26238
rect 31836 25452 31892 25508
rect 31276 23100 31332 23156
rect 31500 25004 31556 25060
rect 31724 25004 31780 25060
rect 31724 24668 31780 24724
rect 31836 24556 31892 24612
rect 31948 25228 32004 25284
rect 31612 23938 31668 23940
rect 31612 23886 31614 23938
rect 31614 23886 31666 23938
rect 31666 23886 31668 23938
rect 31612 23884 31668 23886
rect 31052 22146 31108 22148
rect 31052 22094 31054 22146
rect 31054 22094 31106 22146
rect 31106 22094 31108 22146
rect 31052 22092 31108 22094
rect 31276 21308 31332 21364
rect 30716 20018 30772 20020
rect 30716 19966 30718 20018
rect 30718 19966 30770 20018
rect 30770 19966 30772 20018
rect 30716 19964 30772 19966
rect 31500 22370 31556 22372
rect 31500 22318 31502 22370
rect 31502 22318 31554 22370
rect 31554 22318 31556 22370
rect 31500 22316 31556 22318
rect 32508 30156 32564 30212
rect 32172 28364 32228 28420
rect 32172 28140 32228 28196
rect 32172 27468 32228 27524
rect 33068 32732 33124 32788
rect 33516 34188 33572 34244
rect 33292 34018 33348 34020
rect 33292 33966 33294 34018
rect 33294 33966 33346 34018
rect 33346 33966 33348 34018
rect 33292 33964 33348 33966
rect 32956 31948 33012 32004
rect 33180 31778 33236 31780
rect 33180 31726 33182 31778
rect 33182 31726 33234 31778
rect 33234 31726 33236 31778
rect 33180 31724 33236 31726
rect 33516 31666 33572 31668
rect 33516 31614 33518 31666
rect 33518 31614 33570 31666
rect 33570 31614 33572 31666
rect 33516 31612 33572 31614
rect 32844 29372 32900 29428
rect 33852 34802 33908 34804
rect 33852 34750 33854 34802
rect 33854 34750 33906 34802
rect 33906 34750 33908 34802
rect 33852 34748 33908 34750
rect 33740 34242 33796 34244
rect 33740 34190 33742 34242
rect 33742 34190 33794 34242
rect 33794 34190 33796 34242
rect 33740 34188 33796 34190
rect 33404 29596 33460 29652
rect 34636 35532 34692 35588
rect 34860 36988 34916 37044
rect 34860 35420 34916 35476
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 35308 38162 35364 38164
rect 35308 38110 35310 38162
rect 35310 38110 35362 38162
rect 35362 38110 35364 38162
rect 35308 38108 35364 38110
rect 35644 38108 35700 38164
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 36204 42252 36260 42308
rect 37436 45666 37492 45668
rect 37436 45614 37438 45666
rect 37438 45614 37490 45666
rect 37490 45614 37492 45666
rect 37436 45612 37492 45614
rect 37324 45388 37380 45444
rect 38332 46508 38388 46564
rect 38332 45612 38388 45668
rect 38220 45276 38276 45332
rect 38892 51548 38948 51604
rect 38556 51266 38612 51268
rect 38556 51214 38558 51266
rect 38558 51214 38610 51266
rect 38610 51214 38612 51266
rect 38556 51212 38612 51214
rect 38780 51100 38836 51156
rect 38556 49084 38612 49140
rect 39116 51602 39172 51604
rect 39116 51550 39118 51602
rect 39118 51550 39170 51602
rect 39170 51550 39172 51602
rect 39116 51548 39172 51550
rect 39340 53564 39396 53620
rect 39340 52892 39396 52948
rect 40236 55468 40292 55524
rect 39788 54124 39844 54180
rect 39564 53618 39620 53620
rect 39564 53566 39566 53618
rect 39566 53566 39618 53618
rect 39618 53566 39620 53618
rect 39564 53564 39620 53566
rect 38892 49922 38948 49924
rect 38892 49870 38894 49922
rect 38894 49870 38946 49922
rect 38946 49870 38948 49922
rect 38892 49868 38948 49870
rect 39228 49756 39284 49812
rect 39116 49084 39172 49140
rect 38892 48242 38948 48244
rect 38892 48190 38894 48242
rect 38894 48190 38946 48242
rect 38946 48190 38948 48242
rect 38892 48188 38948 48190
rect 38556 47404 38612 47460
rect 39004 46732 39060 46788
rect 38556 45890 38612 45892
rect 38556 45838 38558 45890
rect 38558 45838 38610 45890
rect 38610 45838 38612 45890
rect 38556 45836 38612 45838
rect 38780 45724 38836 45780
rect 38892 45836 38948 45892
rect 38556 45612 38612 45668
rect 37324 43650 37380 43652
rect 37324 43598 37326 43650
rect 37326 43598 37378 43650
rect 37378 43598 37380 43650
rect 37324 43596 37380 43598
rect 37212 43148 37268 43204
rect 37884 43372 37940 43428
rect 36988 42642 37044 42644
rect 36988 42590 36990 42642
rect 36990 42590 37042 42642
rect 37042 42590 37044 42642
rect 36988 42588 37044 42590
rect 36540 42476 36596 42532
rect 36316 41298 36372 41300
rect 36316 41246 36318 41298
rect 36318 41246 36370 41298
rect 36370 41246 36372 41298
rect 36316 41244 36372 41246
rect 37548 42530 37604 42532
rect 37548 42478 37550 42530
rect 37550 42478 37602 42530
rect 37602 42478 37604 42530
rect 37548 42476 37604 42478
rect 37548 42252 37604 42308
rect 36988 42194 37044 42196
rect 36988 42142 36990 42194
rect 36990 42142 37042 42194
rect 37042 42142 37044 42194
rect 36988 42140 37044 42142
rect 36764 40572 36820 40628
rect 37100 41020 37156 41076
rect 35868 38556 35924 38612
rect 37212 39506 37268 39508
rect 37212 39454 37214 39506
rect 37214 39454 37266 39506
rect 37266 39454 37268 39506
rect 37212 39452 37268 39454
rect 38108 41916 38164 41972
rect 37660 40348 37716 40404
rect 38444 43820 38500 43876
rect 39116 45724 39172 45780
rect 38668 44380 38724 44436
rect 38780 43932 38836 43988
rect 38556 41970 38612 41972
rect 38556 41918 38558 41970
rect 38558 41918 38610 41970
rect 38610 41918 38612 41970
rect 38556 41916 38612 41918
rect 38332 41020 38388 41076
rect 38556 40572 38612 40628
rect 38332 40402 38388 40404
rect 38332 40350 38334 40402
rect 38334 40350 38386 40402
rect 38386 40350 38388 40402
rect 38332 40348 38388 40350
rect 38556 40290 38612 40292
rect 38556 40238 38558 40290
rect 38558 40238 38610 40290
rect 38610 40238 38612 40290
rect 38556 40236 38612 40238
rect 38220 39730 38276 39732
rect 38220 39678 38222 39730
rect 38222 39678 38274 39730
rect 38274 39678 38276 39730
rect 38220 39676 38276 39678
rect 36540 38780 36596 38836
rect 36092 38050 36148 38052
rect 36092 37998 36094 38050
rect 36094 37998 36146 38050
rect 36146 37998 36148 38050
rect 36092 37996 36148 37998
rect 37436 38050 37492 38052
rect 37436 37998 37438 38050
rect 37438 37998 37490 38050
rect 37490 37998 37492 38050
rect 37436 37996 37492 37998
rect 35868 36988 35924 37044
rect 35756 36540 35812 36596
rect 36316 36204 36372 36260
rect 36316 35644 36372 35700
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 36428 35420 36484 35476
rect 33180 28812 33236 28868
rect 33292 28924 33348 28980
rect 33292 28642 33348 28644
rect 33292 28590 33294 28642
rect 33294 28590 33346 28642
rect 33346 28590 33348 28642
rect 33292 28588 33348 28590
rect 32844 28140 32900 28196
rect 33180 28140 33236 28196
rect 32732 27244 32788 27300
rect 33068 27468 33124 27524
rect 32620 27132 32676 27188
rect 32844 27132 32900 27188
rect 32172 26908 32228 26964
rect 32172 26402 32228 26404
rect 32172 26350 32174 26402
rect 32174 26350 32226 26402
rect 32226 26350 32228 26402
rect 32172 26348 32228 26350
rect 32172 25452 32228 25508
rect 32172 25282 32228 25284
rect 32172 25230 32174 25282
rect 32174 25230 32226 25282
rect 32226 25230 32228 25282
rect 32172 25228 32228 25230
rect 33068 26572 33124 26628
rect 34300 33740 34356 33796
rect 34412 33458 34468 33460
rect 34412 33406 34414 33458
rect 34414 33406 34466 33458
rect 34466 33406 34468 33458
rect 34412 33404 34468 33406
rect 35196 34802 35252 34804
rect 35196 34750 35198 34802
rect 35198 34750 35250 34802
rect 35250 34750 35252 34802
rect 35196 34748 35252 34750
rect 34972 34636 35028 34692
rect 35420 34354 35476 34356
rect 35420 34302 35422 34354
rect 35422 34302 35474 34354
rect 35474 34302 35476 34354
rect 35420 34300 35476 34302
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 33964 33068 34020 33124
rect 34188 31836 34244 31892
rect 33852 31778 33908 31780
rect 33852 31726 33854 31778
rect 33854 31726 33906 31778
rect 33906 31726 33908 31778
rect 33852 31724 33908 31726
rect 34076 31724 34132 31780
rect 34076 31554 34132 31556
rect 34076 31502 34078 31554
rect 34078 31502 34130 31554
rect 34130 31502 34132 31554
rect 34076 31500 34132 31502
rect 34972 33122 35028 33124
rect 34972 33070 34974 33122
rect 34974 33070 35026 33122
rect 35026 33070 35028 33122
rect 34972 33068 35028 33070
rect 34524 31836 34580 31892
rect 33852 30940 33908 30996
rect 34300 31276 34356 31332
rect 33740 29260 33796 29316
rect 33852 30716 33908 30772
rect 34188 31106 34244 31108
rect 34188 31054 34190 31106
rect 34190 31054 34242 31106
rect 34242 31054 34244 31106
rect 34188 31052 34244 31054
rect 34076 30994 34132 30996
rect 34076 30942 34078 30994
rect 34078 30942 34130 30994
rect 34130 30942 34132 30994
rect 34076 30940 34132 30942
rect 33964 30380 34020 30436
rect 34300 29986 34356 29988
rect 34300 29934 34302 29986
rect 34302 29934 34354 29986
rect 34354 29934 34356 29986
rect 34300 29932 34356 29934
rect 33516 27468 33572 27524
rect 33628 28082 33684 28084
rect 33628 28030 33630 28082
rect 33630 28030 33682 28082
rect 33682 28030 33684 28082
rect 33628 28028 33684 28030
rect 33964 29484 34020 29540
rect 34748 30828 34804 30884
rect 34860 32396 34916 32452
rect 35644 33516 35700 33572
rect 35980 34690 36036 34692
rect 35980 34638 35982 34690
rect 35982 34638 36034 34690
rect 36034 34638 36036 34690
rect 35980 34636 36036 34638
rect 35756 33292 35812 33348
rect 35868 33234 35924 33236
rect 35868 33182 35870 33234
rect 35870 33182 35922 33234
rect 35922 33182 35924 33234
rect 35868 33180 35924 33182
rect 35756 33122 35812 33124
rect 35756 33070 35758 33122
rect 35758 33070 35810 33122
rect 35810 33070 35812 33122
rect 35756 33068 35812 33070
rect 35196 32396 35252 32452
rect 35868 32956 35924 33012
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35308 31948 35364 32004
rect 35532 31836 35588 31892
rect 35196 31106 35252 31108
rect 35196 31054 35198 31106
rect 35198 31054 35250 31106
rect 35250 31054 35252 31106
rect 35196 31052 35252 31054
rect 35532 31052 35588 31108
rect 35980 31276 36036 31332
rect 36204 31052 36260 31108
rect 35308 30716 35364 30772
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 34524 29148 34580 29204
rect 34524 28476 34580 28532
rect 33404 27244 33460 27300
rect 33964 27074 34020 27076
rect 33964 27022 33966 27074
rect 33966 27022 34018 27074
rect 34018 27022 34020 27074
rect 33964 27020 34020 27022
rect 32508 25564 32564 25620
rect 33068 25900 33124 25956
rect 32620 25340 32676 25396
rect 32844 25340 32900 25396
rect 32508 24946 32564 24948
rect 32508 24894 32510 24946
rect 32510 24894 32562 24946
rect 32562 24894 32564 24946
rect 32508 24892 32564 24894
rect 32284 24780 32340 24836
rect 32060 23324 32116 23380
rect 32172 24556 32228 24612
rect 31724 22370 31780 22372
rect 31724 22318 31726 22370
rect 31726 22318 31778 22370
rect 31778 22318 31780 22370
rect 31724 22316 31780 22318
rect 32956 24780 33012 24836
rect 33852 26850 33908 26852
rect 33852 26798 33854 26850
rect 33854 26798 33906 26850
rect 33906 26798 33908 26850
rect 33852 26796 33908 26798
rect 33516 26402 33572 26404
rect 33516 26350 33518 26402
rect 33518 26350 33570 26402
rect 33570 26350 33572 26402
rect 33516 26348 33572 26350
rect 33404 26236 33460 26292
rect 33292 25564 33348 25620
rect 33404 25506 33460 25508
rect 33404 25454 33406 25506
rect 33406 25454 33458 25506
rect 33458 25454 33460 25506
rect 33404 25452 33460 25454
rect 33180 25394 33236 25396
rect 33180 25342 33182 25394
rect 33182 25342 33234 25394
rect 33234 25342 33236 25394
rect 33180 25340 33236 25342
rect 33292 23714 33348 23716
rect 33292 23662 33294 23714
rect 33294 23662 33346 23714
rect 33346 23662 33348 23714
rect 33292 23660 33348 23662
rect 33180 23548 33236 23604
rect 32172 21644 32228 21700
rect 32620 21644 32676 21700
rect 31724 20690 31780 20692
rect 31724 20638 31726 20690
rect 31726 20638 31778 20690
rect 31778 20638 31780 20690
rect 31724 20636 31780 20638
rect 30828 19404 30884 19460
rect 31612 20130 31668 20132
rect 31612 20078 31614 20130
rect 31614 20078 31666 20130
rect 31666 20078 31668 20130
rect 31612 20076 31668 20078
rect 31500 19516 31556 19572
rect 30044 18508 30100 18564
rect 29708 16658 29764 16660
rect 29708 16606 29710 16658
rect 29710 16606 29762 16658
rect 29762 16606 29764 16658
rect 29708 16604 29764 16606
rect 30604 18450 30660 18452
rect 30604 18398 30606 18450
rect 30606 18398 30658 18450
rect 30658 18398 30660 18450
rect 30604 18396 30660 18398
rect 31724 19628 31780 19684
rect 31612 19234 31668 19236
rect 31612 19182 31614 19234
rect 31614 19182 31666 19234
rect 31666 19182 31668 19234
rect 31612 19180 31668 19182
rect 31500 19122 31556 19124
rect 31500 19070 31502 19122
rect 31502 19070 31554 19122
rect 31554 19070 31556 19122
rect 31500 19068 31556 19070
rect 31500 18674 31556 18676
rect 31500 18622 31502 18674
rect 31502 18622 31554 18674
rect 31554 18622 31556 18674
rect 31500 18620 31556 18622
rect 31052 18284 31108 18340
rect 30380 17500 30436 17556
rect 30604 17724 30660 17780
rect 30156 16716 30212 16772
rect 29260 16268 29316 16324
rect 29148 15596 29204 15652
rect 28364 14530 28420 14532
rect 28364 14478 28366 14530
rect 28366 14478 28418 14530
rect 28418 14478 28420 14530
rect 28364 14476 28420 14478
rect 28252 13858 28308 13860
rect 28252 13806 28254 13858
rect 28254 13806 28306 13858
rect 28306 13806 28308 13858
rect 28252 13804 28308 13806
rect 28028 13468 28084 13524
rect 28028 12178 28084 12180
rect 28028 12126 28030 12178
rect 28030 12126 28082 12178
rect 28082 12126 28084 12178
rect 28028 12124 28084 12126
rect 28028 11676 28084 11732
rect 28028 11282 28084 11284
rect 28028 11230 28030 11282
rect 28030 11230 28082 11282
rect 28082 11230 28084 11282
rect 28028 11228 28084 11230
rect 28700 14252 28756 14308
rect 29484 14306 29540 14308
rect 29484 14254 29486 14306
rect 29486 14254 29538 14306
rect 29538 14254 29540 14306
rect 29484 14252 29540 14254
rect 28924 14140 28980 14196
rect 28588 13074 28644 13076
rect 28588 13022 28590 13074
rect 28590 13022 28642 13074
rect 28642 13022 28644 13074
rect 28588 13020 28644 13022
rect 28588 12684 28644 12740
rect 27580 9772 27636 9828
rect 27356 9660 27412 9716
rect 28140 10386 28196 10388
rect 28140 10334 28142 10386
rect 28142 10334 28194 10386
rect 28194 10334 28196 10386
rect 28140 10332 28196 10334
rect 27916 9884 27972 9940
rect 27692 9266 27748 9268
rect 27692 9214 27694 9266
rect 27694 9214 27746 9266
rect 27746 9214 27748 9266
rect 27692 9212 27748 9214
rect 27244 7474 27300 7476
rect 27244 7422 27246 7474
rect 27246 7422 27298 7474
rect 27298 7422 27300 7474
rect 27244 7420 27300 7422
rect 27020 7308 27076 7364
rect 26348 6748 26404 6804
rect 25340 6412 25396 6468
rect 28364 9884 28420 9940
rect 29484 12850 29540 12852
rect 29484 12798 29486 12850
rect 29486 12798 29538 12850
rect 29538 12798 29540 12850
rect 29484 12796 29540 12798
rect 29260 11788 29316 11844
rect 29372 10332 29428 10388
rect 29260 9938 29316 9940
rect 29260 9886 29262 9938
rect 29262 9886 29314 9938
rect 29314 9886 29316 9938
rect 29260 9884 29316 9886
rect 28588 9714 28644 9716
rect 28588 9662 28590 9714
rect 28590 9662 28642 9714
rect 28642 9662 28644 9714
rect 28588 9660 28644 9662
rect 28476 9212 28532 9268
rect 28476 8316 28532 8372
rect 28364 8258 28420 8260
rect 28364 8206 28366 8258
rect 28366 8206 28418 8258
rect 28418 8206 28420 8258
rect 28364 8204 28420 8206
rect 29148 9660 29204 9716
rect 29148 8146 29204 8148
rect 29148 8094 29150 8146
rect 29150 8094 29202 8146
rect 29202 8094 29204 8146
rect 29148 8092 29204 8094
rect 28028 7644 28084 7700
rect 27804 7586 27860 7588
rect 27804 7534 27806 7586
rect 27806 7534 27858 7586
rect 27858 7534 27860 7586
rect 27804 7532 27860 7534
rect 27692 7308 27748 7364
rect 28140 7420 28196 7476
rect 28588 5180 28644 5236
rect 28364 5122 28420 5124
rect 28364 5070 28366 5122
rect 28366 5070 28418 5122
rect 28418 5070 28420 5122
rect 28364 5068 28420 5070
rect 28700 4844 28756 4900
rect 28364 3442 28420 3444
rect 28364 3390 28366 3442
rect 28366 3390 28418 3442
rect 28418 3390 28420 3442
rect 28364 3388 28420 3390
rect 28476 4060 28532 4116
rect 29148 7474 29204 7476
rect 29148 7422 29150 7474
rect 29150 7422 29202 7474
rect 29202 7422 29204 7474
rect 29148 7420 29204 7422
rect 28924 7362 28980 7364
rect 28924 7310 28926 7362
rect 28926 7310 28978 7362
rect 28978 7310 28980 7362
rect 28924 7308 28980 7310
rect 29484 8652 29540 8708
rect 29372 8370 29428 8372
rect 29372 8318 29374 8370
rect 29374 8318 29426 8370
rect 29426 8318 29428 8370
rect 29372 8316 29428 8318
rect 28924 6748 28980 6804
rect 29708 15314 29764 15316
rect 29708 15262 29710 15314
rect 29710 15262 29762 15314
rect 29762 15262 29764 15314
rect 29708 15260 29764 15262
rect 30380 15874 30436 15876
rect 30380 15822 30382 15874
rect 30382 15822 30434 15874
rect 30434 15822 30436 15874
rect 30380 15820 30436 15822
rect 30492 15148 30548 15204
rect 29708 15036 29764 15092
rect 29708 14530 29764 14532
rect 29708 14478 29710 14530
rect 29710 14478 29762 14530
rect 29762 14478 29764 14530
rect 29708 14476 29764 14478
rect 30268 14530 30324 14532
rect 30268 14478 30270 14530
rect 30270 14478 30322 14530
rect 30322 14478 30324 14530
rect 30268 14476 30324 14478
rect 30044 14364 30100 14420
rect 30380 14252 30436 14308
rect 30268 12796 30324 12852
rect 30716 17612 30772 17668
rect 31052 17500 31108 17556
rect 31388 18284 31444 18340
rect 31388 17052 31444 17108
rect 31500 16828 31556 16884
rect 31836 18956 31892 19012
rect 31724 18620 31780 18676
rect 32060 19964 32116 20020
rect 32172 18620 32228 18676
rect 31836 18338 31892 18340
rect 31836 18286 31838 18338
rect 31838 18286 31890 18338
rect 31890 18286 31892 18338
rect 31836 18284 31892 18286
rect 30940 15314 30996 15316
rect 30940 15262 30942 15314
rect 30942 15262 30994 15314
rect 30994 15262 30996 15314
rect 30940 15260 30996 15262
rect 31276 15314 31332 15316
rect 31276 15262 31278 15314
rect 31278 15262 31330 15314
rect 31330 15262 31332 15314
rect 31276 15260 31332 15262
rect 31276 14530 31332 14532
rect 31276 14478 31278 14530
rect 31278 14478 31330 14530
rect 31330 14478 31332 14530
rect 31276 14476 31332 14478
rect 32060 16828 32116 16884
rect 31836 15820 31892 15876
rect 31612 15148 31668 15204
rect 31500 14476 31556 14532
rect 30380 11788 30436 11844
rect 29820 8316 29876 8372
rect 30716 9436 30772 9492
rect 30492 8316 30548 8372
rect 30268 8204 30324 8260
rect 30828 9266 30884 9268
rect 30828 9214 30830 9266
rect 30830 9214 30882 9266
rect 30882 9214 30884 9266
rect 30828 9212 30884 9214
rect 30604 8204 30660 8260
rect 30604 7474 30660 7476
rect 30604 7422 30606 7474
rect 30606 7422 30658 7474
rect 30658 7422 30660 7474
rect 30604 7420 30660 7422
rect 30268 7308 30324 7364
rect 32172 11788 32228 11844
rect 31948 10498 32004 10500
rect 31948 10446 31950 10498
rect 31950 10446 32002 10498
rect 32002 10446 32004 10498
rect 31948 10444 32004 10446
rect 32508 20914 32564 20916
rect 32508 20862 32510 20914
rect 32510 20862 32562 20914
rect 32562 20862 32564 20914
rect 32508 20860 32564 20862
rect 32732 21420 32788 21476
rect 32844 21756 32900 21812
rect 32620 20636 32676 20692
rect 33180 21810 33236 21812
rect 33180 21758 33182 21810
rect 33182 21758 33234 21810
rect 33234 21758 33236 21810
rect 33180 21756 33236 21758
rect 32844 20188 32900 20244
rect 33292 20018 33348 20020
rect 33292 19966 33294 20018
rect 33294 19966 33346 20018
rect 33346 19966 33348 20018
rect 33292 19964 33348 19966
rect 32732 19234 32788 19236
rect 32732 19182 32734 19234
rect 32734 19182 32786 19234
rect 32786 19182 32788 19234
rect 32732 19180 32788 19182
rect 32508 19122 32564 19124
rect 32508 19070 32510 19122
rect 32510 19070 32562 19122
rect 32562 19070 32564 19122
rect 32508 19068 32564 19070
rect 32732 18956 32788 19012
rect 33292 18674 33348 18676
rect 33292 18622 33294 18674
rect 33294 18622 33346 18674
rect 33346 18622 33348 18674
rect 33292 18620 33348 18622
rect 33628 23996 33684 24052
rect 33740 25340 33796 25396
rect 34076 26290 34132 26292
rect 34076 26238 34078 26290
rect 34078 26238 34130 26290
rect 34130 26238 34132 26290
rect 34076 26236 34132 26238
rect 33964 25676 34020 25732
rect 34076 26012 34132 26068
rect 34524 27692 34580 27748
rect 34748 28700 34804 28756
rect 34748 28418 34804 28420
rect 34748 28366 34750 28418
rect 34750 28366 34802 28418
rect 34802 28366 34804 28418
rect 34748 28364 34804 28366
rect 34636 27468 34692 27524
rect 34748 27804 34804 27860
rect 34524 27356 34580 27412
rect 34748 27244 34804 27300
rect 34972 30098 35028 30100
rect 34972 30046 34974 30098
rect 34974 30046 35026 30098
rect 35026 30046 35028 30098
rect 34972 30044 35028 30046
rect 35308 30210 35364 30212
rect 35308 30158 35310 30210
rect 35310 30158 35362 30210
rect 35362 30158 35364 30210
rect 35308 30156 35364 30158
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35420 28812 35476 28868
rect 34972 28530 35028 28532
rect 34972 28478 34974 28530
rect 34974 28478 35026 28530
rect 35026 28478 35028 28530
rect 34972 28476 35028 28478
rect 34972 28140 35028 28196
rect 35084 27804 35140 27860
rect 36876 34690 36932 34692
rect 36876 34638 36878 34690
rect 36878 34638 36930 34690
rect 36930 34638 36932 34690
rect 36876 34636 36932 34638
rect 36652 33628 36708 33684
rect 36428 33068 36484 33124
rect 36540 33180 36596 33236
rect 36428 31778 36484 31780
rect 36428 31726 36430 31778
rect 36430 31726 36482 31778
rect 36482 31726 36484 31778
rect 36428 31724 36484 31726
rect 36428 31276 36484 31332
rect 37660 38834 37716 38836
rect 37660 38782 37662 38834
rect 37662 38782 37714 38834
rect 37714 38782 37716 38834
rect 37660 38780 37716 38782
rect 37212 37266 37268 37268
rect 37212 37214 37214 37266
rect 37214 37214 37266 37266
rect 37266 37214 37268 37266
rect 37212 37212 37268 37214
rect 37436 37266 37492 37268
rect 37436 37214 37438 37266
rect 37438 37214 37490 37266
rect 37490 37214 37492 37266
rect 37436 37212 37492 37214
rect 37772 37100 37828 37156
rect 37660 36988 37716 37044
rect 37548 35644 37604 35700
rect 37100 35420 37156 35476
rect 37660 35420 37716 35476
rect 37212 35084 37268 35140
rect 38220 37826 38276 37828
rect 38220 37774 38222 37826
rect 38222 37774 38274 37826
rect 38274 37774 38276 37826
rect 38220 37772 38276 37774
rect 39004 43820 39060 43876
rect 39452 52668 39508 52724
rect 40124 54572 40180 54628
rect 40012 53788 40068 53844
rect 40460 55074 40516 55076
rect 40460 55022 40462 55074
rect 40462 55022 40514 55074
rect 40514 55022 40516 55074
rect 40460 55020 40516 55022
rect 40236 53900 40292 53956
rect 39788 52668 39844 52724
rect 39900 53452 39956 53508
rect 39452 52108 39508 52164
rect 39564 52050 39620 52052
rect 39564 51998 39566 52050
rect 39566 51998 39618 52050
rect 39618 51998 39620 52050
rect 39564 51996 39620 51998
rect 39452 49196 39508 49252
rect 39564 49756 39620 49812
rect 39452 48524 39508 48580
rect 39452 47404 39508 47460
rect 39564 47068 39620 47124
rect 39564 45836 39620 45892
rect 40124 52946 40180 52948
rect 40124 52894 40126 52946
rect 40126 52894 40178 52946
rect 40178 52894 40180 52946
rect 40124 52892 40180 52894
rect 40012 52220 40068 52276
rect 39900 51548 39956 51604
rect 39788 51212 39844 51268
rect 40348 50594 40404 50596
rect 40348 50542 40350 50594
rect 40350 50542 40402 50594
rect 40402 50542 40404 50594
rect 40348 50540 40404 50542
rect 41020 56306 41076 56308
rect 41020 56254 41022 56306
rect 41022 56254 41074 56306
rect 41074 56254 41076 56306
rect 41020 56252 41076 56254
rect 43036 56306 43092 56308
rect 43036 56254 43038 56306
rect 43038 56254 43090 56306
rect 43090 56254 43092 56306
rect 43036 56252 43092 56254
rect 50556 56474 50612 56476
rect 50556 56422 50558 56474
rect 50558 56422 50610 56474
rect 50610 56422 50612 56474
rect 50556 56420 50612 56422
rect 50660 56474 50716 56476
rect 50660 56422 50662 56474
rect 50662 56422 50714 56474
rect 50714 56422 50716 56474
rect 50660 56420 50716 56422
rect 50764 56474 50820 56476
rect 50764 56422 50766 56474
rect 50766 56422 50818 56474
rect 50818 56422 50820 56474
rect 50764 56420 50820 56422
rect 41020 55298 41076 55300
rect 41020 55246 41022 55298
rect 41022 55246 41074 55298
rect 41074 55246 41076 55298
rect 41020 55244 41076 55246
rect 41020 54626 41076 54628
rect 41020 54574 41022 54626
rect 41022 54574 41074 54626
rect 41074 54574 41076 54626
rect 41020 54572 41076 54574
rect 41580 56140 41636 56196
rect 43708 56194 43764 56196
rect 43708 56142 43710 56194
rect 43710 56142 43762 56194
rect 43762 56142 43764 56194
rect 43708 56140 43764 56142
rect 42588 56082 42644 56084
rect 42588 56030 42590 56082
rect 42590 56030 42642 56082
rect 42642 56030 42644 56082
rect 42588 56028 42644 56030
rect 42140 55970 42196 55972
rect 42140 55918 42142 55970
rect 42142 55918 42194 55970
rect 42194 55918 42196 55970
rect 42140 55916 42196 55918
rect 42028 55410 42084 55412
rect 42028 55358 42030 55410
rect 42030 55358 42082 55410
rect 42082 55358 42084 55410
rect 42028 55356 42084 55358
rect 42476 55298 42532 55300
rect 42476 55246 42478 55298
rect 42478 55246 42530 55298
rect 42530 55246 42532 55298
rect 42476 55244 42532 55246
rect 41580 55186 41636 55188
rect 41580 55134 41582 55186
rect 41582 55134 41634 55186
rect 41634 55134 41636 55186
rect 41580 55132 41636 55134
rect 41356 54012 41412 54068
rect 42588 53618 42644 53620
rect 42588 53566 42590 53618
rect 42590 53566 42642 53618
rect 42642 53566 42644 53618
rect 42588 53564 42644 53566
rect 42700 53506 42756 53508
rect 42700 53454 42702 53506
rect 42702 53454 42754 53506
rect 42754 53454 42756 53506
rect 42700 53452 42756 53454
rect 42364 53340 42420 53396
rect 41020 53170 41076 53172
rect 41020 53118 41022 53170
rect 41022 53118 41074 53170
rect 41074 53118 41076 53170
rect 41020 53116 41076 53118
rect 41132 53058 41188 53060
rect 41132 53006 41134 53058
rect 41134 53006 41186 53058
rect 41186 53006 41188 53058
rect 41132 53004 41188 53006
rect 40908 52946 40964 52948
rect 40908 52894 40910 52946
rect 40910 52894 40962 52946
rect 40962 52894 40964 52946
rect 40908 52892 40964 52894
rect 41132 52332 41188 52388
rect 40124 48636 40180 48692
rect 40124 46956 40180 47012
rect 40012 46786 40068 46788
rect 40012 46734 40014 46786
rect 40014 46734 40066 46786
rect 40066 46734 40068 46786
rect 40012 46732 40068 46734
rect 40236 46844 40292 46900
rect 40348 46508 40404 46564
rect 40684 48636 40740 48692
rect 42812 52892 42868 52948
rect 41356 52780 41412 52836
rect 42028 52834 42084 52836
rect 42028 52782 42030 52834
rect 42030 52782 42082 52834
rect 42082 52782 42084 52834
rect 42028 52780 42084 52782
rect 42924 52780 42980 52836
rect 42700 52332 42756 52388
rect 41356 52220 41412 52276
rect 41132 52162 41188 52164
rect 41132 52110 41134 52162
rect 41134 52110 41186 52162
rect 41186 52110 41188 52162
rect 41132 52108 41188 52110
rect 41132 51266 41188 51268
rect 41132 51214 41134 51266
rect 41134 51214 41186 51266
rect 41186 51214 41188 51266
rect 41132 51212 41188 51214
rect 41244 51100 41300 51156
rect 41468 48972 41524 49028
rect 41132 46956 41188 47012
rect 40572 46060 40628 46116
rect 41244 46620 41300 46676
rect 39788 45948 39844 46004
rect 40908 45890 40964 45892
rect 40908 45838 40910 45890
rect 40910 45838 40962 45890
rect 40962 45838 40964 45890
rect 40908 45836 40964 45838
rect 40572 45724 40628 45780
rect 39452 43932 39508 43988
rect 39340 43596 39396 43652
rect 39004 43148 39060 43204
rect 38892 42812 38948 42868
rect 40796 45778 40852 45780
rect 40796 45726 40798 45778
rect 40798 45726 40850 45778
rect 40850 45726 40852 45778
rect 40796 45724 40852 45726
rect 40460 44434 40516 44436
rect 40460 44382 40462 44434
rect 40462 44382 40514 44434
rect 40514 44382 40516 44434
rect 40460 44380 40516 44382
rect 41804 51378 41860 51380
rect 41804 51326 41806 51378
rect 41806 51326 41858 51378
rect 41858 51326 41860 51378
rect 41804 51324 41860 51326
rect 42588 52162 42644 52164
rect 42588 52110 42590 52162
rect 42590 52110 42642 52162
rect 42642 52110 42644 52162
rect 42588 52108 42644 52110
rect 43372 53340 43428 53396
rect 44380 53452 44436 53508
rect 43372 52946 43428 52948
rect 43372 52894 43374 52946
rect 43374 52894 43426 52946
rect 43426 52894 43428 52946
rect 43372 52892 43428 52894
rect 43596 52834 43652 52836
rect 43596 52782 43598 52834
rect 43598 52782 43650 52834
rect 43650 52782 43652 52834
rect 43596 52780 43652 52782
rect 43260 51772 43316 51828
rect 43596 52332 43652 52388
rect 42588 51548 42644 51604
rect 42476 51436 42532 51492
rect 41916 51212 41972 51268
rect 42924 51602 42980 51604
rect 42924 51550 42926 51602
rect 42926 51550 42978 51602
rect 42978 51550 42980 51602
rect 42924 51548 42980 51550
rect 43036 51378 43092 51380
rect 43036 51326 43038 51378
rect 43038 51326 43090 51378
rect 43090 51326 43092 51378
rect 43036 51324 43092 51326
rect 42476 50764 42532 50820
rect 41692 48636 41748 48692
rect 42028 48242 42084 48244
rect 42028 48190 42030 48242
rect 42030 48190 42082 48242
rect 42082 48190 42084 48242
rect 42028 48188 42084 48190
rect 41468 47068 41524 47124
rect 42140 46844 42196 46900
rect 41468 46732 41524 46788
rect 41804 46674 41860 46676
rect 41804 46622 41806 46674
rect 41806 46622 41858 46674
rect 41858 46622 41860 46674
rect 41804 46620 41860 46622
rect 41356 45948 41412 46004
rect 42028 46508 42084 46564
rect 41468 45388 41524 45444
rect 42252 44716 42308 44772
rect 40572 43596 40628 43652
rect 39788 43314 39844 43316
rect 39788 43262 39790 43314
rect 39790 43262 39842 43314
rect 39842 43262 39844 43314
rect 39788 43260 39844 43262
rect 40012 43148 40068 43204
rect 39788 42252 39844 42308
rect 39564 41970 39620 41972
rect 39564 41918 39566 41970
rect 39566 41918 39618 41970
rect 39618 41918 39620 41970
rect 39564 41916 39620 41918
rect 39228 41244 39284 41300
rect 39340 41074 39396 41076
rect 39340 41022 39342 41074
rect 39342 41022 39394 41074
rect 39394 41022 39396 41074
rect 39340 41020 39396 41022
rect 39452 39676 39508 39732
rect 40124 42194 40180 42196
rect 40124 42142 40126 42194
rect 40126 42142 40178 42194
rect 40178 42142 40180 42194
rect 40124 42140 40180 42142
rect 40124 41916 40180 41972
rect 40572 43260 40628 43316
rect 41692 43762 41748 43764
rect 41692 43710 41694 43762
rect 41694 43710 41746 43762
rect 41746 43710 41748 43762
rect 41692 43708 41748 43710
rect 42588 50034 42644 50036
rect 42588 49982 42590 50034
rect 42590 49982 42642 50034
rect 42642 49982 42644 50034
rect 42588 49980 42644 49982
rect 43484 51378 43540 51380
rect 43484 51326 43486 51378
rect 43486 51326 43538 51378
rect 43538 51326 43540 51378
rect 43484 51324 43540 51326
rect 43932 51996 43988 52052
rect 43820 51548 43876 51604
rect 43484 50764 43540 50820
rect 44156 51436 44212 51492
rect 43820 50092 43876 50148
rect 43932 49980 43988 50036
rect 43260 49810 43316 49812
rect 43260 49758 43262 49810
rect 43262 49758 43314 49810
rect 43314 49758 43316 49810
rect 43260 49756 43316 49758
rect 43708 48524 43764 48580
rect 43148 47458 43204 47460
rect 43148 47406 43150 47458
rect 43150 47406 43202 47458
rect 43202 47406 43204 47458
rect 43148 47404 43204 47406
rect 42924 46674 42980 46676
rect 42924 46622 42926 46674
rect 42926 46622 42978 46674
rect 42978 46622 42980 46674
rect 42924 46620 42980 46622
rect 43260 46450 43316 46452
rect 43260 46398 43262 46450
rect 43262 46398 43314 46450
rect 43314 46398 43316 46450
rect 43260 46396 43316 46398
rect 43820 47346 43876 47348
rect 43820 47294 43822 47346
rect 43822 47294 43874 47346
rect 43874 47294 43876 47346
rect 43820 47292 43876 47294
rect 47852 53618 47908 53620
rect 47852 53566 47854 53618
rect 47854 53566 47906 53618
rect 47906 53566 47908 53618
rect 47852 53564 47908 53566
rect 44492 53116 44548 53172
rect 46284 53116 46340 53172
rect 44940 51996 44996 52052
rect 44828 51436 44884 51492
rect 44492 50316 44548 50372
rect 45500 51548 45556 51604
rect 45612 51490 45668 51492
rect 45612 51438 45614 51490
rect 45614 51438 45666 51490
rect 45666 51438 45668 51490
rect 45612 51436 45668 51438
rect 45388 51212 45444 51268
rect 44492 49980 44548 50036
rect 46956 51996 47012 52052
rect 46956 51490 47012 51492
rect 46956 51438 46958 51490
rect 46958 51438 47010 51490
rect 47010 51438 47012 51490
rect 46956 51436 47012 51438
rect 46508 51378 46564 51380
rect 46508 51326 46510 51378
rect 46510 51326 46562 51378
rect 46562 51326 46564 51378
rect 46508 51324 46564 51326
rect 46620 51212 46676 51268
rect 47180 51100 47236 51156
rect 46060 50540 46116 50596
rect 46620 50540 46676 50596
rect 45612 50482 45668 50484
rect 45612 50430 45614 50482
rect 45614 50430 45666 50482
rect 45666 50430 45668 50482
rect 45612 50428 45668 50430
rect 45164 50316 45220 50372
rect 44940 50092 44996 50148
rect 44044 48860 44100 48916
rect 46956 50428 47012 50484
rect 47852 51378 47908 51380
rect 47852 51326 47854 51378
rect 47854 51326 47906 51378
rect 47906 51326 47908 51378
rect 47852 51324 47908 51326
rect 48188 53340 48244 53396
rect 48188 52220 48244 52276
rect 48412 52162 48468 52164
rect 48412 52110 48414 52162
rect 48414 52110 48466 52162
rect 48466 52110 48468 52162
rect 48412 52108 48468 52110
rect 49084 52332 49140 52388
rect 48636 52050 48692 52052
rect 48636 51998 48638 52050
rect 48638 51998 48690 52050
rect 48690 51998 48692 52050
rect 48636 51996 48692 51998
rect 49644 52332 49700 52388
rect 50556 54906 50612 54908
rect 50556 54854 50558 54906
rect 50558 54854 50610 54906
rect 50610 54854 50612 54906
rect 50556 54852 50612 54854
rect 50660 54906 50716 54908
rect 50660 54854 50662 54906
rect 50662 54854 50714 54906
rect 50714 54854 50716 54906
rect 50660 54852 50716 54854
rect 50764 54906 50820 54908
rect 50764 54854 50766 54906
rect 50766 54854 50818 54906
rect 50818 54854 50820 54906
rect 50764 54852 50820 54854
rect 50556 53338 50612 53340
rect 50556 53286 50558 53338
rect 50558 53286 50610 53338
rect 50610 53286 50612 53338
rect 50556 53284 50612 53286
rect 50660 53338 50716 53340
rect 50660 53286 50662 53338
rect 50662 53286 50714 53338
rect 50714 53286 50716 53338
rect 50660 53284 50716 53286
rect 50764 53338 50820 53340
rect 50764 53286 50766 53338
rect 50766 53286 50818 53338
rect 50818 53286 50820 53338
rect 50764 53284 50820 53286
rect 50316 52220 50372 52276
rect 49308 52162 49364 52164
rect 49308 52110 49310 52162
rect 49310 52110 49362 52162
rect 49362 52110 49364 52162
rect 49308 52108 49364 52110
rect 50876 52332 50932 52388
rect 50988 52108 51044 52164
rect 49196 51996 49252 52052
rect 48748 51378 48804 51380
rect 48748 51326 48750 51378
rect 48750 51326 48802 51378
rect 48802 51326 48804 51378
rect 48748 51324 48804 51326
rect 48076 50988 48132 51044
rect 47404 50316 47460 50372
rect 46844 48914 46900 48916
rect 46844 48862 46846 48914
rect 46846 48862 46898 48914
rect 46898 48862 46900 48914
rect 46844 48860 46900 48862
rect 44940 48748 44996 48804
rect 45276 48636 45332 48692
rect 44044 48076 44100 48132
rect 43932 46844 43988 46900
rect 44268 48130 44324 48132
rect 44268 48078 44270 48130
rect 44270 48078 44322 48130
rect 44322 48078 44324 48130
rect 44268 48076 44324 48078
rect 46172 48636 46228 48692
rect 45052 46396 45108 46452
rect 43596 45612 43652 45668
rect 43036 45052 43092 45108
rect 42252 43596 42308 43652
rect 41020 43148 41076 43204
rect 41468 42140 41524 42196
rect 40348 40236 40404 40292
rect 39116 39228 39172 39284
rect 38780 38108 38836 38164
rect 40908 40626 40964 40628
rect 40908 40574 40910 40626
rect 40910 40574 40962 40626
rect 40962 40574 40964 40626
rect 40908 40572 40964 40574
rect 40572 39730 40628 39732
rect 40572 39678 40574 39730
rect 40574 39678 40626 39730
rect 40626 39678 40628 39730
rect 40572 39676 40628 39678
rect 40684 40460 40740 40516
rect 40348 38780 40404 38836
rect 40236 38050 40292 38052
rect 40236 37998 40238 38050
rect 40238 37998 40290 38050
rect 40290 37998 40292 38050
rect 40236 37996 40292 37998
rect 39788 37772 39844 37828
rect 38220 37212 38276 37268
rect 38332 37100 38388 37156
rect 38220 36988 38276 37044
rect 38220 36482 38276 36484
rect 38220 36430 38222 36482
rect 38222 36430 38274 36482
rect 38274 36430 38276 36482
rect 38220 36428 38276 36430
rect 38108 36258 38164 36260
rect 38108 36206 38110 36258
rect 38110 36206 38162 36258
rect 38162 36206 38164 36258
rect 38108 36204 38164 36206
rect 38668 36258 38724 36260
rect 38668 36206 38670 36258
rect 38670 36206 38722 36258
rect 38722 36206 38724 36258
rect 38668 36204 38724 36206
rect 38892 37154 38948 37156
rect 38892 37102 38894 37154
rect 38894 37102 38946 37154
rect 38946 37102 38948 37154
rect 38892 37100 38948 37102
rect 40460 37436 40516 37492
rect 39452 36428 39508 36484
rect 37996 35868 38052 35924
rect 38332 35868 38388 35924
rect 37884 35756 37940 35812
rect 38220 35810 38276 35812
rect 38220 35758 38222 35810
rect 38222 35758 38274 35810
rect 38274 35758 38276 35810
rect 38220 35756 38276 35758
rect 38780 35756 38836 35812
rect 38556 35698 38612 35700
rect 38556 35646 38558 35698
rect 38558 35646 38610 35698
rect 38610 35646 38612 35698
rect 38556 35644 38612 35646
rect 38220 35586 38276 35588
rect 38220 35534 38222 35586
rect 38222 35534 38274 35586
rect 38274 35534 38276 35586
rect 38220 35532 38276 35534
rect 38108 35084 38164 35140
rect 37772 34972 37828 35028
rect 38444 34972 38500 35028
rect 37660 34188 37716 34244
rect 38220 34188 38276 34244
rect 37212 33628 37268 33684
rect 37996 33628 38052 33684
rect 37100 33516 37156 33572
rect 37100 31778 37156 31780
rect 37100 31726 37102 31778
rect 37102 31726 37154 31778
rect 37154 31726 37156 31778
rect 37100 31724 37156 31726
rect 36988 30940 37044 30996
rect 36540 30492 36596 30548
rect 36316 30210 36372 30212
rect 36316 30158 36318 30210
rect 36318 30158 36370 30210
rect 36370 30158 36372 30210
rect 36316 30156 36372 30158
rect 36652 30044 36708 30100
rect 35756 29484 35812 29540
rect 36204 29426 36260 29428
rect 36204 29374 36206 29426
rect 36206 29374 36258 29426
rect 36258 29374 36260 29426
rect 36204 29372 36260 29374
rect 35980 29260 36036 29316
rect 35196 28700 35252 28756
rect 35980 28812 36036 28868
rect 35308 28028 35364 28084
rect 35420 28252 35476 28308
rect 35196 27692 35252 27748
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 34524 26236 34580 26292
rect 34524 25900 34580 25956
rect 35196 27132 35252 27188
rect 35196 26012 35252 26068
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 34300 24892 34356 24948
rect 34524 25564 34580 25620
rect 34188 24556 34244 24612
rect 34412 24220 34468 24276
rect 34860 25004 34916 25060
rect 34636 24892 34692 24948
rect 34748 24444 34804 24500
rect 35196 25394 35252 25396
rect 35196 25342 35198 25394
rect 35198 25342 35250 25394
rect 35250 25342 35252 25394
rect 35196 25340 35252 25342
rect 35084 25116 35140 25172
rect 35868 28418 35924 28420
rect 35868 28366 35870 28418
rect 35870 28366 35922 28418
rect 35922 28366 35924 28418
rect 35868 28364 35924 28366
rect 36092 28252 36148 28308
rect 35980 28140 36036 28196
rect 35868 28028 35924 28084
rect 35756 26460 35812 26516
rect 36652 29372 36708 29428
rect 36428 29148 36484 29204
rect 37324 32844 37380 32900
rect 38332 33234 38388 33236
rect 38332 33182 38334 33234
rect 38334 33182 38386 33234
rect 38386 33182 38388 33234
rect 38332 33180 38388 33182
rect 37772 31164 37828 31220
rect 37324 30994 37380 30996
rect 37324 30942 37326 30994
rect 37326 30942 37378 30994
rect 37378 30942 37380 30994
rect 37324 30940 37380 30942
rect 37660 30770 37716 30772
rect 37660 30718 37662 30770
rect 37662 30718 37714 30770
rect 37714 30718 37716 30770
rect 37660 30716 37716 30718
rect 37212 30380 37268 30436
rect 37436 30268 37492 30324
rect 36988 29260 37044 29316
rect 37324 29538 37380 29540
rect 37324 29486 37326 29538
rect 37326 29486 37378 29538
rect 37378 29486 37380 29538
rect 37324 29484 37380 29486
rect 38556 34188 38612 34244
rect 38556 33346 38612 33348
rect 38556 33294 38558 33346
rect 38558 33294 38610 33346
rect 38610 33294 38612 33346
rect 38556 33292 38612 33294
rect 39676 35922 39732 35924
rect 39676 35870 39678 35922
rect 39678 35870 39730 35922
rect 39730 35870 39732 35922
rect 39676 35868 39732 35870
rect 40012 37042 40068 37044
rect 40012 36990 40014 37042
rect 40014 36990 40066 37042
rect 40066 36990 40068 37042
rect 40012 36988 40068 36990
rect 40012 36540 40068 36596
rect 40572 36988 40628 37044
rect 40236 36482 40292 36484
rect 40236 36430 40238 36482
rect 40238 36430 40290 36482
rect 40290 36430 40292 36482
rect 40236 36428 40292 36430
rect 40012 35922 40068 35924
rect 40012 35870 40014 35922
rect 40014 35870 40066 35922
rect 40066 35870 40068 35922
rect 40012 35868 40068 35870
rect 42588 43260 42644 43316
rect 42364 42252 42420 42308
rect 43036 43708 43092 43764
rect 43372 45388 43428 45444
rect 44940 45836 44996 45892
rect 44828 45778 44884 45780
rect 44828 45726 44830 45778
rect 44830 45726 44882 45778
rect 44882 45726 44884 45778
rect 44828 45724 44884 45726
rect 46844 48636 46900 48692
rect 47292 48636 47348 48692
rect 48748 50428 48804 50484
rect 49084 51212 49140 51268
rect 49084 50988 49140 51044
rect 48636 48972 48692 49028
rect 50556 51770 50612 51772
rect 50556 51718 50558 51770
rect 50558 51718 50610 51770
rect 50610 51718 50612 51770
rect 50556 51716 50612 51718
rect 50660 51770 50716 51772
rect 50660 51718 50662 51770
rect 50662 51718 50714 51770
rect 50714 51718 50716 51770
rect 50660 51716 50716 51718
rect 50764 51770 50820 51772
rect 50764 51718 50766 51770
rect 50766 51718 50818 51770
rect 50818 51718 50820 51770
rect 50764 51716 50820 51718
rect 49532 51266 49588 51268
rect 49532 51214 49534 51266
rect 49534 51214 49586 51266
rect 49586 51214 49588 51266
rect 49532 51212 49588 51214
rect 49756 51154 49812 51156
rect 49756 51102 49758 51154
rect 49758 51102 49810 51154
rect 49810 51102 49812 51154
rect 49756 51100 49812 51102
rect 49532 50594 49588 50596
rect 49532 50542 49534 50594
rect 49534 50542 49586 50594
rect 49586 50542 49588 50594
rect 49532 50540 49588 50542
rect 50092 51100 50148 51156
rect 50092 50706 50148 50708
rect 50092 50654 50094 50706
rect 50094 50654 50146 50706
rect 50146 50654 50148 50706
rect 50092 50652 50148 50654
rect 49980 50316 50036 50372
rect 51548 51996 51604 52052
rect 51884 51490 51940 51492
rect 51884 51438 51886 51490
rect 51886 51438 51938 51490
rect 51938 51438 51940 51490
rect 51884 51436 51940 51438
rect 52668 51436 52724 51492
rect 51100 51266 51156 51268
rect 51100 51214 51102 51266
rect 51102 51214 51154 51266
rect 51154 51214 51156 51266
rect 51100 51212 51156 51214
rect 51884 50652 51940 50708
rect 50556 50202 50612 50204
rect 50556 50150 50558 50202
rect 50558 50150 50610 50202
rect 50610 50150 50612 50202
rect 50556 50148 50612 50150
rect 50660 50202 50716 50204
rect 50660 50150 50662 50202
rect 50662 50150 50714 50202
rect 50714 50150 50716 50202
rect 50660 50148 50716 50150
rect 50764 50202 50820 50204
rect 50764 50150 50766 50202
rect 50766 50150 50818 50202
rect 50818 50150 50820 50202
rect 50764 50148 50820 50150
rect 50428 49980 50484 50036
rect 49532 49420 49588 49476
rect 50316 49420 50372 49476
rect 49532 49250 49588 49252
rect 49532 49198 49534 49250
rect 49534 49198 49586 49250
rect 49586 49198 49588 49250
rect 49532 49196 49588 49198
rect 50428 49196 50484 49252
rect 50428 48972 50484 49028
rect 47852 48524 47908 48580
rect 50556 48634 50612 48636
rect 50556 48582 50558 48634
rect 50558 48582 50610 48634
rect 50610 48582 50612 48634
rect 50556 48580 50612 48582
rect 50660 48634 50716 48636
rect 50660 48582 50662 48634
rect 50662 48582 50714 48634
rect 50714 48582 50716 48634
rect 50660 48580 50716 48582
rect 50764 48634 50820 48636
rect 50764 48582 50766 48634
rect 50766 48582 50818 48634
rect 50818 48582 50820 48634
rect 50764 48580 50820 48582
rect 51436 50370 51492 50372
rect 51436 50318 51438 50370
rect 51438 50318 51490 50370
rect 51490 50318 51492 50370
rect 51436 50316 51492 50318
rect 52444 50316 52500 50372
rect 52108 49980 52164 50036
rect 51100 48972 51156 49028
rect 50764 48412 50820 48468
rect 43932 44940 43988 44996
rect 43932 44380 43988 44436
rect 43932 44156 43988 44212
rect 43708 43596 43764 43652
rect 42700 41916 42756 41972
rect 43708 42812 43764 42868
rect 43596 42700 43652 42756
rect 43484 41916 43540 41972
rect 44156 43260 44212 43316
rect 45388 45388 45444 45444
rect 45052 45276 45108 45332
rect 44940 45106 44996 45108
rect 44940 45054 44942 45106
rect 44942 45054 44994 45106
rect 44994 45054 44996 45106
rect 44940 45052 44996 45054
rect 45276 44716 45332 44772
rect 44492 44156 44548 44212
rect 45500 45052 45556 45108
rect 45052 44156 45108 44212
rect 46060 46898 46116 46900
rect 46060 46846 46062 46898
rect 46062 46846 46114 46898
rect 46114 46846 46116 46898
rect 46060 46844 46116 46846
rect 50988 48354 51044 48356
rect 50988 48302 50990 48354
rect 50990 48302 51042 48354
rect 51042 48302 51044 48354
rect 50988 48300 51044 48302
rect 49308 47516 49364 47572
rect 52332 49420 52388 49476
rect 52444 48748 52500 48804
rect 51436 48412 51492 48468
rect 51212 47570 51268 47572
rect 51212 47518 51214 47570
rect 51214 47518 51266 47570
rect 51266 47518 51268 47570
rect 51212 47516 51268 47518
rect 51324 48300 51380 48356
rect 47964 46956 48020 47012
rect 48188 46786 48244 46788
rect 48188 46734 48190 46786
rect 48190 46734 48242 46786
rect 48242 46734 48244 46786
rect 48188 46732 48244 46734
rect 47852 46508 47908 46564
rect 46396 45948 46452 46004
rect 47628 45948 47684 46004
rect 46172 45778 46228 45780
rect 46172 45726 46174 45778
rect 46174 45726 46226 45778
rect 46226 45726 46228 45778
rect 46172 45724 46228 45726
rect 47516 45778 47572 45780
rect 47516 45726 47518 45778
rect 47518 45726 47570 45778
rect 47570 45726 47572 45778
rect 47516 45724 47572 45726
rect 45836 45666 45892 45668
rect 45836 45614 45838 45666
rect 45838 45614 45890 45666
rect 45890 45614 45892 45666
rect 45836 45612 45892 45614
rect 45836 45330 45892 45332
rect 45836 45278 45838 45330
rect 45838 45278 45890 45330
rect 45890 45278 45892 45330
rect 45836 45276 45892 45278
rect 46732 45276 46788 45332
rect 46284 44994 46340 44996
rect 46284 44942 46286 44994
rect 46286 44942 46338 44994
rect 46338 44942 46340 44994
rect 46284 44940 46340 44942
rect 46844 44940 46900 44996
rect 45612 44156 45668 44212
rect 46060 44380 46116 44436
rect 44940 42140 44996 42196
rect 44268 42028 44324 42084
rect 46732 43650 46788 43652
rect 46732 43598 46734 43650
rect 46734 43598 46786 43650
rect 46786 43598 46788 43650
rect 46732 43596 46788 43598
rect 46396 43260 46452 43316
rect 45388 42754 45444 42756
rect 45388 42702 45390 42754
rect 45390 42702 45442 42754
rect 45442 42702 45444 42754
rect 45388 42700 45444 42702
rect 45500 42028 45556 42084
rect 45388 41970 45444 41972
rect 45388 41918 45390 41970
rect 45390 41918 45442 41970
rect 45442 41918 45444 41970
rect 45388 41916 45444 41918
rect 42588 41186 42644 41188
rect 42588 41134 42590 41186
rect 42590 41134 42642 41186
rect 42642 41134 42644 41186
rect 42588 41132 42644 41134
rect 43260 40684 43316 40740
rect 42028 40460 42084 40516
rect 42476 40514 42532 40516
rect 42476 40462 42478 40514
rect 42478 40462 42530 40514
rect 42530 40462 42532 40514
rect 42476 40460 42532 40462
rect 41468 40402 41524 40404
rect 41468 40350 41470 40402
rect 41470 40350 41522 40402
rect 41522 40350 41524 40402
rect 41468 40348 41524 40350
rect 43036 40348 43092 40404
rect 41804 39564 41860 39620
rect 41244 38834 41300 38836
rect 41244 38782 41246 38834
rect 41246 38782 41298 38834
rect 41298 38782 41300 38834
rect 41244 38780 41300 38782
rect 40908 37996 40964 38052
rect 41692 36988 41748 37044
rect 41356 36482 41412 36484
rect 41356 36430 41358 36482
rect 41358 36430 41410 36482
rect 41410 36430 41412 36482
rect 41356 36428 41412 36430
rect 40684 35868 40740 35924
rect 39900 35644 39956 35700
rect 39116 35084 39172 35140
rect 39676 35196 39732 35252
rect 39452 35026 39508 35028
rect 39452 34974 39454 35026
rect 39454 34974 39506 35026
rect 39506 34974 39508 35026
rect 39452 34972 39508 34974
rect 40012 34972 40068 35028
rect 39676 34524 39732 34580
rect 40236 34188 40292 34244
rect 39228 34018 39284 34020
rect 39228 33966 39230 34018
rect 39230 33966 39282 34018
rect 39282 33966 39284 34018
rect 39228 33964 39284 33966
rect 40124 34018 40180 34020
rect 40124 33966 40126 34018
rect 40126 33966 40178 34018
rect 40178 33966 40180 34018
rect 40124 33964 40180 33966
rect 40124 33516 40180 33572
rect 41132 35698 41188 35700
rect 41132 35646 41134 35698
rect 41134 35646 41186 35698
rect 41186 35646 41188 35698
rect 41132 35644 41188 35646
rect 41804 35698 41860 35700
rect 41804 35646 41806 35698
rect 41806 35646 41858 35698
rect 41858 35646 41860 35698
rect 41804 35644 41860 35646
rect 41132 34972 41188 35028
rect 41804 35026 41860 35028
rect 41804 34974 41806 35026
rect 41806 34974 41858 35026
rect 41858 34974 41860 35026
rect 41804 34972 41860 34974
rect 42812 37436 42868 37492
rect 42700 35644 42756 35700
rect 43372 40402 43428 40404
rect 43372 40350 43374 40402
rect 43374 40350 43426 40402
rect 43426 40350 43428 40402
rect 43372 40348 43428 40350
rect 43596 40402 43652 40404
rect 43596 40350 43598 40402
rect 43598 40350 43650 40402
rect 43650 40350 43652 40402
rect 43596 40348 43652 40350
rect 43484 39564 43540 39620
rect 43708 39004 43764 39060
rect 43484 38892 43540 38948
rect 44940 41186 44996 41188
rect 44940 41134 44942 41186
rect 44942 41134 44994 41186
rect 44994 41134 44996 41186
rect 44940 41132 44996 41134
rect 44828 40684 44884 40740
rect 44492 38946 44548 38948
rect 44492 38894 44494 38946
rect 44494 38894 44546 38946
rect 44546 38894 44548 38946
rect 44492 38892 44548 38894
rect 43596 38834 43652 38836
rect 43596 38782 43598 38834
rect 43598 38782 43650 38834
rect 43650 38782 43652 38834
rect 43596 38780 43652 38782
rect 46172 41858 46228 41860
rect 46172 41806 46174 41858
rect 46174 41806 46226 41858
rect 46226 41806 46228 41858
rect 46172 41804 46228 41806
rect 45948 40236 46004 40292
rect 45612 39228 45668 39284
rect 45836 39058 45892 39060
rect 45836 39006 45838 39058
rect 45838 39006 45890 39058
rect 45890 39006 45892 39058
rect 45836 39004 45892 39006
rect 44940 38108 44996 38164
rect 46284 38834 46340 38836
rect 46284 38782 46286 38834
rect 46286 38782 46338 38834
rect 46338 38782 46340 38834
rect 46284 38780 46340 38782
rect 46956 44210 47012 44212
rect 46956 44158 46958 44210
rect 46958 44158 47010 44210
rect 47010 44158 47012 44210
rect 46956 44156 47012 44158
rect 47404 42476 47460 42532
rect 46956 41804 47012 41860
rect 47404 41580 47460 41636
rect 48188 45948 48244 46004
rect 47964 45724 48020 45780
rect 48748 45890 48804 45892
rect 48748 45838 48750 45890
rect 48750 45838 48802 45890
rect 48802 45838 48804 45890
rect 48748 45836 48804 45838
rect 48188 44156 48244 44212
rect 49084 44994 49140 44996
rect 49084 44942 49086 44994
rect 49086 44942 49138 44994
rect 49138 44942 49140 44994
rect 49084 44940 49140 44942
rect 49196 44156 49252 44212
rect 50556 47066 50612 47068
rect 50556 47014 50558 47066
rect 50558 47014 50610 47066
rect 50610 47014 50612 47066
rect 50556 47012 50612 47014
rect 50660 47066 50716 47068
rect 50660 47014 50662 47066
rect 50662 47014 50714 47066
rect 50714 47014 50716 47066
rect 50660 47012 50716 47014
rect 50764 47066 50820 47068
rect 50764 47014 50766 47066
rect 50766 47014 50818 47066
rect 50818 47014 50820 47066
rect 50764 47012 50820 47014
rect 50428 46786 50484 46788
rect 50428 46734 50430 46786
rect 50430 46734 50482 46786
rect 50482 46734 50484 46786
rect 50428 46732 50484 46734
rect 49756 44940 49812 44996
rect 49196 43314 49252 43316
rect 49196 43262 49198 43314
rect 49198 43262 49250 43314
rect 49250 43262 49252 43314
rect 49196 43260 49252 43262
rect 48972 42700 49028 42756
rect 47964 41580 48020 41636
rect 48300 40572 48356 40628
rect 47180 40290 47236 40292
rect 47180 40238 47182 40290
rect 47182 40238 47234 40290
rect 47234 40238 47236 40290
rect 47180 40236 47236 40238
rect 48748 40236 48804 40292
rect 48188 39676 48244 39732
rect 46620 39618 46676 39620
rect 46620 39566 46622 39618
rect 46622 39566 46674 39618
rect 46674 39566 46676 39618
rect 46620 39564 46676 39566
rect 46844 39004 46900 39060
rect 47180 38050 47236 38052
rect 47180 37998 47182 38050
rect 47182 37998 47234 38050
rect 47234 37998 47236 38050
rect 47180 37996 47236 37998
rect 45612 37212 45668 37268
rect 46732 37266 46788 37268
rect 46732 37214 46734 37266
rect 46734 37214 46786 37266
rect 46786 37214 46788 37266
rect 46732 37212 46788 37214
rect 41580 34636 41636 34692
rect 41132 34242 41188 34244
rect 41132 34190 41134 34242
rect 41134 34190 41186 34242
rect 41186 34190 41188 34242
rect 41132 34188 41188 34190
rect 41020 34076 41076 34132
rect 41020 33570 41076 33572
rect 41020 33518 41022 33570
rect 41022 33518 41074 33570
rect 41074 33518 41076 33570
rect 41020 33516 41076 33518
rect 42588 34524 42644 34580
rect 42140 34242 42196 34244
rect 42140 34190 42142 34242
rect 42142 34190 42194 34242
rect 42194 34190 42196 34242
rect 42140 34188 42196 34190
rect 41804 34130 41860 34132
rect 41804 34078 41806 34130
rect 41806 34078 41858 34130
rect 41858 34078 41860 34130
rect 41804 34076 41860 34078
rect 43372 36540 43428 36596
rect 46172 37154 46228 37156
rect 46172 37102 46174 37154
rect 46174 37102 46226 37154
rect 46226 37102 46228 37154
rect 46172 37100 46228 37102
rect 45612 36988 45668 37044
rect 44044 36594 44100 36596
rect 44044 36542 44046 36594
rect 44046 36542 44098 36594
rect 44098 36542 44100 36594
rect 44044 36540 44100 36542
rect 45612 36540 45668 36596
rect 45948 36876 46004 36932
rect 46956 36876 47012 36932
rect 47964 38220 48020 38276
rect 48076 39340 48132 39396
rect 47964 38050 48020 38052
rect 47964 37998 47966 38050
rect 47966 37998 48018 38050
rect 48018 37998 48020 38050
rect 47964 37996 48020 37998
rect 47628 37884 47684 37940
rect 47516 37266 47572 37268
rect 47516 37214 47518 37266
rect 47518 37214 47570 37266
rect 47570 37214 47572 37266
rect 47516 37212 47572 37214
rect 48188 38162 48244 38164
rect 48188 38110 48190 38162
rect 48190 38110 48242 38162
rect 48242 38110 48244 38162
rect 48188 38108 48244 38110
rect 48972 41916 49028 41972
rect 49308 41692 49364 41748
rect 49084 40460 49140 40516
rect 48860 39788 48916 39844
rect 48972 39676 49028 39732
rect 48748 39394 48804 39396
rect 48748 39342 48750 39394
rect 48750 39342 48802 39394
rect 48802 39342 48804 39394
rect 48748 39340 48804 39342
rect 48860 39228 48916 39284
rect 49308 39618 49364 39620
rect 49308 39566 49310 39618
rect 49310 39566 49362 39618
rect 49362 39566 49364 39618
rect 49308 39564 49364 39566
rect 49756 43260 49812 43316
rect 49532 41858 49588 41860
rect 49532 41806 49534 41858
rect 49534 41806 49586 41858
rect 49586 41806 49588 41858
rect 49532 41804 49588 41806
rect 50316 46508 50372 46564
rect 50092 44882 50148 44884
rect 50092 44830 50094 44882
rect 50094 44830 50146 44882
rect 50146 44830 50148 44882
rect 50092 44828 50148 44830
rect 49980 42700 50036 42756
rect 52780 50316 52836 50372
rect 52780 49980 52836 50036
rect 53228 50316 53284 50372
rect 53676 49980 53732 50036
rect 51436 46898 51492 46900
rect 51436 46846 51438 46898
rect 51438 46846 51490 46898
rect 51490 46846 51492 46898
rect 51436 46844 51492 46846
rect 50988 45778 51044 45780
rect 50988 45726 50990 45778
rect 50990 45726 51042 45778
rect 51042 45726 51044 45778
rect 50988 45724 51044 45726
rect 50556 45498 50612 45500
rect 50556 45446 50558 45498
rect 50558 45446 50610 45498
rect 50610 45446 50612 45498
rect 50556 45444 50612 45446
rect 50660 45498 50716 45500
rect 50660 45446 50662 45498
rect 50662 45446 50714 45498
rect 50714 45446 50716 45498
rect 50660 45444 50716 45446
rect 50764 45498 50820 45500
rect 50764 45446 50766 45498
rect 50766 45446 50818 45498
rect 50818 45446 50820 45498
rect 50764 45444 50820 45446
rect 50652 44828 50708 44884
rect 50764 44210 50820 44212
rect 50764 44158 50766 44210
rect 50766 44158 50818 44210
rect 50818 44158 50820 44210
rect 50764 44156 50820 44158
rect 50556 43930 50612 43932
rect 50556 43878 50558 43930
rect 50558 43878 50610 43930
rect 50610 43878 50612 43930
rect 50556 43876 50612 43878
rect 50660 43930 50716 43932
rect 50660 43878 50662 43930
rect 50662 43878 50714 43930
rect 50714 43878 50716 43930
rect 50660 43876 50716 43878
rect 50764 43930 50820 43932
rect 50764 43878 50766 43930
rect 50766 43878 50818 43930
rect 50818 43878 50820 43930
rect 50764 43876 50820 43878
rect 51548 46508 51604 46564
rect 51436 46450 51492 46452
rect 51436 46398 51438 46450
rect 51438 46398 51490 46450
rect 51490 46398 51492 46450
rect 51436 46396 51492 46398
rect 53116 49250 53172 49252
rect 53116 49198 53118 49250
rect 53118 49198 53170 49250
rect 53170 49198 53172 49250
rect 53116 49196 53172 49198
rect 52780 47516 52836 47572
rect 53116 48466 53172 48468
rect 53116 48414 53118 48466
rect 53118 48414 53170 48466
rect 53170 48414 53172 48466
rect 53116 48412 53172 48414
rect 53900 49196 53956 49252
rect 52780 46114 52836 46116
rect 52780 46062 52782 46114
rect 52782 46062 52834 46114
rect 52834 46062 52836 46114
rect 52780 46060 52836 46062
rect 51548 44828 51604 44884
rect 51660 44322 51716 44324
rect 51660 44270 51662 44322
rect 51662 44270 51714 44322
rect 51714 44270 51716 44322
rect 51660 44268 51716 44270
rect 52444 45164 52500 45220
rect 51884 44210 51940 44212
rect 51884 44158 51886 44210
rect 51886 44158 51938 44210
rect 51938 44158 51940 44210
rect 51884 44156 51940 44158
rect 51996 45052 52052 45108
rect 51100 43708 51156 43764
rect 52556 45052 52612 45108
rect 52444 44268 52500 44324
rect 49868 41916 49924 41972
rect 49756 41804 49812 41860
rect 49756 41580 49812 41636
rect 51548 43372 51604 43428
rect 50428 42530 50484 42532
rect 50428 42478 50430 42530
rect 50430 42478 50482 42530
rect 50482 42478 50484 42530
rect 50428 42476 50484 42478
rect 50556 42362 50612 42364
rect 50556 42310 50558 42362
rect 50558 42310 50610 42362
rect 50610 42310 50612 42362
rect 50556 42308 50612 42310
rect 50660 42362 50716 42364
rect 50660 42310 50662 42362
rect 50662 42310 50714 42362
rect 50714 42310 50716 42362
rect 50660 42308 50716 42310
rect 50764 42362 50820 42364
rect 50764 42310 50766 42362
rect 50766 42310 50818 42362
rect 50818 42310 50820 42362
rect 50764 42308 50820 42310
rect 51436 41804 51492 41860
rect 50316 41468 50372 41524
rect 51996 43708 52052 43764
rect 50428 41186 50484 41188
rect 50428 41134 50430 41186
rect 50430 41134 50482 41186
rect 50482 41134 50484 41186
rect 50428 41132 50484 41134
rect 50556 40794 50612 40796
rect 50556 40742 50558 40794
rect 50558 40742 50610 40794
rect 50610 40742 50612 40794
rect 50556 40740 50612 40742
rect 50660 40794 50716 40796
rect 50660 40742 50662 40794
rect 50662 40742 50714 40794
rect 50714 40742 50716 40794
rect 50660 40740 50716 40742
rect 50764 40794 50820 40796
rect 50764 40742 50766 40794
rect 50766 40742 50818 40794
rect 50818 40742 50820 40794
rect 50764 40740 50820 40742
rect 50652 40626 50708 40628
rect 50652 40574 50654 40626
rect 50654 40574 50706 40626
rect 50706 40574 50708 40626
rect 50652 40572 50708 40574
rect 52780 45778 52836 45780
rect 52780 45726 52782 45778
rect 52782 45726 52834 45778
rect 52834 45726 52836 45778
rect 52780 45724 52836 45726
rect 54124 47516 54180 47572
rect 53228 46844 53284 46900
rect 54124 46844 54180 46900
rect 52892 45164 52948 45220
rect 53004 45106 53060 45108
rect 53004 45054 53006 45106
rect 53006 45054 53058 45106
rect 53058 45054 53060 45106
rect 53004 45052 53060 45054
rect 53788 46396 53844 46452
rect 53788 45106 53844 45108
rect 53788 45054 53790 45106
rect 53790 45054 53842 45106
rect 53842 45054 53844 45106
rect 53788 45052 53844 45054
rect 54124 45052 54180 45108
rect 53228 43426 53284 43428
rect 53228 43374 53230 43426
rect 53230 43374 53282 43426
rect 53282 43374 53284 43426
rect 53228 43372 53284 43374
rect 54460 46396 54516 46452
rect 54348 46060 54404 46116
rect 54572 45106 54628 45108
rect 54572 45054 54574 45106
rect 54574 45054 54626 45106
rect 54626 45054 54628 45106
rect 54572 45052 54628 45054
rect 54124 43708 54180 43764
rect 55244 43762 55300 43764
rect 55244 43710 55246 43762
rect 55246 43710 55298 43762
rect 55298 43710 55300 43762
rect 55244 43708 55300 43710
rect 52444 41970 52500 41972
rect 52444 41918 52446 41970
rect 52446 41918 52498 41970
rect 52498 41918 52500 41970
rect 52444 41916 52500 41918
rect 51996 41804 52052 41860
rect 52780 42530 52836 42532
rect 52780 42478 52782 42530
rect 52782 42478 52834 42530
rect 52834 42478 52836 42530
rect 52780 42476 52836 42478
rect 52780 42028 52836 42084
rect 51772 41132 51828 41188
rect 49308 38834 49364 38836
rect 49308 38782 49310 38834
rect 49310 38782 49362 38834
rect 49362 38782 49364 38834
rect 49308 38780 49364 38782
rect 48300 37938 48356 37940
rect 48300 37886 48302 37938
rect 48302 37886 48354 37938
rect 48354 37886 48356 37938
rect 48300 37884 48356 37886
rect 43596 35196 43652 35252
rect 43036 34860 43092 34916
rect 42812 34188 42868 34244
rect 41804 33570 41860 33572
rect 41804 33518 41806 33570
rect 41806 33518 41858 33570
rect 41858 33518 41860 33570
rect 41804 33516 41860 33518
rect 43036 34242 43092 34244
rect 43036 34190 43038 34242
rect 43038 34190 43090 34242
rect 43090 34190 43092 34242
rect 43036 34188 43092 34190
rect 43484 34354 43540 34356
rect 43484 34302 43486 34354
rect 43486 34302 43538 34354
rect 43538 34302 43540 34354
rect 43484 34300 43540 34302
rect 43820 34914 43876 34916
rect 43820 34862 43822 34914
rect 43822 34862 43874 34914
rect 43874 34862 43876 34914
rect 43820 34860 43876 34862
rect 44268 35756 44324 35812
rect 44044 34860 44100 34916
rect 45276 35810 45332 35812
rect 45276 35758 45278 35810
rect 45278 35758 45330 35810
rect 45330 35758 45332 35810
rect 45276 35756 45332 35758
rect 45276 35196 45332 35252
rect 43932 34690 43988 34692
rect 43932 34638 43934 34690
rect 43934 34638 43986 34690
rect 43986 34638 43988 34690
rect 43932 34636 43988 34638
rect 41916 33346 41972 33348
rect 41916 33294 41918 33346
rect 41918 33294 41970 33346
rect 41970 33294 41972 33346
rect 41916 33292 41972 33294
rect 42700 33346 42756 33348
rect 42700 33294 42702 33346
rect 42702 33294 42754 33346
rect 42754 33294 42756 33346
rect 42700 33292 42756 33294
rect 43708 33964 43764 34020
rect 40460 33180 40516 33236
rect 38892 32732 38948 32788
rect 40684 32732 40740 32788
rect 38556 32620 38612 32676
rect 38332 31724 38388 31780
rect 38332 31164 38388 31220
rect 39564 31724 39620 31780
rect 38444 30994 38500 30996
rect 38444 30942 38446 30994
rect 38446 30942 38498 30994
rect 38498 30942 38500 30994
rect 38444 30940 38500 30942
rect 37996 30322 38052 30324
rect 37996 30270 37998 30322
rect 37998 30270 38050 30322
rect 38050 30270 38052 30322
rect 37996 30268 38052 30270
rect 37324 28530 37380 28532
rect 37324 28478 37326 28530
rect 37326 28478 37378 28530
rect 37378 28478 37380 28530
rect 37324 28476 37380 28478
rect 36652 27916 36708 27972
rect 37100 28364 37156 28420
rect 37660 28642 37716 28644
rect 37660 28590 37662 28642
rect 37662 28590 37714 28642
rect 37714 28590 37716 28642
rect 37660 28588 37716 28590
rect 38220 30492 38276 30548
rect 39228 31388 39284 31444
rect 39116 30994 39172 30996
rect 39116 30942 39118 30994
rect 39118 30942 39170 30994
rect 39170 30942 39172 30994
rect 39116 30940 39172 30942
rect 38556 30380 38612 30436
rect 40348 31778 40404 31780
rect 40348 31726 40350 31778
rect 40350 31726 40402 31778
rect 40402 31726 40404 31778
rect 40348 31724 40404 31726
rect 39900 31388 39956 31444
rect 39676 30882 39732 30884
rect 39676 30830 39678 30882
rect 39678 30830 39730 30882
rect 39730 30830 39732 30882
rect 39676 30828 39732 30830
rect 40572 30380 40628 30436
rect 40348 29820 40404 29876
rect 40012 29596 40068 29652
rect 39900 29314 39956 29316
rect 39900 29262 39902 29314
rect 39902 29262 39954 29314
rect 39954 29262 39956 29314
rect 39900 29260 39956 29262
rect 37884 28476 37940 28532
rect 36316 26908 36372 26964
rect 37884 28028 37940 28084
rect 38444 27970 38500 27972
rect 38444 27918 38446 27970
rect 38446 27918 38498 27970
rect 38498 27918 38500 27970
rect 38444 27916 38500 27918
rect 38892 28700 38948 28756
rect 38780 28476 38836 28532
rect 38780 28140 38836 28196
rect 38556 27580 38612 27636
rect 39900 28700 39956 28756
rect 39004 28476 39060 28532
rect 39340 28530 39396 28532
rect 39340 28478 39342 28530
rect 39342 28478 39394 28530
rect 39394 28478 39396 28530
rect 39340 28476 39396 28478
rect 39004 28252 39060 28308
rect 39116 28418 39172 28420
rect 39116 28366 39118 28418
rect 39118 28366 39170 28418
rect 39170 28366 39172 28418
rect 39116 28364 39172 28366
rect 39228 28252 39284 28308
rect 42700 32732 42756 32788
rect 42028 31948 42084 32004
rect 41020 30492 41076 30548
rect 41580 29932 41636 29988
rect 40796 29650 40852 29652
rect 40796 29598 40798 29650
rect 40798 29598 40850 29650
rect 40850 29598 40852 29650
rect 40796 29596 40852 29598
rect 40908 29260 40964 29316
rect 39900 27916 39956 27972
rect 40124 27916 40180 27972
rect 38892 27020 38948 27076
rect 39452 27858 39508 27860
rect 39452 27806 39454 27858
rect 39454 27806 39506 27858
rect 39506 27806 39508 27858
rect 39452 27804 39508 27806
rect 37100 26572 37156 26628
rect 36204 25452 36260 25508
rect 35420 24946 35476 24948
rect 35420 24894 35422 24946
rect 35422 24894 35474 24946
rect 35474 24894 35476 24946
rect 35420 24892 35476 24894
rect 37996 25506 38052 25508
rect 37996 25454 37998 25506
rect 37998 25454 38050 25506
rect 38050 25454 38052 25506
rect 37996 25452 38052 25454
rect 37436 25394 37492 25396
rect 37436 25342 37438 25394
rect 37438 25342 37490 25394
rect 37490 25342 37492 25394
rect 37436 25340 37492 25342
rect 37100 25228 37156 25284
rect 34748 23884 34804 23940
rect 34412 23826 34468 23828
rect 34412 23774 34414 23826
rect 34414 23774 34466 23826
rect 34466 23774 34468 23826
rect 34412 23772 34468 23774
rect 34300 23100 34356 23156
rect 34748 23212 34804 23268
rect 34076 22764 34132 22820
rect 34636 23154 34692 23156
rect 34636 23102 34638 23154
rect 34638 23102 34690 23154
rect 34690 23102 34692 23154
rect 34636 23100 34692 23102
rect 34524 23042 34580 23044
rect 34524 22990 34526 23042
rect 34526 22990 34578 23042
rect 34578 22990 34580 23042
rect 34524 22988 34580 22990
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 35756 24834 35812 24836
rect 35756 24782 35758 24834
rect 35758 24782 35810 24834
rect 35810 24782 35812 24834
rect 35756 24780 35812 24782
rect 36316 24780 36372 24836
rect 35644 24722 35700 24724
rect 35644 24670 35646 24722
rect 35646 24670 35698 24722
rect 35698 24670 35700 24722
rect 35644 24668 35700 24670
rect 37100 24780 37156 24836
rect 35532 23772 35588 23828
rect 35980 23714 36036 23716
rect 35980 23662 35982 23714
rect 35982 23662 36034 23714
rect 36034 23662 36036 23714
rect 35980 23660 36036 23662
rect 35308 23548 35364 23604
rect 36988 24444 37044 24500
rect 36316 23548 36372 23604
rect 36428 23996 36484 24052
rect 35196 22876 35252 22932
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 33852 22092 33908 22148
rect 36204 22540 36260 22596
rect 34412 22204 34468 22260
rect 34300 22146 34356 22148
rect 34300 22094 34302 22146
rect 34302 22094 34354 22146
rect 34354 22094 34356 22146
rect 34300 22092 34356 22094
rect 34524 21980 34580 22036
rect 33516 21644 33572 21700
rect 34412 21586 34468 21588
rect 34412 21534 34414 21586
rect 34414 21534 34466 21586
rect 34466 21534 34468 21586
rect 34412 21532 34468 21534
rect 34412 20076 34468 20132
rect 33628 19794 33684 19796
rect 33628 19742 33630 19794
rect 33630 19742 33682 19794
rect 33682 19742 33684 19794
rect 33628 19740 33684 19742
rect 33852 19404 33908 19460
rect 33068 17666 33124 17668
rect 33068 17614 33070 17666
rect 33070 17614 33122 17666
rect 33122 17614 33124 17666
rect 33068 17612 33124 17614
rect 34524 18172 34580 18228
rect 33516 17666 33572 17668
rect 33516 17614 33518 17666
rect 33518 17614 33570 17666
rect 33570 17614 33572 17666
rect 33516 17612 33572 17614
rect 35196 22370 35252 22372
rect 35196 22318 35198 22370
rect 35198 22318 35250 22370
rect 35250 22318 35252 22370
rect 35196 22316 35252 22318
rect 34972 22258 35028 22260
rect 34972 22206 34974 22258
rect 34974 22206 35026 22258
rect 35026 22206 35028 22258
rect 34972 22204 35028 22206
rect 38332 25676 38388 25732
rect 39900 27746 39956 27748
rect 39900 27694 39902 27746
rect 39902 27694 39954 27746
rect 39954 27694 39956 27746
rect 39900 27692 39956 27694
rect 41020 28642 41076 28644
rect 41020 28590 41022 28642
rect 41022 28590 41074 28642
rect 41074 28590 41076 28642
rect 41020 28588 41076 28590
rect 42476 31106 42532 31108
rect 42476 31054 42478 31106
rect 42478 31054 42530 31106
rect 42530 31054 42532 31106
rect 42476 31052 42532 31054
rect 42924 32674 42980 32676
rect 42924 32622 42926 32674
rect 42926 32622 42978 32674
rect 42978 32622 42980 32674
rect 42924 32620 42980 32622
rect 45724 35196 45780 35252
rect 45724 34914 45780 34916
rect 45724 34862 45726 34914
rect 45726 34862 45778 34914
rect 45778 34862 45780 34914
rect 45724 34860 45780 34862
rect 45388 34636 45444 34692
rect 45164 34300 45220 34356
rect 44156 34130 44212 34132
rect 44156 34078 44158 34130
rect 44158 34078 44210 34130
rect 44210 34078 44212 34130
rect 44156 34076 44212 34078
rect 44268 33964 44324 34020
rect 44716 34076 44772 34132
rect 43932 33516 43988 33572
rect 43820 32620 43876 32676
rect 43932 32844 43988 32900
rect 46284 34690 46340 34692
rect 46284 34638 46286 34690
rect 46286 34638 46338 34690
rect 46338 34638 46340 34690
rect 46284 34636 46340 34638
rect 47292 35756 47348 35812
rect 47180 35644 47236 35700
rect 47068 35196 47124 35252
rect 47180 34972 47236 35028
rect 48076 35308 48132 35364
rect 46508 34690 46564 34692
rect 46508 34638 46510 34690
rect 46510 34638 46562 34690
rect 46562 34638 46564 34690
rect 46508 34636 46564 34638
rect 47516 34636 47572 34692
rect 46620 34524 46676 34580
rect 45612 34354 45668 34356
rect 45612 34302 45614 34354
rect 45614 34302 45666 34354
rect 45666 34302 45668 34354
rect 45612 34300 45668 34302
rect 45948 34130 46004 34132
rect 45948 34078 45950 34130
rect 45950 34078 46002 34130
rect 46002 34078 46004 34130
rect 45948 34076 46004 34078
rect 44828 33234 44884 33236
rect 44828 33182 44830 33234
rect 44830 33182 44882 33234
rect 44882 33182 44884 33234
rect 44828 33180 44884 33182
rect 45276 32844 45332 32900
rect 45052 32508 45108 32564
rect 45836 32562 45892 32564
rect 45836 32510 45838 32562
rect 45838 32510 45890 32562
rect 45890 32510 45892 32562
rect 45836 32508 45892 32510
rect 46060 33234 46116 33236
rect 46060 33182 46062 33234
rect 46062 33182 46114 33234
rect 46114 33182 46116 33234
rect 46060 33180 46116 33182
rect 45500 31948 45556 32004
rect 46620 33068 46676 33124
rect 48524 34914 48580 34916
rect 48524 34862 48526 34914
rect 48526 34862 48578 34914
rect 48578 34862 48580 34914
rect 48524 34860 48580 34862
rect 48972 35308 49028 35364
rect 49084 34860 49140 34916
rect 48412 34524 48468 34580
rect 50092 37938 50148 37940
rect 50092 37886 50094 37938
rect 50094 37886 50146 37938
rect 50146 37886 50148 37938
rect 50092 37884 50148 37886
rect 51100 39564 51156 39620
rect 50556 39226 50612 39228
rect 50556 39174 50558 39226
rect 50558 39174 50610 39226
rect 50610 39174 50612 39226
rect 50556 39172 50612 39174
rect 50660 39226 50716 39228
rect 50660 39174 50662 39226
rect 50662 39174 50714 39226
rect 50714 39174 50716 39226
rect 50660 39172 50716 39174
rect 50764 39226 50820 39228
rect 50764 39174 50766 39226
rect 50766 39174 50818 39226
rect 50818 39174 50820 39226
rect 50764 39172 50820 39174
rect 51100 38780 51156 38836
rect 50876 38556 50932 38612
rect 50556 37658 50612 37660
rect 50556 37606 50558 37658
rect 50558 37606 50610 37658
rect 50610 37606 50612 37658
rect 50556 37604 50612 37606
rect 50660 37658 50716 37660
rect 50660 37606 50662 37658
rect 50662 37606 50714 37658
rect 50714 37606 50716 37658
rect 50660 37604 50716 37606
rect 50764 37658 50820 37660
rect 50764 37606 50766 37658
rect 50766 37606 50818 37658
rect 50818 37606 50820 37658
rect 50764 37604 50820 37606
rect 49868 37212 49924 37268
rect 49644 36876 49700 36932
rect 49644 35420 49700 35476
rect 49308 34636 49364 34692
rect 49308 34354 49364 34356
rect 49308 34302 49310 34354
rect 49310 34302 49362 34354
rect 49362 34302 49364 34354
rect 49308 34300 49364 34302
rect 49868 35810 49924 35812
rect 49868 35758 49870 35810
rect 49870 35758 49922 35810
rect 49922 35758 49924 35810
rect 49868 35756 49924 35758
rect 50764 37266 50820 37268
rect 50764 37214 50766 37266
rect 50766 37214 50818 37266
rect 50818 37214 50820 37266
rect 50764 37212 50820 37214
rect 49868 34972 49924 35028
rect 49980 34914 50036 34916
rect 49980 34862 49982 34914
rect 49982 34862 50034 34914
rect 50034 34862 50036 34914
rect 49980 34860 50036 34862
rect 49868 34690 49924 34692
rect 49868 34638 49870 34690
rect 49870 34638 49922 34690
rect 49922 34638 49924 34690
rect 49868 34636 49924 34638
rect 49756 34524 49812 34580
rect 49868 34076 49924 34132
rect 49532 33180 49588 33236
rect 46620 31948 46676 32004
rect 46732 32620 46788 32676
rect 45164 31612 45220 31668
rect 46060 31666 46116 31668
rect 46060 31614 46062 31666
rect 46062 31614 46114 31666
rect 46114 31614 46116 31666
rect 46060 31612 46116 31614
rect 47068 31666 47124 31668
rect 47068 31614 47070 31666
rect 47070 31614 47122 31666
rect 47122 31614 47124 31666
rect 47068 31612 47124 31614
rect 49308 33122 49364 33124
rect 49308 33070 49310 33122
rect 49310 33070 49362 33122
rect 49362 33070 49364 33122
rect 49308 33068 49364 33070
rect 49308 32844 49364 32900
rect 47964 31890 48020 31892
rect 47964 31838 47966 31890
rect 47966 31838 48018 31890
rect 48018 31838 48020 31890
rect 47964 31836 48020 31838
rect 48300 31836 48356 31892
rect 44940 31276 44996 31332
rect 42252 30156 42308 30212
rect 41916 29820 41972 29876
rect 42812 30716 42868 30772
rect 42924 30044 42980 30100
rect 43036 29986 43092 29988
rect 43036 29934 43038 29986
rect 43038 29934 43090 29986
rect 43090 29934 43092 29986
rect 43036 29932 43092 29934
rect 43596 31052 43652 31108
rect 44492 31106 44548 31108
rect 44492 31054 44494 31106
rect 44494 31054 44546 31106
rect 44546 31054 44548 31106
rect 44492 31052 44548 31054
rect 43932 30322 43988 30324
rect 43932 30270 43934 30322
rect 43934 30270 43986 30322
rect 43986 30270 43988 30322
rect 43932 30268 43988 30270
rect 43372 30156 43428 30212
rect 44268 30210 44324 30212
rect 44268 30158 44270 30210
rect 44270 30158 44322 30210
rect 44322 30158 44324 30210
rect 44268 30156 44324 30158
rect 44604 30044 44660 30100
rect 44044 29986 44100 29988
rect 44044 29934 44046 29986
rect 44046 29934 44098 29986
rect 44098 29934 44100 29986
rect 44044 29932 44100 29934
rect 43148 29820 43204 29876
rect 44716 29932 44772 29988
rect 45276 30770 45332 30772
rect 45276 30718 45278 30770
rect 45278 30718 45330 30770
rect 45330 30718 45332 30770
rect 45276 30716 45332 30718
rect 45612 30770 45668 30772
rect 45612 30718 45614 30770
rect 45614 30718 45666 30770
rect 45666 30718 45668 30770
rect 45612 30716 45668 30718
rect 45164 30156 45220 30212
rect 45052 29596 45108 29652
rect 44492 29372 44548 29428
rect 40348 27916 40404 27972
rect 41692 28418 41748 28420
rect 41692 28366 41694 28418
rect 41694 28366 41746 28418
rect 41746 28366 41748 28418
rect 41692 28364 41748 28366
rect 43148 28530 43204 28532
rect 43148 28478 43150 28530
rect 43150 28478 43202 28530
rect 43202 28478 43204 28530
rect 43148 28476 43204 28478
rect 43820 28476 43876 28532
rect 42364 28418 42420 28420
rect 42364 28366 42366 28418
rect 42366 28366 42418 28418
rect 42418 28366 42420 28418
rect 42364 28364 42420 28366
rect 42140 28252 42196 28308
rect 41020 27692 41076 27748
rect 41916 27580 41972 27636
rect 40348 26684 40404 26740
rect 41020 26684 41076 26740
rect 41804 26514 41860 26516
rect 41804 26462 41806 26514
rect 41806 26462 41858 26514
rect 41858 26462 41860 26514
rect 41804 26460 41860 26462
rect 46844 31500 46900 31556
rect 47628 31554 47684 31556
rect 47628 31502 47630 31554
rect 47630 31502 47682 31554
rect 47682 31502 47684 31554
rect 47628 31500 47684 31502
rect 46284 30828 46340 30884
rect 46396 30716 46452 30772
rect 48748 31164 48804 31220
rect 49084 31778 49140 31780
rect 49084 31726 49086 31778
rect 49086 31726 49138 31778
rect 49138 31726 49140 31778
rect 49084 31724 49140 31726
rect 50540 36652 50596 36708
rect 52668 41468 52724 41524
rect 51996 40962 52052 40964
rect 51996 40910 51998 40962
rect 51998 40910 52050 40962
rect 52050 40910 52052 40962
rect 51996 40908 52052 40910
rect 51996 40460 52052 40516
rect 51884 39506 51940 39508
rect 51884 39454 51886 39506
rect 51886 39454 51938 39506
rect 51938 39454 51940 39506
rect 51884 39452 51940 39454
rect 52220 40460 52276 40516
rect 52332 39452 52388 39508
rect 51996 39004 52052 39060
rect 52220 39116 52276 39172
rect 51884 38556 51940 38612
rect 51548 37212 51604 37268
rect 51436 36428 51492 36484
rect 50556 36090 50612 36092
rect 50556 36038 50558 36090
rect 50558 36038 50610 36090
rect 50610 36038 50612 36090
rect 50556 36036 50612 36038
rect 50660 36090 50716 36092
rect 50660 36038 50662 36090
rect 50662 36038 50714 36090
rect 50714 36038 50716 36090
rect 50660 36036 50716 36038
rect 50764 36090 50820 36092
rect 50764 36038 50766 36090
rect 50766 36038 50818 36090
rect 50818 36038 50820 36090
rect 50764 36036 50820 36038
rect 52220 36988 52276 37044
rect 52444 39058 52500 39060
rect 52444 39006 52446 39058
rect 52446 39006 52498 39058
rect 52498 39006 52500 39058
rect 52444 39004 52500 39006
rect 52892 41692 52948 41748
rect 54348 42082 54404 42084
rect 54348 42030 54350 42082
rect 54350 42030 54402 42082
rect 54402 42030 54404 42082
rect 54348 42028 54404 42030
rect 54236 41804 54292 41860
rect 53004 40572 53060 40628
rect 53004 39506 53060 39508
rect 53004 39454 53006 39506
rect 53006 39454 53058 39506
rect 53058 39454 53060 39506
rect 53004 39452 53060 39454
rect 54124 40572 54180 40628
rect 53228 40460 53284 40516
rect 53340 40348 53396 40404
rect 54012 40402 54068 40404
rect 54012 40350 54014 40402
rect 54014 40350 54066 40402
rect 54066 40350 54068 40402
rect 54012 40348 54068 40350
rect 53116 39116 53172 39172
rect 53452 39564 53508 39620
rect 53004 36706 53060 36708
rect 53004 36654 53006 36706
rect 53006 36654 53058 36706
rect 53058 36654 53060 36706
rect 53004 36652 53060 36654
rect 53228 36482 53284 36484
rect 53228 36430 53230 36482
rect 53230 36430 53282 36482
rect 53282 36430 53284 36482
rect 53228 36428 53284 36430
rect 52332 35756 52388 35812
rect 51884 34914 51940 34916
rect 51884 34862 51886 34914
rect 51886 34862 51938 34914
rect 51938 34862 51940 34914
rect 51884 34860 51940 34862
rect 51996 35420 52052 35476
rect 52108 34972 52164 35028
rect 50556 34522 50612 34524
rect 50556 34470 50558 34522
rect 50558 34470 50610 34522
rect 50610 34470 50612 34522
rect 50556 34468 50612 34470
rect 50660 34522 50716 34524
rect 50660 34470 50662 34522
rect 50662 34470 50714 34522
rect 50714 34470 50716 34522
rect 50660 34468 50716 34470
rect 50764 34522 50820 34524
rect 50764 34470 50766 34522
rect 50766 34470 50818 34522
rect 50818 34470 50820 34522
rect 50764 34468 50820 34470
rect 50316 34188 50372 34244
rect 51324 34188 51380 34244
rect 50652 34130 50708 34132
rect 50652 34078 50654 34130
rect 50654 34078 50706 34130
rect 50706 34078 50708 34130
rect 50652 34076 50708 34078
rect 51996 34242 52052 34244
rect 51996 34190 51998 34242
rect 51998 34190 52050 34242
rect 52050 34190 52052 34242
rect 51996 34188 52052 34190
rect 51548 33628 51604 33684
rect 50764 33234 50820 33236
rect 50764 33182 50766 33234
rect 50766 33182 50818 33234
rect 50818 33182 50820 33234
rect 50764 33180 50820 33182
rect 50556 32954 50612 32956
rect 50556 32902 50558 32954
rect 50558 32902 50610 32954
rect 50610 32902 50612 32954
rect 50556 32900 50612 32902
rect 50660 32954 50716 32956
rect 50660 32902 50662 32954
rect 50662 32902 50714 32954
rect 50714 32902 50716 32954
rect 50660 32900 50716 32902
rect 50764 32954 50820 32956
rect 50764 32902 50766 32954
rect 50766 32902 50818 32954
rect 50818 32902 50820 32954
rect 50764 32900 50820 32902
rect 51660 33068 51716 33124
rect 53564 39058 53620 39060
rect 53564 39006 53566 39058
rect 53566 39006 53618 39058
rect 53618 39006 53620 39058
rect 53564 39004 53620 39006
rect 53452 38556 53508 38612
rect 52668 35026 52724 35028
rect 52668 34974 52670 35026
rect 52670 34974 52722 35026
rect 52722 34974 52724 35026
rect 52668 34972 52724 34974
rect 52780 34860 52836 34916
rect 52444 34130 52500 34132
rect 52444 34078 52446 34130
rect 52446 34078 52498 34130
rect 52498 34078 52500 34130
rect 52444 34076 52500 34078
rect 52668 34188 52724 34244
rect 52332 33180 52388 33236
rect 53116 34636 53172 34692
rect 53452 34914 53508 34916
rect 53452 34862 53454 34914
rect 53454 34862 53506 34914
rect 53506 34862 53508 34914
rect 53452 34860 53508 34862
rect 53340 34242 53396 34244
rect 53340 34190 53342 34242
rect 53342 34190 53394 34242
rect 53394 34190 53396 34242
rect 53340 34188 53396 34190
rect 53004 33628 53060 33684
rect 49756 31724 49812 31780
rect 49756 31388 49812 31444
rect 49532 31164 49588 31220
rect 51548 31890 51604 31892
rect 51548 31838 51550 31890
rect 51550 31838 51602 31890
rect 51602 31838 51604 31890
rect 51548 31836 51604 31838
rect 52108 32562 52164 32564
rect 52108 32510 52110 32562
rect 52110 32510 52162 32562
rect 52162 32510 52164 32562
rect 52108 32508 52164 32510
rect 51996 31836 52052 31892
rect 52332 31948 52388 32004
rect 49868 31052 49924 31108
rect 46620 30716 46676 30772
rect 47180 30882 47236 30884
rect 47180 30830 47182 30882
rect 47182 30830 47234 30882
rect 47234 30830 47236 30882
rect 47180 30828 47236 30830
rect 45612 29820 45668 29876
rect 45836 29650 45892 29652
rect 45836 29598 45838 29650
rect 45838 29598 45890 29650
rect 45890 29598 45892 29650
rect 45836 29596 45892 29598
rect 46284 30210 46340 30212
rect 46284 30158 46286 30210
rect 46286 30158 46338 30210
rect 46338 30158 46340 30210
rect 46284 30156 46340 30158
rect 47740 30716 47796 30772
rect 48972 30604 49028 30660
rect 46396 29986 46452 29988
rect 46396 29934 46398 29986
rect 46398 29934 46450 29986
rect 46450 29934 46452 29986
rect 46396 29932 46452 29934
rect 46172 29820 46228 29876
rect 50204 31500 50260 31556
rect 50556 31386 50612 31388
rect 50556 31334 50558 31386
rect 50558 31334 50610 31386
rect 50610 31334 50612 31386
rect 50556 31332 50612 31334
rect 50660 31386 50716 31388
rect 50660 31334 50662 31386
rect 50662 31334 50714 31386
rect 50714 31334 50716 31386
rect 50660 31332 50716 31334
rect 50764 31386 50820 31388
rect 50764 31334 50766 31386
rect 50766 31334 50818 31386
rect 50818 31334 50820 31386
rect 50764 31332 50820 31334
rect 51100 31106 51156 31108
rect 51100 31054 51102 31106
rect 51102 31054 51154 31106
rect 51154 31054 51156 31106
rect 51100 31052 51156 31054
rect 52780 31948 52836 32004
rect 55356 43314 55412 43316
rect 55356 43262 55358 43314
rect 55358 43262 55410 43314
rect 55410 43262 55412 43314
rect 55356 43260 55412 43262
rect 54684 42700 54740 42756
rect 54908 42140 54964 42196
rect 57148 43260 57204 43316
rect 56700 42754 56756 42756
rect 56700 42702 56702 42754
rect 56702 42702 56754 42754
rect 56754 42702 56756 42754
rect 56700 42700 56756 42702
rect 55692 42140 55748 42196
rect 54684 40908 54740 40964
rect 55244 40908 55300 40964
rect 55132 40572 55188 40628
rect 55468 40460 55524 40516
rect 54236 37212 54292 37268
rect 53900 34914 53956 34916
rect 53900 34862 53902 34914
rect 53902 34862 53954 34914
rect 53954 34862 53956 34914
rect 53900 34860 53956 34862
rect 54124 36988 54180 37044
rect 54572 36988 54628 37044
rect 53676 34690 53732 34692
rect 53676 34638 53678 34690
rect 53678 34638 53730 34690
rect 53730 34638 53732 34690
rect 53676 34636 53732 34638
rect 53676 33292 53732 33348
rect 54460 36428 54516 36484
rect 55468 37212 55524 37268
rect 55244 36988 55300 37044
rect 57820 37378 57876 37380
rect 57820 37326 57822 37378
rect 57822 37326 57874 37378
rect 57874 37326 57876 37378
rect 57820 37324 57876 37326
rect 54124 33628 54180 33684
rect 55244 36482 55300 36484
rect 55244 36430 55246 36482
rect 55246 36430 55298 36482
rect 55298 36430 55300 36482
rect 55244 36428 55300 36430
rect 57596 36988 57652 37044
rect 58156 36988 58212 37044
rect 55468 35810 55524 35812
rect 55468 35758 55470 35810
rect 55470 35758 55522 35810
rect 55522 35758 55524 35810
rect 55468 35756 55524 35758
rect 57820 35868 57876 35924
rect 57932 35756 57988 35812
rect 55580 35532 55636 35588
rect 58156 34972 58212 35028
rect 54572 33346 54628 33348
rect 54572 33294 54574 33346
rect 54574 33294 54626 33346
rect 54626 33294 54628 33346
rect 54572 33292 54628 33294
rect 53564 33234 53620 33236
rect 53564 33182 53566 33234
rect 53566 33182 53618 33234
rect 53618 33182 53620 33234
rect 53564 33180 53620 33182
rect 53228 33122 53284 33124
rect 53228 33070 53230 33122
rect 53230 33070 53282 33122
rect 53282 33070 53284 33122
rect 53228 33068 53284 33070
rect 53228 32674 53284 32676
rect 53228 32622 53230 32674
rect 53230 32622 53282 32674
rect 53282 32622 53284 32674
rect 53228 32620 53284 32622
rect 53452 32508 53508 32564
rect 52556 31612 52612 31668
rect 52892 31554 52948 31556
rect 52892 31502 52894 31554
rect 52894 31502 52946 31554
rect 52946 31502 52948 31554
rect 52892 31500 52948 31502
rect 52444 31164 52500 31220
rect 51884 31052 51940 31108
rect 50988 30940 51044 30996
rect 51660 30940 51716 30996
rect 52556 30770 52612 30772
rect 52556 30718 52558 30770
rect 52558 30718 52610 30770
rect 52610 30718 52612 30770
rect 52556 30716 52612 30718
rect 51212 30322 51268 30324
rect 51212 30270 51214 30322
rect 51214 30270 51266 30322
rect 51266 30270 51268 30322
rect 51212 30268 51268 30270
rect 54124 32508 54180 32564
rect 57148 33628 57204 33684
rect 55580 32732 55636 32788
rect 54684 32620 54740 32676
rect 54124 31836 54180 31892
rect 54684 31836 54740 31892
rect 53676 31164 53732 31220
rect 53004 30994 53060 30996
rect 53004 30942 53006 30994
rect 53006 30942 53058 30994
rect 53058 30942 53060 30994
rect 53004 30940 53060 30942
rect 54348 31164 54404 31220
rect 54124 30994 54180 30996
rect 54124 30942 54126 30994
rect 54126 30942 54178 30994
rect 54178 30942 54180 30994
rect 54124 30940 54180 30942
rect 52668 30322 52724 30324
rect 52668 30270 52670 30322
rect 52670 30270 52722 30322
rect 52722 30270 52724 30322
rect 52668 30268 52724 30270
rect 53340 30716 53396 30772
rect 56588 32562 56644 32564
rect 56588 32510 56590 32562
rect 56590 32510 56642 32562
rect 56642 32510 56644 32562
rect 56588 32508 56644 32510
rect 55580 31778 55636 31780
rect 55580 31726 55582 31778
rect 55582 31726 55634 31778
rect 55634 31726 55636 31778
rect 55580 31724 55636 31726
rect 57260 33068 57316 33124
rect 56700 30940 56756 30996
rect 57932 32284 57988 32340
rect 57820 30940 57876 30996
rect 57932 31612 57988 31668
rect 55020 30770 55076 30772
rect 55020 30718 55022 30770
rect 55022 30718 55074 30770
rect 55074 30718 55076 30770
rect 55020 30716 55076 30718
rect 48972 29986 49028 29988
rect 48972 29934 48974 29986
rect 48974 29934 49026 29986
rect 49026 29934 49028 29986
rect 48972 29932 49028 29934
rect 47068 29820 47124 29876
rect 50556 29818 50612 29820
rect 50556 29766 50558 29818
rect 50558 29766 50610 29818
rect 50610 29766 50612 29818
rect 50556 29764 50612 29766
rect 50660 29818 50716 29820
rect 50660 29766 50662 29818
rect 50662 29766 50714 29818
rect 50714 29766 50716 29818
rect 50660 29764 50716 29766
rect 50764 29818 50820 29820
rect 50764 29766 50766 29818
rect 50766 29766 50818 29818
rect 50818 29766 50820 29818
rect 50764 29764 50820 29766
rect 55580 29708 55636 29764
rect 46620 29484 46676 29540
rect 49756 28812 49812 28868
rect 48748 28140 48804 28196
rect 43260 27580 43316 27636
rect 43148 27186 43204 27188
rect 43148 27134 43150 27186
rect 43150 27134 43202 27186
rect 43202 27134 43204 27186
rect 43148 27132 43204 27134
rect 42812 26796 42868 26852
rect 43148 26460 43204 26516
rect 45276 26908 45332 26964
rect 39900 25788 39956 25844
rect 39452 25564 39508 25620
rect 38332 25452 38388 25508
rect 40236 25506 40292 25508
rect 40236 25454 40238 25506
rect 40238 25454 40290 25506
rect 40290 25454 40292 25506
rect 40236 25452 40292 25454
rect 40684 25506 40740 25508
rect 40684 25454 40686 25506
rect 40686 25454 40738 25506
rect 40738 25454 40740 25506
rect 40684 25452 40740 25454
rect 39004 25340 39060 25396
rect 39452 25282 39508 25284
rect 39452 25230 39454 25282
rect 39454 25230 39506 25282
rect 39506 25230 39508 25282
rect 39452 25228 39508 25230
rect 39900 25282 39956 25284
rect 39900 25230 39902 25282
rect 39902 25230 39954 25282
rect 39954 25230 39956 25282
rect 39900 25228 39956 25230
rect 39228 24780 39284 24836
rect 37660 23884 37716 23940
rect 38108 23884 38164 23940
rect 37436 23714 37492 23716
rect 37436 23662 37438 23714
rect 37438 23662 37490 23714
rect 37490 23662 37492 23714
rect 37436 23660 37492 23662
rect 37100 23100 37156 23156
rect 36540 22370 36596 22372
rect 36540 22318 36542 22370
rect 36542 22318 36594 22370
rect 36594 22318 36596 22370
rect 36540 22316 36596 22318
rect 36988 22092 37044 22148
rect 39340 23826 39396 23828
rect 39340 23774 39342 23826
rect 39342 23774 39394 23826
rect 39394 23774 39396 23826
rect 39340 23772 39396 23774
rect 38556 23436 38612 23492
rect 38668 23100 38724 23156
rect 37436 22370 37492 22372
rect 37436 22318 37438 22370
rect 37438 22318 37490 22370
rect 37490 22318 37492 22370
rect 37436 22316 37492 22318
rect 35980 21698 36036 21700
rect 35980 21646 35982 21698
rect 35982 21646 36034 21698
rect 36034 21646 36036 21698
rect 35980 21644 36036 21646
rect 35868 21420 35924 21476
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 35084 20860 35140 20916
rect 35644 20636 35700 20692
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 36204 21532 36260 21588
rect 36428 21474 36484 21476
rect 36428 21422 36430 21474
rect 36430 21422 36482 21474
rect 36482 21422 36484 21474
rect 36428 21420 36484 21422
rect 36204 19516 36260 19572
rect 34972 18508 35028 18564
rect 35084 18396 35140 18452
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 35980 18284 36036 18340
rect 35868 18226 35924 18228
rect 35868 18174 35870 18226
rect 35870 18174 35922 18226
rect 35922 18174 35924 18226
rect 35868 18172 35924 18174
rect 35644 17666 35700 17668
rect 35644 17614 35646 17666
rect 35646 17614 35698 17666
rect 35698 17614 35700 17666
rect 35644 17612 35700 17614
rect 34300 16044 34356 16100
rect 33404 15986 33460 15988
rect 33404 15934 33406 15986
rect 33406 15934 33458 15986
rect 33458 15934 33460 15986
rect 33404 15932 33460 15934
rect 33068 15260 33124 15316
rect 34188 15372 34244 15428
rect 33740 15314 33796 15316
rect 33740 15262 33742 15314
rect 33742 15262 33794 15314
rect 33794 15262 33796 15314
rect 33740 15260 33796 15262
rect 32732 14306 32788 14308
rect 32732 14254 32734 14306
rect 32734 14254 32786 14306
rect 32786 14254 32788 14306
rect 32732 14252 32788 14254
rect 32508 13970 32564 13972
rect 32508 13918 32510 13970
rect 32510 13918 32562 13970
rect 32562 13918 32564 13970
rect 32508 13916 32564 13918
rect 33180 13580 33236 13636
rect 33628 14252 33684 14308
rect 34412 16380 34468 16436
rect 34636 15932 34692 15988
rect 35756 17442 35812 17444
rect 35756 17390 35758 17442
rect 35758 17390 35810 17442
rect 35810 17390 35812 17442
rect 35756 17388 35812 17390
rect 35532 17052 35588 17108
rect 34972 16716 35028 16772
rect 34972 16380 35028 16436
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 35308 16268 35364 16324
rect 35084 15820 35140 15876
rect 34860 15596 34916 15652
rect 34860 15426 34916 15428
rect 34860 15374 34862 15426
rect 34862 15374 34914 15426
rect 34914 15374 34916 15426
rect 34860 15372 34916 15374
rect 34860 15036 34916 15092
rect 34524 14530 34580 14532
rect 34524 14478 34526 14530
rect 34526 14478 34578 14530
rect 34578 14478 34580 14530
rect 34524 14476 34580 14478
rect 34076 13580 34132 13636
rect 34188 13804 34244 13860
rect 33628 13468 33684 13524
rect 32508 10722 32564 10724
rect 32508 10670 32510 10722
rect 32510 10670 32562 10722
rect 32562 10670 32564 10722
rect 32508 10668 32564 10670
rect 32284 9772 32340 9828
rect 32172 9660 32228 9716
rect 31164 9436 31220 9492
rect 31052 9324 31108 9380
rect 32060 9324 32116 9380
rect 32284 9602 32340 9604
rect 32284 9550 32286 9602
rect 32286 9550 32338 9602
rect 32338 9550 32340 9602
rect 32284 9548 32340 9550
rect 32956 9996 33012 10052
rect 33068 10444 33124 10500
rect 32172 9212 32228 9268
rect 31388 8818 31444 8820
rect 31388 8766 31390 8818
rect 31390 8766 31442 8818
rect 31442 8766 31444 8818
rect 31388 8764 31444 8766
rect 31388 8204 31444 8260
rect 30940 6636 30996 6692
rect 30492 6578 30548 6580
rect 30492 6526 30494 6578
rect 30494 6526 30546 6578
rect 30546 6526 30548 6578
rect 30492 6524 30548 6526
rect 31388 7532 31444 7588
rect 32284 8764 32340 8820
rect 31836 8316 31892 8372
rect 31948 7474 32004 7476
rect 31948 7422 31950 7474
rect 31950 7422 32002 7474
rect 32002 7422 32004 7474
rect 31948 7420 32004 7422
rect 31052 6300 31108 6356
rect 30044 5404 30100 5460
rect 29260 5068 29316 5124
rect 29708 5122 29764 5124
rect 29708 5070 29710 5122
rect 29710 5070 29762 5122
rect 29762 5070 29764 5122
rect 29708 5068 29764 5070
rect 30044 5068 30100 5124
rect 30940 5906 30996 5908
rect 30940 5854 30942 5906
rect 30942 5854 30994 5906
rect 30994 5854 30996 5906
rect 30940 5852 30996 5854
rect 30940 5516 30996 5572
rect 30492 4956 30548 5012
rect 29260 4732 29316 4788
rect 30380 4898 30436 4900
rect 30380 4846 30382 4898
rect 30382 4846 30434 4898
rect 30434 4846 30436 4898
rect 30380 4844 30436 4846
rect 29484 4114 29540 4116
rect 29484 4062 29486 4114
rect 29486 4062 29538 4114
rect 29538 4062 29540 4114
rect 29484 4060 29540 4062
rect 30268 3612 30324 3668
rect 32060 6300 32116 6356
rect 31836 5628 31892 5684
rect 32396 6690 32452 6692
rect 32396 6638 32398 6690
rect 32398 6638 32450 6690
rect 32450 6638 32452 6690
rect 32396 6636 32452 6638
rect 32172 5740 32228 5796
rect 32172 5404 32228 5460
rect 31500 5180 31556 5236
rect 31612 5122 31668 5124
rect 31612 5070 31614 5122
rect 31614 5070 31666 5122
rect 31666 5070 31668 5122
rect 31612 5068 31668 5070
rect 31724 4844 31780 4900
rect 31948 5180 32004 5236
rect 32060 5068 32116 5124
rect 32172 4508 32228 4564
rect 32284 5180 32340 5236
rect 31612 3500 31668 3556
rect 30940 3388 30996 3444
rect 32172 3164 32228 3220
rect 32732 9660 32788 9716
rect 32620 9324 32676 9380
rect 33404 9884 33460 9940
rect 33068 7586 33124 7588
rect 33068 7534 33070 7586
rect 33070 7534 33122 7586
rect 33122 7534 33124 7586
rect 33068 7532 33124 7534
rect 34748 13804 34804 13860
rect 33852 11788 33908 11844
rect 33628 8652 33684 8708
rect 33740 9548 33796 9604
rect 33740 8428 33796 8484
rect 33740 8204 33796 8260
rect 33292 7474 33348 7476
rect 33292 7422 33294 7474
rect 33294 7422 33346 7474
rect 33346 7422 33348 7474
rect 33292 7420 33348 7422
rect 33516 7250 33572 7252
rect 33516 7198 33518 7250
rect 33518 7198 33570 7250
rect 33570 7198 33572 7250
rect 33516 7196 33572 7198
rect 32732 6524 32788 6580
rect 33516 6076 33572 6132
rect 32396 3666 32452 3668
rect 32396 3614 32398 3666
rect 32398 3614 32450 3666
rect 32450 3614 32452 3666
rect 32396 3612 32452 3614
rect 35532 16098 35588 16100
rect 35532 16046 35534 16098
rect 35534 16046 35586 16098
rect 35586 16046 35588 16098
rect 35532 16044 35588 16046
rect 35868 15986 35924 15988
rect 35868 15934 35870 15986
rect 35870 15934 35922 15986
rect 35922 15934 35924 15986
rect 35868 15932 35924 15934
rect 35756 15820 35812 15876
rect 36092 16716 36148 16772
rect 36204 16098 36260 16100
rect 36204 16046 36206 16098
rect 36206 16046 36258 16098
rect 36258 16046 36260 16098
rect 36204 16044 36260 16046
rect 35980 15036 36036 15092
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 35644 14476 35700 14532
rect 35196 14364 35252 14420
rect 34972 13916 35028 13972
rect 35532 14306 35588 14308
rect 35532 14254 35534 14306
rect 35534 14254 35586 14306
rect 35586 14254 35588 14306
rect 35532 14252 35588 14254
rect 37884 21756 37940 21812
rect 37324 21420 37380 21476
rect 37100 20076 37156 20132
rect 37772 20130 37828 20132
rect 37772 20078 37774 20130
rect 37774 20078 37826 20130
rect 37826 20078 37828 20130
rect 37772 20076 37828 20078
rect 37324 19404 37380 19460
rect 39340 21868 39396 21924
rect 38556 21308 38612 21364
rect 39004 21756 39060 21812
rect 40012 24220 40068 24276
rect 42588 26236 42644 26292
rect 41020 25228 41076 25284
rect 41132 24722 41188 24724
rect 41132 24670 41134 24722
rect 41134 24670 41186 24722
rect 41186 24670 41188 24722
rect 41132 24668 41188 24670
rect 41580 25506 41636 25508
rect 41580 25454 41582 25506
rect 41582 25454 41634 25506
rect 41634 25454 41636 25506
rect 41580 25452 41636 25454
rect 43260 26290 43316 26292
rect 43260 26238 43262 26290
rect 43262 26238 43314 26290
rect 43314 26238 43316 26290
rect 43260 26236 43316 26238
rect 44492 26290 44548 26292
rect 44492 26238 44494 26290
rect 44494 26238 44546 26290
rect 44546 26238 44548 26290
rect 44492 26236 44548 26238
rect 43708 26178 43764 26180
rect 43708 26126 43710 26178
rect 43710 26126 43762 26178
rect 43762 26126 43764 26178
rect 43708 26124 43764 26126
rect 44380 26178 44436 26180
rect 44380 26126 44382 26178
rect 44382 26126 44434 26178
rect 44434 26126 44436 26178
rect 44380 26124 44436 26126
rect 42476 24722 42532 24724
rect 42476 24670 42478 24722
rect 42478 24670 42530 24722
rect 42530 24670 42532 24722
rect 42476 24668 42532 24670
rect 41020 23378 41076 23380
rect 41020 23326 41022 23378
rect 41022 23326 41074 23378
rect 41074 23326 41076 23378
rect 41020 23324 41076 23326
rect 42140 24220 42196 24276
rect 40908 23154 40964 23156
rect 40908 23102 40910 23154
rect 40910 23102 40962 23154
rect 40962 23102 40964 23154
rect 40908 23100 40964 23102
rect 40236 22988 40292 23044
rect 40012 22092 40068 22148
rect 44044 24220 44100 24276
rect 42140 23378 42196 23380
rect 42140 23326 42142 23378
rect 42142 23326 42194 23378
rect 42194 23326 42196 23378
rect 42140 23324 42196 23326
rect 43036 23772 43092 23828
rect 43932 23826 43988 23828
rect 43932 23774 43934 23826
rect 43934 23774 43986 23826
rect 43986 23774 43988 23826
rect 43932 23772 43988 23774
rect 44156 23996 44212 24052
rect 44940 24220 44996 24276
rect 45948 27244 46004 27300
rect 45612 26962 45668 26964
rect 45612 26910 45614 26962
rect 45614 26910 45666 26962
rect 45666 26910 45668 26962
rect 45612 26908 45668 26910
rect 45612 25452 45668 25508
rect 46508 27020 46564 27076
rect 46284 26012 46340 26068
rect 45388 24892 45444 24948
rect 47628 26796 47684 26852
rect 50556 28250 50612 28252
rect 50556 28198 50558 28250
rect 50558 28198 50610 28250
rect 50610 28198 50612 28250
rect 50556 28196 50612 28198
rect 50660 28250 50716 28252
rect 50660 28198 50662 28250
rect 50662 28198 50714 28250
rect 50714 28198 50716 28250
rect 50660 28196 50716 28198
rect 50764 28250 50820 28252
rect 50764 28198 50766 28250
rect 50766 28198 50818 28250
rect 50818 28198 50820 28250
rect 50764 28196 50820 28198
rect 48076 27074 48132 27076
rect 48076 27022 48078 27074
rect 48078 27022 48130 27074
rect 48130 27022 48132 27074
rect 48076 27020 48132 27022
rect 48748 26962 48804 26964
rect 48748 26910 48750 26962
rect 48750 26910 48802 26962
rect 48802 26910 48804 26962
rect 48748 26908 48804 26910
rect 47852 26796 47908 26852
rect 47404 26066 47460 26068
rect 47404 26014 47406 26066
rect 47406 26014 47458 26066
rect 47458 26014 47460 26066
rect 47404 26012 47460 26014
rect 47404 25564 47460 25620
rect 46284 25340 46340 25396
rect 46060 24946 46116 24948
rect 46060 24894 46062 24946
rect 46062 24894 46114 24946
rect 46114 24894 46116 24946
rect 46060 24892 46116 24894
rect 45388 24220 45444 24276
rect 45052 23996 45108 24052
rect 45836 24050 45892 24052
rect 45836 23998 45838 24050
rect 45838 23998 45890 24050
rect 45890 23998 45892 24050
rect 45836 23996 45892 23998
rect 45276 23548 45332 23604
rect 42812 23042 42868 23044
rect 42812 22990 42814 23042
rect 42814 22990 42866 23042
rect 42866 22990 42868 23042
rect 42812 22988 42868 22990
rect 40460 22204 40516 22260
rect 41244 22258 41300 22260
rect 41244 22206 41246 22258
rect 41246 22206 41298 22258
rect 41298 22206 41300 22258
rect 41244 22204 41300 22206
rect 40908 22092 40964 22148
rect 40124 21868 40180 21924
rect 40236 21308 40292 21364
rect 39564 20860 39620 20916
rect 40012 19964 40068 20020
rect 42588 22370 42644 22372
rect 42588 22318 42590 22370
rect 42590 22318 42642 22370
rect 42642 22318 42644 22370
rect 42588 22316 42644 22318
rect 41916 21810 41972 21812
rect 41916 21758 41918 21810
rect 41918 21758 41970 21810
rect 41970 21758 41972 21810
rect 41916 21756 41972 21758
rect 42476 21308 42532 21364
rect 40796 19964 40852 20020
rect 38668 19516 38724 19572
rect 39900 19516 39956 19572
rect 39004 19404 39060 19460
rect 37324 19180 37380 19236
rect 37212 18732 37268 18788
rect 36988 18562 37044 18564
rect 36988 18510 36990 18562
rect 36990 18510 37042 18562
rect 37042 18510 37044 18562
rect 36988 18508 37044 18510
rect 36540 18396 36596 18452
rect 36428 18338 36484 18340
rect 36428 18286 36430 18338
rect 36430 18286 36482 18338
rect 36482 18286 36484 18338
rect 36428 18284 36484 18286
rect 38780 19234 38836 19236
rect 38780 19182 38782 19234
rect 38782 19182 38834 19234
rect 38834 19182 38836 19234
rect 38780 19180 38836 19182
rect 37884 18562 37940 18564
rect 37884 18510 37886 18562
rect 37886 18510 37938 18562
rect 37938 18510 37940 18562
rect 37884 18508 37940 18510
rect 38892 18508 38948 18564
rect 38332 18450 38388 18452
rect 38332 18398 38334 18450
rect 38334 18398 38386 18450
rect 38386 18398 38388 18450
rect 38332 18396 38388 18398
rect 37884 18338 37940 18340
rect 37884 18286 37886 18338
rect 37886 18286 37938 18338
rect 37938 18286 37940 18338
rect 37884 18284 37940 18286
rect 38556 18284 38612 18340
rect 37548 17890 37604 17892
rect 37548 17838 37550 17890
rect 37550 17838 37602 17890
rect 37602 17838 37604 17890
rect 37548 17836 37604 17838
rect 38780 17666 38836 17668
rect 38780 17614 38782 17666
rect 38782 17614 38834 17666
rect 38834 17614 38836 17666
rect 38780 17612 38836 17614
rect 37100 17442 37156 17444
rect 37100 17390 37102 17442
rect 37102 17390 37154 17442
rect 37154 17390 37156 17442
rect 37100 17388 37156 17390
rect 38332 17500 38388 17556
rect 38108 17388 38164 17444
rect 36540 17052 36596 17108
rect 36764 16882 36820 16884
rect 36764 16830 36766 16882
rect 36766 16830 36818 16882
rect 36818 16830 36820 16882
rect 36764 16828 36820 16830
rect 36428 16268 36484 16324
rect 37324 16098 37380 16100
rect 37324 16046 37326 16098
rect 37326 16046 37378 16098
rect 37378 16046 37380 16098
rect 37324 16044 37380 16046
rect 35420 13804 35476 13860
rect 36204 13916 36260 13972
rect 35084 13692 35140 13748
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35644 13580 35700 13636
rect 35308 12850 35364 12852
rect 35308 12798 35310 12850
rect 35310 12798 35362 12850
rect 35362 12798 35364 12850
rect 35308 12796 35364 12798
rect 36540 14476 36596 14532
rect 36988 15036 37044 15092
rect 36876 14588 36932 14644
rect 36764 14364 36820 14420
rect 37660 15820 37716 15876
rect 37660 15596 37716 15652
rect 37324 15314 37380 15316
rect 37324 15262 37326 15314
rect 37326 15262 37378 15314
rect 37378 15262 37380 15314
rect 37324 15260 37380 15262
rect 37772 15260 37828 15316
rect 38780 17388 38836 17444
rect 38668 16044 38724 16100
rect 38892 15484 38948 15540
rect 39116 18732 39172 18788
rect 39676 18508 39732 18564
rect 40572 19346 40628 19348
rect 40572 19294 40574 19346
rect 40574 19294 40626 19346
rect 40626 19294 40628 19346
rect 40572 19292 40628 19294
rect 40348 18338 40404 18340
rect 40348 18286 40350 18338
rect 40350 18286 40402 18338
rect 40402 18286 40404 18338
rect 40348 18284 40404 18286
rect 41356 20018 41412 20020
rect 41356 19966 41358 20018
rect 41358 19966 41410 20018
rect 41410 19966 41412 20018
rect 41356 19964 41412 19966
rect 41132 19852 41188 19908
rect 41692 19906 41748 19908
rect 41692 19854 41694 19906
rect 41694 19854 41746 19906
rect 41746 19854 41748 19906
rect 41692 19852 41748 19854
rect 42364 19852 42420 19908
rect 42476 19964 42532 20020
rect 41020 19346 41076 19348
rect 41020 19294 41022 19346
rect 41022 19294 41074 19346
rect 41074 19294 41076 19346
rect 41020 19292 41076 19294
rect 42028 19234 42084 19236
rect 42028 19182 42030 19234
rect 42030 19182 42082 19234
rect 42082 19182 42084 19234
rect 42028 19180 42084 19182
rect 42700 20018 42756 20020
rect 42700 19966 42702 20018
rect 42702 19966 42754 20018
rect 42754 19966 42756 20018
rect 42700 19964 42756 19966
rect 42924 19852 42980 19908
rect 43932 23154 43988 23156
rect 43932 23102 43934 23154
rect 43934 23102 43986 23154
rect 43986 23102 43988 23154
rect 43932 23100 43988 23102
rect 43372 21868 43428 21924
rect 44268 22428 44324 22484
rect 44604 22764 44660 22820
rect 44268 21868 44324 21924
rect 44492 21868 44548 21924
rect 43708 21756 43764 21812
rect 43148 20018 43204 20020
rect 43148 19966 43150 20018
rect 43150 19966 43202 20018
rect 43202 19966 43204 20018
rect 43148 19964 43204 19966
rect 43708 20802 43764 20804
rect 43708 20750 43710 20802
rect 43710 20750 43762 20802
rect 43762 20750 43764 20802
rect 43708 20748 43764 20750
rect 43820 20130 43876 20132
rect 43820 20078 43822 20130
rect 43822 20078 43874 20130
rect 43874 20078 43876 20130
rect 43820 20076 43876 20078
rect 43596 20018 43652 20020
rect 43596 19966 43598 20018
rect 43598 19966 43650 20018
rect 43650 19966 43652 20018
rect 43596 19964 43652 19966
rect 43932 19852 43988 19908
rect 42812 19458 42868 19460
rect 42812 19406 42814 19458
rect 42814 19406 42866 19458
rect 42866 19406 42868 19458
rect 42812 19404 42868 19406
rect 43484 19740 43540 19796
rect 44156 19740 44212 19796
rect 43596 19628 43652 19684
rect 41804 19122 41860 19124
rect 41804 19070 41806 19122
rect 41806 19070 41858 19122
rect 41858 19070 41860 19122
rect 41804 19068 41860 19070
rect 43148 19010 43204 19012
rect 43148 18958 43150 19010
rect 43150 18958 43202 19010
rect 43202 18958 43204 19010
rect 43148 18956 43204 18958
rect 41916 18396 41972 18452
rect 41356 18284 41412 18340
rect 39228 17612 39284 17668
rect 40348 17666 40404 17668
rect 40348 17614 40350 17666
rect 40350 17614 40402 17666
rect 40402 17614 40404 17666
rect 40348 17612 40404 17614
rect 39228 17388 39284 17444
rect 39564 16994 39620 16996
rect 39564 16942 39566 16994
rect 39566 16942 39618 16994
rect 39618 16942 39620 16994
rect 39564 16940 39620 16942
rect 39452 15820 39508 15876
rect 39788 16882 39844 16884
rect 39788 16830 39790 16882
rect 39790 16830 39842 16882
rect 39842 16830 39844 16882
rect 39788 16828 39844 16830
rect 40460 16882 40516 16884
rect 40460 16830 40462 16882
rect 40462 16830 40514 16882
rect 40514 16830 40516 16882
rect 40460 16828 40516 16830
rect 39900 16770 39956 16772
rect 39900 16718 39902 16770
rect 39902 16718 39954 16770
rect 39954 16718 39956 16770
rect 39900 16716 39956 16718
rect 38108 14700 38164 14756
rect 38332 14588 38388 14644
rect 37212 14476 37268 14532
rect 37100 13916 37156 13972
rect 36428 12796 36484 12852
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 36428 12178 36484 12180
rect 36428 12126 36430 12178
rect 36430 12126 36482 12178
rect 36482 12126 36484 12178
rect 36428 12124 36484 12126
rect 36316 11564 36372 11620
rect 34076 10668 34132 10724
rect 34300 10556 34356 10612
rect 36540 11282 36596 11284
rect 36540 11230 36542 11282
rect 36542 11230 36594 11282
rect 36594 11230 36596 11282
rect 36540 11228 36596 11230
rect 36316 11170 36372 11172
rect 36316 11118 36318 11170
rect 36318 11118 36370 11170
rect 36370 11118 36372 11170
rect 36316 11116 36372 11118
rect 35420 10780 35476 10836
rect 36428 10610 36484 10612
rect 36428 10558 36430 10610
rect 36430 10558 36482 10610
rect 36482 10558 36484 10610
rect 36428 10556 36484 10558
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 33964 9324 34020 9380
rect 34860 9938 34916 9940
rect 34860 9886 34862 9938
rect 34862 9886 34914 9938
rect 34914 9886 34916 9938
rect 34860 9884 34916 9886
rect 35420 9996 35476 10052
rect 34188 8988 34244 9044
rect 35084 9826 35140 9828
rect 35084 9774 35086 9826
rect 35086 9774 35138 9826
rect 35138 9774 35140 9826
rect 35084 9772 35140 9774
rect 35644 9772 35700 9828
rect 34748 9660 34804 9716
rect 35420 9602 35476 9604
rect 35420 9550 35422 9602
rect 35422 9550 35474 9602
rect 35474 9550 35476 9602
rect 35420 9548 35476 9550
rect 35196 9266 35252 9268
rect 35196 9214 35198 9266
rect 35198 9214 35250 9266
rect 35250 9214 35252 9266
rect 35196 9212 35252 9214
rect 36540 9212 36596 9268
rect 35868 9042 35924 9044
rect 35868 8990 35870 9042
rect 35870 8990 35922 9042
rect 35922 8990 35924 9042
rect 35868 8988 35924 8990
rect 34524 8652 34580 8708
rect 34412 8482 34468 8484
rect 34412 8430 34414 8482
rect 34414 8430 34466 8482
rect 34466 8430 34468 8482
rect 34412 8428 34468 8430
rect 34860 7980 34916 8036
rect 34300 7532 34356 7588
rect 34076 7420 34132 7476
rect 34636 7196 34692 7252
rect 33852 6412 33908 6468
rect 34300 6690 34356 6692
rect 34300 6638 34302 6690
rect 34302 6638 34354 6690
rect 34354 6638 34356 6690
rect 34300 6636 34356 6638
rect 34188 6018 34244 6020
rect 34188 5966 34190 6018
rect 34190 5966 34242 6018
rect 34242 5966 34244 6018
rect 34188 5964 34244 5966
rect 33740 5852 33796 5908
rect 33068 5292 33124 5348
rect 33516 5234 33572 5236
rect 33516 5182 33518 5234
rect 33518 5182 33570 5234
rect 33570 5182 33572 5234
rect 33516 5180 33572 5182
rect 32620 3500 32676 3556
rect 32956 4732 33012 4788
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 36204 8428 36260 8484
rect 36428 8370 36484 8372
rect 36428 8318 36430 8370
rect 36430 8318 36482 8370
rect 36482 8318 36484 8370
rect 36428 8316 36484 8318
rect 35756 8258 35812 8260
rect 35756 8206 35758 8258
rect 35758 8206 35810 8258
rect 35810 8206 35812 8258
rect 35756 8204 35812 8206
rect 35532 7980 35588 8036
rect 35308 7250 35364 7252
rect 35308 7198 35310 7250
rect 35310 7198 35362 7250
rect 35362 7198 35364 7250
rect 35308 7196 35364 7198
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35084 6636 35140 6692
rect 34412 5906 34468 5908
rect 34412 5854 34414 5906
rect 34414 5854 34466 5906
rect 34466 5854 34468 5906
rect 34412 5852 34468 5854
rect 34300 5516 34356 5572
rect 34524 5628 34580 5684
rect 34524 4844 34580 4900
rect 34636 6412 34692 6468
rect 34412 4732 34468 4788
rect 33964 4284 34020 4340
rect 33628 4060 33684 4116
rect 34860 4450 34916 4452
rect 34860 4398 34862 4450
rect 34862 4398 34914 4450
rect 34914 4398 34916 4450
rect 34860 4396 34916 4398
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 35084 4956 35140 5012
rect 34972 3724 35028 3780
rect 34300 2492 34356 2548
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 35308 3554 35364 3556
rect 35308 3502 35310 3554
rect 35310 3502 35362 3554
rect 35362 3502 35364 3554
rect 35308 3500 35364 3502
rect 35644 6524 35700 6580
rect 36316 8034 36372 8036
rect 36316 7982 36318 8034
rect 36318 7982 36370 8034
rect 36370 7982 36372 8034
rect 36316 7980 36372 7982
rect 35868 6748 35924 6804
rect 36204 6300 36260 6356
rect 36428 7420 36484 7476
rect 36540 7196 36596 7252
rect 36428 6466 36484 6468
rect 36428 6414 36430 6466
rect 36430 6414 36482 6466
rect 36482 6414 36484 6466
rect 36428 6412 36484 6414
rect 36316 6076 36372 6132
rect 35756 5292 35812 5348
rect 35868 5740 35924 5796
rect 35756 5122 35812 5124
rect 35756 5070 35758 5122
rect 35758 5070 35810 5122
rect 35810 5070 35812 5122
rect 35756 5068 35812 5070
rect 35980 4898 36036 4900
rect 35980 4846 35982 4898
rect 35982 4846 36034 4898
rect 36034 4846 36036 4898
rect 35980 4844 36036 4846
rect 35532 3164 35588 3220
rect 35644 3612 35700 3668
rect 36204 4898 36260 4900
rect 36204 4846 36206 4898
rect 36206 4846 36258 4898
rect 36258 4846 36260 4898
rect 36204 4844 36260 4846
rect 36764 13244 36820 13300
rect 37772 14252 37828 14308
rect 37548 13746 37604 13748
rect 37548 13694 37550 13746
rect 37550 13694 37602 13746
rect 37602 13694 37604 13746
rect 37548 13692 37604 13694
rect 38668 14418 38724 14420
rect 38668 14366 38670 14418
rect 38670 14366 38722 14418
rect 38722 14366 38724 14418
rect 38668 14364 38724 14366
rect 38332 13692 38388 13748
rect 37212 13468 37268 13524
rect 38220 13468 38276 13524
rect 38444 13804 38500 13860
rect 37100 12572 37156 12628
rect 38108 12684 38164 12740
rect 37660 12460 37716 12516
rect 37100 12178 37156 12180
rect 37100 12126 37102 12178
rect 37102 12126 37154 12178
rect 37154 12126 37156 12178
rect 37100 12124 37156 12126
rect 36764 12012 36820 12068
rect 37548 11788 37604 11844
rect 38556 12850 38612 12852
rect 38556 12798 38558 12850
rect 38558 12798 38610 12850
rect 38610 12798 38612 12850
rect 38556 12796 38612 12798
rect 38780 12738 38836 12740
rect 38780 12686 38782 12738
rect 38782 12686 38834 12738
rect 38834 12686 38836 12738
rect 38780 12684 38836 12686
rect 36764 11564 36820 11620
rect 36428 5180 36484 5236
rect 36316 4508 36372 4564
rect 35980 3276 36036 3332
rect 36316 3836 36372 3892
rect 37324 11282 37380 11284
rect 37324 11230 37326 11282
rect 37326 11230 37378 11282
rect 37378 11230 37380 11282
rect 37324 11228 37380 11230
rect 37436 10780 37492 10836
rect 37884 10668 37940 10724
rect 38332 12290 38388 12292
rect 38332 12238 38334 12290
rect 38334 12238 38386 12290
rect 38386 12238 38388 12290
rect 38332 12236 38388 12238
rect 38892 12290 38948 12292
rect 38892 12238 38894 12290
rect 38894 12238 38946 12290
rect 38946 12238 38948 12290
rect 38892 12236 38948 12238
rect 38444 12178 38500 12180
rect 38444 12126 38446 12178
rect 38446 12126 38498 12178
rect 38498 12126 38500 12178
rect 38444 12124 38500 12126
rect 37996 11116 38052 11172
rect 37772 10444 37828 10500
rect 38892 11394 38948 11396
rect 38892 11342 38894 11394
rect 38894 11342 38946 11394
rect 38946 11342 38948 11394
rect 38892 11340 38948 11342
rect 38220 10780 38276 10836
rect 37996 10108 38052 10164
rect 37548 9826 37604 9828
rect 37548 9774 37550 9826
rect 37550 9774 37602 9826
rect 37602 9774 37604 9826
rect 37548 9772 37604 9774
rect 37100 9660 37156 9716
rect 37884 9714 37940 9716
rect 37884 9662 37886 9714
rect 37886 9662 37938 9714
rect 37938 9662 37940 9714
rect 37884 9660 37940 9662
rect 37212 9154 37268 9156
rect 37212 9102 37214 9154
rect 37214 9102 37266 9154
rect 37266 9102 37268 9154
rect 37212 9100 37268 9102
rect 37100 8370 37156 8372
rect 37100 8318 37102 8370
rect 37102 8318 37154 8370
rect 37154 8318 37156 8370
rect 37100 8316 37156 8318
rect 37324 8316 37380 8372
rect 37884 9212 37940 9268
rect 37772 9154 37828 9156
rect 37772 9102 37774 9154
rect 37774 9102 37826 9154
rect 37826 9102 37828 9154
rect 37772 9100 37828 9102
rect 37772 8204 37828 8260
rect 36988 7420 37044 7476
rect 37548 7474 37604 7476
rect 37548 7422 37550 7474
rect 37550 7422 37602 7474
rect 37602 7422 37604 7474
rect 37548 7420 37604 7422
rect 37436 6914 37492 6916
rect 37436 6862 37438 6914
rect 37438 6862 37490 6914
rect 37490 6862 37492 6914
rect 37436 6860 37492 6862
rect 37212 6802 37268 6804
rect 37212 6750 37214 6802
rect 37214 6750 37266 6802
rect 37266 6750 37268 6802
rect 37212 6748 37268 6750
rect 37100 6188 37156 6244
rect 38108 8428 38164 8484
rect 38220 9826 38276 9828
rect 38220 9774 38222 9826
rect 38222 9774 38274 9826
rect 38274 9774 38276 9826
rect 38220 9772 38276 9774
rect 38556 10220 38612 10276
rect 38444 10108 38500 10164
rect 38892 9938 38948 9940
rect 38892 9886 38894 9938
rect 38894 9886 38946 9938
rect 38946 9886 38948 9938
rect 38892 9884 38948 9886
rect 38668 9212 38724 9268
rect 39004 9602 39060 9604
rect 39004 9550 39006 9602
rect 39006 9550 39058 9602
rect 39058 9550 39060 9602
rect 39004 9548 39060 9550
rect 39004 9154 39060 9156
rect 39004 9102 39006 9154
rect 39006 9102 39058 9154
rect 39058 9102 39060 9154
rect 39004 9100 39060 9102
rect 38444 7196 38500 7252
rect 38220 7084 38276 7140
rect 38556 6972 38612 7028
rect 38668 6860 38724 6916
rect 39004 7420 39060 7476
rect 39788 16098 39844 16100
rect 39788 16046 39790 16098
rect 39790 16046 39842 16098
rect 39842 16046 39844 16098
rect 39788 16044 39844 16046
rect 39900 15538 39956 15540
rect 39900 15486 39902 15538
rect 39902 15486 39954 15538
rect 39954 15486 39956 15538
rect 39900 15484 39956 15486
rect 41132 15484 41188 15540
rect 41692 18338 41748 18340
rect 41692 18286 41694 18338
rect 41694 18286 41746 18338
rect 41746 18286 41748 18338
rect 41692 18284 41748 18286
rect 41468 16044 41524 16100
rect 41804 16156 41860 16212
rect 42812 18396 42868 18452
rect 42252 18284 42308 18340
rect 42476 17666 42532 17668
rect 42476 17614 42478 17666
rect 42478 17614 42530 17666
rect 42530 17614 42532 17666
rect 42476 17612 42532 17614
rect 42140 17052 42196 17108
rect 42028 16716 42084 16772
rect 41692 15372 41748 15428
rect 42028 15260 42084 15316
rect 39564 13746 39620 13748
rect 39564 13694 39566 13746
rect 39566 13694 39618 13746
rect 39618 13694 39620 13746
rect 39564 13692 39620 13694
rect 41132 13692 41188 13748
rect 40124 13634 40180 13636
rect 40124 13582 40126 13634
rect 40126 13582 40178 13634
rect 40178 13582 40180 13634
rect 40124 13580 40180 13582
rect 39788 13522 39844 13524
rect 39788 13470 39790 13522
rect 39790 13470 39842 13522
rect 39842 13470 39844 13522
rect 39788 13468 39844 13470
rect 39676 12850 39732 12852
rect 39676 12798 39678 12850
rect 39678 12798 39730 12850
rect 39730 12798 39732 12850
rect 39676 12796 39732 12798
rect 39340 12348 39396 12404
rect 40012 12572 40068 12628
rect 40460 12460 40516 12516
rect 40012 11452 40068 11508
rect 40236 12178 40292 12180
rect 40236 12126 40238 12178
rect 40238 12126 40290 12178
rect 40290 12126 40292 12178
rect 40236 12124 40292 12126
rect 40348 11394 40404 11396
rect 40348 11342 40350 11394
rect 40350 11342 40402 11394
rect 40402 11342 40404 11394
rect 40348 11340 40404 11342
rect 39228 9660 39284 9716
rect 39340 9100 39396 9156
rect 40012 9212 40068 9268
rect 39788 9100 39844 9156
rect 40348 9154 40404 9156
rect 40348 9102 40350 9154
rect 40350 9102 40402 9154
rect 40402 9102 40404 9154
rect 40348 9100 40404 9102
rect 40124 8876 40180 8932
rect 39452 8482 39508 8484
rect 39452 8430 39454 8482
rect 39454 8430 39506 8482
rect 39506 8430 39508 8482
rect 39452 8428 39508 8430
rect 39788 7756 39844 7812
rect 39116 6636 39172 6692
rect 39452 7474 39508 7476
rect 39452 7422 39454 7474
rect 39454 7422 39506 7474
rect 39506 7422 39508 7474
rect 39452 7420 39508 7422
rect 39228 6076 39284 6132
rect 39452 6636 39508 6692
rect 36764 5180 36820 5236
rect 36652 5068 36708 5124
rect 36988 4338 37044 4340
rect 36988 4286 36990 4338
rect 36990 4286 37042 4338
rect 37042 4286 37044 4338
rect 36988 4284 37044 4286
rect 36988 3666 37044 3668
rect 36988 3614 36990 3666
rect 36990 3614 37042 3666
rect 37042 3614 37044 3666
rect 36988 3612 37044 3614
rect 39340 5404 39396 5460
rect 39004 5292 39060 5348
rect 38892 5068 38948 5124
rect 37660 3948 37716 4004
rect 38332 3500 38388 3556
rect 39228 5180 39284 5236
rect 39004 3612 39060 3668
rect 39116 4732 39172 4788
rect 39228 4508 39284 4564
rect 40012 8204 40068 8260
rect 39900 7474 39956 7476
rect 39900 7422 39902 7474
rect 39902 7422 39954 7474
rect 39954 7422 39956 7474
rect 39900 7420 39956 7422
rect 41468 13634 41524 13636
rect 41468 13582 41470 13634
rect 41470 13582 41522 13634
rect 41522 13582 41524 13634
rect 41468 13580 41524 13582
rect 41468 13132 41524 13188
rect 41580 12684 41636 12740
rect 41468 12236 41524 12292
rect 41244 11676 41300 11732
rect 40572 10668 40628 10724
rect 41804 13468 41860 13524
rect 41916 12796 41972 12852
rect 41916 11676 41972 11732
rect 41132 9884 41188 9940
rect 41020 9042 41076 9044
rect 41020 8990 41022 9042
rect 41022 8990 41074 9042
rect 41074 8990 41076 9042
rect 41020 8988 41076 8990
rect 41468 10444 41524 10500
rect 41244 9100 41300 9156
rect 40908 8876 40964 8932
rect 41580 9884 41636 9940
rect 40796 8316 40852 8372
rect 41132 8258 41188 8260
rect 41132 8206 41134 8258
rect 41134 8206 41186 8258
rect 41186 8206 41188 8258
rect 41132 8204 41188 8206
rect 40460 7756 40516 7812
rect 41132 7644 41188 7700
rect 40236 7532 40292 7588
rect 40236 6972 40292 7028
rect 41468 7308 41524 7364
rect 40684 7196 40740 7252
rect 39788 5964 39844 6020
rect 39452 5122 39508 5124
rect 39452 5070 39454 5122
rect 39454 5070 39506 5122
rect 39506 5070 39508 5122
rect 39452 5068 39508 5070
rect 39564 5794 39620 5796
rect 39564 5742 39566 5794
rect 39566 5742 39618 5794
rect 39618 5742 39620 5794
rect 39564 5740 39620 5742
rect 40236 5292 40292 5348
rect 40348 5068 40404 5124
rect 41020 6578 41076 6580
rect 41020 6526 41022 6578
rect 41022 6526 41074 6578
rect 41074 6526 41076 6578
rect 41020 6524 41076 6526
rect 41356 6188 41412 6244
rect 40908 6076 40964 6132
rect 40572 5122 40628 5124
rect 40572 5070 40574 5122
rect 40574 5070 40626 5122
rect 40626 5070 40628 5122
rect 40572 5068 40628 5070
rect 40908 4450 40964 4452
rect 40908 4398 40910 4450
rect 40910 4398 40962 4450
rect 40962 4398 40964 4450
rect 40908 4396 40964 4398
rect 42028 8092 42084 8148
rect 41804 7980 41860 8036
rect 42252 16940 42308 16996
rect 43036 16994 43092 16996
rect 43036 16942 43038 16994
rect 43038 16942 43090 16994
rect 43090 16942 43092 16994
rect 43036 16940 43092 16942
rect 42252 16156 42308 16212
rect 43708 19234 43764 19236
rect 43708 19182 43710 19234
rect 43710 19182 43762 19234
rect 43762 19182 43764 19234
rect 43708 19180 43764 19182
rect 43820 19122 43876 19124
rect 43820 19070 43822 19122
rect 43822 19070 43874 19122
rect 43874 19070 43876 19122
rect 43820 19068 43876 19070
rect 44268 19122 44324 19124
rect 44268 19070 44270 19122
rect 44270 19070 44322 19122
rect 44322 19070 44324 19122
rect 44268 19068 44324 19070
rect 44268 18844 44324 18900
rect 44156 18562 44212 18564
rect 44156 18510 44158 18562
rect 44158 18510 44210 18562
rect 44210 18510 44212 18562
rect 44156 18508 44212 18510
rect 45276 22540 45332 22596
rect 45388 23100 45444 23156
rect 45164 22482 45220 22484
rect 45164 22430 45166 22482
rect 45166 22430 45218 22482
rect 45218 22430 45220 22482
rect 45164 22428 45220 22430
rect 44828 22370 44884 22372
rect 44828 22318 44830 22370
rect 44830 22318 44882 22370
rect 44882 22318 44884 22370
rect 44828 22316 44884 22318
rect 46284 22764 46340 22820
rect 46396 22988 46452 23044
rect 46284 22370 46340 22372
rect 46284 22318 46286 22370
rect 46286 22318 46338 22370
rect 46338 22318 46340 22370
rect 46284 22316 46340 22318
rect 45948 21868 46004 21924
rect 47180 25506 47236 25508
rect 47180 25454 47182 25506
rect 47182 25454 47234 25506
rect 47234 25454 47236 25506
rect 47180 25452 47236 25454
rect 47740 26290 47796 26292
rect 47740 26238 47742 26290
rect 47742 26238 47794 26290
rect 47794 26238 47796 26290
rect 47740 26236 47796 26238
rect 47404 25394 47460 25396
rect 47404 25342 47406 25394
rect 47406 25342 47458 25394
rect 47458 25342 47460 25394
rect 47404 25340 47460 25342
rect 49196 26962 49252 26964
rect 49196 26910 49198 26962
rect 49198 26910 49250 26962
rect 49250 26910 49252 26962
rect 49196 26908 49252 26910
rect 50316 27804 50372 27860
rect 51100 28642 51156 28644
rect 51100 28590 51102 28642
rect 51102 28590 51154 28642
rect 51154 28590 51156 28642
rect 51100 28588 51156 28590
rect 51772 28140 51828 28196
rect 51212 27858 51268 27860
rect 51212 27806 51214 27858
rect 51214 27806 51266 27858
rect 51266 27806 51268 27858
rect 51212 27804 51268 27806
rect 55580 28642 55636 28644
rect 55580 28590 55582 28642
rect 55582 28590 55634 28642
rect 55634 28590 55636 28642
rect 55580 28588 55636 28590
rect 57932 28252 57988 28308
rect 52780 28140 52836 28196
rect 52668 28082 52724 28084
rect 52668 28030 52670 28082
rect 52670 28030 52722 28082
rect 52722 28030 52724 28082
rect 52668 28028 52724 28030
rect 52108 27804 52164 27860
rect 50556 26682 50612 26684
rect 50556 26630 50558 26682
rect 50558 26630 50610 26682
rect 50610 26630 50612 26682
rect 50556 26628 50612 26630
rect 50660 26682 50716 26684
rect 50660 26630 50662 26682
rect 50662 26630 50714 26682
rect 50714 26630 50716 26682
rect 50660 26628 50716 26630
rect 50764 26682 50820 26684
rect 50764 26630 50766 26682
rect 50766 26630 50818 26682
rect 50818 26630 50820 26682
rect 50764 26628 50820 26630
rect 49420 25900 49476 25956
rect 47964 25564 48020 25620
rect 48636 25506 48692 25508
rect 48636 25454 48638 25506
rect 48638 25454 48690 25506
rect 48690 25454 48692 25506
rect 48636 25452 48692 25454
rect 49644 25676 49700 25732
rect 49756 26012 49812 26068
rect 48412 25340 48468 25396
rect 47740 24556 47796 24612
rect 46732 23660 46788 23716
rect 47516 23660 47572 23716
rect 49644 25340 49700 25396
rect 48860 25282 48916 25284
rect 48860 25230 48862 25282
rect 48862 25230 48914 25282
rect 48914 25230 48916 25282
rect 48860 25228 48916 25230
rect 50316 26402 50372 26404
rect 50316 26350 50318 26402
rect 50318 26350 50370 26402
rect 50370 26350 50372 26402
rect 50316 26348 50372 26350
rect 50092 26290 50148 26292
rect 50092 26238 50094 26290
rect 50094 26238 50146 26290
rect 50146 26238 50148 26290
rect 50092 26236 50148 26238
rect 50316 25676 50372 25732
rect 49756 25228 49812 25284
rect 49868 25452 49924 25508
rect 50204 25506 50260 25508
rect 50204 25454 50206 25506
rect 50206 25454 50258 25506
rect 50258 25454 50260 25506
rect 50204 25452 50260 25454
rect 51996 26402 52052 26404
rect 51996 26350 51998 26402
rect 51998 26350 52050 26402
rect 52050 26350 52052 26402
rect 51996 26348 52052 26350
rect 52444 26796 52500 26852
rect 53228 28140 53284 28196
rect 53116 27858 53172 27860
rect 53116 27806 53118 27858
rect 53118 27806 53170 27858
rect 53170 27806 53172 27858
rect 53116 27804 53172 27806
rect 53564 26908 53620 26964
rect 52892 26796 52948 26852
rect 54460 26962 54516 26964
rect 54460 26910 54462 26962
rect 54462 26910 54514 26962
rect 54514 26910 54516 26962
rect 54460 26908 54516 26910
rect 54124 26402 54180 26404
rect 54124 26350 54126 26402
rect 54126 26350 54178 26402
rect 54178 26350 54180 26402
rect 54124 26348 54180 26350
rect 53564 26236 53620 26292
rect 53116 26012 53172 26068
rect 51884 25676 51940 25732
rect 52780 25730 52836 25732
rect 52780 25678 52782 25730
rect 52782 25678 52834 25730
rect 52834 25678 52836 25730
rect 52780 25676 52836 25678
rect 52108 25564 52164 25620
rect 50652 25506 50708 25508
rect 50652 25454 50654 25506
rect 50654 25454 50706 25506
rect 50706 25454 50708 25506
rect 50652 25452 50708 25454
rect 51548 25452 51604 25508
rect 50428 25340 50484 25396
rect 49980 25228 50036 25284
rect 50540 25282 50596 25284
rect 50540 25230 50542 25282
rect 50542 25230 50594 25282
rect 50594 25230 50596 25282
rect 50540 25228 50596 25230
rect 49084 24722 49140 24724
rect 49084 24670 49086 24722
rect 49086 24670 49138 24722
rect 49138 24670 49140 24722
rect 49084 24668 49140 24670
rect 49980 24722 50036 24724
rect 49980 24670 49982 24722
rect 49982 24670 50034 24722
rect 50034 24670 50036 24722
rect 49980 24668 50036 24670
rect 47740 23548 47796 23604
rect 48076 23378 48132 23380
rect 48076 23326 48078 23378
rect 48078 23326 48130 23378
rect 48130 23326 48132 23378
rect 48076 23324 48132 23326
rect 47068 22764 47124 22820
rect 47516 22370 47572 22372
rect 47516 22318 47518 22370
rect 47518 22318 47570 22370
rect 47570 22318 47572 22370
rect 47516 22316 47572 22318
rect 47404 22092 47460 22148
rect 46620 21868 46676 21924
rect 47180 21644 47236 21700
rect 45052 20748 45108 20804
rect 45276 20636 45332 20692
rect 45948 20690 46004 20692
rect 45948 20638 45950 20690
rect 45950 20638 46002 20690
rect 46002 20638 46004 20690
rect 45948 20636 46004 20638
rect 46732 20690 46788 20692
rect 46732 20638 46734 20690
rect 46734 20638 46786 20690
rect 46786 20638 46788 20690
rect 46732 20636 46788 20638
rect 45612 19292 45668 19348
rect 45052 19068 45108 19124
rect 45388 19010 45444 19012
rect 45388 18958 45390 19010
rect 45390 18958 45442 19010
rect 45442 18958 45444 19010
rect 45388 18956 45444 18958
rect 45164 18844 45220 18900
rect 43820 18396 43876 18452
rect 44156 18226 44212 18228
rect 44156 18174 44158 18226
rect 44158 18174 44210 18226
rect 44210 18174 44212 18226
rect 44156 18172 44212 18174
rect 43148 15372 43204 15428
rect 42924 15314 42980 15316
rect 42924 15262 42926 15314
rect 42926 15262 42978 15314
rect 42978 15262 42980 15314
rect 42924 15260 42980 15262
rect 42364 13186 42420 13188
rect 42364 13134 42366 13186
rect 42366 13134 42418 13186
rect 42418 13134 42420 13186
rect 42364 13132 42420 13134
rect 43036 14418 43092 14420
rect 43036 14366 43038 14418
rect 43038 14366 43090 14418
rect 43090 14366 43092 14418
rect 43036 14364 43092 14366
rect 43036 13692 43092 13748
rect 43372 15986 43428 15988
rect 43372 15934 43374 15986
rect 43374 15934 43426 15986
rect 43426 15934 43428 15986
rect 43372 15932 43428 15934
rect 43484 15874 43540 15876
rect 43484 15822 43486 15874
rect 43486 15822 43538 15874
rect 43538 15822 43540 15874
rect 43484 15820 43540 15822
rect 45276 18450 45332 18452
rect 45276 18398 45278 18450
rect 45278 18398 45330 18450
rect 45330 18398 45332 18450
rect 45276 18396 45332 18398
rect 45276 17612 45332 17668
rect 44940 15986 44996 15988
rect 44940 15934 44942 15986
rect 44942 15934 44994 15986
rect 44994 15934 44996 15986
rect 44940 15932 44996 15934
rect 44156 15820 44212 15876
rect 43596 15260 43652 15316
rect 43260 13804 43316 13860
rect 43708 14530 43764 14532
rect 43708 14478 43710 14530
rect 43710 14478 43762 14530
rect 43762 14478 43764 14530
rect 43708 14476 43764 14478
rect 43596 13858 43652 13860
rect 43596 13806 43598 13858
rect 43598 13806 43650 13858
rect 43650 13806 43652 13858
rect 43596 13804 43652 13806
rect 44044 14364 44100 14420
rect 43932 13468 43988 13524
rect 44940 14530 44996 14532
rect 44940 14478 44942 14530
rect 44942 14478 44994 14530
rect 44994 14478 44996 14530
rect 44940 14476 44996 14478
rect 44380 14364 44436 14420
rect 42588 12738 42644 12740
rect 42588 12686 42590 12738
rect 42590 12686 42642 12738
rect 42642 12686 42644 12738
rect 42588 12684 42644 12686
rect 42700 12402 42756 12404
rect 42700 12350 42702 12402
rect 42702 12350 42754 12402
rect 42754 12350 42756 12402
rect 42700 12348 42756 12350
rect 43372 12402 43428 12404
rect 43372 12350 43374 12402
rect 43374 12350 43426 12402
rect 43426 12350 43428 12402
rect 43372 12348 43428 12350
rect 44380 12290 44436 12292
rect 44380 12238 44382 12290
rect 44382 12238 44434 12290
rect 44434 12238 44436 12290
rect 44380 12236 44436 12238
rect 44828 12850 44884 12852
rect 44828 12798 44830 12850
rect 44830 12798 44882 12850
rect 44882 12798 44884 12850
rect 44828 12796 44884 12798
rect 42924 12012 42980 12068
rect 43820 12012 43876 12068
rect 43708 11564 43764 11620
rect 42476 10722 42532 10724
rect 42476 10670 42478 10722
rect 42478 10670 42530 10722
rect 42530 10670 42532 10722
rect 42476 10668 42532 10670
rect 43372 10556 43428 10612
rect 43148 9938 43204 9940
rect 43148 9886 43150 9938
rect 43150 9886 43202 9938
rect 43202 9886 43204 9938
rect 43148 9884 43204 9886
rect 43036 9772 43092 9828
rect 43484 9826 43540 9828
rect 43484 9774 43486 9826
rect 43486 9774 43538 9826
rect 43538 9774 43540 9826
rect 43484 9772 43540 9774
rect 43932 11282 43988 11284
rect 43932 11230 43934 11282
rect 43934 11230 43986 11282
rect 43986 11230 43988 11282
rect 43932 11228 43988 11230
rect 44156 11394 44212 11396
rect 44156 11342 44158 11394
rect 44158 11342 44210 11394
rect 44210 11342 44212 11394
rect 44156 11340 44212 11342
rect 44716 11340 44772 11396
rect 44828 11228 44884 11284
rect 44156 9884 44212 9940
rect 43260 9042 43316 9044
rect 43260 8990 43262 9042
rect 43262 8990 43314 9042
rect 43314 8990 43316 9042
rect 43260 8988 43316 8990
rect 43484 9042 43540 9044
rect 43484 8990 43486 9042
rect 43486 8990 43538 9042
rect 43538 8990 43540 9042
rect 43484 8988 43540 8990
rect 43148 8428 43204 8484
rect 42924 8370 42980 8372
rect 42924 8318 42926 8370
rect 42926 8318 42978 8370
rect 42978 8318 42980 8370
rect 42924 8316 42980 8318
rect 42588 8204 42644 8260
rect 42700 7980 42756 8036
rect 42140 7308 42196 7364
rect 42252 7532 42308 7588
rect 42252 7196 42308 7252
rect 42140 6412 42196 6468
rect 41132 5740 41188 5796
rect 41132 4060 41188 4116
rect 41916 5852 41972 5908
rect 41468 5068 41524 5124
rect 42028 4226 42084 4228
rect 42028 4174 42030 4226
rect 42030 4174 42082 4226
rect 42082 4174 42084 4226
rect 42028 4172 42084 4174
rect 42700 6748 42756 6804
rect 42924 7196 42980 7252
rect 42924 6300 42980 6356
rect 42588 5964 42644 6020
rect 42476 5794 42532 5796
rect 42476 5742 42478 5794
rect 42478 5742 42530 5794
rect 42530 5742 42532 5794
rect 42476 5740 42532 5742
rect 43484 8258 43540 8260
rect 43484 8206 43486 8258
rect 43486 8206 43538 8258
rect 43538 8206 43540 8258
rect 43484 8204 43540 8206
rect 43372 7644 43428 7700
rect 43148 6636 43204 6692
rect 43708 8146 43764 8148
rect 43708 8094 43710 8146
rect 43710 8094 43762 8146
rect 43762 8094 43764 8146
rect 43708 8092 43764 8094
rect 43820 7980 43876 8036
rect 43932 7474 43988 7476
rect 43932 7422 43934 7474
rect 43934 7422 43986 7474
rect 43986 7422 43988 7474
rect 43932 7420 43988 7422
rect 43820 7308 43876 7364
rect 43596 5964 43652 6020
rect 43820 5628 43876 5684
rect 43932 6860 43988 6916
rect 45500 15986 45556 15988
rect 45500 15934 45502 15986
rect 45502 15934 45554 15986
rect 45554 15934 45556 15986
rect 45500 15932 45556 15934
rect 45388 13804 45444 13860
rect 45276 11228 45332 11284
rect 45500 10668 45556 10724
rect 44940 10610 44996 10612
rect 44940 10558 44942 10610
rect 44942 10558 44994 10610
rect 44994 10558 44996 10610
rect 44940 10556 44996 10558
rect 44828 8652 44884 8708
rect 44940 8988 44996 9044
rect 45276 8428 45332 8484
rect 45276 8258 45332 8260
rect 45276 8206 45278 8258
rect 45278 8206 45330 8258
rect 45330 8206 45332 8258
rect 45276 8204 45332 8206
rect 45052 8092 45108 8148
rect 44716 7980 44772 8036
rect 44380 7644 44436 7700
rect 46844 18956 46900 19012
rect 46620 18338 46676 18340
rect 46620 18286 46622 18338
rect 46622 18286 46674 18338
rect 46674 18286 46676 18338
rect 46620 18284 46676 18286
rect 46172 18172 46228 18228
rect 47852 22316 47908 22372
rect 47740 22092 47796 22148
rect 49868 23938 49924 23940
rect 49868 23886 49870 23938
rect 49870 23886 49922 23938
rect 49922 23886 49924 23938
rect 49868 23884 49924 23886
rect 49756 23660 49812 23716
rect 49980 23324 50036 23380
rect 49756 22092 49812 22148
rect 49644 21756 49700 21812
rect 47628 20188 47684 20244
rect 48524 20578 48580 20580
rect 48524 20526 48526 20578
rect 48526 20526 48578 20578
rect 48578 20526 48580 20578
rect 48524 20524 48580 20526
rect 48412 20076 48468 20132
rect 48524 20300 48580 20356
rect 47516 19458 47572 19460
rect 47516 19406 47518 19458
rect 47518 19406 47570 19458
rect 47570 19406 47572 19458
rect 47516 19404 47572 19406
rect 48748 20188 48804 20244
rect 49084 20076 49140 20132
rect 49308 20300 49364 20356
rect 48860 19404 48916 19460
rect 47404 19010 47460 19012
rect 47404 18958 47406 19010
rect 47406 18958 47458 19010
rect 47458 18958 47460 19010
rect 47404 18956 47460 18958
rect 47292 18620 47348 18676
rect 47404 18450 47460 18452
rect 47404 18398 47406 18450
rect 47406 18398 47458 18450
rect 47458 18398 47460 18450
rect 47404 18396 47460 18398
rect 46844 18172 46900 18228
rect 45948 16940 46004 16996
rect 47292 18284 47348 18340
rect 47740 18284 47796 18340
rect 47852 18396 47908 18452
rect 45724 15314 45780 15316
rect 45724 15262 45726 15314
rect 45726 15262 45778 15314
rect 45778 15262 45780 15314
rect 45724 15260 45780 15262
rect 46172 15260 46228 15316
rect 46844 16492 46900 16548
rect 46620 15932 46676 15988
rect 48524 18732 48580 18788
rect 48412 17612 48468 17668
rect 48524 17778 48580 17780
rect 48524 17726 48526 17778
rect 48526 17726 48578 17778
rect 48578 17726 48580 17778
rect 48524 17724 48580 17726
rect 47516 15314 47572 15316
rect 47516 15262 47518 15314
rect 47518 15262 47570 15314
rect 47570 15262 47572 15314
rect 47516 15260 47572 15262
rect 47852 15260 47908 15316
rect 47068 14700 47124 14756
rect 46508 14476 46564 14532
rect 45724 13692 45780 13748
rect 45836 11452 45892 11508
rect 45724 8316 45780 8372
rect 45724 8092 45780 8148
rect 45724 7698 45780 7700
rect 45724 7646 45726 7698
rect 45726 7646 45778 7698
rect 45778 7646 45780 7698
rect 45724 7644 45780 7646
rect 46060 10722 46116 10724
rect 46060 10670 46062 10722
rect 46062 10670 46114 10722
rect 46114 10670 46116 10722
rect 46060 10668 46116 10670
rect 46060 9154 46116 9156
rect 46060 9102 46062 9154
rect 46062 9102 46114 9154
rect 46114 9102 46116 9154
rect 46060 9100 46116 9102
rect 46396 11788 46452 11844
rect 47068 11788 47124 11844
rect 46732 11340 46788 11396
rect 47628 14924 47684 14980
rect 47516 14530 47572 14532
rect 47516 14478 47518 14530
rect 47518 14478 47570 14530
rect 47570 14478 47572 14530
rect 47516 14476 47572 14478
rect 47292 13746 47348 13748
rect 47292 13694 47294 13746
rect 47294 13694 47346 13746
rect 47346 13694 47348 13746
rect 47292 13692 47348 13694
rect 49084 18338 49140 18340
rect 49084 18286 49086 18338
rect 49086 18286 49138 18338
rect 49138 18286 49140 18338
rect 49084 18284 49140 18286
rect 49420 19180 49476 19236
rect 50556 25114 50612 25116
rect 50556 25062 50558 25114
rect 50558 25062 50610 25114
rect 50610 25062 50612 25114
rect 50556 25060 50612 25062
rect 50660 25114 50716 25116
rect 50660 25062 50662 25114
rect 50662 25062 50714 25114
rect 50714 25062 50716 25114
rect 50660 25060 50716 25062
rect 50764 25114 50820 25116
rect 50764 25062 50766 25114
rect 50766 25062 50818 25114
rect 50818 25062 50820 25114
rect 50764 25060 50820 25062
rect 50316 23772 50372 23828
rect 50988 23884 51044 23940
rect 51212 23826 51268 23828
rect 51212 23774 51214 23826
rect 51214 23774 51266 23826
rect 51266 23774 51268 23826
rect 51212 23772 51268 23774
rect 50556 23546 50612 23548
rect 50556 23494 50558 23546
rect 50558 23494 50610 23546
rect 50610 23494 50612 23546
rect 50556 23492 50612 23494
rect 50660 23546 50716 23548
rect 50660 23494 50662 23546
rect 50662 23494 50714 23546
rect 50714 23494 50716 23546
rect 50660 23492 50716 23494
rect 50764 23546 50820 23548
rect 50764 23494 50766 23546
rect 50766 23494 50818 23546
rect 50818 23494 50820 23546
rect 50764 23492 50820 23494
rect 50428 23154 50484 23156
rect 50428 23102 50430 23154
rect 50430 23102 50482 23154
rect 50482 23102 50484 23154
rect 50428 23100 50484 23102
rect 50540 22482 50596 22484
rect 50540 22430 50542 22482
rect 50542 22430 50594 22482
rect 50594 22430 50596 22482
rect 50540 22428 50596 22430
rect 50428 22316 50484 22372
rect 50204 21756 50260 21812
rect 51436 22316 51492 22372
rect 51100 22204 51156 22260
rect 50556 21978 50612 21980
rect 50556 21926 50558 21978
rect 50558 21926 50610 21978
rect 50610 21926 50612 21978
rect 50556 21924 50612 21926
rect 50660 21978 50716 21980
rect 50660 21926 50662 21978
rect 50662 21926 50714 21978
rect 50714 21926 50716 21978
rect 50660 21924 50716 21926
rect 50764 21978 50820 21980
rect 50764 21926 50766 21978
rect 50766 21926 50818 21978
rect 50818 21926 50820 21978
rect 50764 21924 50820 21926
rect 51324 21868 51380 21924
rect 52108 25282 52164 25284
rect 52108 25230 52110 25282
rect 52110 25230 52162 25282
rect 52162 25230 52164 25282
rect 52108 25228 52164 25230
rect 51996 24668 52052 24724
rect 52780 25394 52836 25396
rect 52780 25342 52782 25394
rect 52782 25342 52834 25394
rect 52834 25342 52836 25394
rect 52780 25340 52836 25342
rect 53788 26178 53844 26180
rect 53788 26126 53790 26178
rect 53790 26126 53842 26178
rect 53842 26126 53844 26178
rect 53788 26124 53844 26126
rect 53116 25340 53172 25396
rect 55580 27074 55636 27076
rect 55580 27022 55582 27074
rect 55582 27022 55634 27074
rect 55634 27022 55636 27074
rect 55580 27020 55636 27022
rect 57932 27580 57988 27636
rect 57484 26796 57540 26852
rect 54908 26460 54964 26516
rect 55580 26514 55636 26516
rect 55580 26462 55582 26514
rect 55582 26462 55634 26514
rect 55634 26462 55636 26514
rect 55580 26460 55636 26462
rect 53676 25228 53732 25284
rect 51884 23772 51940 23828
rect 51996 23714 52052 23716
rect 51996 23662 51998 23714
rect 51998 23662 52050 23714
rect 52050 23662 52052 23714
rect 51996 23660 52052 23662
rect 51660 22988 51716 23044
rect 51884 22370 51940 22372
rect 51884 22318 51886 22370
rect 51886 22318 51938 22370
rect 51938 22318 51940 22370
rect 51884 22316 51940 22318
rect 51548 22092 51604 22148
rect 52108 23042 52164 23044
rect 52108 22990 52110 23042
rect 52110 22990 52162 23042
rect 52162 22990 52164 23042
rect 52108 22988 52164 22990
rect 51884 22092 51940 22148
rect 50988 21810 51044 21812
rect 50988 21758 50990 21810
rect 50990 21758 51042 21810
rect 51042 21758 51044 21810
rect 50988 21756 51044 21758
rect 50316 20578 50372 20580
rect 50316 20526 50318 20578
rect 50318 20526 50370 20578
rect 50370 20526 50372 20578
rect 50316 20524 50372 20526
rect 51436 21756 51492 21812
rect 51996 21868 52052 21924
rect 51884 21698 51940 21700
rect 51884 21646 51886 21698
rect 51886 21646 51938 21698
rect 51938 21646 51940 21698
rect 51884 21644 51940 21646
rect 50988 20690 51044 20692
rect 50988 20638 50990 20690
rect 50990 20638 51042 20690
rect 51042 20638 51044 20690
rect 50988 20636 51044 20638
rect 50556 20410 50612 20412
rect 50556 20358 50558 20410
rect 50558 20358 50610 20410
rect 50610 20358 50612 20410
rect 50556 20356 50612 20358
rect 50660 20410 50716 20412
rect 50660 20358 50662 20410
rect 50662 20358 50714 20410
rect 50714 20358 50716 20410
rect 50660 20356 50716 20358
rect 50764 20410 50820 20412
rect 50764 20358 50766 20410
rect 50766 20358 50818 20410
rect 50818 20358 50820 20410
rect 50764 20356 50820 20358
rect 50092 19964 50148 20020
rect 51212 19852 51268 19908
rect 49532 18956 49588 19012
rect 51548 20018 51604 20020
rect 51548 19966 51550 20018
rect 51550 19966 51602 20018
rect 51602 19966 51604 20018
rect 51548 19964 51604 19966
rect 49644 18732 49700 18788
rect 49644 18508 49700 18564
rect 49308 18172 49364 18228
rect 50556 18842 50612 18844
rect 50556 18790 50558 18842
rect 50558 18790 50610 18842
rect 50610 18790 50612 18842
rect 50556 18788 50612 18790
rect 50660 18842 50716 18844
rect 50660 18790 50662 18842
rect 50662 18790 50714 18842
rect 50714 18790 50716 18842
rect 50660 18788 50716 18790
rect 50764 18842 50820 18844
rect 50764 18790 50766 18842
rect 50766 18790 50818 18842
rect 50818 18790 50820 18842
rect 50764 18788 50820 18790
rect 49084 17724 49140 17780
rect 50316 17554 50372 17556
rect 50316 17502 50318 17554
rect 50318 17502 50370 17554
rect 50370 17502 50372 17554
rect 50316 17500 50372 17502
rect 50428 18620 50484 18676
rect 50764 18620 50820 18676
rect 50540 18226 50596 18228
rect 50540 18174 50542 18226
rect 50542 18174 50594 18226
rect 50594 18174 50596 18226
rect 50540 18172 50596 18174
rect 50876 18284 50932 18340
rect 50988 18508 51044 18564
rect 50556 17274 50612 17276
rect 50556 17222 50558 17274
rect 50558 17222 50610 17274
rect 50610 17222 50612 17274
rect 50556 17220 50612 17222
rect 50660 17274 50716 17276
rect 50660 17222 50662 17274
rect 50662 17222 50714 17274
rect 50714 17222 50716 17274
rect 50660 17220 50716 17222
rect 50764 17274 50820 17276
rect 50764 17222 50766 17274
rect 50766 17222 50818 17274
rect 50818 17222 50820 17274
rect 50764 17220 50820 17222
rect 53452 23996 53508 24052
rect 53676 23996 53732 24052
rect 53452 23826 53508 23828
rect 53452 23774 53454 23826
rect 53454 23774 53506 23826
rect 53506 23774 53508 23826
rect 53452 23772 53508 23774
rect 55356 26290 55412 26292
rect 55356 26238 55358 26290
rect 55358 26238 55410 26290
rect 55410 26238 55412 26290
rect 55356 26236 55412 26238
rect 55020 25452 55076 25508
rect 55020 23884 55076 23940
rect 54796 23548 54852 23604
rect 53004 23324 53060 23380
rect 53900 23378 53956 23380
rect 53900 23326 53902 23378
rect 53902 23326 53954 23378
rect 53954 23326 53956 23378
rect 53900 23324 53956 23326
rect 53340 23100 53396 23156
rect 53004 22428 53060 22484
rect 52556 22204 52612 22260
rect 52668 21868 52724 21924
rect 53004 21756 53060 21812
rect 52444 19964 52500 20020
rect 52108 18396 52164 18452
rect 51212 17442 51268 17444
rect 51212 17390 51214 17442
rect 51214 17390 51266 17442
rect 51266 17390 51268 17442
rect 51212 17388 51268 17390
rect 52108 17388 52164 17444
rect 52220 17500 52276 17556
rect 51660 16770 51716 16772
rect 51660 16718 51662 16770
rect 51662 16718 51714 16770
rect 51714 16718 51716 16770
rect 51660 16716 51716 16718
rect 49084 16492 49140 16548
rect 48972 15986 49028 15988
rect 48972 15934 48974 15986
rect 48974 15934 49026 15986
rect 49026 15934 49028 15986
rect 48972 15932 49028 15934
rect 48748 15314 48804 15316
rect 48748 15262 48750 15314
rect 48750 15262 48802 15314
rect 48802 15262 48804 15314
rect 48748 15260 48804 15262
rect 50204 16268 50260 16324
rect 49980 16044 50036 16100
rect 49308 15932 49364 15988
rect 48524 14754 48580 14756
rect 48524 14702 48526 14754
rect 48526 14702 48578 14754
rect 48578 14702 48580 14754
rect 48524 14700 48580 14702
rect 48300 14476 48356 14532
rect 49196 15260 49252 15316
rect 48972 13746 49028 13748
rect 48972 13694 48974 13746
rect 48974 13694 49026 13746
rect 49026 13694 49028 13746
rect 48972 13692 49028 13694
rect 47852 12738 47908 12740
rect 47852 12686 47854 12738
rect 47854 12686 47906 12738
rect 47906 12686 47908 12738
rect 47852 12684 47908 12686
rect 48076 12572 48132 12628
rect 47628 12124 47684 12180
rect 47964 12178 48020 12180
rect 47964 12126 47966 12178
rect 47966 12126 48018 12178
rect 48018 12126 48020 12178
rect 47964 12124 48020 12126
rect 48188 12290 48244 12292
rect 48188 12238 48190 12290
rect 48190 12238 48242 12290
rect 48242 12238 48244 12290
rect 48188 12236 48244 12238
rect 48748 12572 48804 12628
rect 49084 12572 49140 12628
rect 49868 15932 49924 15988
rect 50764 16098 50820 16100
rect 50764 16046 50766 16098
rect 50766 16046 50818 16098
rect 50818 16046 50820 16098
rect 50764 16044 50820 16046
rect 50204 15484 50260 15540
rect 49420 15090 49476 15092
rect 49420 15038 49422 15090
rect 49422 15038 49474 15090
rect 49474 15038 49476 15090
rect 49420 15036 49476 15038
rect 49420 12850 49476 12852
rect 49420 12798 49422 12850
rect 49422 12798 49474 12850
rect 49474 12798 49476 12850
rect 49420 12796 49476 12798
rect 50988 15986 51044 15988
rect 50988 15934 50990 15986
rect 50990 15934 51042 15986
rect 51042 15934 51044 15986
rect 50988 15932 51044 15934
rect 50556 15706 50612 15708
rect 50556 15654 50558 15706
rect 50558 15654 50610 15706
rect 50610 15654 50612 15706
rect 50556 15652 50612 15654
rect 50660 15706 50716 15708
rect 50660 15654 50662 15706
rect 50662 15654 50714 15706
rect 50714 15654 50716 15706
rect 50660 15652 50716 15654
rect 50764 15706 50820 15708
rect 50764 15654 50766 15706
rect 50766 15654 50818 15706
rect 50818 15654 50820 15706
rect 50764 15652 50820 15654
rect 50540 15538 50596 15540
rect 50540 15486 50542 15538
rect 50542 15486 50594 15538
rect 50594 15486 50596 15538
rect 50540 15484 50596 15486
rect 50428 14924 50484 14980
rect 50764 15036 50820 15092
rect 50428 14530 50484 14532
rect 50428 14478 50430 14530
rect 50430 14478 50482 14530
rect 50482 14478 50484 14530
rect 50428 14476 50484 14478
rect 50556 14138 50612 14140
rect 50556 14086 50558 14138
rect 50558 14086 50610 14138
rect 50610 14086 50612 14138
rect 50556 14084 50612 14086
rect 50660 14138 50716 14140
rect 50660 14086 50662 14138
rect 50662 14086 50714 14138
rect 50714 14086 50716 14138
rect 50660 14084 50716 14086
rect 50764 14138 50820 14140
rect 50764 14086 50766 14138
rect 50766 14086 50818 14138
rect 50818 14086 50820 14138
rect 50764 14084 50820 14086
rect 50988 14812 51044 14868
rect 50764 13858 50820 13860
rect 50764 13806 50766 13858
rect 50766 13806 50818 13858
rect 50818 13806 50820 13858
rect 50764 13804 50820 13806
rect 50988 12962 51044 12964
rect 50988 12910 50990 12962
rect 50990 12910 51042 12962
rect 51042 12910 51044 12962
rect 50988 12908 51044 12910
rect 49868 12796 49924 12852
rect 52892 20636 52948 20692
rect 53452 22258 53508 22260
rect 53452 22206 53454 22258
rect 53454 22206 53506 22258
rect 53506 22206 53508 22258
rect 53452 22204 53508 22206
rect 55020 23266 55076 23268
rect 55020 23214 55022 23266
rect 55022 23214 55074 23266
rect 55074 23214 55076 23266
rect 55020 23212 55076 23214
rect 54684 23154 54740 23156
rect 54684 23102 54686 23154
rect 54686 23102 54738 23154
rect 54738 23102 54740 23154
rect 54684 23100 54740 23102
rect 55692 26124 55748 26180
rect 55580 25788 55636 25844
rect 55468 25452 55524 25508
rect 55356 24220 55412 24276
rect 55244 23660 55300 23716
rect 55580 24780 55636 24836
rect 55580 24108 55636 24164
rect 55692 23772 55748 23828
rect 55468 23436 55524 23492
rect 54348 22146 54404 22148
rect 54348 22094 54350 22146
rect 54350 22094 54402 22146
rect 54402 22094 54404 22146
rect 54348 22092 54404 22094
rect 54348 21810 54404 21812
rect 54348 21758 54350 21810
rect 54350 21758 54402 21810
rect 54402 21758 54404 21810
rect 54348 21756 54404 21758
rect 54796 21532 54852 21588
rect 54124 19964 54180 20020
rect 53788 19906 53844 19908
rect 53788 19854 53790 19906
rect 53790 19854 53842 19906
rect 53842 19854 53844 19906
rect 53788 19852 53844 19854
rect 55244 22316 55300 22372
rect 55468 22258 55524 22260
rect 55468 22206 55470 22258
rect 55470 22206 55522 22258
rect 55522 22206 55524 22258
rect 55468 22204 55524 22206
rect 55916 25452 55972 25508
rect 55804 23436 55860 23492
rect 56140 23996 56196 24052
rect 55804 23266 55860 23268
rect 55804 23214 55806 23266
rect 55806 23214 55858 23266
rect 55858 23214 55860 23266
rect 55804 23212 55860 23214
rect 55356 21980 55412 22036
rect 55804 21868 55860 21924
rect 56700 25900 56756 25956
rect 57372 25788 57428 25844
rect 57820 25340 57876 25396
rect 57932 24892 57988 24948
rect 56700 23884 56756 23940
rect 56812 23548 56868 23604
rect 55916 21698 55972 21700
rect 55916 21646 55918 21698
rect 55918 21646 55970 21698
rect 55970 21646 55972 21698
rect 55916 21644 55972 21646
rect 55020 20636 55076 20692
rect 55804 20690 55860 20692
rect 55804 20638 55806 20690
rect 55806 20638 55858 20690
rect 55858 20638 55860 20690
rect 55804 20636 55860 20638
rect 56812 21644 56868 21700
rect 56588 21586 56644 21588
rect 56588 21534 56590 21586
rect 56590 21534 56642 21586
rect 56642 21534 56644 21586
rect 56588 21532 56644 21534
rect 58044 24108 58100 24164
rect 57372 23660 57428 23716
rect 57148 22092 57204 22148
rect 58156 23548 58212 23604
rect 57260 22204 57316 22260
rect 56924 21868 56980 21924
rect 58156 21532 58212 21588
rect 57820 21308 57876 21364
rect 53564 19404 53620 19460
rect 53116 19180 53172 19236
rect 53340 18508 53396 18564
rect 53564 19122 53620 19124
rect 53564 19070 53566 19122
rect 53566 19070 53618 19122
rect 53618 19070 53620 19122
rect 53564 19068 53620 19070
rect 53564 18450 53620 18452
rect 53564 18398 53566 18450
rect 53566 18398 53618 18450
rect 53618 18398 53620 18450
rect 53564 18396 53620 18398
rect 53452 18338 53508 18340
rect 53452 18286 53454 18338
rect 53454 18286 53506 18338
rect 53506 18286 53508 18338
rect 53452 18284 53508 18286
rect 52444 17052 52500 17108
rect 53228 17052 53284 17108
rect 54460 19346 54516 19348
rect 54460 19294 54462 19346
rect 54462 19294 54514 19346
rect 54514 19294 54516 19346
rect 54460 19292 54516 19294
rect 53900 19234 53956 19236
rect 53900 19182 53902 19234
rect 53902 19182 53954 19234
rect 53954 19182 53956 19234
rect 53900 19180 53956 19182
rect 54124 18562 54180 18564
rect 54124 18510 54126 18562
rect 54126 18510 54178 18562
rect 54178 18510 54180 18562
rect 54124 18508 54180 18510
rect 55020 19122 55076 19124
rect 55020 19070 55022 19122
rect 55022 19070 55074 19122
rect 55074 19070 55076 19122
rect 55020 19068 55076 19070
rect 54796 18508 54852 18564
rect 55132 18396 55188 18452
rect 54572 18284 54628 18340
rect 55020 18338 55076 18340
rect 55020 18286 55022 18338
rect 55022 18286 55074 18338
rect 55074 18286 55076 18338
rect 55020 18284 55076 18286
rect 53340 16716 53396 16772
rect 53228 16268 53284 16324
rect 55804 19458 55860 19460
rect 55804 19406 55806 19458
rect 55806 19406 55858 19458
rect 55858 19406 55860 19458
rect 55804 19404 55860 19406
rect 56700 19292 56756 19348
rect 55580 18396 55636 18452
rect 51548 14588 51604 14644
rect 52892 14642 52948 14644
rect 52892 14590 52894 14642
rect 52894 14590 52946 14642
rect 52946 14590 52948 14642
rect 52892 14588 52948 14590
rect 51660 13468 51716 13524
rect 53004 13468 53060 13524
rect 49532 12684 49588 12740
rect 50556 12570 50612 12572
rect 50556 12518 50558 12570
rect 50558 12518 50610 12570
rect 50610 12518 50612 12570
rect 50556 12516 50612 12518
rect 50660 12570 50716 12572
rect 50660 12518 50662 12570
rect 50662 12518 50714 12570
rect 50714 12518 50716 12570
rect 50660 12516 50716 12518
rect 50764 12570 50820 12572
rect 50764 12518 50766 12570
rect 50766 12518 50818 12570
rect 50818 12518 50820 12570
rect 50764 12516 50820 12518
rect 51884 12402 51940 12404
rect 51884 12350 51886 12402
rect 51886 12350 51938 12402
rect 51938 12350 51940 12402
rect 51884 12348 51940 12350
rect 51660 12290 51716 12292
rect 51660 12238 51662 12290
rect 51662 12238 51714 12290
rect 51714 12238 51716 12290
rect 51660 12236 51716 12238
rect 53676 16268 53732 16324
rect 54572 16268 54628 16324
rect 55916 18284 55972 18340
rect 56140 17666 56196 17668
rect 56140 17614 56142 17666
rect 56142 17614 56194 17666
rect 56194 17614 56196 17666
rect 56140 17612 56196 17614
rect 55916 17052 55972 17108
rect 54348 15874 54404 15876
rect 54348 15822 54350 15874
rect 54350 15822 54402 15874
rect 54402 15822 54404 15874
rect 54348 15820 54404 15822
rect 55580 16940 55636 16996
rect 55468 16882 55524 16884
rect 55468 16830 55470 16882
rect 55470 16830 55522 16882
rect 55522 16830 55524 16882
rect 55468 16828 55524 16830
rect 55020 16268 55076 16324
rect 55132 16716 55188 16772
rect 53228 13804 53284 13860
rect 53676 13746 53732 13748
rect 53676 13694 53678 13746
rect 53678 13694 53730 13746
rect 53730 13694 53732 13746
rect 53676 13692 53732 13694
rect 53340 13522 53396 13524
rect 53340 13470 53342 13522
rect 53342 13470 53394 13522
rect 53394 13470 53396 13522
rect 53340 13468 53396 13470
rect 54236 13692 54292 13748
rect 54460 14252 54516 14308
rect 55804 16044 55860 16100
rect 55804 15820 55860 15876
rect 55132 15036 55188 15092
rect 57484 19292 57540 19348
rect 57484 17612 57540 17668
rect 57372 16994 57428 16996
rect 57372 16942 57374 16994
rect 57374 16942 57426 16994
rect 57426 16942 57428 16994
rect 57372 16940 57428 16942
rect 56812 16828 56868 16884
rect 56028 16044 56084 16100
rect 56476 16098 56532 16100
rect 56476 16046 56478 16098
rect 56478 16046 56530 16098
rect 56530 16046 56532 16098
rect 56476 16044 56532 16046
rect 56588 15820 56644 15876
rect 57036 15148 57092 15204
rect 55692 14252 55748 14308
rect 54796 13804 54852 13860
rect 54572 13746 54628 13748
rect 54572 13694 54574 13746
rect 54574 13694 54626 13746
rect 54626 13694 54628 13746
rect 54572 13692 54628 13694
rect 54348 13468 54404 13524
rect 54572 13468 54628 13524
rect 49644 12178 49700 12180
rect 49644 12126 49646 12178
rect 49646 12126 49698 12178
rect 49698 12126 49700 12178
rect 49644 12124 49700 12126
rect 50204 12178 50260 12180
rect 50204 12126 50206 12178
rect 50206 12126 50258 12178
rect 50258 12126 50260 12178
rect 50204 12124 50260 12126
rect 50876 12124 50932 12180
rect 49532 12066 49588 12068
rect 49532 12014 49534 12066
rect 49534 12014 49586 12066
rect 49586 12014 49588 12066
rect 49532 12012 49588 12014
rect 47628 11394 47684 11396
rect 47628 11342 47630 11394
rect 47630 11342 47682 11394
rect 47682 11342 47684 11394
rect 47628 11340 47684 11342
rect 47852 10834 47908 10836
rect 47852 10782 47854 10834
rect 47854 10782 47906 10834
rect 47906 10782 47908 10834
rect 47852 10780 47908 10782
rect 47404 10668 47460 10724
rect 50428 12066 50484 12068
rect 50428 12014 50430 12066
rect 50430 12014 50482 12066
rect 50482 12014 50484 12066
rect 50428 12012 50484 12014
rect 49868 11340 49924 11396
rect 49868 10780 49924 10836
rect 47852 10610 47908 10612
rect 47852 10558 47854 10610
rect 47854 10558 47906 10610
rect 47906 10558 47908 10610
rect 47852 10556 47908 10558
rect 46396 8652 46452 8708
rect 46844 8428 46900 8484
rect 47180 9154 47236 9156
rect 47180 9102 47182 9154
rect 47182 9102 47234 9154
rect 47234 9102 47236 9154
rect 47180 9100 47236 9102
rect 47404 8764 47460 8820
rect 47292 8258 47348 8260
rect 47292 8206 47294 8258
rect 47294 8206 47346 8258
rect 47346 8206 47348 8258
rect 47292 8204 47348 8206
rect 44940 6802 44996 6804
rect 44940 6750 44942 6802
rect 44942 6750 44994 6802
rect 44994 6750 44996 6802
rect 44940 6748 44996 6750
rect 44156 6636 44212 6692
rect 44044 5906 44100 5908
rect 44044 5854 44046 5906
rect 44046 5854 44098 5906
rect 44098 5854 44100 5906
rect 44044 5852 44100 5854
rect 44604 5964 44660 6020
rect 45388 6636 45444 6692
rect 43708 5516 43764 5572
rect 43484 5292 43540 5348
rect 43932 5404 43988 5460
rect 43820 5068 43876 5124
rect 43260 4898 43316 4900
rect 43260 4846 43262 4898
rect 43262 4846 43314 4898
rect 43314 4846 43316 4898
rect 43260 4844 43316 4846
rect 43036 4732 43092 4788
rect 42924 4508 42980 4564
rect 42700 4338 42756 4340
rect 42700 4286 42702 4338
rect 42702 4286 42754 4338
rect 42754 4286 42756 4338
rect 42700 4284 42756 4286
rect 42140 3724 42196 3780
rect 41804 3666 41860 3668
rect 41804 3614 41806 3666
rect 41806 3614 41858 3666
rect 41858 3614 41860 3666
rect 41804 3612 41860 3614
rect 39004 3388 39060 3444
rect 43148 4338 43204 4340
rect 43148 4286 43150 4338
rect 43150 4286 43202 4338
rect 43202 4286 43204 4338
rect 43148 4284 43204 4286
rect 43372 4172 43428 4228
rect 43820 4844 43876 4900
rect 43148 3612 43204 3668
rect 42700 3164 42756 3220
rect 39676 2604 39732 2660
rect 43596 4508 43652 4564
rect 43932 3724 43988 3780
rect 43484 3276 43540 3332
rect 44380 5628 44436 5684
rect 44156 5180 44212 5236
rect 44268 5010 44324 5012
rect 44268 4958 44270 5010
rect 44270 4958 44322 5010
rect 44322 4958 44324 5010
rect 44268 4956 44324 4958
rect 44828 5122 44884 5124
rect 44828 5070 44830 5122
rect 44830 5070 44882 5122
rect 44882 5070 44884 5122
rect 44828 5068 44884 5070
rect 44940 3948 44996 4004
rect 44492 3836 44548 3892
rect 45612 6466 45668 6468
rect 45612 6414 45614 6466
rect 45614 6414 45666 6466
rect 45666 6414 45668 6466
rect 45612 6412 45668 6414
rect 45164 5794 45220 5796
rect 45164 5742 45166 5794
rect 45166 5742 45218 5794
rect 45218 5742 45220 5794
rect 45164 5740 45220 5742
rect 45164 5292 45220 5348
rect 45612 4956 45668 5012
rect 45388 4732 45444 4788
rect 45612 4338 45668 4340
rect 45612 4286 45614 4338
rect 45614 4286 45666 4338
rect 45666 4286 45668 4338
rect 45612 4284 45668 4286
rect 45164 3554 45220 3556
rect 45164 3502 45166 3554
rect 45166 3502 45218 3554
rect 45218 3502 45220 3554
rect 45164 3500 45220 3502
rect 46060 7308 46116 7364
rect 46844 7474 46900 7476
rect 46844 7422 46846 7474
rect 46846 7422 46898 7474
rect 46898 7422 46900 7474
rect 46844 7420 46900 7422
rect 46060 6412 46116 6468
rect 47068 7644 47124 7700
rect 47292 6690 47348 6692
rect 47292 6638 47294 6690
rect 47294 6638 47346 6690
rect 47346 6638 47348 6690
rect 47292 6636 47348 6638
rect 47068 6412 47124 6468
rect 50764 11394 50820 11396
rect 50764 11342 50766 11394
rect 50766 11342 50818 11394
rect 50818 11342 50820 11394
rect 50764 11340 50820 11342
rect 51548 12178 51604 12180
rect 51548 12126 51550 12178
rect 51550 12126 51602 12178
rect 51602 12126 51604 12178
rect 51548 12124 51604 12126
rect 50556 11002 50612 11004
rect 50556 10950 50558 11002
rect 50558 10950 50610 11002
rect 50610 10950 50612 11002
rect 50556 10948 50612 10950
rect 50660 11002 50716 11004
rect 50660 10950 50662 11002
rect 50662 10950 50714 11002
rect 50714 10950 50716 11002
rect 50660 10948 50716 10950
rect 50764 11002 50820 11004
rect 50764 10950 50766 11002
rect 50766 10950 50818 11002
rect 50818 10950 50820 11002
rect 50764 10948 50820 10950
rect 50092 9772 50148 9828
rect 51212 9884 51268 9940
rect 50556 9434 50612 9436
rect 50556 9382 50558 9434
rect 50558 9382 50610 9434
rect 50610 9382 50612 9434
rect 50556 9380 50612 9382
rect 50660 9434 50716 9436
rect 50660 9382 50662 9434
rect 50662 9382 50714 9434
rect 50714 9382 50716 9434
rect 50660 9380 50716 9382
rect 50764 9434 50820 9436
rect 50764 9382 50766 9434
rect 50766 9382 50818 9434
rect 50818 9382 50820 9434
rect 50764 9380 50820 9382
rect 48188 9212 48244 9268
rect 48860 9266 48916 9268
rect 48860 9214 48862 9266
rect 48862 9214 48914 9266
rect 48914 9214 48916 9266
rect 48860 9212 48916 9214
rect 48300 8316 48356 8372
rect 48300 7868 48356 7924
rect 47628 7698 47684 7700
rect 47628 7646 47630 7698
rect 47630 7646 47682 7698
rect 47682 7646 47684 7698
rect 47628 7644 47684 7646
rect 49644 8876 49700 8932
rect 48972 8818 49028 8820
rect 48972 8766 48974 8818
rect 48974 8766 49026 8818
rect 49026 8766 49028 8818
rect 48972 8764 49028 8766
rect 49196 8540 49252 8596
rect 49532 8428 49588 8484
rect 48860 7868 48916 7924
rect 48972 7980 49028 8036
rect 48748 7644 48804 7700
rect 48076 7420 48132 7476
rect 49756 8428 49812 8484
rect 49980 8764 50036 8820
rect 50428 8818 50484 8820
rect 50428 8766 50430 8818
rect 50430 8766 50482 8818
rect 50482 8766 50484 8818
rect 50428 8764 50484 8766
rect 49756 7980 49812 8036
rect 49980 8540 50036 8596
rect 49420 7474 49476 7476
rect 49420 7422 49422 7474
rect 49422 7422 49474 7474
rect 49474 7422 49476 7474
rect 49420 7420 49476 7422
rect 50876 8258 50932 8260
rect 50876 8206 50878 8258
rect 50878 8206 50930 8258
rect 50930 8206 50932 8258
rect 50876 8204 50932 8206
rect 50556 7866 50612 7868
rect 50556 7814 50558 7866
rect 50558 7814 50610 7866
rect 50610 7814 50612 7866
rect 50556 7812 50612 7814
rect 50660 7866 50716 7868
rect 50660 7814 50662 7866
rect 50662 7814 50714 7866
rect 50714 7814 50716 7866
rect 50660 7812 50716 7814
rect 50764 7866 50820 7868
rect 50764 7814 50766 7866
rect 50766 7814 50818 7866
rect 50818 7814 50820 7866
rect 50764 7812 50820 7814
rect 50764 7644 50820 7700
rect 50204 7586 50260 7588
rect 50204 7534 50206 7586
rect 50206 7534 50258 7586
rect 50258 7534 50260 7586
rect 50204 7532 50260 7534
rect 47964 7308 48020 7364
rect 47516 6524 47572 6580
rect 49308 6636 49364 6692
rect 46396 5740 46452 5796
rect 45948 5628 46004 5684
rect 45836 5516 45892 5572
rect 45948 5068 46004 5124
rect 46620 5628 46676 5684
rect 46396 4450 46452 4452
rect 46396 4398 46398 4450
rect 46398 4398 46450 4450
rect 46450 4398 46452 4450
rect 46396 4396 46452 4398
rect 46284 4284 46340 4340
rect 45948 4172 46004 4228
rect 46844 3724 46900 3780
rect 48972 5906 49028 5908
rect 48972 5854 48974 5906
rect 48974 5854 49026 5906
rect 49026 5854 49028 5906
rect 48972 5852 49028 5854
rect 48860 5682 48916 5684
rect 48860 5630 48862 5682
rect 48862 5630 48914 5682
rect 48914 5630 48916 5682
rect 48860 5628 48916 5630
rect 47964 5292 48020 5348
rect 47180 5122 47236 5124
rect 47180 5070 47182 5122
rect 47182 5070 47234 5122
rect 47234 5070 47236 5122
rect 47180 5068 47236 5070
rect 50428 6636 50484 6692
rect 49532 6578 49588 6580
rect 49532 6526 49534 6578
rect 49534 6526 49586 6578
rect 49586 6526 49588 6578
rect 49532 6524 49588 6526
rect 49084 5292 49140 5348
rect 48076 5068 48132 5124
rect 48412 5068 48468 5124
rect 47404 4396 47460 4452
rect 47292 3948 47348 4004
rect 47292 3500 47348 3556
rect 45948 3276 46004 3332
rect 48188 4226 48244 4228
rect 48188 4174 48190 4226
rect 48190 4174 48242 4226
rect 48242 4174 48244 4226
rect 48188 4172 48244 4174
rect 47740 3836 47796 3892
rect 47628 3612 47684 3668
rect 48188 3554 48244 3556
rect 48188 3502 48190 3554
rect 48190 3502 48242 3554
rect 48242 3502 48244 3554
rect 48188 3500 48244 3502
rect 50316 6578 50372 6580
rect 50316 6526 50318 6578
rect 50318 6526 50370 6578
rect 50370 6526 50372 6578
rect 50316 6524 50372 6526
rect 49868 6076 49924 6132
rect 49868 5740 49924 5796
rect 49980 5628 50036 5684
rect 50204 5852 50260 5908
rect 49980 5122 50036 5124
rect 49980 5070 49982 5122
rect 49982 5070 50034 5122
rect 50034 5070 50036 5122
rect 49980 5068 50036 5070
rect 49308 3666 49364 3668
rect 49308 3614 49310 3666
rect 49310 3614 49362 3666
rect 49362 3614 49364 3666
rect 49308 3612 49364 3614
rect 48860 3500 48916 3556
rect 48748 3388 48804 3444
rect 46508 2604 46564 2660
rect 43932 2492 43988 2548
rect 50540 6412 50596 6468
rect 52668 12124 52724 12180
rect 53228 12012 53284 12068
rect 53564 12348 53620 12404
rect 53788 12066 53844 12068
rect 53788 12014 53790 12066
rect 53790 12014 53842 12066
rect 53842 12014 53844 12066
rect 53788 12012 53844 12014
rect 56476 14252 56532 14308
rect 55356 13858 55412 13860
rect 55356 13806 55358 13858
rect 55358 13806 55410 13858
rect 55410 13806 55412 13858
rect 55356 13804 55412 13806
rect 55132 13468 55188 13524
rect 54908 12290 54964 12292
rect 54908 12238 54910 12290
rect 54910 12238 54962 12290
rect 54962 12238 54964 12290
rect 54908 12236 54964 12238
rect 52892 10668 52948 10724
rect 51100 7644 51156 7700
rect 51884 9212 51940 9268
rect 51548 9042 51604 9044
rect 51548 8990 51550 9042
rect 51550 8990 51602 9042
rect 51602 8990 51604 9042
rect 51548 8988 51604 8990
rect 51436 8316 51492 8372
rect 51772 8204 51828 8260
rect 51436 7420 51492 7476
rect 50876 6860 50932 6916
rect 51436 6690 51492 6692
rect 51436 6638 51438 6690
rect 51438 6638 51490 6690
rect 51490 6638 51492 6690
rect 51436 6636 51492 6638
rect 50556 6298 50612 6300
rect 50556 6246 50558 6298
rect 50558 6246 50610 6298
rect 50610 6246 50612 6298
rect 50556 6244 50612 6246
rect 50660 6298 50716 6300
rect 50660 6246 50662 6298
rect 50662 6246 50714 6298
rect 50714 6246 50716 6298
rect 50660 6244 50716 6246
rect 50764 6298 50820 6300
rect 50764 6246 50766 6298
rect 50766 6246 50818 6298
rect 50818 6246 50820 6298
rect 50764 6244 50820 6246
rect 52556 9772 52612 9828
rect 52108 9154 52164 9156
rect 52108 9102 52110 9154
rect 52110 9102 52162 9154
rect 52162 9102 52164 9154
rect 52108 9100 52164 9102
rect 53228 10834 53284 10836
rect 53228 10782 53230 10834
rect 53230 10782 53282 10834
rect 53282 10782 53284 10834
rect 53228 10780 53284 10782
rect 54012 10780 54068 10836
rect 53788 10722 53844 10724
rect 53788 10670 53790 10722
rect 53790 10670 53842 10722
rect 53842 10670 53844 10722
rect 53788 10668 53844 10670
rect 53452 10386 53508 10388
rect 53452 10334 53454 10386
rect 53454 10334 53506 10386
rect 53506 10334 53508 10386
rect 53452 10332 53508 10334
rect 54012 10332 54068 10388
rect 53676 9884 53732 9940
rect 53116 9826 53172 9828
rect 53116 9774 53118 9826
rect 53118 9774 53170 9826
rect 53170 9774 53172 9826
rect 53116 9772 53172 9774
rect 52892 9042 52948 9044
rect 52892 8990 52894 9042
rect 52894 8990 52946 9042
rect 52946 8990 52948 9042
rect 52892 8988 52948 8990
rect 52556 8652 52612 8708
rect 52556 8370 52612 8372
rect 52556 8318 52558 8370
rect 52558 8318 52610 8370
rect 52610 8318 52612 8370
rect 52556 8316 52612 8318
rect 52444 7532 52500 7588
rect 53004 8092 53060 8148
rect 52892 7980 52948 8036
rect 53004 6860 53060 6916
rect 54684 9884 54740 9940
rect 53228 9212 53284 9268
rect 54124 9826 54180 9828
rect 54124 9774 54126 9826
rect 54126 9774 54178 9826
rect 54178 9774 54180 9826
rect 54124 9772 54180 9774
rect 53900 9212 53956 9268
rect 53340 8652 53396 8708
rect 53228 7980 53284 8036
rect 53452 8316 53508 8372
rect 54012 8316 54068 8372
rect 53900 8258 53956 8260
rect 53900 8206 53902 8258
rect 53902 8206 53954 8258
rect 53954 8206 53956 8258
rect 53900 8204 53956 8206
rect 54236 8146 54292 8148
rect 54236 8094 54238 8146
rect 54238 8094 54290 8146
rect 54290 8094 54292 8146
rect 54236 8092 54292 8094
rect 53788 8034 53844 8036
rect 53788 7982 53790 8034
rect 53790 7982 53842 8034
rect 53842 7982 53844 8034
rect 53788 7980 53844 7982
rect 53452 6860 53508 6916
rect 52220 6076 52276 6132
rect 51324 5906 51380 5908
rect 51324 5854 51326 5906
rect 51326 5854 51378 5906
rect 51378 5854 51380 5906
rect 51324 5852 51380 5854
rect 50316 5628 50372 5684
rect 52668 6130 52724 6132
rect 52668 6078 52670 6130
rect 52670 6078 52722 6130
rect 52722 6078 52724 6130
rect 52668 6076 52724 6078
rect 52108 5628 52164 5684
rect 50556 4730 50612 4732
rect 50556 4678 50558 4730
rect 50558 4678 50610 4730
rect 50610 4678 50612 4730
rect 50556 4676 50612 4678
rect 50660 4730 50716 4732
rect 50660 4678 50662 4730
rect 50662 4678 50714 4730
rect 50714 4678 50716 4730
rect 50660 4676 50716 4678
rect 50764 4730 50820 4732
rect 50764 4678 50766 4730
rect 50766 4678 50818 4730
rect 50818 4678 50820 4730
rect 50764 4676 50820 4678
rect 50556 3162 50612 3164
rect 50556 3110 50558 3162
rect 50558 3110 50610 3162
rect 50610 3110 50612 3162
rect 50556 3108 50612 3110
rect 50660 3162 50716 3164
rect 50660 3110 50662 3162
rect 50662 3110 50714 3162
rect 50714 3110 50716 3162
rect 50660 3108 50716 3110
rect 50764 3162 50820 3164
rect 50764 3110 50766 3162
rect 50766 3110 50818 3162
rect 50818 3110 50820 3162
rect 50764 3108 50820 3110
<< metal3 >>
rect 19826 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20110 56476
rect 50546 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50830 56476
rect 31602 56252 31612 56308
rect 31668 56252 33180 56308
rect 33236 56252 33246 56308
rect 36306 56252 36316 56308
rect 36372 56252 41020 56308
rect 41076 56252 43036 56308
rect 43092 56252 43102 56308
rect 36978 56140 36988 56196
rect 37044 56140 41580 56196
rect 41636 56140 43708 56196
rect 43764 56140 43774 56196
rect 39218 56028 39228 56084
rect 39284 56028 42588 56084
rect 42644 56028 42654 56084
rect 27570 55916 27580 55972
rect 27636 55916 28588 55972
rect 28644 55916 28654 55972
rect 34290 55916 34300 55972
rect 34356 55916 36204 55972
rect 36260 55916 36270 55972
rect 38546 55916 38556 55972
rect 38612 55916 42140 55972
rect 42196 55916 42206 55972
rect 4466 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4750 55692
rect 35186 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35470 55692
rect 28914 55468 28924 55524
rect 28980 55468 28990 55524
rect 40226 55468 40236 55524
rect 40292 55468 40302 55524
rect 28924 55412 28980 55468
rect 40236 55412 40292 55468
rect 27458 55356 27468 55412
rect 27524 55356 28140 55412
rect 28196 55356 28206 55412
rect 28476 55356 28980 55412
rect 32274 55356 32284 55412
rect 32340 55356 33516 55412
rect 33572 55356 33582 55412
rect 33730 55356 33740 55412
rect 33796 55356 35532 55412
rect 35588 55356 35598 55412
rect 36082 55356 36092 55412
rect 36148 55356 37212 55412
rect 37268 55356 37278 55412
rect 40236 55356 42028 55412
rect 42084 55356 42094 55412
rect 28476 55300 28532 55356
rect 28466 55244 28476 55300
rect 28532 55244 28542 55300
rect 34962 55244 34972 55300
rect 35028 55244 39228 55300
rect 39284 55244 39294 55300
rect 41010 55244 41020 55300
rect 41076 55244 42476 55300
rect 42532 55244 42542 55300
rect 35746 55132 35756 55188
rect 35812 55132 36428 55188
rect 36484 55132 36494 55188
rect 39442 55132 39452 55188
rect 39508 55132 41580 55188
rect 41636 55132 41646 55188
rect 35970 55020 35980 55076
rect 36036 55020 36764 55076
rect 36820 55020 36830 55076
rect 38770 55020 38780 55076
rect 38836 55020 40460 55076
rect 40516 55020 40526 55076
rect 19826 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20110 54908
rect 50546 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50830 54908
rect 29138 54796 29148 54852
rect 29204 54796 29708 54852
rect 29764 54796 29774 54852
rect 32946 54684 32956 54740
rect 33012 54684 34188 54740
rect 34244 54684 34254 54740
rect 28466 54572 28476 54628
rect 28532 54572 29148 54628
rect 29204 54572 29214 54628
rect 31714 54572 31724 54628
rect 31780 54572 32396 54628
rect 32452 54572 32462 54628
rect 37650 54572 37660 54628
rect 37716 54572 40124 54628
rect 40180 54572 41020 54628
rect 41076 54572 41086 54628
rect 32498 54460 32508 54516
rect 32564 54460 33180 54516
rect 33236 54460 33246 54516
rect 31266 54348 31276 54404
rect 31332 54348 31836 54404
rect 31892 54348 31902 54404
rect 32610 54348 32620 54404
rect 32676 54348 35644 54404
rect 35700 54348 35710 54404
rect 35532 54124 36876 54180
rect 36932 54124 39788 54180
rect 39844 54124 39854 54180
rect 4466 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4750 54124
rect 35186 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35470 54124
rect 35532 53956 35588 54124
rect 37426 54012 37436 54068
rect 37492 54012 41356 54068
rect 41412 54012 41422 54068
rect 30594 53900 30604 53956
rect 30660 53900 30670 53956
rect 32386 53900 32396 53956
rect 32452 53900 35420 53956
rect 35476 53900 35588 53956
rect 36194 53900 36204 53956
rect 36260 53900 40236 53956
rect 40292 53900 40302 53956
rect 30604 53732 30660 53900
rect 36754 53788 36764 53844
rect 36820 53788 40012 53844
rect 40068 53788 40078 53844
rect 28802 53676 28812 53732
rect 28868 53676 31612 53732
rect 31668 53676 31678 53732
rect 23874 53564 23884 53620
rect 23940 53564 25228 53620
rect 25284 53564 25294 53620
rect 31154 53564 31164 53620
rect 31220 53564 32396 53620
rect 32452 53564 32462 53620
rect 37090 53564 37100 53620
rect 37156 53564 39340 53620
rect 39396 53564 39564 53620
rect 39620 53564 39630 53620
rect 42578 53564 42588 53620
rect 42644 53564 47852 53620
rect 47908 53564 47918 53620
rect 24322 53452 24332 53508
rect 24388 53452 25676 53508
rect 25732 53452 25742 53508
rect 29922 53452 29932 53508
rect 29988 53452 30268 53508
rect 30324 53452 30334 53508
rect 38546 53452 38556 53508
rect 38612 53396 38668 53508
rect 39890 53452 39900 53508
rect 39956 53452 42700 53508
rect 42756 53452 44380 53508
rect 44436 53452 44446 53508
rect 38612 53340 42364 53396
rect 42420 53340 42430 53396
rect 43362 53340 43372 53396
rect 43428 53340 48188 53396
rect 48244 53340 48254 53396
rect 19826 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20110 53340
rect 50546 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50830 53340
rect 27682 53116 27692 53172
rect 27748 53116 29148 53172
rect 29204 53116 29988 53172
rect 41010 53116 41020 53172
rect 41076 53116 44492 53172
rect 44548 53116 46284 53172
rect 46340 53116 46350 53172
rect 29932 53060 29988 53116
rect 14914 53004 14924 53060
rect 14980 53004 15596 53060
rect 15652 53004 16156 53060
rect 16212 53004 16222 53060
rect 21522 53004 21532 53060
rect 21588 53004 22652 53060
rect 22708 53004 23660 53060
rect 23716 53004 23726 53060
rect 29922 53004 29932 53060
rect 29988 53004 29998 53060
rect 31602 53004 31612 53060
rect 31668 53004 32844 53060
rect 32900 53004 33404 53060
rect 33460 53004 33470 53060
rect 36082 53004 36092 53060
rect 36148 53004 36988 53060
rect 37044 53004 37054 53060
rect 37986 53004 37996 53060
rect 38052 53004 38780 53060
rect 38836 53004 41132 53060
rect 41188 53004 41198 53060
rect 12450 52892 12460 52948
rect 12516 52892 13468 52948
rect 13524 52892 13534 52948
rect 19618 52892 19628 52948
rect 19684 52892 20636 52948
rect 20692 52892 20702 52948
rect 32386 52892 32396 52948
rect 32452 52892 33852 52948
rect 33908 52892 33918 52948
rect 38882 52892 38892 52948
rect 38948 52892 39340 52948
rect 39396 52892 39406 52948
rect 40114 52892 40124 52948
rect 40180 52892 40908 52948
rect 40964 52892 40974 52948
rect 42802 52892 42812 52948
rect 42868 52892 43372 52948
rect 43428 52892 43438 52948
rect 18386 52780 18396 52836
rect 18452 52780 19180 52836
rect 19236 52780 20748 52836
rect 20804 52780 21308 52836
rect 21364 52780 21374 52836
rect 23426 52780 23436 52836
rect 23492 52780 23996 52836
rect 24052 52780 24556 52836
rect 24612 52780 25340 52836
rect 25396 52780 25406 52836
rect 29698 52780 29708 52836
rect 29764 52780 30492 52836
rect 30548 52780 31388 52836
rect 31444 52780 35308 52836
rect 35364 52780 36316 52836
rect 36372 52780 36382 52836
rect 41346 52780 41356 52836
rect 41412 52780 42028 52836
rect 42084 52780 42094 52836
rect 42914 52780 42924 52836
rect 42980 52780 43596 52836
rect 43652 52780 43662 52836
rect 39442 52668 39452 52724
rect 39508 52668 39788 52724
rect 39844 52668 39854 52724
rect 22306 52556 22316 52612
rect 22372 52556 23884 52612
rect 23940 52556 23950 52612
rect 4466 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4750 52556
rect 35186 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35470 52556
rect 20066 52444 20076 52500
rect 20132 52444 21308 52500
rect 21364 52444 21374 52500
rect 30594 52444 30604 52500
rect 30660 52444 31164 52500
rect 31220 52444 31230 52500
rect 10994 52332 11004 52388
rect 11060 52332 12460 52388
rect 12516 52332 12526 52388
rect 17266 52332 17276 52388
rect 17332 52332 18060 52388
rect 18116 52332 20188 52388
rect 24658 52332 24668 52388
rect 24724 52332 26012 52388
rect 26068 52332 26460 52388
rect 26516 52332 26526 52388
rect 33730 52332 33740 52388
rect 33796 52332 35532 52388
rect 35588 52332 35980 52388
rect 36036 52332 36046 52388
rect 41122 52332 41132 52388
rect 41188 52332 42700 52388
rect 42756 52332 42766 52388
rect 43586 52332 43596 52388
rect 43652 52332 49084 52388
rect 49140 52332 49644 52388
rect 49700 52332 50876 52388
rect 50932 52332 50942 52388
rect 12562 52220 12572 52276
rect 12628 52220 13244 52276
rect 13300 52220 14588 52276
rect 14644 52220 15260 52276
rect 15316 52220 15326 52276
rect 16594 52220 16604 52276
rect 16660 52220 17948 52276
rect 18004 52220 18620 52276
rect 18676 52220 19740 52276
rect 19796 52220 19806 52276
rect 11106 52108 11116 52164
rect 11172 52108 11788 52164
rect 11844 52108 11854 52164
rect 12338 52108 12348 52164
rect 12404 52108 15148 52164
rect 15204 52108 16380 52164
rect 16436 52108 16446 52164
rect 20132 52108 20188 52332
rect 21970 52220 21980 52276
rect 22036 52220 22046 52276
rect 29698 52220 29708 52276
rect 29764 52220 30268 52276
rect 30324 52220 32060 52276
rect 32116 52220 35196 52276
rect 35252 52220 35262 52276
rect 40002 52220 40012 52276
rect 40068 52220 41356 52276
rect 41412 52220 41422 52276
rect 48178 52220 48188 52276
rect 48244 52220 50316 52276
rect 50372 52220 50382 52276
rect 21980 52164 22036 52220
rect 20244 52108 20254 52164
rect 21420 52108 24556 52164
rect 24612 52108 24622 52164
rect 26338 52108 26348 52164
rect 26404 52108 27076 52164
rect 29922 52108 29932 52164
rect 29988 52108 31052 52164
rect 31108 52108 31118 52164
rect 32386 52108 32396 52164
rect 32452 52108 33964 52164
rect 34020 52108 34030 52164
rect 37426 52108 37436 52164
rect 37492 52108 39452 52164
rect 39508 52108 39518 52164
rect 41122 52108 41132 52164
rect 41188 52108 42588 52164
rect 42644 52108 42654 52164
rect 48402 52108 48412 52164
rect 48468 52108 49308 52164
rect 49364 52108 50988 52164
rect 51044 52108 51054 52164
rect 21420 52052 21476 52108
rect 27020 52052 27076 52108
rect 12226 51996 12236 52052
rect 12292 51996 12796 52052
rect 12852 51996 12862 52052
rect 21186 51996 21196 52052
rect 21252 51996 21476 52052
rect 21634 51996 21644 52052
rect 21700 51996 21980 52052
rect 22036 51996 22046 52052
rect 27010 51996 27020 52052
rect 27076 51996 27086 52052
rect 30146 51996 30156 52052
rect 30212 51996 30492 52052
rect 30548 51996 30558 52052
rect 36530 51996 36540 52052
rect 36596 51996 39564 52052
rect 39620 51996 39630 52052
rect 43922 51996 43932 52052
rect 43988 51996 44940 52052
rect 44996 51996 45006 52052
rect 46946 51996 46956 52052
rect 47012 51996 48636 52052
rect 48692 51996 48702 52052
rect 49186 51996 49196 52052
rect 49252 51996 51548 52052
rect 51604 51996 51614 52052
rect 21522 51884 21532 51940
rect 21588 51884 22540 51940
rect 22596 51884 23100 51940
rect 23156 51884 23166 51940
rect 31714 51884 31724 51940
rect 31780 51884 32172 51940
rect 32228 51884 32238 51940
rect 36418 51884 36428 51940
rect 36484 51884 37324 51940
rect 37380 51884 37390 51940
rect 37538 51884 37548 51940
rect 37604 51884 37884 51940
rect 37940 51884 38444 51940
rect 38500 51884 38510 51940
rect 21532 51772 21868 51828
rect 21924 51772 21934 51828
rect 34626 51772 34636 51828
rect 34692 51772 36316 51828
rect 36372 51772 38668 51828
rect 38724 51772 43260 51828
rect 43316 51772 43326 51828
rect 19826 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20110 51772
rect 21532 51716 21588 51772
rect 50546 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50830 51772
rect 21522 51660 21532 51716
rect 21588 51660 21598 51716
rect 20626 51548 20636 51604
rect 20692 51548 21644 51604
rect 21700 51548 21710 51604
rect 31892 51548 33180 51604
rect 33236 51548 36316 51604
rect 36372 51548 36876 51604
rect 36932 51548 36942 51604
rect 38882 51548 38892 51604
rect 38948 51548 39116 51604
rect 39172 51548 39900 51604
rect 39956 51548 39966 51604
rect 41244 51548 42588 51604
rect 42644 51548 42654 51604
rect 42914 51548 42924 51604
rect 42980 51548 43820 51604
rect 43876 51548 45500 51604
rect 45556 51548 45566 51604
rect 31892 51492 31948 51548
rect 41244 51492 41300 51548
rect 8306 51436 8316 51492
rect 8372 51436 10332 51492
rect 10388 51436 10836 51492
rect 15474 51436 15484 51492
rect 15540 51436 20076 51492
rect 20132 51436 20860 51492
rect 20916 51436 20926 51492
rect 24770 51436 24780 51492
rect 24836 51436 25564 51492
rect 25620 51436 27356 51492
rect 27412 51436 27422 51492
rect 31602 51436 31612 51492
rect 31668 51436 31948 51492
rect 32498 51436 32508 51492
rect 32564 51436 34076 51492
rect 34132 51436 35532 51492
rect 35588 51436 35598 51492
rect 36418 51436 36428 51492
rect 36484 51436 37436 51492
rect 37492 51436 38332 51492
rect 38388 51436 41300 51492
rect 42466 51436 42476 51492
rect 42532 51436 44156 51492
rect 44212 51436 44828 51492
rect 44884 51436 44894 51492
rect 45602 51436 45612 51492
rect 45668 51436 46956 51492
rect 47012 51436 47022 51492
rect 51874 51436 51884 51492
rect 51940 51436 52668 51492
rect 52724 51436 52734 51492
rect 10780 51380 10836 51436
rect 10770 51324 10780 51380
rect 10836 51324 10846 51380
rect 11218 51324 11228 51380
rect 11284 51324 12348 51380
rect 12404 51324 14476 51380
rect 14532 51324 14542 51380
rect 33058 51324 33068 51380
rect 33124 51324 34860 51380
rect 34916 51324 34926 51380
rect 37314 51324 37324 51380
rect 37380 51324 37772 51380
rect 37828 51324 37838 51380
rect 41794 51324 41804 51380
rect 41860 51324 43036 51380
rect 43092 51324 43484 51380
rect 43540 51324 43550 51380
rect 46498 51324 46508 51380
rect 46564 51324 47852 51380
rect 47908 51324 48748 51380
rect 48804 51324 48814 51380
rect 30594 51212 30604 51268
rect 30660 51212 34524 51268
rect 34580 51212 34590 51268
rect 38546 51212 38556 51268
rect 38612 51212 39788 51268
rect 39844 51212 41132 51268
rect 41188 51212 41916 51268
rect 41972 51212 41982 51268
rect 45378 51212 45388 51268
rect 45444 51212 46620 51268
rect 46676 51212 46686 51268
rect 49074 51212 49084 51268
rect 49140 51212 49532 51268
rect 49588 51212 51100 51268
rect 51156 51212 51166 51268
rect 12450 51100 12460 51156
rect 12516 51100 13692 51156
rect 13748 51100 13758 51156
rect 25554 51100 25564 51156
rect 25620 51100 27020 51156
rect 27076 51100 27086 51156
rect 37762 51100 37772 51156
rect 37828 51100 38780 51156
rect 38836 51100 41244 51156
rect 41300 51100 41310 51156
rect 47170 51100 47180 51156
rect 47236 51100 49756 51156
rect 49812 51100 50092 51156
rect 50148 51100 50158 51156
rect 5954 50988 5964 51044
rect 6020 50988 10108 51044
rect 10164 50988 15484 51044
rect 15540 50988 15550 51044
rect 48066 50988 48076 51044
rect 48132 50988 49084 51044
rect 49140 50988 49150 51044
rect 4466 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4750 50988
rect 35186 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35470 50988
rect 34402 50764 34412 50820
rect 34468 50764 35420 50820
rect 35476 50764 37548 50820
rect 37604 50764 37614 50820
rect 42466 50764 42476 50820
rect 42532 50764 43484 50820
rect 43540 50764 43550 50820
rect 8754 50652 8764 50708
rect 8820 50652 12012 50708
rect 12068 50652 12078 50708
rect 21186 50652 21196 50708
rect 21252 50652 26012 50708
rect 26068 50652 26078 50708
rect 32834 50652 32844 50708
rect 32900 50652 34692 50708
rect 50082 50652 50092 50708
rect 50148 50652 51884 50708
rect 51940 50652 51950 50708
rect 34636 50596 34692 50652
rect 7186 50540 7196 50596
rect 7252 50540 9212 50596
rect 9268 50540 9278 50596
rect 13906 50540 13916 50596
rect 13972 50540 16828 50596
rect 16884 50540 16894 50596
rect 20132 50540 20300 50596
rect 20356 50540 22652 50596
rect 22708 50540 25676 50596
rect 25732 50540 25742 50596
rect 31042 50540 31052 50596
rect 31108 50540 34188 50596
rect 34244 50540 34254 50596
rect 34626 50540 34636 50596
rect 34692 50540 35756 50596
rect 35812 50540 35822 50596
rect 37762 50540 37772 50596
rect 37828 50540 38332 50596
rect 38388 50540 40348 50596
rect 40404 50540 40414 50596
rect 46050 50540 46060 50596
rect 46116 50540 46620 50596
rect 46676 50540 49532 50596
rect 49588 50540 49598 50596
rect 0 50484 800 50512
rect 20132 50484 20188 50540
rect 0 50428 1708 50484
rect 1764 50428 2940 50484
rect 2996 50428 3006 50484
rect 15698 50428 15708 50484
rect 15764 50428 18508 50484
rect 18564 50428 20188 50484
rect 24546 50428 24556 50484
rect 24612 50428 25788 50484
rect 25844 50428 25854 50484
rect 31154 50428 31164 50484
rect 31220 50428 31724 50484
rect 31780 50428 32956 50484
rect 33012 50428 33022 50484
rect 34850 50428 34860 50484
rect 34916 50428 35532 50484
rect 35588 50428 35598 50484
rect 45602 50428 45612 50484
rect 45668 50428 46956 50484
rect 47012 50428 48748 50484
rect 48804 50428 48814 50484
rect 0 50400 800 50428
rect 2034 50316 2044 50372
rect 2100 50316 4844 50372
rect 4900 50316 5628 50372
rect 5684 50316 5694 50372
rect 44482 50316 44492 50372
rect 44548 50316 45164 50372
rect 45220 50316 47404 50372
rect 47460 50316 47470 50372
rect 49970 50316 49980 50372
rect 50036 50316 51436 50372
rect 51492 50316 51502 50372
rect 52434 50316 52444 50372
rect 52500 50316 52780 50372
rect 52836 50316 53228 50372
rect 53284 50316 53294 50372
rect 19826 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20110 50204
rect 50546 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50830 50204
rect 14130 50092 14140 50148
rect 14196 50092 14700 50148
rect 14756 50092 14766 50148
rect 26450 50092 26460 50148
rect 26516 50092 27916 50148
rect 27972 50092 27982 50148
rect 43810 50092 43820 50148
rect 43876 50092 44940 50148
rect 44996 50092 45006 50148
rect 30370 49980 30380 50036
rect 30436 49980 30828 50036
rect 30884 49980 30894 50036
rect 32162 49980 32172 50036
rect 32228 49980 34748 50036
rect 34804 49980 34814 50036
rect 42578 49980 42588 50036
rect 42644 49980 43932 50036
rect 43988 49980 44492 50036
rect 44548 49980 44558 50036
rect 50418 49980 50428 50036
rect 50484 49980 52108 50036
rect 52164 49980 52780 50036
rect 52836 49980 53676 50036
rect 53732 49980 53742 50036
rect 7634 49868 7644 49924
rect 7700 49868 8204 49924
rect 8260 49868 8270 49924
rect 11666 49868 11676 49924
rect 11732 49868 13580 49924
rect 13636 49868 14028 49924
rect 14084 49868 14094 49924
rect 20178 49868 20188 49924
rect 20244 49868 21532 49924
rect 21588 49868 22652 49924
rect 22708 49868 22718 49924
rect 35634 49868 35644 49924
rect 35700 49868 36204 49924
rect 36260 49868 36876 49924
rect 36932 49868 37772 49924
rect 37828 49868 37838 49924
rect 38098 49868 38108 49924
rect 38164 49868 38892 49924
rect 38948 49868 38958 49924
rect 19282 49756 19292 49812
rect 19348 49756 20524 49812
rect 20580 49756 20590 49812
rect 25778 49756 25788 49812
rect 25844 49756 27244 49812
rect 27300 49756 27310 49812
rect 29698 49756 29708 49812
rect 29764 49756 30380 49812
rect 30436 49756 30446 49812
rect 39218 49756 39228 49812
rect 39284 49756 39564 49812
rect 39620 49756 43260 49812
rect 43316 49756 43326 49812
rect 2790 49644 2828 49700
rect 2884 49644 2894 49700
rect 6850 49644 6860 49700
rect 6916 49644 7756 49700
rect 7812 49644 7822 49700
rect 12898 49644 12908 49700
rect 12964 49644 15148 49700
rect 15204 49644 15214 49700
rect 25890 49644 25900 49700
rect 25956 49644 26796 49700
rect 26852 49644 26862 49700
rect 28578 49644 28588 49700
rect 28644 49644 29932 49700
rect 29988 49644 29998 49700
rect 31490 49644 31500 49700
rect 31556 49644 37324 49700
rect 37380 49644 38332 49700
rect 38388 49644 38398 49700
rect 35970 49420 35980 49476
rect 36036 49420 36764 49476
rect 36820 49420 37212 49476
rect 37268 49420 37660 49476
rect 37716 49420 37726 49476
rect 49522 49420 49532 49476
rect 49588 49420 50316 49476
rect 50372 49420 52332 49476
rect 52388 49420 52398 49476
rect 4466 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4750 49420
rect 35186 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35470 49420
rect 1698 49308 1708 49364
rect 1764 49308 3948 49364
rect 4004 49308 4014 49364
rect 29362 49308 29372 49364
rect 29428 49308 31500 49364
rect 31556 49308 31566 49364
rect 2482 49196 2492 49252
rect 2548 49196 3388 49252
rect 3444 49196 3454 49252
rect 29810 49196 29820 49252
rect 29876 49196 29886 49252
rect 35858 49196 35868 49252
rect 35924 49196 39452 49252
rect 39508 49196 39518 49252
rect 49522 49196 49532 49252
rect 49588 49196 50428 49252
rect 50484 49196 50494 49252
rect 53106 49196 53116 49252
rect 53172 49196 53900 49252
rect 53956 49196 53966 49252
rect 3378 49084 3388 49140
rect 3444 49084 3948 49140
rect 4004 49084 4844 49140
rect 4900 49084 4910 49140
rect 6962 49084 6972 49140
rect 7028 49084 14700 49140
rect 14756 49084 15372 49140
rect 15428 49084 15438 49140
rect 19394 49084 19404 49140
rect 19460 49084 21980 49140
rect 22036 49084 22988 49140
rect 23044 49084 23054 49140
rect 2370 48972 2380 49028
rect 2436 48972 2446 49028
rect 3266 48972 3276 49028
rect 3332 48972 4172 49028
rect 4228 48972 4238 49028
rect 4722 48972 4732 49028
rect 4788 48972 6300 49028
rect 6356 48972 6636 49028
rect 6692 48972 6702 49028
rect 2380 48916 2436 48972
rect 3836 48916 3892 48972
rect 6972 48916 7028 49084
rect 29820 49028 29876 49196
rect 32834 49084 32844 49140
rect 32900 49084 34524 49140
rect 34580 49084 37548 49140
rect 37604 49084 37614 49140
rect 38546 49084 38556 49140
rect 38612 49084 39116 49140
rect 39172 49084 39182 49140
rect 15092 48972 16380 49028
rect 16436 48972 16446 49028
rect 21858 48972 21868 49028
rect 21924 48972 22876 49028
rect 22932 48972 22942 49028
rect 27906 48972 27916 49028
rect 27972 48972 28588 49028
rect 28644 48972 28654 49028
rect 29820 48972 31052 49028
rect 31108 48972 32172 49028
rect 32228 48972 32238 49028
rect 35186 48972 35196 49028
rect 35252 48972 36092 49028
rect 36148 48972 36988 49028
rect 37044 48972 37054 49028
rect 38322 48972 38332 49028
rect 38388 48972 41468 49028
rect 41524 48972 41534 49028
rect 48626 48972 48636 49028
rect 48692 48972 50428 49028
rect 50484 48972 51100 49028
rect 51156 48972 51166 49028
rect 15092 48916 15148 48972
rect 2380 48860 3500 48916
rect 3556 48860 3566 48916
rect 3798 48860 3836 48916
rect 3892 48860 3902 48916
rect 4946 48860 4956 48916
rect 5012 48860 5796 48916
rect 6066 48860 6076 48916
rect 6132 48860 7028 48916
rect 8306 48860 8316 48916
rect 8372 48860 9212 48916
rect 9268 48860 9278 48916
rect 14690 48860 14700 48916
rect 14756 48860 15148 48916
rect 17042 48860 17052 48916
rect 17108 48860 19516 48916
rect 19572 48860 20188 48916
rect 20244 48860 20254 48916
rect 27234 48860 27244 48916
rect 27300 48860 28476 48916
rect 28532 48860 28542 48916
rect 29586 48860 29596 48916
rect 29652 48860 31164 48916
rect 31220 48860 33180 48916
rect 33236 48860 36764 48916
rect 36820 48860 36830 48916
rect 37762 48860 37772 48916
rect 37828 48860 37996 48916
rect 38052 48860 38062 48916
rect 44034 48860 44044 48916
rect 44100 48860 46844 48916
rect 46900 48860 46910 48916
rect 5740 48804 5796 48860
rect 6636 48804 6692 48860
rect 1474 48748 1484 48804
rect 1540 48748 2044 48804
rect 2100 48748 2110 48804
rect 5730 48748 5740 48804
rect 5796 48748 5806 48804
rect 6626 48748 6636 48804
rect 6692 48748 6702 48804
rect 10546 48748 10556 48804
rect 10612 48748 12348 48804
rect 12404 48748 12414 48804
rect 18722 48748 18732 48804
rect 18788 48748 19404 48804
rect 19460 48748 20524 48804
rect 20580 48748 20590 48804
rect 20962 48748 20972 48804
rect 21028 48748 21420 48804
rect 21476 48748 21486 48804
rect 24882 48748 24892 48804
rect 24948 48748 26012 48804
rect 26068 48748 26852 48804
rect 33282 48748 33292 48804
rect 33348 48748 33516 48804
rect 33572 48748 34300 48804
rect 34356 48748 34366 48804
rect 36082 48748 36092 48804
rect 36148 48748 37436 48804
rect 37492 48748 37502 48804
rect 44930 48748 44940 48804
rect 44996 48748 52444 48804
rect 52500 48748 52510 48804
rect 20524 48692 20580 48748
rect 3602 48636 3612 48692
rect 3668 48636 3948 48692
rect 4004 48636 4014 48692
rect 11778 48636 11788 48692
rect 11844 48636 13692 48692
rect 13748 48636 13758 48692
rect 20524 48636 22204 48692
rect 22260 48636 22270 48692
rect 19826 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20110 48636
rect 26796 48580 26852 48748
rect 35410 48636 35420 48692
rect 35476 48636 35756 48692
rect 35812 48636 35822 48692
rect 40114 48636 40124 48692
rect 40180 48636 40684 48692
rect 40740 48636 41692 48692
rect 41748 48636 41758 48692
rect 45266 48636 45276 48692
rect 45332 48636 46172 48692
rect 46228 48636 46844 48692
rect 46900 48636 47292 48692
rect 47348 48636 47358 48692
rect 1698 48524 1708 48580
rect 1764 48524 4508 48580
rect 4564 48524 4574 48580
rect 26786 48524 26796 48580
rect 26852 48524 26862 48580
rect 37090 48524 37100 48580
rect 37156 48524 39452 48580
rect 39508 48524 39518 48580
rect 43698 48524 43708 48580
rect 43764 48524 47852 48580
rect 47908 48524 47918 48580
rect 2706 48412 2716 48468
rect 2772 48412 3388 48468
rect 3444 48412 3454 48468
rect 3948 48356 4004 48524
rect 50428 48468 50484 48748
rect 50546 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50830 48636
rect 11554 48412 11564 48468
rect 11620 48412 11900 48468
rect 11956 48412 11966 48468
rect 15922 48412 15932 48468
rect 15988 48412 17388 48468
rect 17444 48412 17454 48468
rect 19282 48412 19292 48468
rect 19348 48412 19852 48468
rect 19908 48412 19918 48468
rect 20850 48412 20860 48468
rect 20916 48412 21196 48468
rect 21252 48412 21262 48468
rect 22642 48412 22652 48468
rect 22708 48412 25676 48468
rect 25732 48412 25742 48468
rect 50428 48412 50764 48468
rect 50820 48412 50830 48468
rect 51426 48412 51436 48468
rect 51492 48412 53116 48468
rect 53172 48412 53182 48468
rect 2146 48300 2156 48356
rect 2212 48300 3276 48356
rect 3332 48300 3342 48356
rect 3836 48300 4004 48356
rect 9090 48300 9100 48356
rect 9156 48300 9884 48356
rect 9940 48300 13916 48356
rect 13972 48300 13982 48356
rect 32386 48300 32396 48356
rect 32452 48300 35644 48356
rect 35700 48300 35710 48356
rect 50978 48300 50988 48356
rect 51044 48300 51324 48356
rect 51380 48300 51390 48356
rect 2594 48188 2604 48244
rect 2660 48188 3052 48244
rect 3108 48188 3118 48244
rect 3378 48076 3388 48132
rect 3444 48076 3500 48132
rect 3556 48076 3566 48132
rect 3836 47908 3892 48300
rect 8978 48188 8988 48244
rect 9044 48188 11900 48244
rect 11956 48188 12796 48244
rect 12852 48188 12862 48244
rect 19618 48188 19628 48244
rect 19684 48188 19964 48244
rect 20020 48188 20030 48244
rect 25666 48188 25676 48244
rect 25732 48188 26236 48244
rect 26292 48188 26302 48244
rect 32834 48188 32844 48244
rect 32900 48188 33740 48244
rect 33796 48188 33806 48244
rect 34850 48188 34860 48244
rect 34916 48188 37100 48244
rect 37156 48188 37166 48244
rect 38882 48188 38892 48244
rect 38948 48188 42028 48244
rect 42084 48188 42094 48244
rect 4050 48076 4060 48132
rect 4116 48076 4508 48132
rect 4564 48076 5628 48132
rect 5684 48076 5694 48132
rect 5954 48076 5964 48132
rect 6020 48076 7532 48132
rect 7588 48076 7598 48132
rect 31154 48076 31164 48132
rect 31220 48076 33068 48132
rect 33124 48076 33134 48132
rect 44034 48076 44044 48132
rect 44100 48076 44268 48132
rect 44324 48076 44334 48132
rect 25778 47964 25788 48020
rect 25844 47964 27020 48020
rect 27076 47964 27086 48020
rect 30146 47964 30156 48020
rect 30212 47964 33292 48020
rect 33348 47964 33516 48020
rect 33572 47964 33582 48020
rect 3836 47852 4228 47908
rect 4172 47572 4228 47852
rect 4466 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4750 47852
rect 35186 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35470 47852
rect 13906 47740 13916 47796
rect 13972 47740 16380 47796
rect 16436 47740 16446 47796
rect 14130 47628 14140 47684
rect 14196 47628 17724 47684
rect 17780 47628 17790 47684
rect 25890 47628 25900 47684
rect 25956 47628 26236 47684
rect 26292 47628 26302 47684
rect 31714 47628 31724 47684
rect 31780 47628 32284 47684
rect 32340 47628 32350 47684
rect 3164 47516 3724 47572
rect 3780 47516 3790 47572
rect 4162 47516 4172 47572
rect 4228 47516 4238 47572
rect 7522 47516 7532 47572
rect 7588 47516 7980 47572
rect 8036 47516 8046 47572
rect 8306 47516 8316 47572
rect 8372 47516 9772 47572
rect 9828 47516 9838 47572
rect 14578 47516 14588 47572
rect 14644 47516 15932 47572
rect 15988 47516 15998 47572
rect 16370 47516 16380 47572
rect 16436 47516 18508 47572
rect 18564 47516 18574 47572
rect 30594 47516 30604 47572
rect 30660 47516 31388 47572
rect 31444 47516 34636 47572
rect 34692 47516 34702 47572
rect 49298 47516 49308 47572
rect 49364 47516 51212 47572
rect 51268 47516 51278 47572
rect 52770 47516 52780 47572
rect 52836 47516 54124 47572
rect 54180 47516 54190 47572
rect 3164 47460 3220 47516
rect 2482 47404 2492 47460
rect 2548 47404 3052 47460
rect 3108 47404 3220 47460
rect 3378 47404 3388 47460
rect 3444 47404 5068 47460
rect 5124 47404 5134 47460
rect 17266 47404 17276 47460
rect 17332 47404 21196 47460
rect 21252 47404 21262 47460
rect 38098 47404 38108 47460
rect 38164 47404 38556 47460
rect 38612 47404 38622 47460
rect 39442 47404 39452 47460
rect 39508 47404 43148 47460
rect 43204 47404 43214 47460
rect 3266 47292 3276 47348
rect 3332 47292 6300 47348
rect 6356 47292 6366 47348
rect 8866 47292 8876 47348
rect 8932 47292 9548 47348
rect 9604 47292 10332 47348
rect 10388 47292 10398 47348
rect 14690 47292 14700 47348
rect 14756 47292 17500 47348
rect 17556 47292 17948 47348
rect 18004 47292 18014 47348
rect 18610 47292 18620 47348
rect 18676 47292 19292 47348
rect 19348 47292 19852 47348
rect 19908 47292 19918 47348
rect 20290 47292 20300 47348
rect 20356 47292 21532 47348
rect 21588 47292 21598 47348
rect 41468 47292 43820 47348
rect 43876 47292 43886 47348
rect 2034 47180 2044 47236
rect 2100 47180 9212 47236
rect 9268 47180 9278 47236
rect 15026 47180 15036 47236
rect 15092 47180 15596 47236
rect 15652 47180 15662 47236
rect 19058 47180 19068 47236
rect 19124 47180 19740 47236
rect 19796 47180 19806 47236
rect 21970 47180 21980 47236
rect 22036 47180 22652 47236
rect 22708 47180 22718 47236
rect 31266 47180 31276 47236
rect 31332 47180 31612 47236
rect 31668 47180 31678 47236
rect 41468 47124 41524 47292
rect 3042 47068 3052 47124
rect 3108 47068 3836 47124
rect 3892 47068 5404 47124
rect 5460 47068 5470 47124
rect 31378 47068 31388 47124
rect 31444 47068 35084 47124
rect 35140 47068 35150 47124
rect 35522 47068 35532 47124
rect 35588 47068 39564 47124
rect 39620 47068 41468 47124
rect 41524 47068 41534 47124
rect 19826 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20110 47068
rect 50546 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50830 47068
rect 32050 46956 32060 47012
rect 32116 46956 33292 47012
rect 33348 46956 33358 47012
rect 40114 46956 40124 47012
rect 40180 46956 41132 47012
rect 41188 46956 47964 47012
rect 48020 46956 48030 47012
rect 47964 46900 48020 46956
rect 19404 46844 20300 46900
rect 20356 46844 20366 46900
rect 22530 46844 22540 46900
rect 22596 46844 22606 46900
rect 40226 46844 40236 46900
rect 40292 46844 42140 46900
rect 42196 46844 42206 46900
rect 43922 46844 43932 46900
rect 43988 46844 46060 46900
rect 46116 46844 46126 46900
rect 47964 46844 51436 46900
rect 51492 46844 51502 46900
rect 53218 46844 53228 46900
rect 53284 46844 54124 46900
rect 54180 46844 54190 46900
rect 19404 46788 19460 46844
rect 1810 46732 1820 46788
rect 1876 46732 2268 46788
rect 2324 46732 2334 46788
rect 16706 46732 16716 46788
rect 16772 46732 19404 46788
rect 19460 46732 19470 46788
rect 19618 46732 19628 46788
rect 19684 46732 20748 46788
rect 20804 46732 20814 46788
rect 22540 46676 22596 46844
rect 30930 46732 30940 46788
rect 30996 46732 31948 46788
rect 32004 46732 32732 46788
rect 32788 46732 32798 46788
rect 38994 46732 39004 46788
rect 39060 46732 40012 46788
rect 40068 46732 41468 46788
rect 41524 46732 41534 46788
rect 48178 46732 48188 46788
rect 48244 46732 50428 46788
rect 50484 46732 50494 46788
rect 3042 46620 3052 46676
rect 3108 46620 3948 46676
rect 4004 46620 4014 46676
rect 6850 46620 6860 46676
rect 6916 46620 7644 46676
rect 7700 46620 7710 46676
rect 10210 46620 10220 46676
rect 10276 46620 11228 46676
rect 11284 46620 12124 46676
rect 12180 46620 12190 46676
rect 16594 46620 16604 46676
rect 16660 46620 17724 46676
rect 17780 46620 17790 46676
rect 20178 46620 20188 46676
rect 20244 46620 20524 46676
rect 20580 46620 20590 46676
rect 20850 46620 20860 46676
rect 20916 46620 22204 46676
rect 22260 46620 23324 46676
rect 23380 46620 23390 46676
rect 26114 46620 26124 46676
rect 26180 46620 26908 46676
rect 26964 46620 26974 46676
rect 32274 46620 32284 46676
rect 32340 46620 33068 46676
rect 33124 46620 33134 46676
rect 33506 46620 33516 46676
rect 33572 46620 36988 46676
rect 37044 46620 37054 46676
rect 41234 46620 41244 46676
rect 41300 46620 41804 46676
rect 41860 46620 42924 46676
rect 42980 46620 42990 46676
rect 22418 46508 22428 46564
rect 22484 46508 23660 46564
rect 23716 46508 23726 46564
rect 31826 46508 31836 46564
rect 31892 46508 34860 46564
rect 34916 46508 34926 46564
rect 38322 46508 38332 46564
rect 38388 46508 40348 46564
rect 40404 46508 42028 46564
rect 42084 46508 42094 46564
rect 47842 46508 47852 46564
rect 47908 46508 50316 46564
rect 50372 46508 51548 46564
rect 51604 46508 51614 46564
rect 23426 46396 23436 46452
rect 23492 46396 27020 46452
rect 27076 46396 27086 46452
rect 43250 46396 43260 46452
rect 43316 46396 45052 46452
rect 45108 46396 45118 46452
rect 51426 46396 51436 46452
rect 51492 46396 53788 46452
rect 53844 46396 54460 46452
rect 54516 46396 54526 46452
rect 27794 46284 27804 46340
rect 27860 46284 29372 46340
rect 29428 46284 29438 46340
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 5618 46060 5628 46116
rect 5684 46060 6300 46116
rect 6356 46060 8540 46116
rect 8596 46060 9660 46116
rect 9716 46060 9726 46116
rect 31042 46060 31052 46116
rect 31108 46060 31948 46116
rect 32004 46060 32014 46116
rect 35298 46060 35308 46116
rect 35364 46060 36316 46116
rect 36372 46060 40572 46116
rect 40628 46060 40638 46116
rect 52770 46060 52780 46116
rect 52836 46060 54348 46116
rect 54404 46060 54414 46116
rect 4162 45948 4172 46004
rect 4228 45948 4238 46004
rect 14802 45948 14812 46004
rect 14868 45948 15484 46004
rect 15540 45948 15550 46004
rect 39778 45948 39788 46004
rect 39844 45948 41356 46004
rect 41412 45948 41422 46004
rect 46386 45948 46396 46004
rect 46452 45948 47628 46004
rect 47684 45948 48188 46004
rect 48244 45948 48254 46004
rect 3154 45836 3164 45892
rect 3220 45836 3724 45892
rect 3780 45836 3790 45892
rect 4172 45668 4228 45948
rect 38546 45836 38556 45892
rect 38612 45836 38892 45892
rect 38948 45836 39564 45892
rect 39620 45836 40908 45892
rect 40964 45836 40974 45892
rect 44930 45836 44940 45892
rect 44996 45836 48748 45892
rect 48804 45836 48814 45892
rect 6402 45724 6412 45780
rect 6468 45724 8652 45780
rect 8708 45724 8718 45780
rect 12786 45724 12796 45780
rect 12852 45724 13804 45780
rect 13860 45724 13870 45780
rect 15922 45724 15932 45780
rect 15988 45724 16716 45780
rect 16772 45724 18732 45780
rect 18788 45724 18798 45780
rect 36418 45724 36428 45780
rect 36484 45724 38780 45780
rect 38836 45724 39116 45780
rect 39172 45724 40572 45780
rect 40628 45724 40638 45780
rect 40786 45724 40796 45780
rect 40852 45724 44828 45780
rect 44884 45724 44894 45780
rect 46162 45724 46172 45780
rect 46228 45724 47516 45780
rect 47572 45724 47964 45780
rect 48020 45724 50988 45780
rect 51044 45724 52780 45780
rect 52836 45724 52846 45780
rect 4172 45612 4620 45668
rect 4676 45612 4686 45668
rect 9762 45612 9772 45668
rect 9828 45612 11340 45668
rect 11396 45612 11900 45668
rect 11956 45612 13580 45668
rect 13636 45612 13646 45668
rect 19058 45612 19068 45668
rect 19124 45612 22316 45668
rect 22372 45612 26124 45668
rect 26180 45612 26190 45668
rect 27234 45612 27244 45668
rect 27300 45612 28252 45668
rect 28308 45612 28318 45668
rect 36082 45612 36092 45668
rect 36148 45612 37100 45668
rect 37156 45612 37166 45668
rect 37426 45612 37436 45668
rect 37492 45612 38332 45668
rect 38388 45612 38556 45668
rect 38612 45612 38622 45668
rect 43586 45612 43596 45668
rect 43652 45612 45836 45668
rect 45892 45612 45902 45668
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 50546 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50830 45500
rect 10434 45388 10444 45444
rect 10500 45388 15932 45444
rect 15988 45388 15998 45444
rect 20514 45388 20524 45444
rect 20580 45388 21532 45444
rect 21588 45388 21598 45444
rect 36194 45388 36204 45444
rect 36260 45388 36270 45444
rect 37314 45388 37324 45444
rect 37380 45388 41468 45444
rect 41524 45388 41534 45444
rect 43362 45388 43372 45444
rect 43428 45388 45388 45444
rect 45444 45388 45454 45444
rect 36204 45332 36260 45388
rect 2146 45276 2156 45332
rect 2212 45276 3388 45332
rect 3444 45276 3454 45332
rect 4722 45276 4732 45332
rect 4788 45276 6412 45332
rect 6468 45276 6478 45332
rect 9762 45276 9772 45332
rect 9828 45276 11116 45332
rect 11172 45276 11182 45332
rect 12002 45276 12012 45332
rect 12068 45276 13916 45332
rect 13972 45276 14364 45332
rect 14420 45276 14430 45332
rect 16370 45276 16380 45332
rect 16436 45276 17724 45332
rect 17780 45276 17790 45332
rect 21858 45276 21868 45332
rect 21924 45276 24332 45332
rect 24388 45276 24398 45332
rect 36204 45276 36764 45332
rect 36820 45276 38220 45332
rect 38276 45276 38286 45332
rect 45042 45276 45052 45332
rect 45108 45276 45836 45332
rect 45892 45276 46732 45332
rect 46788 45276 46798 45332
rect 3388 45220 3444 45276
rect 3388 45164 5124 45220
rect 8978 45164 8988 45220
rect 9044 45164 12348 45220
rect 12404 45164 12414 45220
rect 12562 45164 12572 45220
rect 12628 45164 14140 45220
rect 14196 45164 15820 45220
rect 15876 45164 15886 45220
rect 17602 45164 17612 45220
rect 17668 45164 18956 45220
rect 19012 45164 19022 45220
rect 26562 45164 26572 45220
rect 26628 45164 27132 45220
rect 27188 45164 27580 45220
rect 27636 45164 27646 45220
rect 34850 45164 34860 45220
rect 34916 45164 35308 45220
rect 35364 45164 35374 45220
rect 52434 45164 52444 45220
rect 52500 45164 52892 45220
rect 52948 45164 52958 45220
rect 0 45108 800 45136
rect 5068 45108 5124 45164
rect 0 45052 3500 45108
rect 3556 45052 3566 45108
rect 5058 45052 5068 45108
rect 5124 45052 5134 45108
rect 5842 45052 5852 45108
rect 5908 45052 7196 45108
rect 7252 45052 7262 45108
rect 9202 45052 9212 45108
rect 9268 45052 15148 45108
rect 24770 45052 24780 45108
rect 24836 45052 26796 45108
rect 26852 45052 27468 45108
rect 27524 45052 27534 45108
rect 33730 45052 33740 45108
rect 33796 45052 34972 45108
rect 35028 45052 35038 45108
rect 43026 45052 43036 45108
rect 43092 45052 44940 45108
rect 44996 45052 45500 45108
rect 45556 45052 45566 45108
rect 51986 45052 51996 45108
rect 52052 45052 52556 45108
rect 52612 45052 53004 45108
rect 53060 45052 53070 45108
rect 53778 45052 53788 45108
rect 53844 45052 54124 45108
rect 54180 45052 54572 45108
rect 54628 45052 54638 45108
rect 0 45024 800 45052
rect 3042 44940 3052 44996
rect 3108 44940 5628 44996
rect 5684 44940 5694 44996
rect 9650 44940 9660 44996
rect 9716 44940 12124 44996
rect 12180 44940 12190 44996
rect 15092 44884 15148 45052
rect 33506 44940 33516 44996
rect 33572 44940 35644 44996
rect 35700 44940 35710 44996
rect 43922 44940 43932 44996
rect 43988 44940 46284 44996
rect 46340 44940 46844 44996
rect 46900 44940 49084 44996
rect 49140 44940 49756 44996
rect 49812 44940 49822 44996
rect 3378 44828 3388 44884
rect 3444 44828 3948 44884
rect 4004 44828 5964 44884
rect 6020 44828 6636 44884
rect 6692 44828 6702 44884
rect 9986 44828 9996 44884
rect 10052 44828 11340 44884
rect 11396 44828 11406 44884
rect 15092 44828 16604 44884
rect 16660 44828 16670 44884
rect 32284 44828 35532 44884
rect 35588 44828 35598 44884
rect 50082 44828 50092 44884
rect 50148 44828 50652 44884
rect 50708 44828 51548 44884
rect 51604 44828 51614 44884
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 2706 44604 2716 44660
rect 2772 44604 3220 44660
rect 924 44492 1932 44548
rect 1988 44492 1998 44548
rect 0 44436 800 44464
rect 924 44436 980 44492
rect 0 44380 980 44436
rect 1362 44380 1372 44436
rect 1428 44380 2380 44436
rect 2436 44380 2716 44436
rect 2772 44380 2782 44436
rect 0 44352 800 44380
rect 1586 44268 1596 44324
rect 1652 44268 1662 44324
rect 2146 44268 2156 44324
rect 2212 44268 2940 44324
rect 2996 44268 3006 44324
rect 1596 44212 1652 44268
rect 3164 44212 3220 44604
rect 17826 44492 17836 44548
rect 17892 44492 19404 44548
rect 19460 44492 20412 44548
rect 20468 44492 20478 44548
rect 32284 44436 32340 44828
rect 42242 44716 42252 44772
rect 42308 44716 45276 44772
rect 45332 44716 45342 44772
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 5058 44380 5068 44436
rect 5124 44380 7644 44436
rect 7700 44380 7710 44436
rect 32274 44380 32284 44436
rect 32340 44380 32350 44436
rect 34962 44380 34972 44436
rect 35028 44380 35532 44436
rect 35588 44380 35598 44436
rect 38658 44380 38668 44436
rect 38724 44380 40460 44436
rect 40516 44380 40526 44436
rect 43922 44380 43932 44436
rect 43988 44380 46060 44436
rect 46116 44380 46126 44436
rect 4610 44268 4620 44324
rect 4676 44268 6860 44324
rect 6916 44268 6926 44324
rect 7522 44268 7532 44324
rect 7588 44268 9548 44324
rect 9604 44268 9614 44324
rect 12338 44268 12348 44324
rect 12404 44268 13468 44324
rect 13524 44268 13534 44324
rect 19954 44268 19964 44324
rect 20020 44268 21308 44324
rect 21364 44268 21374 44324
rect 51650 44268 51660 44324
rect 51716 44268 52444 44324
rect 52500 44268 52510 44324
rect 924 44156 1652 44212
rect 2818 44156 2828 44212
rect 2884 44156 6300 44212
rect 6356 44156 6366 44212
rect 8418 44156 8428 44212
rect 8484 44156 9436 44212
rect 9492 44156 9502 44212
rect 33506 44156 33516 44212
rect 33572 44156 34412 44212
rect 34468 44156 34478 44212
rect 43922 44156 43932 44212
rect 43988 44156 44492 44212
rect 44548 44156 45052 44212
rect 45108 44156 45612 44212
rect 45668 44156 45678 44212
rect 46946 44156 46956 44212
rect 47012 44156 48188 44212
rect 48244 44156 49196 44212
rect 49252 44156 49262 44212
rect 50754 44156 50764 44212
rect 50820 44156 51884 44212
rect 51940 44156 51950 44212
rect 0 43764 800 43792
rect 924 43764 980 44156
rect 1698 44044 1708 44100
rect 1764 44044 1774 44100
rect 3378 44044 3388 44100
rect 3444 44044 5852 44100
rect 5908 44044 5918 44100
rect 6402 44044 6412 44100
rect 6468 44044 7196 44100
rect 7252 44044 7262 44100
rect 19282 44044 19292 44100
rect 19348 44044 19852 44100
rect 19908 44044 19918 44100
rect 26534 44044 26572 44100
rect 26628 44044 26638 44100
rect 1708 43876 1764 44044
rect 15092 43932 16828 43988
rect 16884 43932 16894 43988
rect 38770 43932 38780 43988
rect 38836 43932 39452 43988
rect 39508 43932 39518 43988
rect 1708 43820 3612 43876
rect 3668 43820 3678 43876
rect 15092 43764 15148 43932
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 50546 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50830 43932
rect 38434 43820 38444 43876
rect 38500 43820 39004 43876
rect 39060 43820 39070 43876
rect 0 43708 980 43764
rect 2034 43708 2044 43764
rect 2100 43708 6860 43764
rect 6916 43708 6926 43764
rect 14018 43708 14028 43764
rect 14084 43708 15148 43764
rect 25106 43708 25116 43764
rect 25172 43708 25620 43764
rect 32050 43708 32060 43764
rect 32116 43708 33628 43764
rect 33684 43708 33694 43764
rect 36194 43708 36204 43764
rect 36260 43708 37100 43764
rect 37156 43708 37166 43764
rect 41682 43708 41692 43764
rect 41748 43708 43036 43764
rect 43092 43708 43102 43764
rect 51090 43708 51100 43764
rect 51156 43708 51996 43764
rect 52052 43708 52062 43764
rect 54114 43708 54124 43764
rect 54180 43708 55244 43764
rect 55300 43708 55310 43764
rect 0 43680 800 43708
rect 25564 43652 25620 43708
rect 2706 43596 2716 43652
rect 2772 43596 4620 43652
rect 4676 43596 5740 43652
rect 5796 43596 5806 43652
rect 19506 43596 19516 43652
rect 19572 43596 20076 43652
rect 20132 43596 22540 43652
rect 22596 43596 22606 43652
rect 24210 43596 24220 43652
rect 24276 43596 25340 43652
rect 25396 43596 25406 43652
rect 25564 43596 27076 43652
rect 27234 43596 27244 43652
rect 27300 43596 28812 43652
rect 28868 43596 29148 43652
rect 29204 43596 29214 43652
rect 34066 43596 34076 43652
rect 34132 43596 36092 43652
rect 36148 43596 37324 43652
rect 37380 43596 39340 43652
rect 39396 43596 39406 43652
rect 40562 43596 40572 43652
rect 40628 43596 42252 43652
rect 42308 43596 42318 43652
rect 43698 43596 43708 43652
rect 43764 43596 46732 43652
rect 46788 43596 46798 43652
rect 27020 43540 27076 43596
rect 3332 43484 4060 43540
rect 4116 43484 4126 43540
rect 4834 43484 4844 43540
rect 4900 43484 6748 43540
rect 6804 43484 7308 43540
rect 7364 43484 7374 43540
rect 14914 43484 14924 43540
rect 14980 43484 15764 43540
rect 24658 43484 24668 43540
rect 24724 43484 25228 43540
rect 25284 43484 25294 43540
rect 26786 43484 26796 43540
rect 3332 43428 3388 43484
rect 15708 43428 15764 43484
rect 26852 43428 26908 43540
rect 27020 43484 27132 43540
rect 27188 43484 27198 43540
rect 28018 43484 28028 43540
rect 28084 43484 28094 43540
rect 28242 43484 28252 43540
rect 28308 43484 28924 43540
rect 28980 43484 28990 43540
rect 33730 43484 33740 43540
rect 33796 43484 36204 43540
rect 36260 43484 36270 43540
rect 28028 43428 28084 43484
rect 2930 43372 2940 43428
rect 2996 43372 3388 43428
rect 3938 43372 3948 43428
rect 4004 43372 5852 43428
rect 5908 43372 5918 43428
rect 11330 43372 11340 43428
rect 11396 43372 12908 43428
rect 12964 43372 14028 43428
rect 14084 43372 14094 43428
rect 15698 43372 15708 43428
rect 15764 43372 17724 43428
rect 17780 43372 17790 43428
rect 18610 43372 18620 43428
rect 18676 43372 19404 43428
rect 19460 43372 19470 43428
rect 19730 43372 19740 43428
rect 19796 43372 20412 43428
rect 20468 43372 20478 43428
rect 26852 43372 28084 43428
rect 36866 43372 36876 43428
rect 36932 43372 37884 43428
rect 37940 43372 37950 43428
rect 51538 43372 51548 43428
rect 51604 43372 53228 43428
rect 53284 43372 53294 43428
rect 3948 43316 4004 43372
rect 3042 43260 3052 43316
rect 3108 43260 4004 43316
rect 4274 43260 4284 43316
rect 4340 43260 8092 43316
rect 8148 43260 17388 43316
rect 17444 43260 17454 43316
rect 26338 43260 26348 43316
rect 26404 43260 26908 43316
rect 26964 43260 26974 43316
rect 27122 43260 27132 43316
rect 27188 43260 28476 43316
rect 28532 43260 28542 43316
rect 34738 43260 34748 43316
rect 34804 43260 35980 43316
rect 36036 43260 36046 43316
rect 39778 43260 39788 43316
rect 39844 43260 40572 43316
rect 40628 43260 40638 43316
rect 42578 43260 42588 43316
rect 42644 43260 44156 43316
rect 44212 43260 46396 43316
rect 46452 43260 46462 43316
rect 49186 43260 49196 43316
rect 49252 43260 49756 43316
rect 49812 43260 49822 43316
rect 55346 43260 55356 43316
rect 55412 43260 57148 43316
rect 57204 43260 57214 43316
rect 5506 43148 5516 43204
rect 5572 43148 11228 43204
rect 11284 43148 11294 43204
rect 25554 43148 25564 43204
rect 25620 43148 26124 43204
rect 26180 43148 26190 43204
rect 30594 43148 30604 43204
rect 30660 43148 31388 43204
rect 31444 43148 33180 43204
rect 33236 43148 33246 43204
rect 35858 43148 35868 43204
rect 35924 43148 37212 43204
rect 37268 43148 37278 43204
rect 38994 43148 39004 43204
rect 39060 43148 40012 43204
rect 40068 43148 41020 43204
rect 41076 43148 41086 43204
rect 0 43092 800 43120
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 0 43036 3388 43092
rect 0 43008 800 43036
rect 3332 42980 3388 43036
rect 15092 43036 22988 43092
rect 23044 43036 23054 43092
rect 15092 42980 15148 43036
rect 3332 42924 15148 42980
rect 25778 42924 25788 42980
rect 25844 42924 26124 42980
rect 26180 42924 26908 42980
rect 28018 42924 28028 42980
rect 28084 42924 29260 42980
rect 29316 42924 29326 42980
rect 26852 42868 26908 42924
rect 2034 42812 2044 42868
rect 2100 42812 2716 42868
rect 2772 42812 4620 42868
rect 4676 42812 4686 42868
rect 26852 42812 27244 42868
rect 27300 42812 27310 42868
rect 33282 42812 33292 42868
rect 33348 42812 34524 42868
rect 34580 42812 34590 42868
rect 34738 42812 34748 42868
rect 34804 42812 38892 42868
rect 38948 42812 43708 42868
rect 43764 42812 43774 42868
rect 21410 42700 21420 42756
rect 21476 42700 22092 42756
rect 22148 42700 22158 42756
rect 23874 42700 23884 42756
rect 23940 42700 25340 42756
rect 25396 42700 25406 42756
rect 43586 42700 43596 42756
rect 43652 42700 45388 42756
rect 45444 42700 45454 42756
rect 48962 42700 48972 42756
rect 49028 42700 49980 42756
rect 50036 42700 50046 42756
rect 54674 42700 54684 42756
rect 54740 42700 56700 42756
rect 56756 42700 56766 42756
rect 16370 42588 16380 42644
rect 16436 42588 18060 42644
rect 18116 42588 19180 42644
rect 19236 42588 19246 42644
rect 20514 42588 20524 42644
rect 20580 42588 21308 42644
rect 21364 42588 21374 42644
rect 27794 42588 27804 42644
rect 27860 42588 29148 42644
rect 29204 42588 29214 42644
rect 30594 42588 30604 42644
rect 30660 42588 31724 42644
rect 31780 42588 31790 42644
rect 34850 42588 34860 42644
rect 34916 42588 35756 42644
rect 35812 42588 36988 42644
rect 37044 42588 37054 42644
rect 9762 42476 9772 42532
rect 9828 42476 10108 42532
rect 10164 42476 10174 42532
rect 12674 42476 12684 42532
rect 12740 42476 13804 42532
rect 13860 42476 13870 42532
rect 17602 42476 17612 42532
rect 17668 42476 18956 42532
rect 19012 42476 19022 42532
rect 20738 42476 20748 42532
rect 20804 42476 21644 42532
rect 21700 42476 21710 42532
rect 26786 42476 26796 42532
rect 26852 42476 27132 42532
rect 27188 42476 27198 42532
rect 36530 42476 36540 42532
rect 36596 42476 37548 42532
rect 37604 42476 37614 42532
rect 47394 42476 47404 42532
rect 47460 42476 50428 42532
rect 50484 42476 52780 42532
rect 52836 42476 52846 42532
rect 0 42420 800 42448
rect 0 42364 1932 42420
rect 1988 42364 1998 42420
rect 22642 42364 22652 42420
rect 22708 42364 22718 42420
rect 0 42336 800 42364
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 22652 42196 22708 42364
rect 50546 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50830 42364
rect 36194 42252 36204 42308
rect 36260 42252 37548 42308
rect 37604 42252 37614 42308
rect 38612 42252 39788 42308
rect 39844 42252 42364 42308
rect 42420 42252 42430 42308
rect 38612 42196 38668 42252
rect 13916 42140 16492 42196
rect 16548 42140 16716 42196
rect 16772 42140 27132 42196
rect 27188 42140 27198 42196
rect 36978 42140 36988 42196
rect 37044 42140 38668 42196
rect 40114 42140 40124 42196
rect 40180 42140 41468 42196
rect 41524 42140 44940 42196
rect 44996 42140 45006 42196
rect 54898 42140 54908 42196
rect 54964 42140 55692 42196
rect 55748 42140 55758 42196
rect 13916 42084 13972 42140
rect 5404 42028 6860 42084
rect 6916 42028 6926 42084
rect 10434 42028 10444 42084
rect 10500 42028 13916 42084
rect 13972 42028 13982 42084
rect 14354 42028 14364 42084
rect 14420 42028 15484 42084
rect 15540 42028 15550 42084
rect 44258 42028 44268 42084
rect 44324 42028 45500 42084
rect 45556 42028 45566 42084
rect 52770 42028 52780 42084
rect 52836 42028 54348 42084
rect 54404 42028 54414 42084
rect 5404 41972 5460 42028
rect 1698 41916 1708 41972
rect 1764 41916 2828 41972
rect 2884 41916 2894 41972
rect 5394 41916 5404 41972
rect 5460 41916 5470 41972
rect 6290 41916 6300 41972
rect 6356 41916 6636 41972
rect 6692 41916 6702 41972
rect 8306 41916 8316 41972
rect 8372 41916 10668 41972
rect 10724 41916 12796 41972
rect 12852 41916 12862 41972
rect 13346 41916 13356 41972
rect 13412 41916 15372 41972
rect 15428 41916 15438 41972
rect 21634 41916 21644 41972
rect 21700 41916 22204 41972
rect 22260 41916 23100 41972
rect 23156 41916 23166 41972
rect 30706 41916 30716 41972
rect 30772 41916 31836 41972
rect 31892 41916 31902 41972
rect 32386 41916 32396 41972
rect 32452 41916 33404 41972
rect 33460 41916 33470 41972
rect 38098 41916 38108 41972
rect 38164 41916 38556 41972
rect 38612 41916 39564 41972
rect 39620 41916 39630 41972
rect 40114 41916 40124 41972
rect 40180 41916 42700 41972
rect 42756 41916 42766 41972
rect 43474 41916 43484 41972
rect 43540 41916 45388 41972
rect 45444 41916 45454 41972
rect 48962 41916 48972 41972
rect 49028 41916 49868 41972
rect 49924 41916 52444 41972
rect 52500 41916 52510 41972
rect 4610 41804 4620 41860
rect 4676 41804 6188 41860
rect 6244 41804 6254 41860
rect 11554 41804 11564 41860
rect 11620 41804 12012 41860
rect 12068 41804 14252 41860
rect 14308 41804 14318 41860
rect 25638 41804 25676 41860
rect 25732 41804 25742 41860
rect 33282 41804 33292 41860
rect 33348 41804 34748 41860
rect 34804 41804 34814 41860
rect 46162 41804 46172 41860
rect 46228 41804 46956 41860
rect 47012 41804 49532 41860
rect 49588 41804 49598 41860
rect 49746 41804 49756 41860
rect 49812 41804 51436 41860
rect 51492 41804 51502 41860
rect 51986 41804 51996 41860
rect 52052 41804 54236 41860
rect 54292 41804 54302 41860
rect 0 41748 800 41776
rect 0 41692 3836 41748
rect 3892 41692 3902 41748
rect 8642 41692 8652 41748
rect 8708 41692 10892 41748
rect 10948 41692 10958 41748
rect 49298 41692 49308 41748
rect 49364 41692 52892 41748
rect 52948 41692 52958 41748
rect 0 41664 800 41692
rect 8082 41580 8092 41636
rect 8148 41580 9324 41636
rect 9380 41580 9660 41636
rect 9716 41580 9726 41636
rect 47394 41580 47404 41636
rect 47460 41580 47964 41636
rect 48020 41580 49756 41636
rect 49812 41580 49822 41636
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 21746 41468 21756 41524
rect 21812 41468 22540 41524
rect 22596 41468 23324 41524
rect 23380 41468 23390 41524
rect 50306 41468 50316 41524
rect 50372 41468 52668 41524
rect 52724 41468 52734 41524
rect 4274 41356 4284 41412
rect 4340 41356 8988 41412
rect 9044 41356 9054 41412
rect 6178 41244 6188 41300
rect 6244 41244 7196 41300
rect 7252 41244 7262 41300
rect 16706 41244 16716 41300
rect 16772 41244 17500 41300
rect 17556 41244 17566 41300
rect 36306 41244 36316 41300
rect 36372 41244 39228 41300
rect 39284 41244 39294 41300
rect 6738 41132 6748 41188
rect 6804 41132 7420 41188
rect 7476 41132 7486 41188
rect 10098 41132 10108 41188
rect 10164 41132 11564 41188
rect 11620 41132 11900 41188
rect 11956 41132 12460 41188
rect 12516 41132 12526 41188
rect 17938 41132 17948 41188
rect 18004 41132 18732 41188
rect 18788 41132 18798 41188
rect 30818 41132 30828 41188
rect 30884 41132 31948 41188
rect 32004 41132 32014 41188
rect 32274 41132 32284 41188
rect 32340 41132 33292 41188
rect 33348 41132 33358 41188
rect 42578 41132 42588 41188
rect 42644 41132 44940 41188
rect 44996 41132 45006 41188
rect 50418 41132 50428 41188
rect 50484 41132 51772 41188
rect 51828 41132 51838 41188
rect 0 41076 800 41104
rect 0 41020 1708 41076
rect 1764 41020 1774 41076
rect 3714 41020 3724 41076
rect 3780 41020 4732 41076
rect 4788 41020 8540 41076
rect 8596 41020 8606 41076
rect 11106 41020 11116 41076
rect 11172 41020 12236 41076
rect 12292 41020 12302 41076
rect 16594 41020 16604 41076
rect 16660 41020 17612 41076
rect 17668 41020 18844 41076
rect 18900 41020 18910 41076
rect 19282 41020 19292 41076
rect 19348 41020 19964 41076
rect 20020 41020 20030 41076
rect 33506 41020 33516 41076
rect 33572 41020 34636 41076
rect 34692 41020 37100 41076
rect 37156 41020 37166 41076
rect 38322 41020 38332 41076
rect 38388 41020 39340 41076
rect 39396 41020 39406 41076
rect 0 40992 800 41020
rect 4946 40908 4956 40964
rect 5012 40908 9884 40964
rect 9940 40908 9950 40964
rect 17826 40908 17836 40964
rect 17892 40908 19068 40964
rect 19124 40908 19134 40964
rect 22082 40908 22092 40964
rect 22148 40908 23772 40964
rect 23828 40908 23838 40964
rect 25330 40908 25340 40964
rect 25396 40908 26012 40964
rect 26068 40908 26684 40964
rect 26740 40908 26750 40964
rect 31826 40908 31836 40964
rect 31892 40908 32508 40964
rect 32564 40908 32574 40964
rect 33842 40908 33852 40964
rect 33908 40908 34412 40964
rect 34468 40908 34478 40964
rect 51986 40908 51996 40964
rect 52052 40908 54684 40964
rect 54740 40908 55244 40964
rect 55300 40908 55310 40964
rect 4274 40796 4284 40852
rect 4340 40796 9100 40852
rect 9156 40796 9166 40852
rect 25890 40796 25900 40852
rect 25956 40796 26460 40852
rect 26516 40796 26526 40852
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 50546 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50830 40796
rect 4162 40684 4172 40740
rect 4228 40684 6860 40740
rect 6916 40684 9324 40740
rect 9380 40684 9390 40740
rect 21298 40684 21308 40740
rect 21364 40684 27244 40740
rect 27300 40684 27310 40740
rect 43250 40684 43260 40740
rect 43316 40684 44828 40740
rect 44884 40684 44894 40740
rect 6626 40572 6636 40628
rect 6692 40572 7196 40628
rect 7252 40572 7262 40628
rect 7410 40572 7420 40628
rect 7476 40572 9212 40628
rect 9268 40572 9278 40628
rect 9436 40572 13356 40628
rect 13412 40572 13422 40628
rect 19058 40572 19068 40628
rect 19124 40572 19852 40628
rect 19908 40572 19918 40628
rect 20514 40572 20524 40628
rect 20580 40572 21756 40628
rect 21812 40572 21822 40628
rect 35410 40572 35420 40628
rect 35476 40572 36764 40628
rect 36820 40572 36830 40628
rect 38546 40572 38556 40628
rect 38612 40572 40908 40628
rect 40964 40572 40974 40628
rect 48290 40572 48300 40628
rect 48356 40572 50652 40628
rect 50708 40572 50718 40628
rect 52994 40572 53004 40628
rect 53060 40572 54124 40628
rect 54180 40572 55132 40628
rect 55188 40572 55198 40628
rect 7420 40516 7476 40572
rect 9436 40516 9492 40572
rect 5058 40460 5068 40516
rect 5124 40460 6300 40516
rect 6356 40460 7476 40516
rect 9090 40460 9100 40516
rect 9156 40460 9492 40516
rect 10658 40460 10668 40516
rect 10724 40460 11788 40516
rect 11844 40460 14028 40516
rect 14084 40460 14094 40516
rect 14578 40460 14588 40516
rect 14644 40460 15148 40516
rect 18274 40460 18284 40516
rect 18340 40460 19292 40516
rect 19348 40460 20412 40516
rect 20468 40460 20478 40516
rect 27122 40460 27132 40516
rect 27188 40460 29148 40516
rect 29204 40460 29214 40516
rect 40674 40460 40684 40516
rect 40740 40460 42028 40516
rect 42084 40460 42094 40516
rect 42466 40460 42476 40516
rect 42532 40460 49084 40516
rect 49140 40460 51996 40516
rect 52052 40460 52062 40516
rect 52210 40460 52220 40516
rect 52276 40460 53228 40516
rect 53284 40460 55468 40516
rect 55524 40460 55534 40516
rect 0 40404 800 40432
rect 15092 40404 15148 40460
rect 0 40348 1932 40404
rect 1988 40348 1998 40404
rect 3602 40348 3612 40404
rect 3668 40348 4060 40404
rect 4116 40348 6076 40404
rect 6132 40348 6142 40404
rect 7522 40348 7532 40404
rect 7588 40348 8316 40404
rect 8372 40348 8382 40404
rect 10882 40348 10892 40404
rect 10948 40348 12460 40404
rect 12516 40348 13244 40404
rect 13300 40348 13310 40404
rect 15092 40348 16156 40404
rect 16212 40348 16222 40404
rect 18834 40348 18844 40404
rect 18900 40348 19740 40404
rect 19796 40348 20188 40404
rect 20244 40348 20254 40404
rect 24434 40348 24444 40404
rect 24500 40348 25116 40404
rect 25172 40348 25564 40404
rect 25620 40348 25630 40404
rect 33282 40348 33292 40404
rect 33348 40348 34076 40404
rect 34132 40348 34142 40404
rect 37650 40348 37660 40404
rect 37716 40348 38332 40404
rect 38388 40348 38398 40404
rect 41458 40348 41468 40404
rect 41524 40348 43036 40404
rect 43092 40348 43102 40404
rect 43362 40348 43372 40404
rect 43428 40348 43596 40404
rect 43652 40348 43662 40404
rect 53330 40348 53340 40404
rect 53396 40348 54012 40404
rect 54068 40348 54078 40404
rect 0 40320 800 40348
rect 4620 40292 4676 40348
rect 4610 40236 4620 40292
rect 4676 40236 4686 40292
rect 16034 40236 16044 40292
rect 16100 40236 17724 40292
rect 17780 40236 17790 40292
rect 32470 40236 32508 40292
rect 32564 40236 32574 40292
rect 34402 40236 34412 40292
rect 34468 40236 35308 40292
rect 35364 40236 35374 40292
rect 38546 40236 38556 40292
rect 38612 40236 40348 40292
rect 40404 40236 40414 40292
rect 45938 40236 45948 40292
rect 46004 40236 47180 40292
rect 47236 40236 48748 40292
rect 48804 40236 48814 40292
rect 3938 40124 3948 40180
rect 4004 40124 4284 40180
rect 4340 40124 4732 40180
rect 4788 40124 4798 40180
rect 8978 40124 8988 40180
rect 9044 40124 13244 40180
rect 13300 40124 13310 40180
rect 17378 40124 17388 40180
rect 17444 40124 20524 40180
rect 20580 40124 20590 40180
rect 5842 40012 5852 40068
rect 5908 40012 20636 40068
rect 20692 40012 20702 40068
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 20402 39900 20412 39956
rect 20468 39900 25900 39956
rect 25956 39900 25966 39956
rect 28690 39788 28700 39844
rect 28756 39788 29260 39844
rect 29316 39788 30156 39844
rect 30212 39788 31052 39844
rect 31108 39788 31118 39844
rect 48822 39788 48860 39844
rect 48916 39788 48926 39844
rect 0 39732 800 39760
rect 0 39676 1932 39732
rect 1988 39676 1998 39732
rect 18162 39676 18172 39732
rect 18228 39676 21588 39732
rect 38210 39676 38220 39732
rect 38276 39676 39452 39732
rect 39508 39676 40572 39732
rect 40628 39676 40638 39732
rect 48178 39676 48188 39732
rect 48244 39676 48972 39732
rect 49028 39676 49038 39732
rect 0 39648 800 39676
rect 21532 39620 21588 39676
rect 2034 39564 2044 39620
rect 2100 39564 5964 39620
rect 6020 39564 6030 39620
rect 9090 39564 9100 39620
rect 9156 39564 11340 39620
rect 11396 39564 11406 39620
rect 16146 39564 16156 39620
rect 16212 39564 16828 39620
rect 16884 39564 16894 39620
rect 17490 39564 17500 39620
rect 17556 39564 18508 39620
rect 18564 39564 19180 39620
rect 19236 39564 19246 39620
rect 21522 39564 21532 39620
rect 21588 39564 23996 39620
rect 24052 39564 24062 39620
rect 41794 39564 41804 39620
rect 41860 39564 43484 39620
rect 43540 39564 43550 39620
rect 46610 39564 46620 39620
rect 46676 39564 49308 39620
rect 49364 39564 49374 39620
rect 51090 39564 51100 39620
rect 51156 39564 53452 39620
rect 53508 39564 53518 39620
rect 8082 39452 8092 39508
rect 8148 39452 11452 39508
rect 11508 39452 12908 39508
rect 12964 39452 12974 39508
rect 16258 39452 16268 39508
rect 16324 39452 17836 39508
rect 17892 39452 17902 39508
rect 19394 39452 19404 39508
rect 19460 39452 20188 39508
rect 20244 39452 21644 39508
rect 21700 39452 21710 39508
rect 26450 39452 26460 39508
rect 26516 39452 27132 39508
rect 27188 39452 27198 39508
rect 37202 39452 37212 39508
rect 37268 39452 38668 39508
rect 51874 39452 51884 39508
rect 51940 39452 52332 39508
rect 52388 39452 53004 39508
rect 53060 39452 53070 39508
rect 1250 39340 1260 39396
rect 1316 39340 2044 39396
rect 2100 39340 2110 39396
rect 9986 39340 9996 39396
rect 10052 39340 10556 39396
rect 10612 39340 10622 39396
rect 18946 39340 18956 39396
rect 19012 39340 21308 39396
rect 21364 39340 21374 39396
rect 25218 39340 25228 39396
rect 25284 39340 25900 39396
rect 25956 39340 25966 39396
rect 38612 39284 38668 39452
rect 48066 39340 48076 39396
rect 48132 39340 48748 39396
rect 48804 39340 48814 39396
rect 38612 39228 39116 39284
rect 39172 39228 45612 39284
rect 45668 39228 48860 39284
rect 48916 39228 48926 39284
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 50546 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50830 39228
rect 52210 39116 52220 39172
rect 52276 39116 53116 39172
rect 53172 39116 53182 39172
rect 0 39060 800 39088
rect 0 39004 5516 39060
rect 5572 39004 9436 39060
rect 9492 39004 9502 39060
rect 12114 39004 12124 39060
rect 12180 39004 13804 39060
rect 13860 39004 13870 39060
rect 17378 39004 17388 39060
rect 17444 39004 18060 39060
rect 18116 39004 18126 39060
rect 23874 39004 23884 39060
rect 23940 39004 24556 39060
rect 24612 39004 24622 39060
rect 29474 39004 29484 39060
rect 29540 39004 30828 39060
rect 30884 39004 31164 39060
rect 31220 39004 32732 39060
rect 32788 39004 32798 39060
rect 41244 39004 43708 39060
rect 43764 39004 43774 39060
rect 45826 39004 45836 39060
rect 45892 39004 46844 39060
rect 46900 39004 46910 39060
rect 51986 39004 51996 39060
rect 52052 39004 52444 39060
rect 52500 39004 53564 39060
rect 53620 39004 53630 39060
rect 0 38976 800 39004
rect 2146 38892 2156 38948
rect 2212 38892 2716 38948
rect 2772 38892 2782 38948
rect 8306 38892 8316 38948
rect 8372 38892 10108 38948
rect 10164 38892 11228 38948
rect 11284 38892 11788 38948
rect 11844 38892 11854 38948
rect 4610 38780 4620 38836
rect 4676 38780 5180 38836
rect 5236 38780 5246 38836
rect 13804 38724 13860 39004
rect 14914 38892 14924 38948
rect 14980 38892 15932 38948
rect 15988 38892 16380 38948
rect 16436 38892 16446 38948
rect 17714 38892 17724 38948
rect 17780 38892 19516 38948
rect 19572 38892 19582 38948
rect 20626 38892 20636 38948
rect 20692 38892 21420 38948
rect 21476 38892 21486 38948
rect 24210 38892 24220 38948
rect 24276 38892 25004 38948
rect 25060 38892 25340 38948
rect 25396 38892 25406 38948
rect 41244 38836 41300 39004
rect 43474 38892 43484 38948
rect 43540 38892 44492 38948
rect 44548 38892 44558 38948
rect 14130 38780 14140 38836
rect 14196 38780 15372 38836
rect 15428 38780 15438 38836
rect 19954 38780 19964 38836
rect 20020 38780 21532 38836
rect 21588 38780 22428 38836
rect 22484 38780 23548 38836
rect 23604 38780 23614 38836
rect 36530 38780 36540 38836
rect 36596 38780 37660 38836
rect 37716 38780 37726 38836
rect 40338 38780 40348 38836
rect 40404 38780 41244 38836
rect 41300 38780 41310 38836
rect 43586 38780 43596 38836
rect 43652 38780 46284 38836
rect 46340 38780 46350 38836
rect 49298 38780 49308 38836
rect 49364 38780 51100 38836
rect 51156 38780 51166 38836
rect 5068 38668 6076 38724
rect 6132 38668 6142 38724
rect 13804 38668 17052 38724
rect 17108 38668 17118 38724
rect 21298 38668 21308 38724
rect 21364 38668 22204 38724
rect 22260 38668 22270 38724
rect 33954 38668 33964 38724
rect 34020 38668 34748 38724
rect 34804 38668 34814 38724
rect 1698 38556 1708 38612
rect 1764 38556 2156 38612
rect 2212 38556 2222 38612
rect 5068 38500 5124 38668
rect 13458 38556 13468 38612
rect 13524 38556 14812 38612
rect 14868 38556 14878 38612
rect 22754 38556 22764 38612
rect 22820 38556 23324 38612
rect 23380 38556 23390 38612
rect 32386 38556 32396 38612
rect 32452 38556 33180 38612
rect 33236 38556 35868 38612
rect 35924 38556 35934 38612
rect 50866 38556 50876 38612
rect 50932 38556 51884 38612
rect 51940 38556 53452 38612
rect 53508 38556 53518 38612
rect 2594 38444 2604 38500
rect 2660 38444 4060 38500
rect 4116 38444 4126 38500
rect 4946 38444 4956 38500
rect 5012 38444 5124 38500
rect 8978 38444 8988 38500
rect 9044 38444 9772 38500
rect 9828 38444 9838 38500
rect 25554 38444 25564 38500
rect 25620 38444 25630 38500
rect 0 38388 800 38416
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 25564 38388 25620 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 0 38332 3388 38388
rect 3444 38332 3454 38388
rect 13906 38332 13916 38388
rect 13972 38332 14252 38388
rect 14308 38332 14318 38388
rect 15092 38332 16940 38388
rect 16996 38332 17006 38388
rect 25330 38332 25340 38388
rect 25396 38332 25620 38388
rect 0 38304 800 38332
rect 15092 38276 15148 38332
rect 4162 38220 4172 38276
rect 4228 38220 5404 38276
rect 5460 38220 15148 38276
rect 25106 38220 25116 38276
rect 25172 38220 25900 38276
rect 25956 38220 26796 38276
rect 26852 38220 26862 38276
rect 47954 38220 47964 38276
rect 48020 38220 48030 38276
rect 47964 38164 48020 38220
rect 2268 38108 5740 38164
rect 5796 38108 5806 38164
rect 6850 38108 6860 38164
rect 6916 38108 13580 38164
rect 13636 38108 13646 38164
rect 14018 38108 14028 38164
rect 14084 38108 17388 38164
rect 17444 38108 17454 38164
rect 28130 38108 28140 38164
rect 28196 38108 28812 38164
rect 28868 38108 28878 38164
rect 34290 38108 34300 38164
rect 34356 38108 35308 38164
rect 35364 38108 35644 38164
rect 35700 38108 38780 38164
rect 38836 38108 38846 38164
rect 44930 38108 44940 38164
rect 44996 38108 48188 38164
rect 48244 38108 48254 38164
rect 2268 38052 2324 38108
rect 2258 37996 2268 38052
rect 2324 37996 2334 38052
rect 2706 37996 2716 38052
rect 2772 37996 4284 38052
rect 4340 37996 4732 38052
rect 4788 37996 6748 38052
rect 6804 37996 6814 38052
rect 13010 37996 13020 38052
rect 13076 37996 18284 38052
rect 18340 37996 19740 38052
rect 19796 37996 19806 38052
rect 25106 37996 25116 38052
rect 25172 37996 25452 38052
rect 25508 37996 25518 38052
rect 25666 37996 25676 38052
rect 25732 37996 26124 38052
rect 26180 37996 26190 38052
rect 36082 37996 36092 38052
rect 36148 37996 37436 38052
rect 37492 37996 37502 38052
rect 40226 37996 40236 38052
rect 40292 37996 40908 38052
rect 40964 37996 40974 38052
rect 47170 37996 47180 38052
rect 47236 37996 47964 38052
rect 48020 37996 48030 38052
rect 7634 37884 7644 37940
rect 7700 37884 9212 37940
rect 9268 37884 9548 37940
rect 9604 37884 9614 37940
rect 14354 37884 14364 37940
rect 14420 37884 15036 37940
rect 15092 37884 15102 37940
rect 27906 37884 27916 37940
rect 27972 37884 29820 37940
rect 29876 37884 29886 37940
rect 47618 37884 47628 37940
rect 47684 37884 48300 37940
rect 48356 37884 50092 37940
rect 50148 37884 50158 37940
rect 9874 37772 9884 37828
rect 9940 37772 10444 37828
rect 10500 37772 10780 37828
rect 10836 37772 10846 37828
rect 12786 37772 12796 37828
rect 12852 37772 15596 37828
rect 15652 37772 15662 37828
rect 17938 37772 17948 37828
rect 18004 37772 18956 37828
rect 19012 37772 19022 37828
rect 29922 37772 29932 37828
rect 29988 37772 30492 37828
rect 30548 37772 30558 37828
rect 38210 37772 38220 37828
rect 38276 37772 39788 37828
rect 39844 37772 39854 37828
rect 0 37716 800 37744
rect 0 37660 3724 37716
rect 3780 37660 3790 37716
rect 13346 37660 13356 37716
rect 13412 37660 17388 37716
rect 17444 37660 17454 37716
rect 25638 37660 25676 37716
rect 25732 37660 25742 37716
rect 26348 37660 26572 37716
rect 26628 37660 26638 37716
rect 0 37632 800 37660
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 2370 37548 2380 37604
rect 2436 37548 2716 37604
rect 2772 37548 2782 37604
rect 4834 37548 4844 37604
rect 4900 37548 5740 37604
rect 5796 37548 5806 37604
rect 15362 37548 15372 37604
rect 15428 37548 18172 37604
rect 18228 37548 18238 37604
rect 18610 37548 18620 37604
rect 18676 37548 19628 37604
rect 19684 37548 19694 37604
rect 24546 37548 24556 37604
rect 24612 37548 25004 37604
rect 25060 37548 25070 37604
rect 11218 37436 11228 37492
rect 11284 37436 12012 37492
rect 12068 37436 13916 37492
rect 13972 37436 14588 37492
rect 14644 37436 15932 37492
rect 15988 37436 15998 37492
rect 2370 37324 2380 37380
rect 2436 37324 3724 37380
rect 3780 37324 4732 37380
rect 4788 37324 4798 37380
rect 9874 37324 9884 37380
rect 9940 37324 14028 37380
rect 14084 37324 16268 37380
rect 16324 37324 16334 37380
rect 20178 37324 20188 37380
rect 20244 37324 21196 37380
rect 21252 37324 21262 37380
rect 26348 37268 26404 37660
rect 50546 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50830 37660
rect 28354 37436 28364 37492
rect 28420 37436 29596 37492
rect 29652 37436 30940 37492
rect 30996 37436 31612 37492
rect 31668 37436 32396 37492
rect 32452 37436 32462 37492
rect 32722 37436 32732 37492
rect 32788 37436 33516 37492
rect 33572 37436 34524 37492
rect 34580 37436 34590 37492
rect 40450 37436 40460 37492
rect 40516 37436 42812 37492
rect 42868 37436 42878 37492
rect 26572 37324 26796 37380
rect 26852 37324 26862 37380
rect 57810 37324 57820 37380
rect 57876 37324 57886 37380
rect 26572 37268 26628 37324
rect 5730 37212 5740 37268
rect 5796 37212 7868 37268
rect 7924 37212 7934 37268
rect 15586 37212 15596 37268
rect 15652 37212 19068 37268
rect 19124 37212 19134 37268
rect 20738 37212 20748 37268
rect 20804 37212 21532 37268
rect 21588 37212 23884 37268
rect 23940 37212 23950 37268
rect 26338 37212 26348 37268
rect 26404 37212 26414 37268
rect 26562 37212 26572 37268
rect 26628 37212 26638 37268
rect 37202 37212 37212 37268
rect 37268 37212 37436 37268
rect 37492 37212 38220 37268
rect 38276 37212 38286 37268
rect 45602 37212 45612 37268
rect 45668 37212 46732 37268
rect 46788 37212 47516 37268
rect 47572 37212 47582 37268
rect 49858 37212 49868 37268
rect 49924 37212 50764 37268
rect 50820 37212 51548 37268
rect 51604 37212 51614 37268
rect 54226 37212 54236 37268
rect 54292 37212 55468 37268
rect 55524 37212 55534 37268
rect 57820 37156 57876 37324
rect 6290 37100 6300 37156
rect 6356 37100 6860 37156
rect 6916 37100 8764 37156
rect 8820 37100 8830 37156
rect 15698 37100 15708 37156
rect 15764 37100 17500 37156
rect 17556 37100 18732 37156
rect 18788 37100 18798 37156
rect 22876 37100 29484 37156
rect 29540 37100 29550 37156
rect 30482 37100 30492 37156
rect 30548 37100 31164 37156
rect 31220 37100 31230 37156
rect 37762 37100 37772 37156
rect 37828 37100 38332 37156
rect 38388 37100 38892 37156
rect 38948 37100 38958 37156
rect 45612 37100 46172 37156
rect 46228 37100 57876 37156
rect 0 37044 800 37072
rect 22876 37044 22932 37100
rect 45612 37044 45668 37100
rect 59200 37044 60000 37072
rect 0 36988 1932 37044
rect 1988 36988 1998 37044
rect 2818 36988 2828 37044
rect 2884 36988 4396 37044
rect 4452 36988 4462 37044
rect 5506 36988 5516 37044
rect 5572 36988 8316 37044
rect 8372 36988 8876 37044
rect 8932 36988 8942 37044
rect 18946 36988 18956 37044
rect 19012 36988 20076 37044
rect 20132 36988 20142 37044
rect 22866 36988 22876 37044
rect 22932 36988 22942 37044
rect 23100 36988 24332 37044
rect 24388 36988 24398 37044
rect 26226 36988 26236 37044
rect 26292 36988 26684 37044
rect 26740 36988 26750 37044
rect 34850 36988 34860 37044
rect 34916 36988 35868 37044
rect 35924 36988 37660 37044
rect 37716 36988 37726 37044
rect 38210 36988 38220 37044
rect 38276 36988 40012 37044
rect 40068 36988 40078 37044
rect 40562 36988 40572 37044
rect 40628 36988 41692 37044
rect 41748 36988 41758 37044
rect 45602 36988 45612 37044
rect 45668 36988 45678 37044
rect 52210 36988 52220 37044
rect 52276 36988 54124 37044
rect 54180 36988 54572 37044
rect 54628 36988 55244 37044
rect 55300 36988 55310 37044
rect 57586 36988 57596 37044
rect 57652 36988 58156 37044
rect 58212 36988 60000 37044
rect 0 36960 800 36988
rect 23100 36932 23156 36988
rect 59200 36960 60000 36988
rect 4834 36876 4844 36932
rect 4900 36876 6524 36932
rect 6580 36876 6590 36932
rect 23090 36876 23100 36932
rect 23156 36876 23166 36932
rect 45938 36876 45948 36932
rect 46004 36876 46956 36932
rect 47012 36876 49644 36932
rect 49700 36876 49710 36932
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 26534 36764 26572 36820
rect 26628 36764 26638 36820
rect 32946 36764 32956 36820
rect 33012 36764 34188 36820
rect 34244 36764 34254 36820
rect 6626 36652 6636 36708
rect 6692 36652 7420 36708
rect 7476 36652 7486 36708
rect 14690 36652 14700 36708
rect 14756 36652 17164 36708
rect 17220 36652 17230 36708
rect 18050 36652 18060 36708
rect 18116 36652 18508 36708
rect 18564 36652 18574 36708
rect 50530 36652 50540 36708
rect 50596 36652 53004 36708
rect 53060 36652 53070 36708
rect 2118 36540 2156 36596
rect 2212 36540 2222 36596
rect 12898 36540 12908 36596
rect 12964 36540 13804 36596
rect 13860 36540 13870 36596
rect 14466 36540 14476 36596
rect 14532 36540 15148 36596
rect 15204 36540 15820 36596
rect 15876 36540 15886 36596
rect 18722 36540 18732 36596
rect 18788 36540 19964 36596
rect 20020 36540 20030 36596
rect 33170 36540 33180 36596
rect 33236 36540 33852 36596
rect 33908 36540 34412 36596
rect 34468 36540 35756 36596
rect 35812 36540 35822 36596
rect 40002 36540 40012 36596
rect 40068 36540 43372 36596
rect 43428 36540 44044 36596
rect 44100 36540 45612 36596
rect 45668 36540 45678 36596
rect 1586 36428 1596 36484
rect 1652 36428 1662 36484
rect 8978 36428 8988 36484
rect 9044 36428 10220 36484
rect 10276 36428 11116 36484
rect 11172 36428 11182 36484
rect 11666 36428 11676 36484
rect 11732 36428 12348 36484
rect 12404 36428 12414 36484
rect 27346 36428 27356 36484
rect 27412 36428 27916 36484
rect 27972 36428 29372 36484
rect 29428 36428 29438 36484
rect 38210 36428 38220 36484
rect 38276 36428 39452 36484
rect 39508 36428 40236 36484
rect 40292 36428 41356 36484
rect 41412 36428 41422 36484
rect 51426 36428 51436 36484
rect 51492 36428 53228 36484
rect 53284 36428 53294 36484
rect 54450 36428 54460 36484
rect 54516 36428 55244 36484
rect 55300 36428 55310 36484
rect 0 36372 800 36400
rect 1596 36372 1652 36428
rect 0 36316 1652 36372
rect 2258 36316 2268 36372
rect 2324 36316 2716 36372
rect 2772 36316 2782 36372
rect 3332 36316 4620 36372
rect 4676 36316 4686 36372
rect 15250 36316 15260 36372
rect 15316 36316 16156 36372
rect 16212 36316 20188 36372
rect 20244 36316 20254 36372
rect 21644 36316 24108 36372
rect 24164 36316 24174 36372
rect 31602 36316 31612 36372
rect 31668 36316 32172 36372
rect 32228 36316 32238 36372
rect 0 36288 800 36316
rect 1810 36204 1820 36260
rect 1876 36204 2940 36260
rect 2996 36204 3006 36260
rect 3332 36148 3388 36316
rect 21644 36260 21700 36316
rect 6514 36204 6524 36260
rect 6580 36204 8204 36260
rect 8260 36204 8270 36260
rect 11778 36204 11788 36260
rect 11844 36204 17612 36260
rect 17668 36204 21644 36260
rect 21700 36204 21710 36260
rect 23090 36204 23100 36260
rect 23156 36204 27692 36260
rect 27748 36204 27758 36260
rect 28130 36204 28140 36260
rect 28196 36204 29148 36260
rect 29204 36204 29214 36260
rect 36306 36204 36316 36260
rect 36372 36204 38108 36260
rect 38164 36204 38668 36260
rect 38724 36204 38734 36260
rect 2146 36092 2156 36148
rect 2212 36092 2492 36148
rect 2548 36092 2558 36148
rect 2706 36092 2716 36148
rect 2772 36092 3388 36148
rect 3826 36092 3836 36148
rect 3892 36092 4284 36148
rect 4340 36092 4350 36148
rect 6962 36092 6972 36148
rect 7028 36092 7756 36148
rect 7812 36092 10724 36148
rect 10668 36036 10724 36092
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 50546 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50830 36092
rect 10658 35980 10668 36036
rect 10724 35980 10734 36036
rect 1698 35868 1708 35924
rect 1764 35868 2604 35924
rect 2660 35868 2670 35924
rect 5282 35868 5292 35924
rect 5348 35868 5964 35924
rect 6020 35868 7196 35924
rect 7252 35868 7262 35924
rect 8642 35868 8652 35924
rect 8708 35868 10892 35924
rect 10948 35868 12348 35924
rect 12404 35868 12414 35924
rect 37986 35868 37996 35924
rect 38052 35868 38332 35924
rect 38388 35868 39676 35924
rect 39732 35868 39742 35924
rect 40002 35868 40012 35924
rect 40068 35868 40684 35924
rect 40740 35868 40750 35924
rect 50372 35868 57820 35924
rect 57876 35868 57886 35924
rect 40012 35812 40068 35868
rect 1708 35756 5404 35812
rect 5460 35756 5470 35812
rect 13682 35756 13692 35812
rect 13748 35756 14476 35812
rect 14532 35756 14542 35812
rect 15474 35756 15484 35812
rect 15540 35756 17388 35812
rect 17444 35756 17454 35812
rect 18834 35756 18844 35812
rect 18900 35756 19180 35812
rect 19236 35756 19246 35812
rect 22978 35756 22988 35812
rect 23044 35756 23660 35812
rect 23716 35756 26124 35812
rect 26180 35756 30268 35812
rect 30324 35756 30334 35812
rect 37874 35756 37884 35812
rect 37940 35756 38220 35812
rect 38276 35756 38780 35812
rect 38836 35756 40068 35812
rect 44258 35756 44268 35812
rect 44324 35756 45276 35812
rect 45332 35756 45342 35812
rect 47282 35756 47292 35812
rect 47348 35756 49868 35812
rect 49924 35756 49934 35812
rect 0 35700 800 35728
rect 1708 35700 1764 35756
rect 50372 35700 50428 35868
rect 52322 35756 52332 35812
rect 52388 35756 55468 35812
rect 55524 35756 55534 35812
rect 57922 35756 57932 35812
rect 57988 35756 57998 35812
rect 0 35644 1764 35700
rect 2268 35644 5628 35700
rect 5684 35644 5694 35700
rect 7746 35644 7756 35700
rect 7812 35644 8652 35700
rect 8708 35644 9548 35700
rect 9604 35644 9614 35700
rect 12674 35644 12684 35700
rect 12740 35644 12908 35700
rect 12964 35644 12974 35700
rect 13794 35644 13804 35700
rect 13860 35644 15372 35700
rect 15428 35644 15438 35700
rect 17154 35644 17164 35700
rect 17220 35644 17948 35700
rect 18004 35644 18014 35700
rect 29586 35644 29596 35700
rect 29652 35644 36316 35700
rect 36372 35644 36382 35700
rect 37538 35644 37548 35700
rect 37604 35644 38556 35700
rect 38612 35644 38622 35700
rect 39890 35644 39900 35700
rect 39956 35644 41132 35700
rect 41188 35644 41198 35700
rect 41794 35644 41804 35700
rect 41860 35644 42700 35700
rect 42756 35644 42766 35700
rect 47170 35644 47180 35700
rect 47236 35644 50428 35700
rect 57932 35700 57988 35756
rect 59200 35700 60000 35728
rect 57932 35644 60000 35700
rect 0 35616 800 35644
rect 2268 35364 2324 35644
rect 59200 35616 60000 35644
rect 4946 35532 4956 35588
rect 5012 35532 6524 35588
rect 6580 35532 6590 35588
rect 17826 35532 17836 35588
rect 17892 35532 23436 35588
rect 23492 35532 23502 35588
rect 25330 35532 25340 35588
rect 25396 35532 25676 35588
rect 25732 35532 25742 35588
rect 27234 35532 27244 35588
rect 27300 35532 28252 35588
rect 28308 35532 29372 35588
rect 29428 35532 29438 35588
rect 34626 35532 34636 35588
rect 34692 35532 38220 35588
rect 38276 35532 38286 35588
rect 38612 35532 55580 35588
rect 55636 35532 55646 35588
rect 38612 35476 38668 35532
rect 3238 35420 3276 35476
rect 3332 35420 3342 35476
rect 4386 35420 4396 35476
rect 4452 35420 6860 35476
rect 6916 35420 7980 35476
rect 8036 35420 8988 35476
rect 9044 35420 9772 35476
rect 9828 35420 9838 35476
rect 26898 35420 26908 35476
rect 26964 35420 29484 35476
rect 29540 35420 29550 35476
rect 34850 35420 34860 35476
rect 34916 35420 36428 35476
rect 36484 35420 36494 35476
rect 37090 35420 37100 35476
rect 37156 35420 37660 35476
rect 37716 35420 38668 35476
rect 49634 35420 49644 35476
rect 49700 35420 51996 35476
rect 52052 35420 52062 35476
rect 27244 35364 27300 35420
rect 1698 35308 1708 35364
rect 1764 35308 2268 35364
rect 2324 35308 2334 35364
rect 2594 35308 2604 35364
rect 2660 35308 4284 35364
rect 4340 35308 4350 35364
rect 4844 35308 6076 35364
rect 6132 35308 9660 35364
rect 9716 35308 9726 35364
rect 27234 35308 27244 35364
rect 27300 35308 27310 35364
rect 27906 35308 27916 35364
rect 27972 35308 28364 35364
rect 28420 35308 28430 35364
rect 33282 35308 33292 35364
rect 33348 35308 33358 35364
rect 48066 35308 48076 35364
rect 48132 35308 48972 35364
rect 49028 35308 49038 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 1922 35196 1932 35252
rect 1988 35196 2156 35252
rect 2212 35196 2222 35252
rect 3490 35196 3500 35252
rect 3556 35196 4060 35252
rect 4116 35196 4126 35252
rect 4844 35140 4900 35308
rect 33292 35252 33348 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 24546 35196 24556 35252
rect 24612 35196 25788 35252
rect 25844 35196 27132 35252
rect 27188 35196 27198 35252
rect 31938 35196 31948 35252
rect 32004 35196 33348 35252
rect 33292 35140 33348 35196
rect 38612 35196 39676 35252
rect 39732 35196 39742 35252
rect 43586 35196 43596 35252
rect 43652 35196 45276 35252
rect 45332 35196 45724 35252
rect 45780 35196 47068 35252
rect 47124 35196 47134 35252
rect 38612 35140 38668 35196
rect 2034 35084 2044 35140
rect 2100 35084 2604 35140
rect 2660 35084 2670 35140
rect 3332 35084 4900 35140
rect 7298 35084 7308 35140
rect 7364 35084 7980 35140
rect 8036 35084 8046 35140
rect 17714 35084 17724 35140
rect 17780 35084 19068 35140
rect 19124 35084 19134 35140
rect 25666 35084 25676 35140
rect 25732 35084 26012 35140
rect 26068 35084 26078 35140
rect 27346 35084 27356 35140
rect 27412 35084 28476 35140
rect 28532 35084 29260 35140
rect 29316 35084 29708 35140
rect 29764 35084 29774 35140
rect 33292 35084 37212 35140
rect 37268 35084 37278 35140
rect 38098 35084 38108 35140
rect 38164 35084 38668 35140
rect 39106 35084 39116 35140
rect 39172 35084 39182 35140
rect 0 35028 800 35056
rect 3332 35028 3388 35084
rect 39116 35028 39172 35084
rect 59200 35028 60000 35056
rect 0 34972 3388 35028
rect 3826 34972 3836 35028
rect 3892 34972 4508 35028
rect 4564 34972 4574 35028
rect 11330 34972 11340 35028
rect 11396 34972 13580 35028
rect 13636 34972 13646 35028
rect 15026 34972 15036 35028
rect 15092 34972 16156 35028
rect 16212 34972 16222 35028
rect 19282 34972 19292 35028
rect 19348 34972 20188 35028
rect 20244 34972 20254 35028
rect 20402 34972 20412 35028
rect 20468 34972 21868 35028
rect 21924 34972 30380 35028
rect 30436 34972 31052 35028
rect 31108 34972 31118 35028
rect 37762 34972 37772 35028
rect 37828 34972 38444 35028
rect 38500 34972 39172 35028
rect 39442 34972 39452 35028
rect 39508 34972 40012 35028
rect 40068 34972 41132 35028
rect 41188 34972 41804 35028
rect 41860 34972 47180 35028
rect 47236 34972 47246 35028
rect 49858 34972 49868 35028
rect 49924 34972 52108 35028
rect 52164 34972 52668 35028
rect 52724 34972 52734 35028
rect 58146 34972 58156 35028
rect 58212 34972 60000 35028
rect 0 34944 800 34972
rect 59200 34944 60000 34972
rect 3266 34860 3276 34916
rect 3332 34860 5068 34916
rect 5124 34860 5134 34916
rect 6962 34860 6972 34916
rect 7028 34860 10332 34916
rect 10388 34860 10556 34916
rect 10612 34860 10622 34916
rect 11442 34860 11452 34916
rect 11508 34860 14140 34916
rect 14196 34860 15148 34916
rect 15204 34860 15214 34916
rect 16034 34860 16044 34916
rect 16100 34860 17164 34916
rect 17220 34860 17230 34916
rect 17490 34860 17500 34916
rect 17556 34860 23996 34916
rect 24052 34860 24062 34916
rect 43026 34860 43036 34916
rect 43092 34860 43820 34916
rect 43876 34860 43886 34916
rect 44034 34860 44044 34916
rect 44100 34860 45724 34916
rect 45780 34860 48524 34916
rect 48580 34860 49084 34916
rect 49140 34860 49150 34916
rect 49970 34860 49980 34916
rect 50036 34860 51884 34916
rect 51940 34860 52780 34916
rect 52836 34860 52846 34916
rect 53442 34860 53452 34916
rect 53508 34860 53900 34916
rect 53956 34860 53966 34916
rect 17500 34804 17556 34860
rect 1362 34748 1372 34804
rect 1428 34748 6300 34804
rect 6356 34748 6366 34804
rect 7746 34748 7756 34804
rect 7812 34748 9212 34804
rect 9268 34748 9278 34804
rect 10658 34748 10668 34804
rect 10724 34748 12796 34804
rect 12852 34748 12862 34804
rect 13010 34748 13020 34804
rect 13076 34748 13916 34804
rect 13972 34748 13982 34804
rect 16370 34748 16380 34804
rect 16436 34748 17556 34804
rect 26226 34748 26236 34804
rect 26292 34748 27244 34804
rect 27300 34748 27310 34804
rect 27906 34748 27916 34804
rect 27972 34748 29372 34804
rect 29428 34748 29438 34804
rect 30594 34748 30604 34804
rect 30660 34748 32060 34804
rect 32116 34748 32126 34804
rect 33842 34748 33852 34804
rect 33908 34748 35196 34804
rect 35252 34748 35262 34804
rect 4050 34636 4060 34692
rect 4116 34636 5852 34692
rect 5908 34636 6188 34692
rect 6244 34636 6254 34692
rect 8642 34636 8652 34692
rect 8708 34636 10108 34692
rect 10164 34636 10174 34692
rect 24434 34636 24444 34692
rect 24500 34636 25676 34692
rect 25732 34636 25742 34692
rect 26674 34636 26684 34692
rect 26740 34636 28140 34692
rect 28196 34636 28206 34692
rect 33282 34636 33292 34692
rect 33348 34636 34972 34692
rect 35028 34636 35038 34692
rect 35970 34636 35980 34692
rect 36036 34636 36876 34692
rect 36932 34636 36942 34692
rect 41570 34636 41580 34692
rect 41636 34636 43932 34692
rect 43988 34636 45388 34692
rect 45444 34636 46284 34692
rect 46340 34636 46350 34692
rect 46498 34636 46508 34692
rect 46564 34636 47516 34692
rect 47572 34636 47582 34692
rect 49298 34636 49308 34692
rect 49364 34636 49868 34692
rect 49924 34636 49934 34692
rect 53106 34636 53116 34692
rect 53172 34636 53676 34692
rect 53732 34636 53742 34692
rect 39666 34524 39676 34580
rect 39732 34524 42588 34580
rect 42644 34524 42654 34580
rect 46610 34524 46620 34580
rect 46676 34524 48412 34580
rect 48468 34524 49756 34580
rect 49812 34524 49822 34580
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 50546 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50830 34524
rect 1474 34412 1484 34468
rect 1540 34412 17276 34468
rect 17332 34412 17342 34468
rect 0 34356 800 34384
rect 0 34300 4956 34356
rect 5012 34300 5022 34356
rect 7186 34300 7196 34356
rect 7252 34300 7644 34356
rect 7700 34300 7710 34356
rect 14466 34300 14476 34356
rect 14532 34300 15596 34356
rect 15652 34300 15662 34356
rect 16930 34300 16940 34356
rect 16996 34300 21756 34356
rect 21812 34300 21822 34356
rect 24322 34300 24332 34356
rect 24388 34300 26012 34356
rect 26068 34300 26078 34356
rect 32162 34300 32172 34356
rect 32228 34300 32956 34356
rect 33012 34300 33022 34356
rect 35410 34300 35420 34356
rect 35476 34300 43484 34356
rect 43540 34300 43550 34356
rect 45154 34300 45164 34356
rect 45220 34300 45612 34356
rect 45668 34300 49308 34356
rect 49364 34300 49374 34356
rect 0 34272 800 34300
rect 45164 34244 45220 34300
rect 3686 34188 3724 34244
rect 3780 34188 3790 34244
rect 9986 34188 9996 34244
rect 10052 34188 10556 34244
rect 10612 34188 10622 34244
rect 13906 34188 13916 34244
rect 13972 34188 15708 34244
rect 15764 34188 15774 34244
rect 19730 34188 19740 34244
rect 19796 34188 20860 34244
rect 20916 34188 20926 34244
rect 31602 34188 31612 34244
rect 31668 34188 33516 34244
rect 33572 34188 33582 34244
rect 33730 34188 33740 34244
rect 33796 34188 37660 34244
rect 37716 34188 37726 34244
rect 38210 34188 38220 34244
rect 38276 34188 38556 34244
rect 38612 34188 40236 34244
rect 40292 34188 41132 34244
rect 41188 34188 41198 34244
rect 42130 34188 42140 34244
rect 42196 34188 42812 34244
rect 42868 34188 42878 34244
rect 43026 34188 43036 34244
rect 43092 34188 45220 34244
rect 50306 34188 50316 34244
rect 50372 34188 51324 34244
rect 51380 34188 51996 34244
rect 52052 34188 52062 34244
rect 52658 34188 52668 34244
rect 52724 34188 53340 34244
rect 53396 34188 53406 34244
rect 1698 34076 1708 34132
rect 1764 34076 3948 34132
rect 4004 34076 4732 34132
rect 4788 34076 4798 34132
rect 8418 34076 8428 34132
rect 8484 34076 9884 34132
rect 9940 34076 11340 34132
rect 11396 34076 11406 34132
rect 20402 34076 20412 34132
rect 20468 34076 21420 34132
rect 21476 34076 23548 34132
rect 23604 34076 24556 34132
rect 24612 34076 25004 34132
rect 25060 34076 25070 34132
rect 31266 34076 31276 34132
rect 31332 34076 32172 34132
rect 32228 34076 32238 34132
rect 2034 33964 2044 34020
rect 2100 33964 5404 34020
rect 5460 33964 5470 34020
rect 9202 33964 9212 34020
rect 9268 33964 11564 34020
rect 11620 33964 11630 34020
rect 17602 33964 17612 34020
rect 17668 33964 19180 34020
rect 19236 33964 19852 34020
rect 19908 33964 19918 34020
rect 23874 33964 23884 34020
rect 23940 33964 25116 34020
rect 25172 33964 25182 34020
rect 32396 33908 32452 34188
rect 32582 34076 32620 34132
rect 32676 34076 32686 34132
rect 41010 34076 41020 34132
rect 41076 34076 41804 34132
rect 41860 34076 41870 34132
rect 42140 34020 42196 34188
rect 44146 34076 44156 34132
rect 44212 34076 44716 34132
rect 44772 34076 45948 34132
rect 46004 34076 46014 34132
rect 49858 34076 49868 34132
rect 49924 34076 50652 34132
rect 50708 34076 52444 34132
rect 52500 34076 52510 34132
rect 33282 33964 33292 34020
rect 33348 33964 39228 34020
rect 39284 33964 39294 34020
rect 40114 33964 40124 34020
rect 40180 33964 42196 34020
rect 43698 33964 43708 34020
rect 43764 33964 44268 34020
rect 44324 33964 44334 34020
rect 1922 33852 1932 33908
rect 1988 33852 1998 33908
rect 3490 33852 3500 33908
rect 3556 33852 3836 33908
rect 3892 33852 3902 33908
rect 4274 33852 4284 33908
rect 4340 33852 9324 33908
rect 9380 33852 9390 33908
rect 26898 33852 26908 33908
rect 26964 33852 31948 33908
rect 32004 33852 32014 33908
rect 32386 33852 32396 33908
rect 32452 33852 32462 33908
rect 0 33684 800 33712
rect 1932 33684 1988 33852
rect 23090 33740 23100 33796
rect 23156 33740 27020 33796
rect 27076 33740 27086 33796
rect 31378 33740 31388 33796
rect 31444 33740 34300 33796
rect 34356 33740 34366 33796
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 0 33628 1988 33684
rect 19506 33628 19516 33684
rect 19572 33628 21084 33684
rect 21140 33628 21150 33684
rect 23202 33628 23212 33684
rect 23268 33628 24668 33684
rect 24724 33628 24734 33684
rect 25442 33628 25452 33684
rect 25508 33628 31948 33684
rect 32004 33628 32014 33684
rect 36642 33628 36652 33684
rect 36708 33628 37212 33684
rect 37268 33628 37996 33684
rect 38052 33628 38062 33684
rect 51538 33628 51548 33684
rect 51604 33628 53004 33684
rect 53060 33628 54124 33684
rect 54180 33628 57148 33684
rect 57204 33628 57214 33684
rect 0 33600 800 33628
rect 3686 33516 3724 33572
rect 3780 33516 3790 33572
rect 5282 33516 5292 33572
rect 5348 33516 6076 33572
rect 6132 33516 6142 33572
rect 9314 33516 9324 33572
rect 9380 33516 21532 33572
rect 21588 33516 21598 33572
rect 35634 33516 35644 33572
rect 35700 33516 37100 33572
rect 37156 33516 37166 33572
rect 40114 33516 40124 33572
rect 40180 33516 41020 33572
rect 41076 33516 41086 33572
rect 41794 33516 41804 33572
rect 41860 33516 43932 33572
rect 43988 33516 43998 33572
rect 6178 33404 6188 33460
rect 6244 33404 8428 33460
rect 8484 33404 8494 33460
rect 9090 33404 9100 33460
rect 9156 33404 9996 33460
rect 10052 33404 10062 33460
rect 10658 33404 10668 33460
rect 10724 33404 11788 33460
rect 11844 33404 11854 33460
rect 12786 33404 12796 33460
rect 12852 33404 14476 33460
rect 14532 33404 14542 33460
rect 17714 33404 17724 33460
rect 17780 33404 20076 33460
rect 20132 33404 21420 33460
rect 21476 33404 21486 33460
rect 27794 33404 27804 33460
rect 27860 33404 29036 33460
rect 29092 33404 29102 33460
rect 30146 33404 30156 33460
rect 30212 33404 34412 33460
rect 34468 33404 34478 33460
rect 2706 33292 2716 33348
rect 2772 33292 5964 33348
rect 6020 33292 6748 33348
rect 6804 33292 6814 33348
rect 7634 33292 7644 33348
rect 7700 33292 9548 33348
rect 9604 33292 9614 33348
rect 21746 33292 21756 33348
rect 21812 33292 22988 33348
rect 23044 33292 23054 33348
rect 35746 33292 35756 33348
rect 35812 33292 38556 33348
rect 38612 33292 38622 33348
rect 41906 33292 41916 33348
rect 41972 33292 42700 33348
rect 42756 33292 42766 33348
rect 53666 33292 53676 33348
rect 53732 33292 54572 33348
rect 54628 33292 54638 33348
rect 5842 33180 5852 33236
rect 5908 33180 7756 33236
rect 7812 33180 7822 33236
rect 20626 33180 20636 33236
rect 20692 33180 20860 33236
rect 20916 33180 22876 33236
rect 22932 33180 22942 33236
rect 25218 33180 25228 33236
rect 25284 33180 30156 33236
rect 30212 33180 31164 33236
rect 31220 33180 31230 33236
rect 35858 33180 35868 33236
rect 35924 33180 36540 33236
rect 36596 33180 36606 33236
rect 38322 33180 38332 33236
rect 38388 33180 40292 33236
rect 40450 33180 40460 33236
rect 40516 33180 44828 33236
rect 44884 33180 46060 33236
rect 46116 33180 46126 33236
rect 49522 33180 49532 33236
rect 49588 33180 50764 33236
rect 50820 33180 50830 33236
rect 52322 33180 52332 33236
rect 52388 33180 53564 33236
rect 53620 33180 53630 33236
rect 25228 33124 25284 33180
rect 1698 33068 1708 33124
rect 1764 33068 2492 33124
rect 2548 33068 2558 33124
rect 17826 33068 17836 33124
rect 17892 33068 18732 33124
rect 18788 33068 25284 33124
rect 25666 33068 25676 33124
rect 25732 33068 28028 33124
rect 28084 33068 28094 33124
rect 31910 33068 31948 33124
rect 32004 33068 32014 33124
rect 32722 33068 32732 33124
rect 32788 33068 33964 33124
rect 34020 33068 34030 33124
rect 34962 33068 34972 33124
rect 35028 33068 35308 33124
rect 35746 33068 35756 33124
rect 35812 33068 36428 33124
rect 36484 33068 36494 33124
rect 0 33012 800 33040
rect 35252 33012 35308 33068
rect 40236 33012 40292 33180
rect 46610 33068 46620 33124
rect 46676 33068 49308 33124
rect 49364 33068 49374 33124
rect 51650 33068 51660 33124
rect 51716 33068 53228 33124
rect 53284 33068 57260 33124
rect 57316 33068 57326 33124
rect 0 32956 1820 33012
rect 1876 32956 1886 33012
rect 6178 32956 6188 33012
rect 6244 32956 7308 33012
rect 7364 32956 8092 33012
rect 8148 32956 17388 33012
rect 17444 32956 17454 33012
rect 23986 32956 23996 33012
rect 24052 32956 25452 33012
rect 25508 32956 25518 33012
rect 26562 32956 26572 33012
rect 26628 32956 27244 33012
rect 27300 32956 27310 33012
rect 35252 32956 35868 33012
rect 35924 32956 35934 33012
rect 40236 32956 49364 33012
rect 0 32928 800 32956
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 49308 32900 49364 32956
rect 50546 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50830 32956
rect 20188 32844 26684 32900
rect 26740 32844 29708 32900
rect 29764 32844 30492 32900
rect 30548 32844 30558 32900
rect 37314 32844 37324 32900
rect 37380 32844 43932 32900
rect 43988 32844 45276 32900
rect 45332 32844 45342 32900
rect 49298 32844 49308 32900
rect 49364 32844 49374 32900
rect 20188 32788 20244 32844
rect 3266 32732 3276 32788
rect 3332 32732 4956 32788
rect 5012 32732 5022 32788
rect 5506 32732 5516 32788
rect 5572 32732 7420 32788
rect 7476 32732 7486 32788
rect 7858 32732 7868 32788
rect 7924 32732 9660 32788
rect 9716 32732 11732 32788
rect 19170 32732 19180 32788
rect 19236 32732 20244 32788
rect 23426 32732 23436 32788
rect 23492 32732 27468 32788
rect 27524 32732 27534 32788
rect 28466 32732 28476 32788
rect 28532 32732 29820 32788
rect 29876 32732 33068 32788
rect 33124 32732 33134 32788
rect 38882 32732 38892 32788
rect 38948 32732 40684 32788
rect 40740 32732 40750 32788
rect 42690 32732 42700 32788
rect 42756 32732 55580 32788
rect 55636 32732 55646 32788
rect 11676 32676 11732 32732
rect 2482 32620 2492 32676
rect 2548 32620 5292 32676
rect 5348 32620 5358 32676
rect 7634 32620 7644 32676
rect 7700 32620 10108 32676
rect 10164 32620 10174 32676
rect 11666 32620 11676 32676
rect 11732 32620 14924 32676
rect 14980 32620 14990 32676
rect 22764 32620 25340 32676
rect 25396 32620 25406 32676
rect 32162 32620 32172 32676
rect 32228 32620 32508 32676
rect 32564 32620 38556 32676
rect 38612 32620 38622 32676
rect 42914 32620 42924 32676
rect 42980 32620 43820 32676
rect 43876 32620 43886 32676
rect 46722 32620 46732 32676
rect 46788 32620 50428 32676
rect 53218 32620 53228 32676
rect 53284 32620 54684 32676
rect 54740 32620 54750 32676
rect 8530 32508 8540 32564
rect 8596 32508 10220 32564
rect 10276 32508 13468 32564
rect 13524 32508 13534 32564
rect 22764 32452 22820 32620
rect 50372 32564 50428 32620
rect 45042 32508 45052 32564
rect 45108 32508 45836 32564
rect 45892 32508 45902 32564
rect 50372 32508 52108 32564
rect 52164 32508 52174 32564
rect 53442 32508 53452 32564
rect 53508 32508 54124 32564
rect 54180 32508 56588 32564
rect 56644 32508 56654 32564
rect 21746 32396 21756 32452
rect 21812 32396 22764 32452
rect 22820 32396 22830 32452
rect 29810 32396 29820 32452
rect 29876 32396 31500 32452
rect 31556 32396 31566 32452
rect 34850 32396 34860 32452
rect 34916 32396 35196 32452
rect 35252 32396 35262 32452
rect 0 32340 800 32368
rect 59200 32340 60000 32368
rect 0 32284 6188 32340
rect 6244 32284 8876 32340
rect 8932 32284 8942 32340
rect 57922 32284 57932 32340
rect 57988 32284 60000 32340
rect 0 32256 800 32284
rect 59200 32256 60000 32284
rect 27906 32172 27916 32228
rect 27972 32172 29036 32228
rect 29092 32172 29596 32228
rect 29652 32172 29662 32228
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 26562 32060 26572 32116
rect 26628 32060 33012 32116
rect 32956 32004 33012 32060
rect 4722 31948 4732 32004
rect 4788 31948 7868 32004
rect 7924 31948 7934 32004
rect 13906 31948 13916 32004
rect 13972 31948 15260 32004
rect 15316 31948 15326 32004
rect 24210 31948 24220 32004
rect 24276 31948 25116 32004
rect 25172 31948 25182 32004
rect 27682 31948 27692 32004
rect 27748 31948 30156 32004
rect 30212 31948 30716 32004
rect 30772 31948 30782 32004
rect 32946 31948 32956 32004
rect 33012 31948 33022 32004
rect 35298 31948 35308 32004
rect 35364 31948 42028 32004
rect 42084 31948 42094 32004
rect 45490 31948 45500 32004
rect 45556 31948 46620 32004
rect 46676 31948 46686 32004
rect 52322 31948 52332 32004
rect 52388 31948 52780 32004
rect 52836 31948 52846 32004
rect 2370 31836 2380 31892
rect 2436 31836 4060 31892
rect 4116 31836 4956 31892
rect 5012 31836 5628 31892
rect 5684 31836 5694 31892
rect 6850 31836 6860 31892
rect 6916 31836 8652 31892
rect 8708 31836 10332 31892
rect 10388 31836 10398 31892
rect 12002 31836 12012 31892
rect 12068 31836 13692 31892
rect 13748 31836 14588 31892
rect 14644 31836 14654 31892
rect 16370 31836 16380 31892
rect 16436 31836 17500 31892
rect 17556 31836 17566 31892
rect 22194 31836 22204 31892
rect 22260 31836 25228 31892
rect 25284 31836 25294 31892
rect 28018 31836 28028 31892
rect 28084 31836 28476 31892
rect 28532 31836 29820 31892
rect 29876 31836 29886 31892
rect 31826 31836 31836 31892
rect 31892 31836 34188 31892
rect 34244 31836 34254 31892
rect 34514 31836 34524 31892
rect 34580 31836 35532 31892
rect 35588 31836 35598 31892
rect 47954 31836 47964 31892
rect 48020 31836 48300 31892
rect 48356 31836 51548 31892
rect 51604 31836 51614 31892
rect 51986 31836 51996 31892
rect 52052 31836 54124 31892
rect 54180 31836 54684 31892
rect 54740 31836 54750 31892
rect 1250 31724 1260 31780
rect 1316 31724 4620 31780
rect 4676 31724 4686 31780
rect 6514 31724 6524 31780
rect 6580 31724 8540 31780
rect 8596 31724 10108 31780
rect 10164 31724 10174 31780
rect 14242 31724 14252 31780
rect 14308 31724 16156 31780
rect 16212 31724 16222 31780
rect 16594 31724 16604 31780
rect 16660 31724 16670 31780
rect 16930 31724 16940 31780
rect 16996 31724 19180 31780
rect 19236 31724 19246 31780
rect 22978 31724 22988 31780
rect 23044 31724 25564 31780
rect 25620 31724 26012 31780
rect 26068 31724 26078 31780
rect 28354 31724 28364 31780
rect 28420 31724 29372 31780
rect 29428 31724 29438 31780
rect 33170 31724 33180 31780
rect 33236 31724 33852 31780
rect 33908 31724 33918 31780
rect 34066 31724 34076 31780
rect 34132 31724 36428 31780
rect 36484 31724 36494 31780
rect 37090 31724 37100 31780
rect 37156 31724 38332 31780
rect 38388 31724 39564 31780
rect 39620 31724 40348 31780
rect 40404 31724 40414 31780
rect 45164 31724 49084 31780
rect 49140 31724 49150 31780
rect 49746 31724 49756 31780
rect 49812 31724 55580 31780
rect 55636 31724 55646 31780
rect 0 31668 800 31696
rect 16604 31668 16660 31724
rect 22988 31668 23044 31724
rect 45164 31668 45220 31724
rect 59200 31668 60000 31696
rect 0 31612 3612 31668
rect 3668 31612 3678 31668
rect 4274 31612 4284 31668
rect 4340 31612 9604 31668
rect 14802 31612 14812 31668
rect 14868 31612 16660 31668
rect 18162 31612 18172 31668
rect 18228 31612 18732 31668
rect 18788 31612 23044 31668
rect 27346 31612 27356 31668
rect 27412 31612 28252 31668
rect 28308 31612 28318 31668
rect 33506 31612 33516 31668
rect 33572 31612 45164 31668
rect 45220 31612 45230 31668
rect 46050 31612 46060 31668
rect 46116 31612 47068 31668
rect 47124 31612 52556 31668
rect 52612 31612 52622 31668
rect 57922 31612 57932 31668
rect 57988 31612 60000 31668
rect 0 31584 800 31612
rect 3042 31500 3052 31556
rect 3108 31500 3500 31556
rect 3556 31500 6524 31556
rect 6580 31500 6590 31556
rect 7298 31500 7308 31556
rect 7364 31500 7374 31556
rect 4162 31388 4172 31444
rect 4228 31388 7084 31444
rect 7140 31388 7150 31444
rect 7308 31332 7364 31500
rect 9548 31444 9604 31612
rect 27356 31556 27412 31612
rect 59200 31584 60000 31612
rect 10210 31500 10220 31556
rect 10276 31500 21084 31556
rect 21140 31500 21150 31556
rect 23650 31500 23660 31556
rect 23716 31500 27020 31556
rect 27076 31500 27412 31556
rect 34066 31500 34076 31556
rect 34132 31500 38668 31556
rect 46834 31500 46844 31556
rect 46900 31500 47628 31556
rect 47684 31500 47694 31556
rect 50194 31500 50204 31556
rect 50260 31500 52892 31556
rect 52948 31500 52958 31556
rect 9548 31388 17388 31444
rect 17444 31388 17454 31444
rect 20738 31388 20748 31444
rect 20804 31388 21308 31444
rect 21364 31388 21374 31444
rect 23314 31388 23324 31444
rect 23380 31388 24444 31444
rect 24500 31388 24510 31444
rect 24770 31388 24780 31444
rect 24836 31388 26012 31444
rect 26068 31388 26078 31444
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 38612 31332 38668 31500
rect 39218 31388 39228 31444
rect 39284 31388 39900 31444
rect 39956 31388 49756 31444
rect 49812 31388 49822 31444
rect 50546 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50830 31388
rect 2706 31276 2716 31332
rect 2772 31276 7364 31332
rect 17042 31276 17052 31332
rect 17108 31276 17948 31332
rect 18004 31276 18014 31332
rect 21186 31276 21196 31332
rect 21252 31276 25452 31332
rect 25508 31276 25518 31332
rect 34290 31276 34300 31332
rect 34356 31276 35980 31332
rect 36036 31276 36428 31332
rect 36484 31276 36494 31332
rect 38612 31276 44940 31332
rect 44996 31276 45006 31332
rect 4946 31164 4956 31220
rect 5012 31164 5852 31220
rect 5908 31164 6636 31220
rect 6692 31164 7140 31220
rect 9426 31164 9436 31220
rect 9492 31164 11452 31220
rect 11508 31164 20636 31220
rect 20692 31164 20702 31220
rect 22306 31164 22316 31220
rect 22372 31164 25228 31220
rect 25284 31164 27468 31220
rect 27524 31164 27534 31220
rect 31490 31164 31500 31220
rect 31556 31164 33292 31220
rect 33348 31164 36484 31220
rect 37762 31164 37772 31220
rect 37828 31164 38332 31220
rect 38388 31164 38398 31220
rect 48738 31164 48748 31220
rect 48804 31164 49532 31220
rect 49588 31164 49598 31220
rect 52434 31164 52444 31220
rect 52500 31164 53676 31220
rect 53732 31164 54348 31220
rect 54404 31164 54414 31220
rect 7084 31108 7140 31164
rect 3714 31052 3724 31108
rect 3780 31052 6076 31108
rect 6132 31052 6412 31108
rect 6468 31052 6748 31108
rect 6804 31052 6814 31108
rect 7074 31052 7084 31108
rect 7140 31052 8148 31108
rect 8866 31052 8876 31108
rect 8932 31052 10220 31108
rect 10276 31052 10286 31108
rect 12450 31052 12460 31108
rect 12516 31052 17724 31108
rect 17780 31052 17790 31108
rect 17938 31052 17948 31108
rect 18004 31052 21756 31108
rect 21812 31052 21822 31108
rect 24546 31052 24556 31108
rect 24612 31052 25340 31108
rect 25396 31052 25406 31108
rect 26002 31052 26012 31108
rect 26068 31052 26572 31108
rect 26628 31052 26638 31108
rect 32386 31052 32396 31108
rect 32452 31052 34188 31108
rect 34244 31052 34254 31108
rect 35186 31052 35196 31108
rect 35252 31052 35532 31108
rect 35588 31052 36204 31108
rect 36260 31052 36270 31108
rect 0 30996 800 31024
rect 8092 30996 8148 31052
rect 0 30940 1932 30996
rect 1988 30940 1998 30996
rect 6514 30940 6524 30996
rect 6580 30940 7532 30996
rect 7588 30940 7868 30996
rect 7924 30940 7934 30996
rect 8092 30940 11788 30996
rect 11844 30940 11854 30996
rect 16594 30940 16604 30996
rect 16660 30940 20188 30996
rect 20244 30940 22988 30996
rect 23044 30940 23054 30996
rect 24658 30940 24668 30996
rect 24724 30940 27244 30996
rect 27300 30940 27310 30996
rect 30706 30940 30716 30996
rect 30772 30940 33852 30996
rect 33908 30940 34076 30996
rect 34132 30940 34142 30996
rect 0 30912 800 30940
rect 3266 30828 3276 30884
rect 3332 30828 5404 30884
rect 5460 30828 5470 30884
rect 13234 30828 13244 30884
rect 13300 30828 15260 30884
rect 15316 30828 15326 30884
rect 20066 30828 20076 30884
rect 20132 30828 22204 30884
rect 22260 30828 22270 30884
rect 26786 30828 26796 30884
rect 26852 30828 31836 30884
rect 31892 30828 34748 30884
rect 34804 30828 34814 30884
rect 16594 30716 16604 30772
rect 16660 30716 17836 30772
rect 17892 30716 17902 30772
rect 20738 30716 20748 30772
rect 20804 30716 31500 30772
rect 31556 30716 31566 30772
rect 33842 30716 33852 30772
rect 33908 30716 35308 30772
rect 35364 30716 35374 30772
rect 36428 30660 36484 31164
rect 42466 31052 42476 31108
rect 42532 31052 43596 31108
rect 43652 31052 44492 31108
rect 44548 31052 44558 31108
rect 49858 31052 49868 31108
rect 49924 31052 51100 31108
rect 51156 31052 51166 31108
rect 51874 31052 51884 31108
rect 51940 31052 54180 31108
rect 54124 30996 54180 31052
rect 59200 30996 60000 31024
rect 36978 30940 36988 30996
rect 37044 30940 37324 30996
rect 37380 30940 37390 30996
rect 38434 30940 38444 30996
rect 38500 30940 39116 30996
rect 39172 30940 39182 30996
rect 50978 30940 50988 30996
rect 51044 30940 51660 30996
rect 51716 30940 53004 30996
rect 53060 30940 53070 30996
rect 54114 30940 54124 30996
rect 54180 30940 56700 30996
rect 56756 30940 56766 30996
rect 57810 30940 57820 30996
rect 57876 30940 60000 30996
rect 37324 30884 37380 30940
rect 59200 30912 60000 30940
rect 37324 30828 39676 30884
rect 39732 30828 39742 30884
rect 46274 30828 46284 30884
rect 46340 30828 47180 30884
rect 47236 30828 47246 30884
rect 37650 30716 37660 30772
rect 37716 30716 38668 30772
rect 42802 30716 42812 30772
rect 42868 30716 45276 30772
rect 45332 30716 45342 30772
rect 45602 30716 45612 30772
rect 45668 30716 46396 30772
rect 46452 30716 46462 30772
rect 46610 30716 46620 30772
rect 46676 30716 47740 30772
rect 47796 30716 52556 30772
rect 52612 30716 52622 30772
rect 53330 30716 53340 30772
rect 53396 30716 55020 30772
rect 55076 30716 55086 30772
rect 38612 30660 38668 30716
rect 2258 30604 2268 30660
rect 2324 30604 3388 30660
rect 3444 30604 3948 30660
rect 4004 30604 4014 30660
rect 36428 30604 38500 30660
rect 38612 30604 48972 30660
rect 49028 30604 49038 30660
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 38444 30548 38500 30604
rect 30818 30492 30828 30548
rect 30884 30492 31500 30548
rect 31556 30492 34244 30548
rect 36530 30492 36540 30548
rect 36596 30492 38220 30548
rect 38276 30492 38286 30548
rect 38444 30492 41020 30548
rect 41076 30492 41086 30548
rect 34188 30436 34244 30492
rect 15250 30380 15260 30436
rect 15316 30380 16044 30436
rect 16100 30380 16110 30436
rect 17378 30380 17388 30436
rect 17444 30380 19404 30436
rect 19460 30380 19470 30436
rect 27346 30380 27356 30436
rect 27412 30380 33964 30436
rect 34020 30380 34030 30436
rect 34188 30380 37212 30436
rect 37268 30380 37278 30436
rect 0 30324 800 30352
rect 0 30268 1708 30324
rect 1764 30268 1774 30324
rect 12450 30268 12460 30324
rect 12516 30268 13916 30324
rect 13972 30268 13982 30324
rect 14690 30268 14700 30324
rect 14756 30268 15372 30324
rect 15428 30268 15438 30324
rect 25778 30268 25788 30324
rect 25844 30268 30772 30324
rect 0 30240 800 30268
rect 8194 30156 8204 30212
rect 8260 30156 8988 30212
rect 9044 30156 9054 30212
rect 10098 30156 10108 30212
rect 10164 30156 11452 30212
rect 11508 30156 11518 30212
rect 14466 30156 14476 30212
rect 14532 30156 15708 30212
rect 15764 30156 15774 30212
rect 20850 30156 20860 30212
rect 20916 30156 21644 30212
rect 21700 30156 24220 30212
rect 24276 30156 24444 30212
rect 24500 30156 24510 30212
rect 26338 30156 26348 30212
rect 26404 30156 27692 30212
rect 27748 30156 27758 30212
rect 28578 30156 28588 30212
rect 28644 30156 30492 30212
rect 30548 30156 30558 30212
rect 30716 30100 30772 30268
rect 32508 30212 32564 30380
rect 37436 30324 37492 30492
rect 38546 30380 38556 30436
rect 38612 30380 40572 30436
rect 40628 30380 40638 30436
rect 37426 30268 37436 30324
rect 37492 30268 37502 30324
rect 37986 30268 37996 30324
rect 38052 30268 43932 30324
rect 43988 30268 43998 30324
rect 51202 30268 51212 30324
rect 51268 30268 52668 30324
rect 52724 30268 52734 30324
rect 32498 30156 32508 30212
rect 32564 30156 32574 30212
rect 35298 30156 35308 30212
rect 35364 30156 36316 30212
rect 36372 30156 38668 30212
rect 42242 30156 42252 30212
rect 42308 30156 43372 30212
rect 43428 30156 43438 30212
rect 44258 30156 44268 30212
rect 44324 30156 45164 30212
rect 45220 30156 46284 30212
rect 46340 30156 46350 30212
rect 38612 30100 38668 30156
rect 43372 30100 43428 30156
rect 8082 30044 8092 30100
rect 8148 30044 10668 30100
rect 10724 30044 10734 30100
rect 18274 30044 18284 30100
rect 18340 30044 19068 30100
rect 19124 30044 19134 30100
rect 25228 30044 27580 30100
rect 27636 30044 27646 30100
rect 28018 30044 28028 30100
rect 28084 30044 29148 30100
rect 29204 30044 29214 30100
rect 30716 30044 34356 30100
rect 34962 30044 34972 30100
rect 35028 30044 36652 30100
rect 36708 30044 36718 30100
rect 38612 30044 42924 30100
rect 42980 30044 42990 30100
rect 43372 30044 44604 30100
rect 44660 30044 44670 30100
rect 25228 29988 25284 30044
rect 34300 29988 34356 30044
rect 4274 29932 4284 29988
rect 4340 29932 13468 29988
rect 13524 29932 13534 29988
rect 20402 29932 20412 29988
rect 20468 29932 25228 29988
rect 25284 29932 25294 29988
rect 27458 29932 27468 29988
rect 27524 29932 28084 29988
rect 29474 29932 29484 29988
rect 29540 29932 30604 29988
rect 30660 29932 31612 29988
rect 31668 29932 31678 29988
rect 34290 29932 34300 29988
rect 34356 29932 34366 29988
rect 41570 29932 41580 29988
rect 41636 29932 43036 29988
rect 43092 29932 43102 29988
rect 44034 29932 44044 29988
rect 44100 29932 44716 29988
rect 44772 29932 46396 29988
rect 46452 29932 48972 29988
rect 49028 29932 49038 29988
rect 6514 29820 6524 29876
rect 6580 29820 7420 29876
rect 7476 29820 8316 29876
rect 8372 29820 8382 29876
rect 26852 29820 27804 29876
rect 27860 29820 27870 29876
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 2818 29708 2828 29764
rect 2884 29708 3388 29764
rect 7746 29708 7756 29764
rect 7812 29708 9660 29764
rect 9716 29708 9726 29764
rect 0 29652 800 29680
rect 3332 29652 3388 29708
rect 26852 29652 26908 29820
rect 28028 29764 28084 29932
rect 29138 29820 29148 29876
rect 29204 29820 30380 29876
rect 30436 29820 31276 29876
rect 31332 29820 31342 29876
rect 35252 29820 40348 29876
rect 40404 29820 41916 29876
rect 41972 29820 41982 29876
rect 43138 29820 43148 29876
rect 43204 29820 43214 29876
rect 45602 29820 45612 29876
rect 45668 29820 46172 29876
rect 46228 29820 47068 29876
rect 47124 29820 47134 29876
rect 35252 29764 35308 29820
rect 28028 29708 30156 29764
rect 30212 29708 30222 29764
rect 31154 29708 31164 29764
rect 31220 29708 34972 29764
rect 35028 29708 35308 29764
rect 43148 29764 43204 29820
rect 50546 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50830 29820
rect 43148 29708 50428 29764
rect 55570 29708 55580 29764
rect 55636 29708 55646 29764
rect 50372 29652 50428 29708
rect 55580 29652 55636 29708
rect 0 29596 2492 29652
rect 2548 29596 2558 29652
rect 3332 29596 20076 29652
rect 20132 29596 21532 29652
rect 21588 29596 21598 29652
rect 25442 29596 25452 29652
rect 25508 29596 26908 29652
rect 28690 29596 28700 29652
rect 28756 29596 30716 29652
rect 30772 29596 30782 29652
rect 31042 29596 31052 29652
rect 31108 29596 31948 29652
rect 32004 29596 32014 29652
rect 32274 29596 32284 29652
rect 32340 29596 33404 29652
rect 33460 29596 33470 29652
rect 40002 29596 40012 29652
rect 40068 29596 40796 29652
rect 40852 29596 40862 29652
rect 45042 29596 45052 29652
rect 45108 29596 45836 29652
rect 45892 29596 45902 29652
rect 50372 29596 55636 29652
rect 0 29568 800 29596
rect 31948 29540 32004 29596
rect 4274 29484 4284 29540
rect 4340 29484 15148 29540
rect 15204 29484 15214 29540
rect 16818 29484 16828 29540
rect 16884 29484 17948 29540
rect 18004 29484 20300 29540
rect 20356 29484 20366 29540
rect 20850 29484 20860 29540
rect 20916 29484 22204 29540
rect 22260 29484 23324 29540
rect 23380 29484 23390 29540
rect 26002 29484 26012 29540
rect 26068 29484 26796 29540
rect 26852 29484 27132 29540
rect 27188 29484 27198 29540
rect 27682 29484 27692 29540
rect 27748 29484 31164 29540
rect 31220 29484 31230 29540
rect 31948 29484 33964 29540
rect 34020 29484 35756 29540
rect 35812 29484 35822 29540
rect 37314 29484 37324 29540
rect 37380 29484 46620 29540
rect 46676 29484 46686 29540
rect 27132 29428 27188 29484
rect 2706 29372 2716 29428
rect 2772 29372 6860 29428
rect 6916 29372 6926 29428
rect 7522 29372 7532 29428
rect 7588 29372 8428 29428
rect 8484 29372 8494 29428
rect 14354 29372 14364 29428
rect 14420 29372 15596 29428
rect 15652 29372 15662 29428
rect 26562 29372 26572 29428
rect 26628 29372 27076 29428
rect 27132 29372 28028 29428
rect 28084 29372 28094 29428
rect 32834 29372 32844 29428
rect 32900 29372 36204 29428
rect 36260 29372 36484 29428
rect 36642 29372 36652 29428
rect 36708 29372 44492 29428
rect 44548 29372 44558 29428
rect 27020 29316 27076 29372
rect 36428 29316 36484 29372
rect 13458 29260 13468 29316
rect 13524 29260 15932 29316
rect 15988 29260 15998 29316
rect 26422 29260 26460 29316
rect 26516 29260 26526 29316
rect 27010 29260 27020 29316
rect 27076 29260 27580 29316
rect 27636 29260 28476 29316
rect 28532 29260 28542 29316
rect 33702 29260 33740 29316
rect 33796 29260 35980 29316
rect 36036 29260 36046 29316
rect 36428 29260 36988 29316
rect 37044 29260 37054 29316
rect 39890 29260 39900 29316
rect 39956 29260 40908 29316
rect 40964 29260 40974 29316
rect 1922 29148 1932 29204
rect 1988 29148 1998 29204
rect 6626 29148 6636 29204
rect 6692 29148 7868 29204
rect 7924 29148 8540 29204
rect 8596 29148 8606 29204
rect 9986 29148 9996 29204
rect 10052 29148 19628 29204
rect 19684 29148 21308 29204
rect 21364 29148 21374 29204
rect 34514 29148 34524 29204
rect 34580 29148 34860 29204
rect 34916 29148 36428 29204
rect 36484 29148 36494 29204
rect 0 28980 800 29008
rect 1932 28980 1988 29148
rect 20738 29036 20748 29092
rect 20804 29036 21420 29092
rect 21476 29036 25116 29092
rect 25172 29036 25182 29092
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 0 28924 1988 28980
rect 15138 28924 15148 28980
rect 15204 28924 17388 28980
rect 17444 28924 17454 28980
rect 25778 28924 25788 28980
rect 25844 28924 33292 28980
rect 33348 28924 33358 28980
rect 0 28896 800 28924
rect 1586 28812 1596 28868
rect 1652 28812 19068 28868
rect 19124 28812 19134 28868
rect 27654 28812 27692 28868
rect 27748 28812 27758 28868
rect 30594 28812 30604 28868
rect 30660 28812 33180 28868
rect 33236 28812 33246 28868
rect 35410 28812 35420 28868
rect 35476 28812 35980 28868
rect 36036 28812 49756 28868
rect 49812 28812 49822 28868
rect 14578 28700 14588 28756
rect 14644 28700 15596 28756
rect 15652 28700 15662 28756
rect 25666 28700 25676 28756
rect 25732 28700 31164 28756
rect 31220 28700 34748 28756
rect 34804 28700 34814 28756
rect 35186 28700 35196 28756
rect 35252 28700 38668 28756
rect 38882 28700 38892 28756
rect 38948 28700 39900 28756
rect 39956 28700 39966 28756
rect 47068 28700 55636 28756
rect 38612 28644 38668 28700
rect 2034 28588 2044 28644
rect 2100 28588 2716 28644
rect 2772 28588 2782 28644
rect 3378 28588 3388 28644
rect 3444 28588 6636 28644
rect 6692 28588 6702 28644
rect 16258 28588 16268 28644
rect 16324 28588 17052 28644
rect 17108 28588 17118 28644
rect 26338 28588 26348 28644
rect 26404 28588 26414 28644
rect 29474 28588 29484 28644
rect 29540 28588 30380 28644
rect 30436 28588 30828 28644
rect 30884 28588 31612 28644
rect 31668 28588 31678 28644
rect 33282 28588 33292 28644
rect 33348 28588 37660 28644
rect 37716 28588 37726 28644
rect 38612 28588 41020 28644
rect 41076 28588 41086 28644
rect 26348 28532 26404 28588
rect 47068 28532 47124 28700
rect 55580 28644 55636 28700
rect 26348 28476 27132 28532
rect 27188 28476 27198 28532
rect 34514 28476 34524 28532
rect 34580 28476 34972 28532
rect 35028 28476 35038 28532
rect 37314 28476 37324 28532
rect 37380 28476 37390 28532
rect 37874 28476 37884 28532
rect 37940 28476 38780 28532
rect 38836 28476 38846 28532
rect 38994 28476 39004 28532
rect 39060 28476 39340 28532
rect 39396 28476 42868 28532
rect 43138 28476 43148 28532
rect 43204 28476 43820 28532
rect 43876 28476 47124 28532
rect 47180 28588 51100 28644
rect 51156 28588 51166 28644
rect 55570 28588 55580 28644
rect 55636 28588 55646 28644
rect 37324 28420 37380 28476
rect 42812 28420 42868 28476
rect 47180 28420 47236 28588
rect 2930 28364 2940 28420
rect 2996 28364 20524 28420
rect 20580 28364 20590 28420
rect 26338 28364 26348 28420
rect 26404 28364 26908 28420
rect 28466 28364 28476 28420
rect 28532 28364 28924 28420
rect 28980 28364 28990 28420
rect 31714 28364 31724 28420
rect 31780 28364 32172 28420
rect 32228 28364 32238 28420
rect 32834 28364 32844 28420
rect 32900 28364 34748 28420
rect 34804 28364 34814 28420
rect 35858 28364 35868 28420
rect 35924 28364 37100 28420
rect 37156 28364 37166 28420
rect 37324 28364 39116 28420
rect 39172 28364 39182 28420
rect 41682 28364 41692 28420
rect 41748 28364 42364 28420
rect 42420 28364 42430 28420
rect 42812 28364 47236 28420
rect 0 28308 800 28336
rect 26852 28308 26908 28364
rect 59200 28308 60000 28336
rect 0 28252 1932 28308
rect 1988 28252 3052 28308
rect 3108 28252 3118 28308
rect 17266 28252 17276 28308
rect 17332 28252 18060 28308
rect 18116 28252 18126 28308
rect 26852 28252 35420 28308
rect 35476 28252 35486 28308
rect 36082 28252 36092 28308
rect 36148 28252 39004 28308
rect 39060 28252 39070 28308
rect 39218 28252 39228 28308
rect 39284 28252 42140 28308
rect 42196 28252 42206 28308
rect 57922 28252 57932 28308
rect 57988 28252 60000 28308
rect 0 28224 800 28252
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 50546 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50830 28252
rect 59200 28224 60000 28252
rect 1250 28140 1260 28196
rect 1316 28140 18172 28196
rect 18228 28140 18508 28196
rect 18564 28140 18574 28196
rect 25330 28140 25340 28196
rect 25396 28140 32172 28196
rect 32228 28140 32238 28196
rect 32834 28140 32844 28196
rect 32900 28140 33180 28196
rect 33236 28140 33246 28196
rect 34962 28140 34972 28196
rect 35028 28140 35980 28196
rect 36036 28140 36046 28196
rect 38770 28140 38780 28196
rect 38836 28140 48748 28196
rect 48804 28140 48814 28196
rect 51762 28140 51772 28196
rect 51828 28140 52780 28196
rect 52836 28140 53228 28196
rect 53284 28140 53294 28196
rect 16370 28028 16380 28084
rect 16436 28028 17948 28084
rect 18004 28028 22092 28084
rect 22148 28028 23548 28084
rect 23604 28028 23614 28084
rect 24658 28028 24668 28084
rect 24724 28028 25564 28084
rect 25620 28028 25630 28084
rect 27346 28028 27356 28084
rect 27412 28028 28140 28084
rect 28196 28028 28206 28084
rect 33618 28028 33628 28084
rect 33684 28028 35308 28084
rect 35364 28028 35374 28084
rect 35858 28028 35868 28084
rect 35924 28028 37884 28084
rect 37940 28028 37950 28084
rect 50372 28028 52668 28084
rect 52724 28028 52734 28084
rect 50372 27972 50428 28028
rect 17602 27916 17612 27972
rect 17668 27916 19068 27972
rect 19124 27916 19134 27972
rect 21634 27916 21644 27972
rect 21700 27916 22204 27972
rect 22260 27916 22270 27972
rect 25228 27916 25788 27972
rect 25844 27916 25854 27972
rect 28690 27916 28700 27972
rect 28756 27916 29372 27972
rect 29428 27916 36652 27972
rect 36708 27916 36718 27972
rect 38434 27916 38444 27972
rect 38500 27916 39900 27972
rect 39956 27916 40124 27972
rect 40180 27916 40190 27972
rect 40338 27916 40348 27972
rect 40404 27916 50428 27972
rect 25228 27860 25284 27916
rect 40348 27860 40404 27916
rect 1810 27804 1820 27860
rect 1876 27804 3612 27860
rect 3668 27804 3678 27860
rect 6626 27804 6636 27860
rect 6692 27804 20188 27860
rect 20244 27804 20254 27860
rect 20514 27804 20524 27860
rect 20580 27804 21756 27860
rect 21812 27804 21822 27860
rect 22082 27804 22092 27860
rect 22148 27804 25284 27860
rect 25666 27804 25676 27860
rect 25732 27804 28364 27860
rect 28420 27804 28430 27860
rect 34738 27804 34748 27860
rect 34804 27804 35084 27860
rect 35140 27804 35150 27860
rect 39442 27804 39452 27860
rect 39508 27804 40404 27860
rect 50306 27804 50316 27860
rect 50372 27804 51212 27860
rect 51268 27804 51278 27860
rect 52098 27804 52108 27860
rect 52164 27804 53116 27860
rect 53172 27804 53182 27860
rect 18050 27692 18060 27748
rect 18116 27692 21196 27748
rect 21252 27692 21262 27748
rect 26786 27692 26796 27748
rect 26852 27692 27692 27748
rect 27748 27692 27758 27748
rect 34514 27692 34524 27748
rect 34580 27692 35196 27748
rect 35252 27692 35262 27748
rect 39890 27692 39900 27748
rect 39956 27692 41020 27748
rect 41076 27692 41086 27748
rect 0 27636 800 27664
rect 59200 27636 60000 27664
rect 0 27580 2380 27636
rect 2436 27580 3164 27636
rect 3220 27580 3230 27636
rect 19954 27580 19964 27636
rect 20020 27580 21308 27636
rect 21364 27580 22652 27636
rect 22708 27580 22718 27636
rect 22978 27580 22988 27636
rect 23044 27580 23660 27636
rect 23716 27580 24220 27636
rect 24276 27580 38556 27636
rect 38612 27580 41916 27636
rect 41972 27580 43260 27636
rect 43316 27580 43326 27636
rect 57922 27580 57932 27636
rect 57988 27580 60000 27636
rect 0 27552 800 27580
rect 59200 27552 60000 27580
rect 25676 27468 26012 27524
rect 26068 27468 26078 27524
rect 26786 27468 26796 27524
rect 26852 27468 27580 27524
rect 27636 27468 27646 27524
rect 32162 27468 32172 27524
rect 32228 27468 33068 27524
rect 33124 27468 33516 27524
rect 33572 27468 33582 27524
rect 34598 27468 34636 27524
rect 34692 27468 34702 27524
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 25676 27412 25732 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 9212 27356 20188 27412
rect 20244 27356 20254 27412
rect 22876 27356 24668 27412
rect 24724 27356 24734 27412
rect 25666 27356 25676 27412
rect 25732 27356 25742 27412
rect 31714 27356 31724 27412
rect 31780 27356 34524 27412
rect 34580 27356 34590 27412
rect 9212 27188 9268 27356
rect 22876 27300 22932 27356
rect 2034 27132 2044 27188
rect 2100 27132 9268 27188
rect 15092 27244 22876 27300
rect 22932 27244 22942 27300
rect 23426 27244 23436 27300
rect 23492 27244 30380 27300
rect 30436 27244 32732 27300
rect 32788 27244 33404 27300
rect 33460 27244 33470 27300
rect 15092 27076 15148 27244
rect 34524 27188 34580 27356
rect 34738 27244 34748 27300
rect 34804 27244 45948 27300
rect 46004 27244 46014 27300
rect 16594 27132 16604 27188
rect 16660 27132 17276 27188
rect 17332 27132 17342 27188
rect 24994 27132 25004 27188
rect 25060 27132 26572 27188
rect 26628 27132 26638 27188
rect 32162 27132 32172 27188
rect 32228 27132 32620 27188
rect 32676 27132 32686 27188
rect 32834 27132 32844 27188
rect 32900 27132 32938 27188
rect 34524 27132 35196 27188
rect 35252 27132 35262 27188
rect 43138 27132 43148 27188
rect 43204 27132 50428 27188
rect 50372 27076 50428 27132
rect 1698 27020 1708 27076
rect 1764 27020 3612 27076
rect 3668 27020 3678 27076
rect 5058 27020 5068 27076
rect 5124 27020 15148 27076
rect 23538 27020 23548 27076
rect 23604 27020 24556 27076
rect 24612 27020 25676 27076
rect 25732 27020 25742 27076
rect 27570 27020 27580 27076
rect 27636 27020 27692 27076
rect 27748 27020 27758 27076
rect 29698 27020 29708 27076
rect 29764 27020 30044 27076
rect 30100 27020 30828 27076
rect 30884 27020 30894 27076
rect 31378 27020 31388 27076
rect 31444 27020 33964 27076
rect 34020 27020 34030 27076
rect 35252 27020 38892 27076
rect 38948 27020 38958 27076
rect 46498 27020 46508 27076
rect 46564 27020 48076 27076
rect 48132 27020 48142 27076
rect 50372 27020 55580 27076
rect 55636 27020 55646 27076
rect 0 26964 800 26992
rect 35252 26964 35308 27020
rect 59200 26964 60000 26992
rect 0 26908 1876 26964
rect 9650 26908 9660 26964
rect 9716 26908 18620 26964
rect 18676 26908 18686 26964
rect 25106 26908 25116 26964
rect 25172 26908 29260 26964
rect 29316 26908 32172 26964
rect 32228 26908 35308 26964
rect 36306 26908 36316 26964
rect 36372 26908 38724 26964
rect 45266 26908 45276 26964
rect 45332 26908 45612 26964
rect 45668 26908 45678 26964
rect 48738 26908 48748 26964
rect 48804 26908 49196 26964
rect 49252 26908 49262 26964
rect 53554 26908 53564 26964
rect 53620 26908 54460 26964
rect 54516 26908 54526 26964
rect 57484 26908 60000 26964
rect 0 26880 800 26908
rect 1820 26404 1876 26908
rect 38668 26852 38724 26908
rect 57484 26852 57540 26908
rect 59200 26880 60000 26908
rect 2482 26796 2492 26852
rect 2548 26796 3164 26852
rect 3220 26796 3230 26852
rect 15138 26796 15148 26852
rect 15204 26796 23436 26852
rect 23492 26796 23502 26852
rect 27794 26796 27804 26852
rect 27860 26796 33852 26852
rect 33908 26796 33918 26852
rect 38668 26796 42812 26852
rect 42868 26796 42878 26852
rect 47618 26796 47628 26852
rect 47684 26796 47852 26852
rect 47908 26796 47918 26852
rect 52434 26796 52444 26852
rect 52500 26796 52892 26852
rect 52948 26796 52958 26852
rect 57474 26796 57484 26852
rect 57540 26796 57550 26852
rect 3378 26684 3388 26740
rect 3444 26684 9996 26740
rect 10052 26684 10062 26740
rect 20514 26684 20524 26740
rect 20580 26684 30604 26740
rect 30660 26684 30670 26740
rect 40338 26684 40348 26740
rect 40404 26684 41020 26740
rect 41076 26684 41086 26740
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 50546 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50830 26684
rect 2706 26572 2716 26628
rect 2772 26572 19068 26628
rect 19124 26572 19134 26628
rect 23846 26572 23884 26628
rect 23940 26572 23950 26628
rect 33058 26572 33068 26628
rect 33124 26572 37100 26628
rect 37156 26572 37166 26628
rect 2034 26460 2044 26516
rect 2100 26460 8036 26516
rect 12674 26460 12684 26516
rect 12740 26460 14364 26516
rect 14420 26460 14430 26516
rect 23202 26460 23212 26516
rect 23268 26460 25564 26516
rect 25620 26460 25630 26516
rect 26422 26460 26460 26516
rect 26516 26460 26526 26516
rect 26674 26460 26684 26516
rect 26740 26460 35756 26516
rect 35812 26460 35822 26516
rect 41794 26460 41804 26516
rect 41860 26460 43148 26516
rect 43204 26460 43214 26516
rect 54898 26460 54908 26516
rect 54964 26460 55580 26516
rect 55636 26460 55646 26516
rect 1782 26348 1820 26404
rect 1876 26348 4732 26404
rect 4788 26348 4798 26404
rect 0 26292 800 26320
rect 0 26236 2492 26292
rect 2548 26236 2558 26292
rect 0 26208 800 26236
rect 7980 26180 8036 26460
rect 9314 26348 9324 26404
rect 9380 26348 9884 26404
rect 9940 26348 11116 26404
rect 11172 26348 13804 26404
rect 13860 26348 13870 26404
rect 14018 26348 14028 26404
rect 14084 26348 20412 26404
rect 20468 26348 20478 26404
rect 29698 26348 29708 26404
rect 29764 26348 30940 26404
rect 30996 26348 31006 26404
rect 31154 26348 31164 26404
rect 31220 26348 31612 26404
rect 31668 26348 31678 26404
rect 32134 26348 32172 26404
rect 32228 26348 33516 26404
rect 33572 26348 33582 26404
rect 50306 26348 50316 26404
rect 8194 26236 8204 26292
rect 8260 26236 10108 26292
rect 10164 26236 10174 26292
rect 11554 26236 11564 26292
rect 11620 26236 12348 26292
rect 12404 26236 13132 26292
rect 13188 26236 13198 26292
rect 15092 26236 18172 26292
rect 18228 26236 18238 26292
rect 23314 26236 23324 26292
rect 23380 26236 27468 26292
rect 27524 26236 27534 26292
rect 30706 26236 30716 26292
rect 30772 26236 31500 26292
rect 31556 26236 31566 26292
rect 31826 26236 31836 26292
rect 31892 26236 33404 26292
rect 33460 26236 33470 26292
rect 34066 26236 34076 26292
rect 34132 26236 34524 26292
rect 34580 26236 34590 26292
rect 42578 26236 42588 26292
rect 42644 26236 43260 26292
rect 43316 26236 44492 26292
rect 44548 26236 44558 26292
rect 47730 26236 47740 26292
rect 47796 26236 50092 26292
rect 50148 26236 50158 26292
rect 15092 26180 15148 26236
rect 1820 26124 3052 26180
rect 3108 26124 3836 26180
rect 3892 26124 3902 26180
rect 4274 26124 4284 26180
rect 4340 26124 4350 26180
rect 7980 26124 15148 26180
rect 20738 26124 20748 26180
rect 20804 26124 24220 26180
rect 24276 26124 24286 26180
rect 24882 26124 24892 26180
rect 24948 26124 26572 26180
rect 26628 26124 26638 26180
rect 43698 26124 43708 26180
rect 43764 26124 44380 26180
rect 44436 26124 44446 26180
rect 0 25620 800 25648
rect 1820 25620 1876 26124
rect 4284 26068 4340 26124
rect 50372 26068 50428 26404
rect 51986 26348 51996 26404
rect 52052 26348 54124 26404
rect 54180 26348 54190 26404
rect 53554 26236 53564 26292
rect 53620 26236 55356 26292
rect 55412 26236 55422 26292
rect 53778 26124 53788 26180
rect 53844 26124 55692 26180
rect 55748 26124 55758 26180
rect 2370 26012 2380 26068
rect 2436 26012 4340 26068
rect 14130 26012 14140 26068
rect 14196 26012 14812 26068
rect 14868 26012 14878 26068
rect 23650 26012 23660 26068
rect 23716 26012 24332 26068
rect 24388 26012 24398 26068
rect 34066 26012 34076 26068
rect 34132 26012 35196 26068
rect 35252 26012 35262 26068
rect 46274 26012 46284 26068
rect 46340 26012 47404 26068
rect 47460 26012 47470 26068
rect 49746 26012 49756 26068
rect 49812 26012 53116 26068
rect 53172 26012 53182 26068
rect 9090 25900 9100 25956
rect 9156 25900 11452 25956
rect 11508 25900 12684 25956
rect 12740 25900 12750 25956
rect 23846 25900 23884 25956
rect 23940 25900 23950 25956
rect 24434 25900 24444 25956
rect 24500 25900 29484 25956
rect 29540 25900 29550 25956
rect 31938 25900 31948 25956
rect 32004 25900 33068 25956
rect 33124 25900 33134 25956
rect 34486 25900 34524 25956
rect 34580 25900 34590 25956
rect 49410 25900 49420 25956
rect 49476 25900 56700 25956
rect 56756 25900 56766 25956
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 5730 25788 5740 25844
rect 5796 25788 6636 25844
rect 6692 25788 6702 25844
rect 15092 25788 19404 25844
rect 19460 25788 19470 25844
rect 39890 25788 39900 25844
rect 39956 25788 55580 25844
rect 55636 25788 57372 25844
rect 57428 25788 57438 25844
rect 4834 25676 4844 25732
rect 4900 25676 5852 25732
rect 5908 25676 5918 25732
rect 15092 25620 15148 25788
rect 22978 25676 22988 25732
rect 23044 25676 33964 25732
rect 34020 25676 34030 25732
rect 34860 25676 38332 25732
rect 38388 25676 38398 25732
rect 49634 25676 49644 25732
rect 49700 25676 50316 25732
rect 50372 25676 50382 25732
rect 51874 25676 51884 25732
rect 51940 25676 52780 25732
rect 52836 25676 52846 25732
rect 0 25564 1876 25620
rect 2034 25564 2044 25620
rect 2100 25564 15148 25620
rect 27010 25564 27020 25620
rect 27076 25564 27468 25620
rect 27524 25564 27534 25620
rect 32498 25564 32508 25620
rect 32564 25564 33292 25620
rect 33348 25564 34524 25620
rect 34580 25564 34590 25620
rect 0 25536 800 25564
rect 34860 25508 34916 25676
rect 37996 25564 39452 25620
rect 39508 25564 39518 25620
rect 47394 25564 47404 25620
rect 47460 25564 47964 25620
rect 48020 25564 52108 25620
rect 52164 25564 52174 25620
rect 37996 25508 38052 25564
rect 4274 25452 4284 25508
rect 4340 25452 4956 25508
rect 5012 25452 5022 25508
rect 5394 25452 5404 25508
rect 5460 25452 6300 25508
rect 6356 25452 7532 25508
rect 7588 25452 7598 25508
rect 7858 25452 7868 25508
rect 7924 25452 8876 25508
rect 8932 25452 9996 25508
rect 10052 25452 10062 25508
rect 14690 25452 14700 25508
rect 14756 25452 18284 25508
rect 18340 25452 18732 25508
rect 18788 25452 18798 25508
rect 28130 25452 28140 25508
rect 28196 25452 31276 25508
rect 31332 25452 31836 25508
rect 31892 25452 31902 25508
rect 32162 25452 32172 25508
rect 32228 25452 32238 25508
rect 32610 25452 32620 25508
rect 32676 25452 33404 25508
rect 33460 25452 34916 25508
rect 36194 25452 36204 25508
rect 36260 25452 37996 25508
rect 38052 25452 38062 25508
rect 38322 25452 38332 25508
rect 38388 25452 40236 25508
rect 40292 25452 40302 25508
rect 40674 25452 40684 25508
rect 40740 25452 41580 25508
rect 41636 25452 41646 25508
rect 45602 25452 45612 25508
rect 45668 25452 47180 25508
rect 47236 25452 48636 25508
rect 48692 25452 49868 25508
rect 49924 25452 49934 25508
rect 50194 25452 50204 25508
rect 50260 25452 50652 25508
rect 50708 25452 51548 25508
rect 51604 25452 51614 25508
rect 55010 25452 55020 25508
rect 55076 25452 55468 25508
rect 55524 25452 55916 25508
rect 55972 25452 55982 25508
rect 32172 25396 32228 25452
rect 4610 25340 4620 25396
rect 4676 25340 5180 25396
rect 5236 25340 5628 25396
rect 5684 25340 5694 25396
rect 5954 25340 5964 25396
rect 6020 25340 7644 25396
rect 7700 25340 7710 25396
rect 7868 25340 8428 25396
rect 8484 25340 9772 25396
rect 9828 25340 9838 25396
rect 10658 25340 10668 25396
rect 10724 25340 10734 25396
rect 15372 25340 23548 25396
rect 23604 25340 23614 25396
rect 30818 25340 30828 25396
rect 30884 25340 32620 25396
rect 32676 25340 32686 25396
rect 32834 25340 32844 25396
rect 32900 25340 33180 25396
rect 33236 25340 33246 25396
rect 33730 25340 33740 25396
rect 33796 25340 34972 25396
rect 35028 25340 35196 25396
rect 35252 25340 35262 25396
rect 37426 25340 37436 25396
rect 37492 25340 39004 25396
rect 39060 25340 39070 25396
rect 46274 25340 46284 25396
rect 46340 25340 47404 25396
rect 47460 25340 48412 25396
rect 48468 25340 48478 25396
rect 49634 25340 49644 25396
rect 49700 25340 50428 25396
rect 50484 25340 50494 25396
rect 52770 25340 52780 25396
rect 52836 25340 53116 25396
rect 53172 25340 53182 25396
rect 57810 25340 57820 25396
rect 57876 25340 57886 25396
rect 7868 25284 7924 25340
rect 5394 25228 5404 25284
rect 5460 25228 7924 25284
rect 8082 25228 8092 25284
rect 8148 25228 9548 25284
rect 9604 25228 9614 25284
rect 10668 25172 10724 25340
rect 15372 25284 15428 25340
rect 57820 25284 57876 25340
rect 10994 25228 11004 25284
rect 11060 25228 15148 25284
rect 15204 25228 15214 25284
rect 15362 25228 15372 25284
rect 15428 25228 15438 25284
rect 15698 25228 15708 25284
rect 15764 25228 18956 25284
rect 19012 25228 19022 25284
rect 20178 25228 20188 25284
rect 20244 25228 23212 25284
rect 23268 25228 23278 25284
rect 31154 25228 31164 25284
rect 31220 25228 31948 25284
rect 32004 25228 32172 25284
rect 32228 25228 32238 25284
rect 37090 25228 37100 25284
rect 37156 25228 39452 25284
rect 39508 25228 39900 25284
rect 39956 25228 41020 25284
rect 41076 25228 41086 25284
rect 48850 25228 48860 25284
rect 48916 25228 49756 25284
rect 49812 25228 49822 25284
rect 49970 25228 49980 25284
rect 50036 25228 50540 25284
rect 50596 25228 50606 25284
rect 52098 25228 52108 25284
rect 52164 25228 53676 25284
rect 53732 25228 53742 25284
rect 54124 25228 57876 25284
rect 9426 25116 9436 25172
rect 9492 25116 10724 25172
rect 11554 25116 11564 25172
rect 11620 25116 12572 25172
rect 12628 25116 12638 25172
rect 12898 25116 12908 25172
rect 12964 25116 14140 25172
rect 14196 25116 14206 25172
rect 34962 25116 34972 25172
rect 35028 25116 35084 25172
rect 35140 25116 35150 25172
rect 10668 25060 10724 25116
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 50546 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50830 25116
rect 10668 25004 13580 25060
rect 13636 25004 13646 25060
rect 30482 25004 30492 25060
rect 30548 25004 31500 25060
rect 31556 25004 31566 25060
rect 31714 25004 31724 25060
rect 31780 25004 33740 25060
rect 33796 25004 33806 25060
rect 34822 25004 34860 25060
rect 34916 25004 34926 25060
rect 0 24948 800 24976
rect 54124 24948 54180 25228
rect 59200 24948 60000 24976
rect 0 24892 1932 24948
rect 1988 24892 1998 24948
rect 7522 24892 7532 24948
rect 7588 24892 8092 24948
rect 8148 24892 8158 24948
rect 21634 24892 21644 24948
rect 21700 24892 22204 24948
rect 22260 24892 23324 24948
rect 23380 24892 24108 24948
rect 24164 24892 24444 24948
rect 24500 24892 24510 24948
rect 25106 24892 25116 24948
rect 25172 24892 26460 24948
rect 26516 24892 26526 24948
rect 26898 24892 26908 24948
rect 26964 24892 27692 24948
rect 27748 24892 27758 24948
rect 29250 24892 29260 24948
rect 29316 24892 32508 24948
rect 32564 24892 32574 24948
rect 34290 24892 34300 24948
rect 34356 24892 34366 24948
rect 34626 24892 34636 24948
rect 34692 24892 35420 24948
rect 35476 24892 35486 24948
rect 45378 24892 45388 24948
rect 45444 24892 46060 24948
rect 46116 24892 54180 24948
rect 57922 24892 57932 24948
rect 57988 24892 60000 24948
rect 0 24864 800 24892
rect 34300 24836 34356 24892
rect 59200 24864 60000 24892
rect 15362 24780 15372 24836
rect 15428 24780 30380 24836
rect 30436 24780 30446 24836
rect 32274 24780 32284 24836
rect 32340 24780 32956 24836
rect 33012 24780 33022 24836
rect 34300 24780 35756 24836
rect 35812 24780 35822 24836
rect 36306 24780 36316 24836
rect 36372 24780 37100 24836
rect 37156 24780 37166 24836
rect 39218 24780 39228 24836
rect 39284 24780 55580 24836
rect 55636 24780 55646 24836
rect 9090 24668 9100 24724
rect 9156 24668 9772 24724
rect 9828 24668 9838 24724
rect 18050 24668 18060 24724
rect 18116 24668 19292 24724
rect 19348 24668 19358 24724
rect 31714 24668 31724 24724
rect 31780 24668 35644 24724
rect 35700 24668 35710 24724
rect 41122 24668 41132 24724
rect 41188 24668 42476 24724
rect 42532 24668 42542 24724
rect 49074 24668 49084 24724
rect 49140 24668 49980 24724
rect 50036 24668 50046 24724
rect 50372 24668 51996 24724
rect 52052 24668 52062 24724
rect 50372 24612 50428 24668
rect 10770 24556 10780 24612
rect 10836 24556 13468 24612
rect 13524 24556 13534 24612
rect 17826 24556 17836 24612
rect 17892 24556 18508 24612
rect 18564 24556 19740 24612
rect 19796 24556 19806 24612
rect 31826 24556 31836 24612
rect 31892 24556 32172 24612
rect 32228 24556 32238 24612
rect 34178 24556 34188 24612
rect 34244 24556 34636 24612
rect 34692 24556 34702 24612
rect 47730 24556 47740 24612
rect 47796 24556 50428 24612
rect 5730 24444 5740 24500
rect 5796 24444 6076 24500
rect 6132 24444 8316 24500
rect 8372 24444 23660 24500
rect 23716 24444 24220 24500
rect 24276 24444 24286 24500
rect 34738 24444 34748 24500
rect 34804 24444 36988 24500
rect 37044 24444 37054 24500
rect 24098 24332 24108 24388
rect 24164 24332 25452 24388
rect 25508 24332 25518 24388
rect 0 24276 800 24304
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 59200 24276 60000 24304
rect 0 24220 2380 24276
rect 2436 24220 2446 24276
rect 30146 24220 30156 24276
rect 30212 24220 34412 24276
rect 34468 24220 34478 24276
rect 40002 24220 40012 24276
rect 40068 24220 42140 24276
rect 42196 24220 44044 24276
rect 44100 24220 44940 24276
rect 44996 24220 45388 24276
rect 45444 24220 45454 24276
rect 55346 24220 55356 24276
rect 55412 24220 60000 24276
rect 0 24192 800 24220
rect 59200 24192 60000 24220
rect 23538 24108 23548 24164
rect 23604 24108 30268 24164
rect 30324 24108 30334 24164
rect 55570 24108 55580 24164
rect 55636 24108 58044 24164
rect 58100 24108 58110 24164
rect 2370 23996 2380 24052
rect 2436 23996 2604 24052
rect 2660 23996 2670 24052
rect 6962 23996 6972 24052
rect 7028 23996 7476 24052
rect 10770 23996 10780 24052
rect 10836 23996 11564 24052
rect 11620 23996 11630 24052
rect 12898 23996 12908 24052
rect 12964 23996 13916 24052
rect 13972 23996 13982 24052
rect 17154 23996 17164 24052
rect 17220 23996 17836 24052
rect 17892 23996 17902 24052
rect 24434 23996 24444 24052
rect 24500 23996 25116 24052
rect 25172 23996 25182 24052
rect 33618 23996 33628 24052
rect 33684 23996 36428 24052
rect 36484 23996 36494 24052
rect 44146 23996 44156 24052
rect 44212 23996 45052 24052
rect 45108 23996 45836 24052
rect 45892 23996 45902 24052
rect 46060 23996 53452 24052
rect 53508 23996 53518 24052
rect 53666 23996 53676 24052
rect 53732 23996 56140 24052
rect 56196 23996 56206 24052
rect 7420 23940 7476 23996
rect 46060 23940 46116 23996
rect 2706 23884 2716 23940
rect 2772 23884 3388 23940
rect 3444 23884 3454 23940
rect 6178 23884 6188 23940
rect 6244 23884 6860 23940
rect 6916 23884 6926 23940
rect 7410 23884 7420 23940
rect 7476 23884 8204 23940
rect 8260 23884 11788 23940
rect 11844 23884 11854 23940
rect 13458 23884 13468 23940
rect 13524 23884 14924 23940
rect 14980 23884 15596 23940
rect 15652 23884 15662 23940
rect 19954 23884 19964 23940
rect 20020 23884 20860 23940
rect 20916 23884 20926 23940
rect 24322 23884 24332 23940
rect 24388 23884 25452 23940
rect 25508 23884 25518 23940
rect 30482 23884 30492 23940
rect 30548 23884 31612 23940
rect 31668 23884 31678 23940
rect 34738 23884 34748 23940
rect 34804 23884 34972 23940
rect 35028 23884 36484 23940
rect 37650 23884 37660 23940
rect 37716 23884 38108 23940
rect 38164 23884 46116 23940
rect 49858 23884 49868 23940
rect 49924 23884 50988 23940
rect 51044 23884 51054 23940
rect 55010 23884 55020 23940
rect 55076 23884 56700 23940
rect 56756 23884 56766 23940
rect 36428 23828 36484 23884
rect 2146 23772 2156 23828
rect 2212 23772 2940 23828
rect 2996 23772 3006 23828
rect 4610 23772 4620 23828
rect 4676 23772 8876 23828
rect 8932 23772 13692 23828
rect 13748 23772 14364 23828
rect 14420 23772 14430 23828
rect 16706 23772 16716 23828
rect 16772 23772 18508 23828
rect 18564 23772 18574 23828
rect 23202 23772 23212 23828
rect 23268 23772 31276 23828
rect 31332 23772 31342 23828
rect 34402 23772 34412 23828
rect 34468 23772 35532 23828
rect 35588 23772 35598 23828
rect 36428 23772 39340 23828
rect 39396 23772 39406 23828
rect 43026 23772 43036 23828
rect 43092 23772 43932 23828
rect 43988 23772 43998 23828
rect 50306 23772 50316 23828
rect 50372 23772 51212 23828
rect 51268 23772 51278 23828
rect 51874 23772 51884 23828
rect 51940 23772 53452 23828
rect 53508 23772 55692 23828
rect 55748 23772 55758 23828
rect 2818 23660 2828 23716
rect 2884 23660 4060 23716
rect 4116 23660 4126 23716
rect 5170 23660 5180 23716
rect 5236 23660 6076 23716
rect 6132 23660 6972 23716
rect 7028 23660 7038 23716
rect 7186 23660 7196 23716
rect 7252 23660 8092 23716
rect 8148 23660 8158 23716
rect 10434 23660 10444 23716
rect 10500 23660 11340 23716
rect 11396 23660 11406 23716
rect 13906 23660 13916 23716
rect 13972 23660 18620 23716
rect 18676 23660 19516 23716
rect 19572 23660 22540 23716
rect 22596 23660 22606 23716
rect 33282 23660 33292 23716
rect 33348 23660 34524 23716
rect 34580 23660 34972 23716
rect 35028 23660 35038 23716
rect 35970 23660 35980 23716
rect 36036 23660 37436 23716
rect 37492 23660 37502 23716
rect 46722 23660 46732 23716
rect 46788 23660 47516 23716
rect 47572 23660 49756 23716
rect 49812 23660 51996 23716
rect 52052 23660 52062 23716
rect 55234 23660 55244 23716
rect 55300 23660 57372 23716
rect 57428 23660 57438 23716
rect 0 23604 800 23632
rect 59200 23604 60000 23632
rect 0 23548 1932 23604
rect 1988 23548 1998 23604
rect 7298 23548 7308 23604
rect 7364 23548 7420 23604
rect 7476 23548 7486 23604
rect 7746 23548 7756 23604
rect 7812 23548 8540 23604
rect 8596 23548 8606 23604
rect 11638 23548 11676 23604
rect 11732 23548 12124 23604
rect 12180 23548 12190 23604
rect 33170 23548 33180 23604
rect 33236 23548 35308 23604
rect 35364 23548 36316 23604
rect 36372 23548 36382 23604
rect 45266 23548 45276 23604
rect 45332 23548 47740 23604
rect 47796 23548 47806 23604
rect 54786 23548 54796 23604
rect 54852 23548 56812 23604
rect 56868 23548 56878 23604
rect 58146 23548 58156 23604
rect 58212 23548 60000 23604
rect 0 23520 800 23548
rect 11676 23492 11732 23548
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 36316 23492 36372 23548
rect 50546 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50830 23548
rect 59200 23520 60000 23548
rect 10098 23436 10108 23492
rect 10164 23436 11732 23492
rect 15362 23436 15372 23492
rect 15428 23436 16492 23492
rect 16548 23436 16558 23492
rect 36316 23436 38556 23492
rect 38612 23436 38622 23492
rect 55458 23436 55468 23492
rect 55524 23436 55804 23492
rect 55860 23436 55870 23492
rect 11666 23324 11676 23380
rect 11732 23324 12572 23380
rect 12628 23324 14476 23380
rect 14532 23324 14542 23380
rect 22306 23324 22316 23380
rect 22372 23324 23436 23380
rect 23492 23324 24444 23380
rect 24500 23324 24510 23380
rect 26226 23324 26236 23380
rect 26292 23324 27468 23380
rect 27524 23324 27534 23380
rect 29362 23324 29372 23380
rect 29428 23324 29708 23380
rect 29764 23324 30828 23380
rect 30884 23324 32060 23380
rect 32116 23324 32126 23380
rect 41010 23324 41020 23380
rect 41076 23324 42140 23380
rect 42196 23324 42206 23380
rect 48066 23324 48076 23380
rect 48132 23324 49980 23380
rect 50036 23324 50428 23380
rect 52994 23324 53004 23380
rect 53060 23324 53900 23380
rect 53956 23324 53966 23380
rect 3332 23212 6860 23268
rect 6916 23212 6926 23268
rect 34710 23212 34748 23268
rect 34804 23212 34814 23268
rect 3332 23156 3388 23212
rect 2258 23100 2268 23156
rect 2324 23100 3164 23156
rect 3220 23100 3388 23156
rect 3602 23100 3612 23156
rect 3668 23100 4844 23156
rect 4900 23100 4910 23156
rect 7074 23100 7084 23156
rect 7140 23100 8204 23156
rect 8260 23100 8652 23156
rect 8708 23100 8718 23156
rect 11218 23100 11228 23156
rect 11284 23100 11900 23156
rect 11956 23100 12684 23156
rect 12740 23100 12750 23156
rect 14802 23100 14812 23156
rect 14868 23100 15036 23156
rect 15092 23100 15102 23156
rect 21298 23100 21308 23156
rect 21364 23100 21980 23156
rect 22036 23100 22540 23156
rect 22596 23100 22606 23156
rect 30818 23100 30828 23156
rect 30884 23100 31276 23156
rect 31332 23100 31342 23156
rect 34290 23100 34300 23156
rect 34356 23100 34636 23156
rect 34692 23100 37100 23156
rect 37156 23100 37166 23156
rect 38658 23100 38668 23156
rect 38724 23100 40908 23156
rect 40964 23100 40974 23156
rect 43922 23100 43932 23156
rect 43988 23100 45388 23156
rect 45444 23100 45454 23156
rect 50372 23100 50428 23324
rect 55010 23212 55020 23268
rect 55076 23212 55804 23268
rect 55860 23212 55870 23268
rect 50484 23100 50494 23156
rect 53330 23100 53340 23156
rect 53396 23100 54684 23156
rect 54740 23100 54750 23156
rect 2818 22988 2828 23044
rect 2884 22988 4172 23044
rect 4228 22988 4238 23044
rect 6412 22988 20412 23044
rect 20468 22988 20478 23044
rect 21746 22988 21756 23044
rect 21812 22988 22652 23044
rect 22708 22988 22718 23044
rect 23734 22988 23772 23044
rect 23828 22988 24668 23044
rect 24724 22988 24734 23044
rect 30930 22988 30940 23044
rect 30996 22988 34524 23044
rect 34580 22988 34590 23044
rect 40226 22988 40236 23044
rect 40292 22988 42812 23044
rect 42868 22988 46396 23044
rect 46452 22988 46462 23044
rect 51650 22988 51660 23044
rect 51716 22988 52108 23044
rect 52164 22988 52174 23044
rect 0 22932 800 22960
rect 6412 22932 6468 22988
rect 0 22876 1708 22932
rect 1764 22876 1774 22932
rect 1932 22876 6468 22932
rect 6626 22876 6636 22932
rect 6692 22876 8764 22932
rect 8820 22876 8830 22932
rect 34850 22876 34860 22932
rect 34916 22876 35196 22932
rect 35252 22876 35262 22932
rect 0 22848 800 22876
rect 1932 22820 1988 22876
rect 1474 22764 1484 22820
rect 1540 22764 1988 22820
rect 2258 22764 2268 22820
rect 2324 22764 2380 22820
rect 2436 22764 2446 22820
rect 34066 22764 34076 22820
rect 34132 22764 34142 22820
rect 44594 22764 44604 22820
rect 44660 22764 46284 22820
rect 46340 22764 47068 22820
rect 47124 22764 47134 22820
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 6066 22652 6076 22708
rect 6132 22652 17500 22708
rect 17556 22652 17566 22708
rect 8978 22540 8988 22596
rect 9044 22540 10108 22596
rect 10164 22540 10174 22596
rect 12898 22540 12908 22596
rect 12964 22540 13804 22596
rect 13860 22540 14812 22596
rect 14868 22540 14878 22596
rect 24546 22540 24556 22596
rect 24612 22540 28028 22596
rect 28084 22540 28094 22596
rect 12226 22428 12236 22484
rect 12292 22428 15820 22484
rect 15876 22428 15886 22484
rect 23650 22428 23660 22484
rect 23716 22428 24220 22484
rect 24276 22428 24286 22484
rect 27906 22428 27916 22484
rect 27972 22428 28700 22484
rect 28756 22428 29260 22484
rect 29316 22428 29326 22484
rect 1474 22316 1484 22372
rect 1540 22316 7084 22372
rect 7140 22316 7150 22372
rect 10658 22316 10668 22372
rect 10724 22316 11452 22372
rect 11508 22316 11518 22372
rect 17826 22316 17836 22372
rect 17892 22316 18396 22372
rect 18452 22316 19068 22372
rect 19124 22316 19134 22372
rect 21858 22316 21868 22372
rect 21924 22316 22652 22372
rect 22708 22316 22876 22372
rect 22932 22316 25564 22372
rect 25620 22316 25630 22372
rect 31490 22316 31500 22372
rect 31556 22316 31724 22372
rect 31780 22316 31790 22372
rect 0 22260 800 22288
rect 0 22204 1764 22260
rect 2706 22204 2716 22260
rect 2772 22204 3724 22260
rect 3780 22204 3790 22260
rect 23202 22204 23212 22260
rect 23268 22204 26348 22260
rect 26404 22204 27356 22260
rect 27412 22204 27422 22260
rect 0 22176 800 22204
rect 1708 22148 1764 22204
rect 34076 22148 34132 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 36194 22540 36204 22596
rect 36260 22540 45276 22596
rect 45332 22540 45342 22596
rect 44258 22428 44268 22484
rect 44324 22428 45164 22484
rect 45220 22428 45230 22484
rect 50530 22428 50540 22484
rect 50596 22428 53004 22484
rect 53060 22428 53070 22484
rect 34738 22316 34748 22372
rect 34804 22316 35196 22372
rect 35252 22316 35262 22372
rect 36530 22316 36540 22372
rect 36596 22316 37436 22372
rect 37492 22316 37502 22372
rect 42578 22316 42588 22372
rect 42644 22316 44828 22372
rect 44884 22316 44894 22372
rect 46274 22316 46284 22372
rect 46340 22316 47516 22372
rect 47572 22316 47582 22372
rect 47842 22316 47852 22372
rect 47908 22316 48020 22372
rect 50418 22316 50428 22372
rect 50484 22316 51436 22372
rect 51492 22316 51502 22372
rect 51874 22316 51884 22372
rect 51940 22316 55244 22372
rect 55300 22316 55310 22372
rect 34402 22204 34412 22260
rect 34468 22204 34972 22260
rect 35028 22204 35038 22260
rect 40450 22204 40460 22260
rect 40516 22204 41244 22260
rect 41300 22204 41310 22260
rect 1708 22092 3500 22148
rect 3556 22092 3566 22148
rect 22082 22092 22092 22148
rect 22148 22092 23660 22148
rect 23716 22092 24780 22148
rect 24836 22092 24846 22148
rect 30482 22092 30492 22148
rect 30548 22092 31052 22148
rect 31108 22092 31118 22148
rect 33842 22092 33852 22148
rect 33908 22092 33918 22148
rect 34076 22092 34300 22148
rect 34356 22092 36988 22148
rect 37044 22092 37054 22148
rect 40002 22092 40012 22148
rect 40068 22092 40908 22148
rect 40964 22092 40974 22148
rect 47394 22092 47404 22148
rect 47460 22092 47740 22148
rect 47796 22092 47806 22148
rect 33852 22036 33908 22092
rect 2594 21980 2604 22036
rect 2660 21980 3612 22036
rect 3668 21980 3678 22036
rect 23538 21980 23548 22036
rect 23604 21980 23772 22036
rect 23828 21980 23838 22036
rect 30146 21980 30156 22036
rect 30212 21980 30716 22036
rect 30772 21980 30782 22036
rect 33852 21980 34524 22036
rect 34580 21980 34590 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 2818 21868 2828 21924
rect 2884 21868 3276 21924
rect 3332 21868 3342 21924
rect 39330 21868 39340 21924
rect 39396 21868 40124 21924
rect 40180 21868 40190 21924
rect 43362 21868 43372 21924
rect 43428 21868 44268 21924
rect 44324 21868 44334 21924
rect 44482 21868 44492 21924
rect 44548 21868 45948 21924
rect 46004 21868 46620 21924
rect 46676 21868 46686 21924
rect 4162 21756 4172 21812
rect 4228 21756 5068 21812
rect 5124 21756 11228 21812
rect 11284 21756 11294 21812
rect 11554 21756 11564 21812
rect 11620 21756 12012 21812
rect 12068 21756 15820 21812
rect 15876 21756 15886 21812
rect 16146 21756 16156 21812
rect 16212 21756 18396 21812
rect 18452 21756 18462 21812
rect 20850 21756 20860 21812
rect 20916 21756 21308 21812
rect 21364 21756 21374 21812
rect 29474 21756 29484 21812
rect 29540 21756 32844 21812
rect 32900 21756 33180 21812
rect 33236 21756 33246 21812
rect 37874 21756 37884 21812
rect 37940 21756 39004 21812
rect 39060 21756 39070 21812
rect 41906 21756 41916 21812
rect 41972 21756 43708 21812
rect 43764 21756 43774 21812
rect 47964 21700 48020 22316
rect 51090 22204 51100 22260
rect 51156 22204 52556 22260
rect 52612 22204 53452 22260
rect 53508 22204 53518 22260
rect 55458 22204 55468 22260
rect 55524 22204 57260 22260
rect 57316 22204 57326 22260
rect 49746 22092 49756 22148
rect 49812 22092 51548 22148
rect 51604 22092 51884 22148
rect 51940 22092 51950 22148
rect 54338 22092 54348 22148
rect 54404 22092 57148 22148
rect 57204 22092 57214 22148
rect 55346 21980 55356 22036
rect 55412 21980 55422 22036
rect 50546 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50830 21980
rect 51314 21868 51324 21924
rect 51380 21868 51996 21924
rect 52052 21868 52668 21924
rect 52724 21868 52734 21924
rect 55356 21812 55412 21980
rect 55794 21868 55804 21924
rect 55860 21868 56924 21924
rect 56980 21868 56990 21924
rect 49634 21756 49644 21812
rect 49700 21756 50204 21812
rect 50260 21756 50988 21812
rect 51044 21756 51054 21812
rect 51426 21756 51436 21812
rect 51492 21756 53004 21812
rect 53060 21756 53070 21812
rect 54338 21756 54348 21812
rect 54404 21756 55412 21812
rect 3266 21644 3276 21700
rect 3332 21644 5684 21700
rect 17938 21644 17948 21700
rect 18004 21644 20300 21700
rect 20356 21644 20366 21700
rect 24322 21644 24332 21700
rect 24388 21644 26012 21700
rect 26068 21644 26684 21700
rect 26740 21644 26750 21700
rect 32162 21644 32172 21700
rect 32228 21644 32238 21700
rect 32610 21644 32620 21700
rect 32676 21644 33516 21700
rect 33572 21644 33582 21700
rect 33740 21644 35980 21700
rect 36036 21644 36046 21700
rect 47170 21644 47180 21700
rect 47236 21644 51884 21700
rect 51940 21644 51950 21700
rect 55906 21644 55916 21700
rect 55972 21644 56812 21700
rect 56868 21644 56878 21700
rect 0 21588 800 21616
rect 5628 21588 5684 21644
rect 32172 21588 32228 21644
rect 33740 21588 33796 21644
rect 59200 21588 60000 21616
rect 0 21532 1932 21588
rect 1988 21532 1998 21588
rect 2706 21532 2716 21588
rect 2772 21532 2782 21588
rect 3276 21532 3612 21588
rect 3668 21532 3678 21588
rect 5618 21532 5628 21588
rect 5684 21532 6524 21588
rect 6580 21532 6590 21588
rect 7186 21532 7196 21588
rect 7252 21532 10444 21588
rect 10500 21532 10510 21588
rect 11218 21532 11228 21588
rect 11284 21532 12124 21588
rect 12180 21532 12190 21588
rect 17602 21532 17612 21588
rect 17668 21532 19068 21588
rect 19124 21532 19134 21588
rect 20402 21532 20412 21588
rect 20468 21532 21756 21588
rect 21812 21532 21822 21588
rect 23538 21532 23548 21588
rect 23604 21532 24556 21588
rect 24612 21532 24622 21588
rect 26338 21532 26348 21588
rect 26404 21532 27132 21588
rect 27188 21532 27468 21588
rect 27524 21532 27534 21588
rect 32172 21532 33796 21588
rect 34402 21532 34412 21588
rect 34468 21532 36204 21588
rect 36260 21532 36270 21588
rect 54786 21532 54796 21588
rect 54852 21532 56588 21588
rect 56644 21532 56654 21588
rect 58146 21532 58156 21588
rect 58212 21532 60000 21588
rect 0 21504 800 21532
rect 2716 21476 2772 21532
rect 3276 21476 3332 21532
rect 2716 21420 3332 21476
rect 12124 21476 12180 21532
rect 59200 21504 60000 21532
rect 12124 21420 12572 21476
rect 12628 21420 13580 21476
rect 13636 21420 13646 21476
rect 18162 21420 18172 21476
rect 18228 21420 19180 21476
rect 19236 21420 19246 21476
rect 28578 21420 28588 21476
rect 28644 21420 29148 21476
rect 29204 21420 32732 21476
rect 32788 21420 32798 21476
rect 35858 21420 35868 21476
rect 35924 21420 36428 21476
rect 36484 21420 37324 21476
rect 37380 21420 37390 21476
rect 2034 21308 2044 21364
rect 2100 21308 12236 21364
rect 12292 21308 12302 21364
rect 28018 21308 28028 21364
rect 28084 21308 31276 21364
rect 31332 21308 31342 21364
rect 38546 21308 38556 21364
rect 38612 21308 40236 21364
rect 40292 21308 42476 21364
rect 42532 21308 57820 21364
rect 57876 21308 57886 21364
rect 3238 21196 3276 21252
rect 3332 21196 3342 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 5170 20972 5180 21028
rect 5236 20972 6412 21028
rect 6468 20972 7196 21028
rect 7252 20972 7262 21028
rect 23090 20972 23100 21028
rect 23156 20972 24444 21028
rect 24500 20972 24510 21028
rect 0 20916 800 20944
rect 0 20860 1820 20916
rect 1876 20860 1886 20916
rect 6290 20860 6300 20916
rect 6356 20860 23548 20916
rect 23604 20860 23614 20916
rect 26002 20860 26012 20916
rect 26068 20860 27692 20916
rect 27748 20860 27758 20916
rect 32498 20860 32508 20916
rect 32564 20860 35084 20916
rect 35140 20860 35150 20916
rect 39554 20860 39564 20916
rect 39620 20860 39630 20916
rect 0 20832 800 20860
rect 1698 20748 1708 20804
rect 1764 20748 2380 20804
rect 2436 20748 2446 20804
rect 6178 20748 6188 20804
rect 6244 20748 6972 20804
rect 7028 20748 7038 20804
rect 7858 20748 7868 20804
rect 7924 20748 8540 20804
rect 8596 20748 9324 20804
rect 9380 20748 9390 20804
rect 16482 20748 16492 20804
rect 16548 20748 17724 20804
rect 17780 20748 19404 20804
rect 19460 20748 19470 20804
rect 39564 20692 39620 20860
rect 43698 20748 43708 20804
rect 43764 20748 45052 20804
rect 45108 20748 46788 20804
rect 46732 20692 46788 20748
rect 3602 20636 3612 20692
rect 3668 20636 3836 20692
rect 3892 20636 4956 20692
rect 5012 20636 5022 20692
rect 8978 20636 8988 20692
rect 9044 20636 9772 20692
rect 9828 20636 10668 20692
rect 10724 20636 11116 20692
rect 11172 20636 11676 20692
rect 11732 20636 11742 20692
rect 12786 20636 12796 20692
rect 12852 20636 14028 20692
rect 14084 20636 14094 20692
rect 31714 20636 31724 20692
rect 31780 20636 32620 20692
rect 32676 20636 32686 20692
rect 35634 20636 35644 20692
rect 35700 20636 39620 20692
rect 45266 20636 45276 20692
rect 45332 20636 45948 20692
rect 46004 20636 46014 20692
rect 46722 20636 46732 20692
rect 46788 20636 46798 20692
rect 50978 20636 50988 20692
rect 51044 20636 52892 20692
rect 52948 20636 55020 20692
rect 55076 20636 55804 20692
rect 55860 20636 55870 20692
rect 2790 20524 2828 20580
rect 2884 20524 2894 20580
rect 3378 20524 3388 20580
rect 3444 20524 4508 20580
rect 4564 20524 4574 20580
rect 4722 20524 4732 20580
rect 4788 20524 4844 20580
rect 4900 20524 4910 20580
rect 8194 20524 8204 20580
rect 8260 20524 8764 20580
rect 8820 20524 9884 20580
rect 9940 20524 9950 20580
rect 11890 20524 11900 20580
rect 11956 20524 23324 20580
rect 23380 20524 23390 20580
rect 29250 20524 29260 20580
rect 29316 20524 29708 20580
rect 29764 20524 29774 20580
rect 48514 20524 48524 20580
rect 48580 20524 50316 20580
rect 50372 20524 50382 20580
rect 4050 20412 4060 20468
rect 4116 20412 4844 20468
rect 4900 20412 8092 20468
rect 8148 20412 8876 20468
rect 8932 20412 10332 20468
rect 10388 20412 10398 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 50546 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50830 20412
rect 3826 20300 3836 20356
rect 3892 20300 5964 20356
rect 6020 20300 7420 20356
rect 7476 20300 7486 20356
rect 48514 20300 48524 20356
rect 48580 20300 49308 20356
rect 49364 20300 49374 20356
rect 0 20244 800 20272
rect 0 20188 1708 20244
rect 1764 20188 1774 20244
rect 5842 20188 5852 20244
rect 5908 20188 6860 20244
rect 6916 20188 6926 20244
rect 15810 20188 15820 20244
rect 15876 20188 16996 20244
rect 19618 20188 19628 20244
rect 19684 20188 20300 20244
rect 20356 20188 20366 20244
rect 21074 20188 21084 20244
rect 21140 20188 26908 20244
rect 32834 20188 32844 20244
rect 32900 20188 33572 20244
rect 47618 20188 47628 20244
rect 47684 20188 48748 20244
rect 48804 20188 48814 20244
rect 0 20160 800 20188
rect 16940 20132 16996 20188
rect 2482 20076 2492 20132
rect 2548 20076 3836 20132
rect 3892 20076 5124 20132
rect 5506 20076 5516 20132
rect 5572 20076 6300 20132
rect 6356 20076 7196 20132
rect 7252 20076 7262 20132
rect 10434 20076 10444 20132
rect 10500 20076 11340 20132
rect 11396 20076 11406 20132
rect 12674 20076 12684 20132
rect 12740 20076 13132 20132
rect 13188 20076 14252 20132
rect 14308 20076 14318 20132
rect 15922 20076 15932 20132
rect 15988 20076 16716 20132
rect 16772 20076 16782 20132
rect 16940 20076 19292 20132
rect 19348 20076 20076 20132
rect 20132 20076 20142 20132
rect 22866 20076 22876 20132
rect 22932 20076 24668 20132
rect 24724 20076 24734 20132
rect 25554 20076 25564 20132
rect 25620 20076 26572 20132
rect 26628 20076 26638 20132
rect 5068 20020 5124 20076
rect 2594 19964 2604 20020
rect 2660 19964 3724 20020
rect 3780 19964 3790 20020
rect 5058 19964 5068 20020
rect 5124 19964 5134 20020
rect 9090 19964 9100 20020
rect 9156 19964 10332 20020
rect 10388 19964 11564 20020
rect 11620 19964 11630 20020
rect 16146 19964 16156 20020
rect 16212 19964 18508 20020
rect 18564 19964 18956 20020
rect 19012 19964 19022 20020
rect 24434 19964 24444 20020
rect 24500 19964 25228 20020
rect 25284 19964 25294 20020
rect 26852 19908 26908 20188
rect 33516 20132 33572 20188
rect 28242 20076 28252 20132
rect 28308 20076 28588 20132
rect 28644 20076 28654 20132
rect 30370 20076 30380 20132
rect 30436 20076 31612 20132
rect 31668 20076 31678 20132
rect 33516 20076 34412 20132
rect 34468 20076 37100 20132
rect 37156 20076 37772 20132
rect 37828 20076 37838 20132
rect 43810 20076 43820 20132
rect 43876 20076 48412 20132
rect 48468 20076 49084 20132
rect 49140 20076 49150 20132
rect 30034 19964 30044 20020
rect 30100 19964 30492 20020
rect 30548 19964 30558 20020
rect 30706 19964 30716 20020
rect 30772 19964 30782 20020
rect 32050 19964 32060 20020
rect 32116 19964 33292 20020
rect 33348 19964 33358 20020
rect 40002 19964 40012 20020
rect 40068 19964 40796 20020
rect 40852 19964 41356 20020
rect 41412 19964 42476 20020
rect 42532 19964 42542 20020
rect 42690 19964 42700 20020
rect 42756 19964 43148 20020
rect 43204 19964 43596 20020
rect 43652 19964 43662 20020
rect 50082 19964 50092 20020
rect 50148 19964 51548 20020
rect 51604 19964 51614 20020
rect 52434 19964 52444 20020
rect 52500 19964 54124 20020
rect 54180 19964 54190 20020
rect 30716 19908 30772 19964
rect 2706 19852 2716 19908
rect 2772 19852 3276 19908
rect 3332 19852 3342 19908
rect 6290 19852 6300 19908
rect 6356 19852 7532 19908
rect 7588 19852 8540 19908
rect 8596 19852 9772 19908
rect 9828 19852 9838 19908
rect 20402 19852 20412 19908
rect 20468 19852 24556 19908
rect 24612 19852 24780 19908
rect 24836 19852 26124 19908
rect 26180 19852 26190 19908
rect 26852 19852 30772 19908
rect 41122 19852 41132 19908
rect 41188 19852 41692 19908
rect 41748 19852 42364 19908
rect 42420 19852 42532 19908
rect 42914 19852 42924 19908
rect 42980 19852 43932 19908
rect 43988 19852 43998 19908
rect 51202 19852 51212 19908
rect 51268 19852 53788 19908
rect 53844 19852 53854 19908
rect 26852 19740 33628 19796
rect 33684 19740 33694 19796
rect 26852 19684 26908 19740
rect 42476 19684 42532 19852
rect 43474 19740 43484 19796
rect 43540 19740 44156 19796
rect 44212 19740 44222 19796
rect 22754 19628 22764 19684
rect 22820 19628 26908 19684
rect 29698 19628 29708 19684
rect 29764 19628 31724 19684
rect 31780 19628 31790 19684
rect 42476 19628 43596 19684
rect 43652 19628 43662 19684
rect 0 19572 800 19600
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 0 19516 1708 19572
rect 1764 19516 1774 19572
rect 15250 19516 15260 19572
rect 15316 19516 20972 19572
rect 21028 19516 21038 19572
rect 29810 19516 29820 19572
rect 29876 19516 31500 19572
rect 31556 19516 31566 19572
rect 36194 19516 36204 19572
rect 36260 19516 38668 19572
rect 38724 19516 39900 19572
rect 39956 19516 39966 19572
rect 0 19488 800 19516
rect 42812 19460 42868 19628
rect 2706 19404 2716 19460
rect 2772 19404 6076 19460
rect 6132 19404 6142 19460
rect 14466 19404 14476 19460
rect 14532 19404 16716 19460
rect 16772 19404 17052 19460
rect 17108 19404 18060 19460
rect 18116 19404 18126 19460
rect 29362 19404 29372 19460
rect 29428 19404 30828 19460
rect 30884 19404 33852 19460
rect 33908 19404 33918 19460
rect 37314 19404 37324 19460
rect 37380 19404 39004 19460
rect 39060 19404 39070 19460
rect 42802 19404 42812 19460
rect 42868 19404 42878 19460
rect 47506 19404 47516 19460
rect 47572 19404 48860 19460
rect 48916 19404 48926 19460
rect 53554 19404 53564 19460
rect 53620 19404 55804 19460
rect 55860 19404 55870 19460
rect 5954 19292 5964 19348
rect 6020 19292 15260 19348
rect 15316 19292 15326 19348
rect 15810 19292 15820 19348
rect 15876 19292 17948 19348
rect 18004 19292 20524 19348
rect 20580 19292 20590 19348
rect 40562 19292 40572 19348
rect 40628 19292 41020 19348
rect 41076 19292 45612 19348
rect 45668 19292 45678 19348
rect 54450 19292 54460 19348
rect 54516 19292 56700 19348
rect 56756 19292 57484 19348
rect 57540 19292 57550 19348
rect 3602 19180 3612 19236
rect 3668 19180 4172 19236
rect 4228 19180 4238 19236
rect 4946 19180 4956 19236
rect 5012 19180 5292 19236
rect 5348 19180 6076 19236
rect 6132 19180 6142 19236
rect 6850 19180 6860 19236
rect 6916 19180 8316 19236
rect 8372 19180 8988 19236
rect 9044 19180 9054 19236
rect 12898 19180 12908 19236
rect 12964 19180 14476 19236
rect 14532 19180 14542 19236
rect 16034 19180 16044 19236
rect 16100 19180 16110 19236
rect 19506 19180 19516 19236
rect 19572 19180 20636 19236
rect 20692 19180 22204 19236
rect 22260 19180 22876 19236
rect 22932 19180 22942 19236
rect 26002 19180 26012 19236
rect 26068 19180 28028 19236
rect 28084 19180 28094 19236
rect 28578 19180 28588 19236
rect 28644 19180 29148 19236
rect 29204 19180 29214 19236
rect 31602 19180 31612 19236
rect 31668 19180 32732 19236
rect 32788 19180 32798 19236
rect 37314 19180 37324 19236
rect 37380 19180 38780 19236
rect 38836 19180 38846 19236
rect 42018 19180 42028 19236
rect 42084 19180 43708 19236
rect 43764 19180 49420 19236
rect 49476 19180 53116 19236
rect 53172 19180 53900 19236
rect 53956 19180 53966 19236
rect 2370 19068 2380 19124
rect 2436 19068 3500 19124
rect 3556 19068 5740 19124
rect 5796 19068 5806 19124
rect 8754 19068 8764 19124
rect 8820 19068 11228 19124
rect 11284 19068 11294 19124
rect 13458 19068 13468 19124
rect 13524 19068 15036 19124
rect 15092 19068 15484 19124
rect 15540 19068 15550 19124
rect 0 18900 800 18928
rect 16044 18900 16100 19180
rect 19730 19068 19740 19124
rect 19796 19068 21420 19124
rect 21476 19068 21756 19124
rect 21812 19068 21822 19124
rect 31490 19068 31500 19124
rect 31556 19068 32508 19124
rect 32564 19068 32574 19124
rect 41794 19068 41804 19124
rect 41860 19068 43820 19124
rect 43876 19068 43886 19124
rect 44258 19068 44268 19124
rect 44324 19068 45052 19124
rect 45108 19068 45118 19124
rect 53554 19068 53564 19124
rect 53620 19068 55020 19124
rect 55076 19068 55086 19124
rect 20402 18956 20412 19012
rect 20468 18956 23436 19012
rect 23492 18956 23502 19012
rect 27010 18956 27020 19012
rect 27076 18956 28812 19012
rect 28868 18956 29260 19012
rect 29316 18956 29326 19012
rect 31826 18956 31836 19012
rect 31892 18956 32732 19012
rect 32788 18956 32798 19012
rect 43138 18956 43148 19012
rect 43204 18956 45388 19012
rect 45444 18956 45454 19012
rect 46834 18956 46844 19012
rect 46900 18956 47404 19012
rect 47460 18956 47470 19012
rect 49522 18956 49532 19012
rect 49588 18956 51044 19012
rect 0 18844 2940 18900
rect 2996 18844 3006 18900
rect 5170 18844 5180 18900
rect 5236 18844 15708 18900
rect 15764 18844 16100 18900
rect 24770 18844 24780 18900
rect 24836 18844 25452 18900
rect 25508 18844 25518 18900
rect 44258 18844 44268 18900
rect 44324 18844 45164 18900
rect 45220 18844 45230 18900
rect 0 18816 800 18844
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 50546 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50830 18844
rect 12114 18732 12124 18788
rect 12180 18732 13468 18788
rect 13524 18732 16604 18788
rect 16660 18732 17500 18788
rect 17556 18732 17566 18788
rect 37202 18732 37212 18788
rect 37268 18732 39116 18788
rect 39172 18732 39182 18788
rect 45276 18732 48524 18788
rect 48580 18732 49644 18788
rect 49700 18732 49710 18788
rect 39116 18676 39172 18732
rect 45276 18676 45332 18732
rect 50988 18676 51044 18956
rect 3266 18620 3276 18676
rect 3332 18620 3724 18676
rect 3780 18620 3790 18676
rect 4022 18620 4060 18676
rect 4116 18620 4126 18676
rect 5842 18620 5852 18676
rect 5908 18620 11900 18676
rect 11956 18620 11966 18676
rect 24546 18620 24556 18676
rect 24612 18620 25228 18676
rect 25284 18620 26572 18676
rect 26628 18620 26638 18676
rect 31490 18620 31500 18676
rect 31556 18620 31724 18676
rect 31780 18620 31790 18676
rect 32162 18620 32172 18676
rect 32228 18620 33292 18676
rect 33348 18620 33358 18676
rect 39116 18620 45332 18676
rect 47282 18620 47292 18676
rect 47348 18620 50428 18676
rect 50484 18620 50494 18676
rect 50754 18620 50764 18676
rect 50820 18620 51044 18676
rect 5058 18508 5068 18564
rect 5124 18508 5516 18564
rect 5572 18508 5582 18564
rect 10882 18508 10892 18564
rect 10948 18508 12236 18564
rect 12292 18508 12302 18564
rect 16034 18508 16044 18564
rect 16100 18508 18060 18564
rect 18116 18508 18126 18564
rect 20514 18508 20524 18564
rect 20580 18508 24444 18564
rect 24500 18508 24510 18564
rect 28242 18508 28252 18564
rect 28308 18508 30044 18564
rect 30100 18508 30110 18564
rect 34962 18508 34972 18564
rect 35028 18508 36988 18564
rect 37044 18508 37884 18564
rect 37940 18508 37950 18564
rect 38882 18508 38892 18564
rect 38948 18508 39676 18564
rect 39732 18508 44156 18564
rect 44212 18508 44222 18564
rect 49634 18508 49644 18564
rect 49700 18508 50988 18564
rect 51044 18508 51054 18564
rect 53330 18508 53340 18564
rect 53396 18508 54124 18564
rect 54180 18508 54796 18564
rect 54852 18508 54862 18564
rect 38892 18452 38948 18508
rect 41916 18452 41972 18508
rect 1474 18396 1484 18452
rect 1540 18396 2716 18452
rect 2772 18396 2782 18452
rect 5842 18396 5852 18452
rect 5908 18396 7756 18452
rect 7812 18396 7822 18452
rect 12002 18396 12012 18452
rect 12068 18396 13356 18452
rect 13412 18396 13804 18452
rect 13860 18396 13870 18452
rect 14588 18396 15372 18452
rect 15428 18396 15438 18452
rect 16482 18396 16492 18452
rect 16548 18396 17388 18452
rect 17444 18396 17454 18452
rect 19618 18396 19628 18452
rect 19684 18396 21084 18452
rect 21140 18396 21150 18452
rect 24770 18396 24780 18452
rect 24836 18396 25340 18452
rect 25396 18396 26796 18452
rect 26852 18396 26862 18452
rect 27346 18396 27356 18452
rect 27412 18396 27692 18452
rect 27748 18396 27758 18452
rect 30594 18396 30604 18452
rect 30660 18396 31108 18452
rect 35074 18396 35084 18452
rect 35140 18396 36540 18452
rect 36596 18396 36606 18452
rect 38322 18396 38332 18452
rect 38388 18396 38948 18452
rect 41906 18396 41916 18452
rect 41972 18396 41982 18452
rect 42802 18396 42812 18452
rect 42868 18396 43820 18452
rect 43876 18396 43886 18452
rect 45266 18396 45276 18452
rect 45332 18396 47404 18452
rect 47460 18396 47852 18452
rect 47908 18396 47918 18452
rect 52098 18396 52108 18452
rect 52164 18396 53564 18452
rect 53620 18396 53630 18452
rect 55122 18396 55132 18452
rect 55188 18396 55580 18452
rect 55636 18396 55646 18452
rect 1810 18284 1820 18340
rect 1876 18284 2492 18340
rect 2548 18284 2558 18340
rect 3798 18284 3836 18340
rect 3892 18284 3902 18340
rect 4498 18284 4508 18340
rect 4564 18284 6300 18340
rect 6356 18284 6366 18340
rect 0 18228 800 18256
rect 14588 18228 14644 18396
rect 15026 18284 15036 18340
rect 15092 18284 15484 18340
rect 15540 18284 15550 18340
rect 16492 18228 16548 18396
rect 31052 18340 31108 18396
rect 19058 18284 19068 18340
rect 19124 18284 20300 18340
rect 20356 18284 20366 18340
rect 25778 18284 25788 18340
rect 25844 18284 26908 18340
rect 26964 18284 27468 18340
rect 27524 18284 27534 18340
rect 31042 18284 31052 18340
rect 31108 18284 31118 18340
rect 31378 18284 31388 18340
rect 31444 18284 31836 18340
rect 31892 18284 31902 18340
rect 35970 18284 35980 18340
rect 36036 18284 36428 18340
rect 36484 18284 36494 18340
rect 37874 18284 37884 18340
rect 37940 18284 38556 18340
rect 38612 18284 38622 18340
rect 40338 18284 40348 18340
rect 40404 18284 41356 18340
rect 41412 18284 41422 18340
rect 41682 18284 41692 18340
rect 41748 18284 42252 18340
rect 42308 18284 42318 18340
rect 46610 18284 46620 18340
rect 46676 18284 47292 18340
rect 47348 18284 47740 18340
rect 47796 18284 47806 18340
rect 49074 18284 49084 18340
rect 49140 18284 50876 18340
rect 50932 18284 50942 18340
rect 53442 18284 53452 18340
rect 53508 18284 54572 18340
rect 54628 18284 54638 18340
rect 55010 18284 55020 18340
rect 55076 18284 55916 18340
rect 55972 18284 55982 18340
rect 0 18172 1204 18228
rect 1362 18172 1372 18228
rect 1428 18172 1820 18228
rect 1876 18172 1886 18228
rect 12562 18172 12572 18228
rect 12628 18172 14588 18228
rect 14644 18172 14654 18228
rect 15138 18172 15148 18228
rect 15204 18172 16548 18228
rect 27346 18172 27356 18228
rect 27412 18172 28364 18228
rect 28420 18172 28430 18228
rect 34514 18172 34524 18228
rect 34580 18172 35868 18228
rect 35924 18172 35934 18228
rect 44146 18172 44156 18228
rect 44212 18172 46172 18228
rect 46228 18172 46844 18228
rect 46900 18172 46910 18228
rect 49298 18172 49308 18228
rect 49364 18172 50540 18228
rect 50596 18172 50606 18228
rect 0 18144 800 18172
rect 1148 18116 1204 18172
rect 1148 18060 2604 18116
rect 2660 18060 2670 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 6962 17948 6972 18004
rect 7028 17948 7644 18004
rect 7700 17948 9436 18004
rect 9492 17948 10108 18004
rect 10164 17948 10174 18004
rect 27234 17948 27244 18004
rect 27300 17948 28476 18004
rect 28532 17948 28542 18004
rect 3378 17836 3388 17892
rect 3444 17836 4396 17892
rect 4452 17836 4462 17892
rect 12114 17836 12124 17892
rect 12180 17836 13692 17892
rect 13748 17836 14532 17892
rect 26002 17836 26012 17892
rect 26068 17836 26796 17892
rect 26852 17836 26862 17892
rect 37538 17836 37548 17892
rect 37604 17836 38668 17892
rect 14476 17780 14532 17836
rect 38612 17780 38668 17836
rect 2930 17724 2940 17780
rect 2996 17724 5740 17780
rect 5796 17724 5806 17780
rect 14466 17724 14476 17780
rect 14532 17724 14542 17780
rect 15474 17724 15484 17780
rect 15540 17724 15932 17780
rect 15988 17724 15998 17780
rect 28802 17724 28812 17780
rect 28868 17724 30604 17780
rect 30660 17724 30670 17780
rect 38612 17724 38836 17780
rect 48514 17724 48524 17780
rect 48580 17724 49084 17780
rect 49140 17724 49150 17780
rect 38780 17668 38836 17724
rect 3378 17612 3388 17668
rect 3444 17612 5180 17668
rect 5236 17612 5246 17668
rect 16370 17612 16380 17668
rect 16436 17612 17164 17668
rect 17220 17612 17230 17668
rect 22194 17612 22204 17668
rect 22260 17612 22876 17668
rect 22932 17612 22942 17668
rect 24322 17612 24332 17668
rect 24388 17612 25004 17668
rect 25060 17612 25788 17668
rect 25844 17612 25854 17668
rect 30706 17612 30716 17668
rect 30772 17612 33068 17668
rect 33124 17612 33134 17668
rect 33506 17612 33516 17668
rect 33572 17612 35644 17668
rect 35700 17612 35710 17668
rect 38770 17612 38780 17668
rect 38836 17612 38846 17668
rect 39218 17612 39228 17668
rect 39284 17612 40348 17668
rect 40404 17612 40414 17668
rect 42466 17612 42476 17668
rect 42532 17612 42542 17668
rect 45266 17612 45276 17668
rect 45332 17612 48412 17668
rect 48468 17612 48478 17668
rect 56130 17612 56140 17668
rect 56196 17612 57484 17668
rect 57540 17612 57550 17668
rect 0 17556 800 17584
rect 42476 17556 42532 17612
rect 0 17500 1820 17556
rect 1876 17500 1886 17556
rect 2034 17500 2044 17556
rect 2100 17500 2138 17556
rect 3574 17500 3612 17556
rect 3668 17500 4508 17556
rect 4564 17500 4574 17556
rect 4806 17500 4844 17556
rect 4900 17500 4910 17556
rect 20402 17500 20412 17556
rect 20468 17500 20972 17556
rect 21028 17500 21038 17556
rect 28354 17500 28364 17556
rect 28420 17500 30380 17556
rect 30436 17500 31052 17556
rect 31108 17500 31118 17556
rect 38322 17500 38332 17556
rect 38388 17500 42532 17556
rect 50306 17500 50316 17556
rect 50372 17500 52220 17556
rect 52276 17500 52286 17556
rect 0 17472 800 17500
rect 1698 17388 1708 17444
rect 1764 17388 1876 17444
rect 4162 17388 4172 17444
rect 4228 17388 7756 17444
rect 7812 17388 12460 17444
rect 12516 17388 13132 17444
rect 13188 17388 13198 17444
rect 14354 17388 14364 17444
rect 14420 17388 15484 17444
rect 15540 17388 16156 17444
rect 16212 17388 16222 17444
rect 34962 17388 34972 17444
rect 35028 17388 35756 17444
rect 35812 17388 37100 17444
rect 37156 17388 38108 17444
rect 38164 17388 38174 17444
rect 38770 17388 38780 17444
rect 38836 17388 39228 17444
rect 39284 17388 39294 17444
rect 51202 17388 51212 17444
rect 51268 17388 52108 17444
rect 52164 17388 52174 17444
rect 1820 17332 1876 17388
rect 1810 17276 1820 17332
rect 1876 17276 6748 17332
rect 6804 17276 6814 17332
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 50546 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50830 17276
rect 2342 17164 2380 17220
rect 2436 17164 2446 17220
rect 1698 17052 1708 17108
rect 1764 17052 6300 17108
rect 6356 17052 6366 17108
rect 20626 17052 20636 17108
rect 20692 17052 22764 17108
rect 22820 17052 22830 17108
rect 28130 17052 28140 17108
rect 28196 17052 28700 17108
rect 28756 17052 28766 17108
rect 28914 17052 28924 17108
rect 28980 17052 31388 17108
rect 31444 17052 31454 17108
rect 35522 17052 35532 17108
rect 35588 17052 36540 17108
rect 36596 17052 42140 17108
rect 42196 17052 42206 17108
rect 52434 17052 52444 17108
rect 52500 17052 53228 17108
rect 53284 17052 55916 17108
rect 55972 17052 55982 17108
rect 1922 16940 1932 16996
rect 1988 16940 2940 16996
rect 2996 16940 3006 16996
rect 4498 16940 4508 16996
rect 4564 16940 5292 16996
rect 5348 16940 5358 16996
rect 20738 16940 20748 16996
rect 20804 16940 21756 16996
rect 21812 16940 24444 16996
rect 24500 16940 24510 16996
rect 39554 16940 39564 16996
rect 39620 16940 42252 16996
rect 42308 16940 42318 16996
rect 43026 16940 43036 16996
rect 43092 16940 45948 16996
rect 46004 16940 46014 16996
rect 55570 16940 55580 16996
rect 55636 16940 57372 16996
rect 57428 16940 57438 16996
rect 0 16884 800 16912
rect 0 16828 3164 16884
rect 3220 16828 3230 16884
rect 3490 16828 3500 16884
rect 3556 16828 3836 16884
rect 3892 16828 3902 16884
rect 14130 16828 14140 16884
rect 14196 16828 15036 16884
rect 15092 16828 16940 16884
rect 16996 16828 17006 16884
rect 20962 16828 20972 16884
rect 21028 16828 22204 16884
rect 22260 16828 22270 16884
rect 26562 16828 26572 16884
rect 26628 16828 26908 16884
rect 26964 16828 26974 16884
rect 27990 16828 28028 16884
rect 28084 16828 28094 16884
rect 31490 16828 31500 16884
rect 31556 16828 32060 16884
rect 32116 16828 32126 16884
rect 36754 16828 36764 16884
rect 36820 16828 39788 16884
rect 39844 16828 40460 16884
rect 40516 16828 40526 16884
rect 55458 16828 55468 16884
rect 55524 16828 56812 16884
rect 56868 16828 56878 16884
rect 0 16800 800 16828
rect 4610 16716 4620 16772
rect 4676 16716 5628 16772
rect 5684 16716 5694 16772
rect 13234 16716 13244 16772
rect 13300 16716 15260 16772
rect 15316 16716 15326 16772
rect 30118 16716 30156 16772
rect 30212 16716 30222 16772
rect 34962 16716 34972 16772
rect 35028 16716 36092 16772
rect 36148 16716 36158 16772
rect 39890 16716 39900 16772
rect 39956 16716 42028 16772
rect 42084 16716 42094 16772
rect 51650 16716 51660 16772
rect 51716 16716 53340 16772
rect 53396 16716 55132 16772
rect 55188 16716 55198 16772
rect 2034 16604 2044 16660
rect 2100 16604 15596 16660
rect 15652 16604 15662 16660
rect 28018 16604 28028 16660
rect 28084 16604 29708 16660
rect 29764 16604 29774 16660
rect 46834 16492 46844 16548
rect 46900 16492 49084 16548
rect 49140 16492 49150 16548
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 34402 16380 34412 16436
rect 34468 16380 34972 16436
rect 35028 16380 35038 16436
rect 6962 16268 6972 16324
rect 7028 16268 8876 16324
rect 8932 16268 8942 16324
rect 28578 16268 28588 16324
rect 28644 16268 29260 16324
rect 29316 16268 29326 16324
rect 35298 16268 35308 16324
rect 35364 16268 36428 16324
rect 36484 16268 50204 16324
rect 50260 16268 53228 16324
rect 53284 16268 53676 16324
rect 53732 16268 54572 16324
rect 54628 16268 55020 16324
rect 55076 16268 55086 16324
rect 0 16212 800 16240
rect 0 16156 1764 16212
rect 3154 16156 3164 16212
rect 3220 16156 4172 16212
rect 4228 16156 7420 16212
rect 7476 16156 7486 16212
rect 16258 16156 16268 16212
rect 16324 16156 18956 16212
rect 19012 16156 19022 16212
rect 41794 16156 41804 16212
rect 41860 16156 42252 16212
rect 42308 16156 42318 16212
rect 0 16128 800 16156
rect 1708 15764 1764 16156
rect 4498 16044 4508 16100
rect 4564 16044 5628 16100
rect 5684 16044 6636 16100
rect 6692 16044 6702 16100
rect 7970 16044 7980 16100
rect 8036 16044 8652 16100
rect 8708 16044 8718 16100
rect 10770 16044 10780 16100
rect 10836 16044 11900 16100
rect 11956 16044 11966 16100
rect 12786 16044 12796 16100
rect 12852 16044 13692 16100
rect 13748 16044 15148 16100
rect 16370 16044 16380 16100
rect 16436 16044 18844 16100
rect 18900 16044 18910 16100
rect 19394 16044 19404 16100
rect 19460 16044 20076 16100
rect 20132 16044 21644 16100
rect 21700 16044 21710 16100
rect 23650 16044 23660 16100
rect 23716 16044 24220 16100
rect 24276 16044 25116 16100
rect 25172 16044 27580 16100
rect 27636 16044 27646 16100
rect 34290 16044 34300 16100
rect 34356 16044 35532 16100
rect 35588 16044 35598 16100
rect 36194 16044 36204 16100
rect 36260 16044 37324 16100
rect 37380 16044 37390 16100
rect 38658 16044 38668 16100
rect 38724 16044 39788 16100
rect 39844 16044 41468 16100
rect 41524 16044 41534 16100
rect 49970 16044 49980 16100
rect 50036 16044 50764 16100
rect 50820 16044 50830 16100
rect 55794 16044 55804 16100
rect 55860 16044 56028 16100
rect 56084 16044 56476 16100
rect 56532 16044 56542 16100
rect 2930 15932 2940 15988
rect 2996 15932 3948 15988
rect 4004 15932 4732 15988
rect 4788 15932 4798 15988
rect 11666 15932 11676 15988
rect 11732 15932 14028 15988
rect 14084 15932 14094 15988
rect 15092 15876 15148 16044
rect 15922 15932 15932 15988
rect 15988 15932 16492 15988
rect 16548 15932 17052 15988
rect 17108 15932 19180 15988
rect 19236 15932 19246 15988
rect 20524 15932 23324 15988
rect 23380 15932 23390 15988
rect 33394 15932 33404 15988
rect 33460 15932 34636 15988
rect 34692 15932 34702 15988
rect 35858 15932 35868 15988
rect 35924 15932 43372 15988
rect 43428 15932 44940 15988
rect 44996 15932 45006 15988
rect 45490 15932 45500 15988
rect 45556 15932 46620 15988
rect 46676 15932 48972 15988
rect 49028 15932 49308 15988
rect 49364 15932 49374 15988
rect 49858 15932 49868 15988
rect 49924 15932 50988 15988
rect 51044 15932 51054 15988
rect 20524 15876 20580 15932
rect 2818 15820 2828 15876
rect 2884 15820 3612 15876
rect 3668 15820 3678 15876
rect 4274 15820 4284 15876
rect 4340 15820 5964 15876
rect 6020 15820 6030 15876
rect 6514 15820 6524 15876
rect 6580 15820 7196 15876
rect 7252 15820 7262 15876
rect 15092 15820 17276 15876
rect 17332 15820 20524 15876
rect 20580 15820 20590 15876
rect 22418 15820 22428 15876
rect 22484 15820 23884 15876
rect 23940 15820 23950 15876
rect 30370 15820 30380 15876
rect 30436 15820 31836 15876
rect 31892 15820 31902 15876
rect 35074 15820 35084 15876
rect 35140 15820 35756 15876
rect 35812 15820 35822 15876
rect 37650 15820 37660 15876
rect 37716 15820 39452 15876
rect 39508 15820 39518 15876
rect 43474 15820 43484 15876
rect 43540 15820 44156 15876
rect 44212 15820 44222 15876
rect 54338 15820 54348 15876
rect 54404 15820 55804 15876
rect 55860 15820 56588 15876
rect 56644 15820 56654 15876
rect 1698 15708 1708 15764
rect 1764 15708 1774 15764
rect 2258 15708 2268 15764
rect 2324 15708 4060 15764
rect 4116 15708 4126 15764
rect 7634 15708 7644 15764
rect 7700 15708 11116 15764
rect 11172 15708 11182 15764
rect 26002 15708 26012 15764
rect 26068 15708 26078 15764
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 26012 15652 26068 15708
rect 50546 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50830 15708
rect 26012 15596 26348 15652
rect 26404 15596 26414 15652
rect 29138 15596 29148 15652
rect 29204 15596 29214 15652
rect 34850 15596 34860 15652
rect 34916 15596 37660 15652
rect 37716 15596 37726 15652
rect 0 15540 800 15568
rect 0 15484 2660 15540
rect 4946 15484 4956 15540
rect 5012 15484 5180 15540
rect 5236 15484 5964 15540
rect 6020 15484 6030 15540
rect 6850 15484 6860 15540
rect 6916 15484 7756 15540
rect 7812 15484 7822 15540
rect 25442 15484 25452 15540
rect 25508 15484 26012 15540
rect 26068 15484 26078 15540
rect 0 15456 800 15484
rect 2604 15428 2660 15484
rect 2594 15372 2604 15428
rect 2660 15372 2670 15428
rect 9202 15372 9212 15428
rect 9268 15372 11676 15428
rect 11732 15372 11742 15428
rect 7522 15260 7532 15316
rect 7588 15260 8540 15316
rect 8596 15260 8606 15316
rect 12898 15260 12908 15316
rect 12964 15260 13580 15316
rect 13636 15260 15148 15316
rect 15204 15260 15214 15316
rect 19282 15260 19292 15316
rect 19348 15260 20300 15316
rect 20356 15260 20366 15316
rect 25554 15260 25564 15316
rect 25620 15260 27244 15316
rect 27300 15260 27310 15316
rect 1698 15148 1708 15204
rect 1764 15148 3052 15204
rect 3108 15148 3118 15204
rect 5506 15148 5516 15204
rect 5572 15148 6636 15204
rect 6692 15148 6702 15204
rect 8754 15148 8764 15204
rect 8820 15148 10556 15204
rect 10612 15148 10622 15204
rect 15698 15148 15708 15204
rect 15764 15148 16380 15204
rect 16436 15148 16446 15204
rect 24658 15148 24668 15204
rect 24724 15148 25900 15204
rect 25956 15148 26460 15204
rect 26516 15148 26526 15204
rect 29148 15092 29204 15596
rect 38882 15484 38892 15540
rect 38948 15484 39900 15540
rect 39956 15484 41132 15540
rect 41188 15484 41198 15540
rect 50194 15484 50204 15540
rect 50260 15484 50540 15540
rect 50596 15484 50606 15540
rect 34178 15372 34188 15428
rect 34244 15372 34860 15428
rect 34916 15372 34926 15428
rect 41682 15372 41692 15428
rect 41748 15372 43148 15428
rect 43204 15372 43652 15428
rect 43596 15316 43652 15372
rect 29698 15260 29708 15316
rect 29764 15260 30940 15316
rect 30996 15260 31276 15316
rect 31332 15260 31342 15316
rect 33058 15260 33068 15316
rect 33124 15260 33740 15316
rect 33796 15260 33806 15316
rect 37314 15260 37324 15316
rect 37380 15260 37772 15316
rect 37828 15260 37838 15316
rect 42018 15260 42028 15316
rect 42084 15260 42924 15316
rect 42980 15260 42990 15316
rect 43586 15260 43596 15316
rect 43652 15260 45724 15316
rect 45780 15260 45790 15316
rect 46162 15260 46172 15316
rect 46228 15260 47516 15316
rect 47572 15260 47582 15316
rect 47842 15260 47852 15316
rect 47908 15260 48748 15316
rect 48804 15260 49196 15316
rect 49252 15260 49262 15316
rect 30482 15148 30492 15204
rect 30548 15148 31612 15204
rect 31668 15148 31678 15204
rect 55132 15148 57036 15204
rect 57092 15148 57102 15204
rect 55132 15092 55188 15148
rect 1922 15036 1932 15092
rect 1988 15036 1998 15092
rect 2482 15036 2492 15092
rect 2548 15036 3836 15092
rect 3892 15036 3902 15092
rect 29148 15036 29708 15092
rect 29764 15036 29774 15092
rect 34822 15036 34860 15092
rect 34916 15036 34926 15092
rect 35970 15036 35980 15092
rect 36036 15036 36988 15092
rect 37044 15036 37054 15092
rect 49410 15036 49420 15092
rect 49476 15036 50764 15092
rect 50820 15036 50830 15092
rect 55122 15036 55132 15092
rect 55188 15036 55198 15092
rect 0 14868 800 14896
rect 1932 14868 1988 15036
rect 22754 14924 22764 14980
rect 22820 14924 23100 14980
rect 23156 14924 23166 14980
rect 27570 14924 27580 14980
rect 27636 14924 28476 14980
rect 28532 14924 28542 14980
rect 47618 14924 47628 14980
rect 47684 14924 50428 14980
rect 50484 14924 50494 14980
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 0 14812 1988 14868
rect 6066 14812 6076 14868
rect 6132 14812 6524 14868
rect 6580 14812 6860 14868
rect 6916 14812 6926 14868
rect 50372 14812 50988 14868
rect 51044 14812 51054 14868
rect 0 14784 800 14812
rect 50372 14756 50428 14812
rect 2034 14700 2044 14756
rect 2100 14700 7644 14756
rect 7700 14700 7710 14756
rect 17938 14700 17948 14756
rect 18004 14700 18844 14756
rect 18900 14700 18910 14756
rect 38098 14700 38108 14756
rect 38164 14700 47068 14756
rect 47124 14700 47134 14756
rect 48514 14700 48524 14756
rect 48580 14700 50428 14756
rect 2594 14588 2604 14644
rect 2660 14588 4956 14644
rect 5012 14588 5022 14644
rect 20066 14588 20076 14644
rect 20132 14588 21308 14644
rect 21364 14588 21374 14644
rect 23538 14588 23548 14644
rect 23604 14588 23884 14644
rect 23940 14588 23950 14644
rect 36866 14588 36876 14644
rect 36932 14588 38332 14644
rect 38388 14588 38398 14644
rect 51538 14588 51548 14644
rect 51604 14588 52892 14644
rect 52948 14588 52958 14644
rect 2818 14476 2828 14532
rect 2884 14476 9660 14532
rect 9716 14476 9726 14532
rect 14914 14476 14924 14532
rect 14980 14476 17724 14532
rect 17780 14476 17790 14532
rect 27234 14476 27244 14532
rect 27300 14476 28364 14532
rect 28420 14476 28430 14532
rect 29698 14476 29708 14532
rect 29764 14476 30268 14532
rect 30324 14476 30334 14532
rect 31266 14476 31276 14532
rect 31332 14476 31500 14532
rect 31556 14476 31566 14532
rect 34514 14476 34524 14532
rect 34580 14476 35644 14532
rect 35700 14476 35710 14532
rect 36530 14476 36540 14532
rect 36596 14476 37212 14532
rect 37268 14476 37278 14532
rect 43698 14476 43708 14532
rect 43764 14476 44940 14532
rect 44996 14476 45006 14532
rect 46498 14476 46508 14532
rect 46564 14476 47516 14532
rect 47572 14476 47582 14532
rect 48290 14476 48300 14532
rect 48356 14476 50428 14532
rect 50484 14476 50494 14532
rect 31276 14420 31332 14476
rect 10322 14364 10332 14420
rect 10388 14364 10780 14420
rect 10836 14364 10846 14420
rect 30034 14364 30044 14420
rect 30100 14364 31332 14420
rect 35186 14364 35196 14420
rect 35252 14364 36764 14420
rect 36820 14364 38668 14420
rect 38724 14364 38734 14420
rect 43026 14364 43036 14420
rect 43092 14364 44044 14420
rect 44100 14364 44380 14420
rect 44436 14364 44446 14420
rect 7298 14252 7308 14308
rect 7364 14252 8092 14308
rect 8148 14252 8158 14308
rect 21410 14252 21420 14308
rect 21476 14252 22540 14308
rect 22596 14252 22606 14308
rect 28690 14252 28700 14308
rect 28756 14252 29484 14308
rect 29540 14252 30380 14308
rect 30436 14252 30446 14308
rect 32722 14252 32732 14308
rect 32788 14252 33628 14308
rect 33684 14252 33694 14308
rect 35522 14252 35532 14308
rect 35588 14252 37772 14308
rect 37828 14252 37838 14308
rect 54450 14252 54460 14308
rect 54516 14252 55692 14308
rect 55748 14252 56476 14308
rect 56532 14252 56542 14308
rect 0 14196 800 14224
rect 0 14140 1876 14196
rect 27346 14140 27356 14196
rect 27412 14140 28924 14196
rect 28980 14140 28990 14196
rect 0 14112 800 14140
rect 1820 13972 1876 14140
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 50546 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50830 14140
rect 8092 14028 8204 14084
rect 8260 14028 8270 14084
rect 1810 13916 1820 13972
rect 1876 13916 3612 13972
rect 3668 13916 3678 13972
rect 8092 13748 8148 14028
rect 32498 13916 32508 13972
rect 32564 13916 34972 13972
rect 35028 13916 35038 13972
rect 36194 13916 36204 13972
rect 36260 13916 37100 13972
rect 37156 13916 37166 13972
rect 8306 13804 8316 13860
rect 8372 13804 10108 13860
rect 10164 13804 10174 13860
rect 26562 13804 26572 13860
rect 26628 13804 28252 13860
rect 28308 13804 28318 13860
rect 34178 13804 34188 13860
rect 34244 13804 34748 13860
rect 34804 13804 35420 13860
rect 35476 13804 38444 13860
rect 38500 13804 38510 13860
rect 43250 13804 43260 13860
rect 43316 13804 43596 13860
rect 43652 13804 45388 13860
rect 45444 13804 45454 13860
rect 50754 13804 50764 13860
rect 50820 13804 53228 13860
rect 53284 13804 53294 13860
rect 54786 13804 54796 13860
rect 54852 13804 55356 13860
rect 55412 13804 55422 13860
rect 2034 13692 2044 13748
rect 2100 13692 2828 13748
rect 2884 13692 2894 13748
rect 7410 13692 7420 13748
rect 7476 13692 8540 13748
rect 8596 13692 8606 13748
rect 8754 13692 8764 13748
rect 8820 13692 9436 13748
rect 9492 13692 9502 13748
rect 23314 13692 23324 13748
rect 23380 13692 24108 13748
rect 24164 13692 24174 13748
rect 35074 13692 35084 13748
rect 35140 13692 37548 13748
rect 37604 13692 37614 13748
rect 38322 13692 38332 13748
rect 38388 13692 39564 13748
rect 39620 13692 39630 13748
rect 41122 13692 41132 13748
rect 41188 13692 43036 13748
rect 43092 13692 43102 13748
rect 45714 13692 45724 13748
rect 45780 13692 47292 13748
rect 47348 13692 48972 13748
rect 49028 13692 49038 13748
rect 53666 13692 53676 13748
rect 53732 13692 54236 13748
rect 54292 13692 54572 13748
rect 54628 13692 54638 13748
rect 8540 13636 8596 13692
rect 3332 13580 4060 13636
rect 4116 13580 4126 13636
rect 8540 13580 9884 13636
rect 9940 13580 9950 13636
rect 20626 13580 20636 13636
rect 20692 13580 22876 13636
rect 22932 13580 23436 13636
rect 23492 13580 23502 13636
rect 33170 13580 33180 13636
rect 33236 13580 34076 13636
rect 34132 13580 35644 13636
rect 35700 13580 35710 13636
rect 40114 13580 40124 13636
rect 40180 13580 41468 13636
rect 41524 13580 41534 13636
rect 0 13524 800 13552
rect 3332 13524 3388 13580
rect 0 13468 2380 13524
rect 2436 13468 3388 13524
rect 22530 13468 22540 13524
rect 22596 13468 23884 13524
rect 23940 13468 23950 13524
rect 27990 13468 28028 13524
rect 28084 13468 28094 13524
rect 33618 13468 33628 13524
rect 33684 13468 36820 13524
rect 37202 13468 37212 13524
rect 37268 13468 38220 13524
rect 38276 13468 39788 13524
rect 39844 13468 39854 13524
rect 41794 13468 41804 13524
rect 41860 13468 43932 13524
rect 43988 13468 43998 13524
rect 51650 13468 51660 13524
rect 51716 13468 53004 13524
rect 53060 13468 53340 13524
rect 53396 13468 54348 13524
rect 54404 13468 54414 13524
rect 54562 13468 54572 13524
rect 54628 13468 55132 13524
rect 55188 13468 55198 13524
rect 0 13440 800 13468
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 36764 13300 36820 13468
rect 36754 13244 36764 13300
rect 36820 13244 36830 13300
rect 21746 13132 21756 13188
rect 21812 13132 23996 13188
rect 24052 13132 24062 13188
rect 41458 13132 41468 13188
rect 41524 13132 42364 13188
rect 42420 13132 42430 13188
rect 6262 13020 6300 13076
rect 6356 13020 6860 13076
rect 6916 13020 6926 13076
rect 28550 13020 28588 13076
rect 28644 13020 28654 13076
rect 4834 12908 4844 12964
rect 4900 12908 5740 12964
rect 5796 12908 5806 12964
rect 6066 12908 6076 12964
rect 6132 12908 6748 12964
rect 6804 12908 6814 12964
rect 19618 12908 19628 12964
rect 19684 12908 20748 12964
rect 20804 12908 21420 12964
rect 21476 12908 21486 12964
rect 50372 12908 50988 12964
rect 51044 12908 51054 12964
rect 0 12852 800 12880
rect 50372 12852 50428 12908
rect 0 12796 1708 12852
rect 1764 12796 3612 12852
rect 3668 12796 3678 12852
rect 9314 12796 9324 12852
rect 9380 12796 12572 12852
rect 12628 12796 12638 12852
rect 18050 12796 18060 12852
rect 18116 12796 19292 12852
rect 19348 12796 19358 12852
rect 19516 12796 20076 12852
rect 20132 12796 21756 12852
rect 21812 12796 21822 12852
rect 26114 12796 26124 12852
rect 26180 12796 29484 12852
rect 29540 12796 30268 12852
rect 30324 12796 30334 12852
rect 35298 12796 35308 12852
rect 35364 12796 36428 12852
rect 36484 12796 36494 12852
rect 38546 12796 38556 12852
rect 38612 12796 39676 12852
rect 39732 12796 39742 12852
rect 41906 12796 41916 12852
rect 41972 12796 44828 12852
rect 44884 12796 44894 12852
rect 49410 12796 49420 12852
rect 49476 12796 49868 12852
rect 49924 12796 50428 12852
rect 0 12768 800 12796
rect 19516 12740 19572 12796
rect 19394 12684 19404 12740
rect 19460 12684 19572 12740
rect 22082 12684 22092 12740
rect 22148 12684 23100 12740
rect 23156 12684 23166 12740
rect 24658 12684 24668 12740
rect 24724 12684 28588 12740
rect 28644 12684 28654 12740
rect 38098 12684 38108 12740
rect 38164 12684 38780 12740
rect 38836 12684 38846 12740
rect 41570 12684 41580 12740
rect 41636 12684 42588 12740
rect 42644 12684 42654 12740
rect 47842 12684 47852 12740
rect 47908 12684 49532 12740
rect 49588 12684 49598 12740
rect 37090 12572 37100 12628
rect 37156 12572 40012 12628
rect 40068 12572 40078 12628
rect 48066 12572 48076 12628
rect 48132 12572 48748 12628
rect 48804 12572 49084 12628
rect 49140 12572 49150 12628
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 50546 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50830 12572
rect 37650 12460 37660 12516
rect 37716 12460 40460 12516
rect 40516 12460 43428 12516
rect 43372 12404 43428 12460
rect 38612 12348 39340 12404
rect 39396 12348 42700 12404
rect 42756 12348 42766 12404
rect 43362 12348 43372 12404
rect 43428 12348 43438 12404
rect 51874 12348 51884 12404
rect 51940 12348 53564 12404
rect 53620 12348 53630 12404
rect 38612 12292 38668 12348
rect 16482 12236 16492 12292
rect 16548 12236 18060 12292
rect 18116 12236 18126 12292
rect 18946 12236 18956 12292
rect 19012 12236 19628 12292
rect 19684 12236 19694 12292
rect 23314 12236 23324 12292
rect 23380 12236 25900 12292
rect 25956 12236 25966 12292
rect 26898 12236 26908 12292
rect 26964 12236 28084 12292
rect 38322 12236 38332 12292
rect 38388 12236 38668 12292
rect 38882 12236 38892 12292
rect 38948 12236 41468 12292
rect 41524 12236 41534 12292
rect 0 12180 800 12208
rect 28028 12180 28084 12236
rect 42700 12180 42756 12348
rect 44370 12236 44380 12292
rect 44436 12236 48188 12292
rect 48244 12236 51660 12292
rect 51716 12236 54908 12292
rect 54964 12236 54974 12292
rect 0 12124 2492 12180
rect 2548 12124 2558 12180
rect 5170 12124 5180 12180
rect 5236 12124 6188 12180
rect 6244 12124 6972 12180
rect 7028 12124 7038 12180
rect 8978 12124 8988 12180
rect 9044 12124 9996 12180
rect 10052 12124 11340 12180
rect 11396 12124 11406 12180
rect 24322 12124 24332 12180
rect 24388 12124 25452 12180
rect 25508 12124 25518 12180
rect 27010 12124 27020 12180
rect 27076 12124 27086 12180
rect 28018 12124 28028 12180
rect 28084 12124 28094 12180
rect 36418 12124 36428 12180
rect 36484 12124 37100 12180
rect 37156 12124 37166 12180
rect 38434 12124 38444 12180
rect 38500 12124 40236 12180
rect 40292 12124 40302 12180
rect 42700 12124 47628 12180
rect 47684 12124 47964 12180
rect 48020 12124 48030 12180
rect 49634 12124 49644 12180
rect 49700 12124 50204 12180
rect 50260 12124 50876 12180
rect 50932 12124 50942 12180
rect 51538 12124 51548 12180
rect 51604 12124 52668 12180
rect 52724 12124 52734 12180
rect 0 12096 800 12124
rect 5954 12012 5964 12068
rect 6020 12012 6748 12068
rect 6804 12012 6814 12068
rect 9650 12012 9660 12068
rect 9716 12012 10220 12068
rect 10276 12012 10286 12068
rect 14578 12012 14588 12068
rect 14644 12012 20972 12068
rect 21028 12012 21038 12068
rect 22978 12012 22988 12068
rect 23044 12012 23996 12068
rect 24052 12012 25340 12068
rect 25396 12012 25406 12068
rect 27020 11956 27076 12124
rect 36754 12012 36764 12068
rect 36820 12012 42924 12068
rect 42980 12012 43820 12068
rect 43876 12012 43886 12068
rect 49522 12012 49532 12068
rect 49588 12012 50428 12068
rect 50484 12012 50494 12068
rect 53218 12012 53228 12068
rect 53284 12012 53788 12068
rect 53844 12012 53854 12068
rect 15026 11900 15036 11956
rect 15092 11900 17836 11956
rect 17892 11900 18508 11956
rect 18564 11900 18574 11956
rect 19618 11900 19628 11956
rect 19684 11900 20412 11956
rect 20468 11900 20478 11956
rect 23090 11900 23100 11956
rect 23156 11900 24332 11956
rect 24388 11900 27076 11956
rect 29148 11788 29260 11844
rect 29316 11788 30380 11844
rect 30436 11788 30446 11844
rect 32162 11788 32172 11844
rect 32228 11788 33852 11844
rect 33908 11788 33918 11844
rect 37538 11788 37548 11844
rect 37604 11788 38668 11844
rect 46386 11788 46396 11844
rect 46452 11788 47068 11844
rect 47124 11788 47134 11844
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 29148 11732 29204 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 5730 11676 5740 11732
rect 5796 11676 8428 11732
rect 8484 11676 10444 11732
rect 10500 11676 10510 11732
rect 21858 11676 21868 11732
rect 21924 11676 26236 11732
rect 26292 11676 26302 11732
rect 28018 11676 28028 11732
rect 28084 11676 29204 11732
rect 38612 11620 38668 11788
rect 41234 11676 41244 11732
rect 41300 11676 41916 11732
rect 41972 11676 41982 11732
rect 11442 11564 11452 11620
rect 11508 11564 11788 11620
rect 11844 11564 12684 11620
rect 12740 11564 12750 11620
rect 36306 11564 36316 11620
rect 36372 11564 36764 11620
rect 36820 11564 36830 11620
rect 38612 11564 43708 11620
rect 43764 11564 43774 11620
rect 0 11508 800 11536
rect 0 11452 1708 11508
rect 1764 11452 2940 11508
rect 2996 11452 3006 11508
rect 6850 11452 6860 11508
rect 6916 11452 8652 11508
rect 8708 11452 8718 11508
rect 14242 11452 14252 11508
rect 14308 11452 15372 11508
rect 15428 11452 15438 11508
rect 40002 11452 40012 11508
rect 40068 11452 45836 11508
rect 45892 11452 45902 11508
rect 0 11424 800 11452
rect 6290 11340 6300 11396
rect 6356 11340 6972 11396
rect 7028 11340 7308 11396
rect 7364 11340 7374 11396
rect 7522 11340 7532 11396
rect 7588 11340 10220 11396
rect 10276 11340 10286 11396
rect 11330 11340 11340 11396
rect 11396 11340 12236 11396
rect 12292 11340 12302 11396
rect 13458 11340 13468 11396
rect 13524 11340 14700 11396
rect 14756 11340 15148 11396
rect 16594 11340 16604 11396
rect 16660 11340 17388 11396
rect 17444 11340 17454 11396
rect 20738 11340 20748 11396
rect 20804 11340 21532 11396
rect 21588 11340 21598 11396
rect 38882 11340 38892 11396
rect 38948 11340 40348 11396
rect 40404 11340 40414 11396
rect 44146 11340 44156 11396
rect 44212 11340 44716 11396
rect 44772 11340 46732 11396
rect 46788 11340 47628 11396
rect 47684 11340 47694 11396
rect 49858 11340 49868 11396
rect 49924 11340 50764 11396
rect 50820 11340 50830 11396
rect 15092 11284 15148 11340
rect 1250 11228 1260 11284
rect 1316 11228 2044 11284
rect 2100 11228 2110 11284
rect 5058 11228 5068 11284
rect 5124 11228 5740 11284
rect 5796 11228 5806 11284
rect 7970 11228 7980 11284
rect 8036 11228 9772 11284
rect 9828 11228 9838 11284
rect 12898 11228 12908 11284
rect 12964 11228 13804 11284
rect 13860 11228 13870 11284
rect 15092 11228 17948 11284
rect 18004 11228 18732 11284
rect 18788 11228 18798 11284
rect 27234 11228 27244 11284
rect 27300 11228 28028 11284
rect 28084 11228 28094 11284
rect 36530 11228 36540 11284
rect 36596 11228 37324 11284
rect 37380 11228 37390 11284
rect 43922 11228 43932 11284
rect 43988 11228 44828 11284
rect 44884 11228 45276 11284
rect 45332 11228 45342 11284
rect 36306 11116 36316 11172
rect 36372 11116 37996 11172
rect 38052 11116 38062 11172
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 50546 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50830 11004
rect 2034 10892 2044 10948
rect 2100 10892 3388 10948
rect 0 10836 800 10864
rect 0 10780 1708 10836
rect 1764 10780 2492 10836
rect 2548 10780 2558 10836
rect 0 10752 800 10780
rect 3332 10724 3388 10892
rect 6066 10780 6076 10836
rect 6132 10780 7644 10836
rect 7700 10780 7710 10836
rect 14242 10780 14252 10836
rect 14308 10780 15036 10836
rect 15092 10780 15102 10836
rect 35410 10780 35420 10836
rect 35476 10780 37436 10836
rect 37492 10780 38220 10836
rect 38276 10780 38286 10836
rect 47842 10780 47852 10836
rect 47908 10780 49868 10836
rect 49924 10780 49934 10836
rect 53218 10780 53228 10836
rect 53284 10780 54012 10836
rect 54068 10780 54078 10836
rect 3332 10668 4844 10724
rect 4900 10668 6188 10724
rect 6244 10668 6254 10724
rect 14914 10668 14924 10724
rect 14980 10668 16604 10724
rect 16660 10668 16670 10724
rect 32498 10668 32508 10724
rect 32564 10668 34076 10724
rect 34132 10668 34142 10724
rect 37874 10668 37884 10724
rect 37940 10668 40572 10724
rect 40628 10668 42476 10724
rect 42532 10668 42542 10724
rect 45490 10668 45500 10724
rect 45556 10668 46060 10724
rect 46116 10668 47404 10724
rect 47460 10668 47470 10724
rect 52882 10668 52892 10724
rect 52948 10668 53788 10724
rect 53844 10668 53854 10724
rect 10098 10556 10108 10612
rect 10164 10556 10892 10612
rect 10948 10556 10958 10612
rect 17042 10556 17052 10612
rect 17108 10556 17836 10612
rect 17892 10556 17902 10612
rect 18274 10556 18284 10612
rect 18340 10556 19404 10612
rect 19460 10556 19470 10612
rect 34290 10556 34300 10612
rect 34356 10556 36428 10612
rect 36484 10556 36494 10612
rect 43362 10556 43372 10612
rect 43428 10556 44940 10612
rect 44996 10556 47852 10612
rect 47908 10556 47918 10612
rect 11554 10444 11564 10500
rect 11620 10444 12124 10500
rect 12180 10444 12190 10500
rect 31938 10444 31948 10500
rect 32004 10444 33068 10500
rect 33124 10444 33134 10500
rect 37762 10444 37772 10500
rect 37828 10444 41468 10500
rect 41524 10444 41534 10500
rect 28130 10332 28140 10388
rect 28196 10332 29372 10388
rect 29428 10332 29438 10388
rect 38546 10220 38556 10276
rect 38612 10220 38668 10444
rect 53442 10332 53452 10388
rect 53508 10332 54012 10388
rect 54068 10332 54078 10388
rect 0 10164 800 10192
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 0 10108 1708 10164
rect 1764 10108 2492 10164
rect 2548 10108 2558 10164
rect 10434 10108 10444 10164
rect 10500 10108 12796 10164
rect 12852 10108 12862 10164
rect 37986 10108 37996 10164
rect 38052 10108 38444 10164
rect 38500 10108 38510 10164
rect 0 10080 800 10108
rect 23986 9996 23996 10052
rect 24052 9996 25452 10052
rect 25508 9996 25900 10052
rect 25956 9996 25966 10052
rect 32946 9996 32956 10052
rect 33012 9996 35420 10052
rect 35476 9996 35486 10052
rect 23426 9884 23436 9940
rect 23492 9884 24108 9940
rect 24164 9884 24780 9940
rect 24836 9884 24846 9940
rect 25900 9884 27916 9940
rect 27972 9884 27982 9940
rect 28354 9884 28364 9940
rect 28420 9884 29260 9940
rect 29316 9884 29326 9940
rect 33394 9884 33404 9940
rect 33460 9884 34860 9940
rect 34916 9884 34926 9940
rect 38882 9884 38892 9940
rect 38948 9884 41132 9940
rect 41188 9884 41198 9940
rect 41570 9884 41580 9940
rect 41636 9884 43148 9940
rect 43204 9884 44156 9940
rect 44212 9884 44222 9940
rect 51202 9884 51212 9940
rect 51268 9884 53676 9940
rect 53732 9884 54684 9940
rect 54740 9884 54750 9940
rect 25900 9828 25956 9884
rect 10770 9772 10780 9828
rect 10836 9772 12796 9828
rect 12852 9772 15148 9828
rect 15204 9772 15214 9828
rect 15362 9772 15372 9828
rect 15428 9772 17052 9828
rect 17108 9772 17118 9828
rect 23650 9772 23660 9828
rect 23716 9772 25900 9828
rect 25956 9772 25966 9828
rect 26898 9772 26908 9828
rect 26964 9772 27580 9828
rect 27636 9772 27646 9828
rect 32274 9772 32284 9828
rect 32340 9772 35084 9828
rect 35140 9772 35150 9828
rect 35634 9772 35644 9828
rect 35700 9772 37548 9828
rect 37604 9772 38220 9828
rect 38276 9772 38286 9828
rect 43026 9772 43036 9828
rect 43092 9772 43484 9828
rect 43540 9772 43550 9828
rect 50082 9772 50092 9828
rect 50148 9772 52556 9828
rect 52612 9772 52622 9828
rect 53106 9772 53116 9828
rect 53172 9772 54124 9828
rect 54180 9772 54190 9828
rect 13682 9660 13692 9716
rect 13748 9660 14476 9716
rect 14532 9660 15484 9716
rect 15540 9660 15550 9716
rect 15810 9660 15820 9716
rect 15876 9660 16940 9716
rect 16996 9660 17006 9716
rect 24322 9660 24332 9716
rect 24388 9660 26236 9716
rect 26292 9660 27356 9716
rect 27412 9660 27422 9716
rect 28578 9660 28588 9716
rect 28644 9660 29148 9716
rect 29204 9660 29214 9716
rect 32162 9660 32172 9716
rect 32228 9660 32732 9716
rect 32788 9660 32798 9716
rect 34738 9660 34748 9716
rect 34804 9660 37100 9716
rect 37156 9660 37166 9716
rect 37874 9660 37884 9716
rect 37940 9660 39228 9716
rect 39284 9660 39294 9716
rect 16370 9548 16380 9604
rect 16436 9548 17724 9604
rect 17780 9548 17790 9604
rect 32274 9548 32284 9604
rect 32340 9548 33740 9604
rect 33796 9548 33806 9604
rect 35410 9548 35420 9604
rect 35476 9548 39004 9604
rect 39060 9548 39070 9604
rect 30706 9436 30716 9492
rect 30772 9436 31164 9492
rect 31220 9436 31230 9492
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 50546 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50830 9436
rect 31042 9324 31052 9380
rect 31108 9324 32060 9380
rect 32116 9324 32452 9380
rect 32610 9324 32620 9380
rect 32676 9324 33964 9380
rect 34020 9324 34030 9380
rect 32396 9268 32452 9324
rect 5618 9212 5628 9268
rect 5684 9212 6300 9268
rect 6356 9212 6748 9268
rect 6804 9212 6814 9268
rect 7970 9212 7980 9268
rect 8036 9212 9100 9268
rect 9156 9212 9548 9268
rect 9604 9212 9614 9268
rect 15250 9212 15260 9268
rect 15316 9212 15820 9268
rect 15876 9212 15886 9268
rect 17826 9212 17836 9268
rect 17892 9212 19180 9268
rect 19236 9212 19246 9268
rect 19506 9212 19516 9268
rect 19572 9212 21532 9268
rect 21588 9212 24892 9268
rect 24948 9212 26012 9268
rect 26068 9212 26078 9268
rect 27682 9212 27692 9268
rect 27748 9212 28476 9268
rect 28532 9212 28542 9268
rect 30818 9212 30828 9268
rect 30884 9212 32172 9268
rect 32228 9212 32238 9268
rect 32396 9212 35196 9268
rect 35252 9212 36540 9268
rect 36596 9212 36606 9268
rect 37874 9212 37884 9268
rect 37940 9212 38668 9268
rect 38724 9212 40012 9268
rect 40068 9212 40078 9268
rect 48178 9212 48188 9268
rect 48244 9212 48860 9268
rect 48916 9212 48926 9268
rect 50372 9212 51884 9268
rect 51940 9212 53228 9268
rect 53284 9212 53900 9268
rect 53956 9212 53966 9268
rect 17836 9156 17892 9212
rect 50372 9156 50428 9212
rect 2034 9100 2044 9156
rect 2100 9100 7084 9156
rect 7140 9100 7644 9156
rect 7700 9100 8652 9156
rect 8708 9100 8718 9156
rect 15138 9100 15148 9156
rect 15204 9100 17892 9156
rect 37202 9100 37212 9156
rect 37268 9100 37772 9156
rect 37828 9100 39004 9156
rect 39060 9100 39340 9156
rect 39396 9100 39788 9156
rect 39844 9100 39854 9156
rect 40338 9100 40348 9156
rect 40404 9100 41244 9156
rect 41300 9100 41310 9156
rect 46050 9100 46060 9156
rect 46116 9100 47180 9156
rect 47236 9100 50428 9156
rect 51212 9100 52108 9156
rect 52164 9100 52174 9156
rect 8866 8988 8876 9044
rect 8932 8988 10108 9044
rect 10164 8988 10174 9044
rect 22082 8988 22092 9044
rect 22148 8988 23660 9044
rect 23716 8988 24220 9044
rect 24276 8988 25228 9044
rect 25284 8988 25294 9044
rect 34178 8988 34188 9044
rect 34244 8988 35868 9044
rect 35924 8988 35934 9044
rect 41010 8988 41020 9044
rect 41076 8988 43260 9044
rect 43316 8988 43326 9044
rect 43474 8988 43484 9044
rect 43540 8988 44940 9044
rect 44996 8988 45006 9044
rect 51212 8932 51268 9100
rect 51538 8988 51548 9044
rect 51604 8988 52892 9044
rect 52948 8988 52958 9044
rect 15922 8876 15932 8932
rect 15988 8876 17500 8932
rect 17556 8876 17566 8932
rect 40114 8876 40124 8932
rect 40180 8876 40908 8932
rect 40964 8876 40974 8932
rect 49634 8876 49644 8932
rect 49700 8876 51268 8932
rect 0 8820 800 8848
rect 0 8764 1708 8820
rect 1764 8764 2492 8820
rect 2548 8764 2558 8820
rect 16706 8764 16716 8820
rect 16772 8764 17948 8820
rect 18004 8764 18014 8820
rect 31378 8764 31388 8820
rect 31444 8764 32284 8820
rect 32340 8764 32350 8820
rect 47394 8764 47404 8820
rect 47460 8764 48972 8820
rect 49028 8764 49980 8820
rect 50036 8764 50428 8820
rect 50484 8764 50494 8820
rect 0 8736 800 8764
rect 29474 8652 29484 8708
rect 29540 8652 33628 8708
rect 33684 8652 34524 8708
rect 34580 8652 34590 8708
rect 44818 8652 44828 8708
rect 44884 8652 46396 8708
rect 46452 8652 50036 8708
rect 52546 8652 52556 8708
rect 52612 8652 53340 8708
rect 53396 8652 53406 8708
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 49980 8596 50036 8652
rect 49186 8540 49196 8596
rect 49252 8540 49262 8596
rect 49970 8540 49980 8596
rect 50036 8540 50046 8596
rect 49196 8484 49252 8540
rect 6178 8428 6188 8484
rect 6244 8428 9212 8484
rect 9268 8428 9278 8484
rect 20066 8428 20076 8484
rect 20132 8428 21868 8484
rect 21924 8428 21934 8484
rect 33730 8428 33740 8484
rect 33796 8428 34412 8484
rect 34468 8428 36204 8484
rect 36260 8428 36270 8484
rect 38098 8428 38108 8484
rect 38164 8428 39452 8484
rect 39508 8428 39518 8484
rect 43138 8428 43148 8484
rect 43204 8428 45276 8484
rect 45332 8428 45342 8484
rect 46834 8428 46844 8484
rect 46900 8428 49532 8484
rect 49588 8428 49756 8484
rect 49812 8428 49822 8484
rect 48300 8372 48356 8428
rect 8642 8316 8652 8372
rect 8708 8316 9548 8372
rect 9604 8316 9614 8372
rect 9986 8316 9996 8372
rect 10052 8316 11228 8372
rect 11284 8316 11294 8372
rect 12338 8316 12348 8372
rect 12404 8316 13020 8372
rect 13076 8316 13804 8372
rect 13860 8316 13870 8372
rect 22866 8316 22876 8372
rect 22932 8316 26572 8372
rect 26628 8316 26638 8372
rect 28466 8316 28476 8372
rect 28532 8316 29372 8372
rect 29428 8316 29820 8372
rect 29876 8316 29886 8372
rect 30482 8316 30492 8372
rect 30548 8316 31836 8372
rect 31892 8316 31902 8372
rect 36418 8316 36428 8372
rect 36484 8316 37100 8372
rect 37156 8316 37166 8372
rect 37314 8316 37324 8372
rect 37380 8316 40796 8372
rect 40852 8316 42924 8372
rect 42980 8316 45724 8372
rect 45780 8316 45790 8372
rect 48290 8316 48300 8372
rect 48356 8316 48366 8372
rect 51426 8316 51436 8372
rect 51492 8316 52556 8372
rect 52612 8316 52622 8372
rect 53442 8316 53452 8372
rect 53508 8316 54012 8372
rect 54068 8316 54078 8372
rect 6962 8204 6972 8260
rect 7028 8204 7644 8260
rect 7700 8204 8764 8260
rect 8820 8204 8830 8260
rect 10994 8204 11004 8260
rect 11060 8204 11788 8260
rect 11844 8204 13580 8260
rect 13636 8204 13646 8260
rect 21746 8204 21756 8260
rect 21812 8204 22428 8260
rect 22484 8204 23436 8260
rect 23492 8204 23502 8260
rect 24434 8204 24444 8260
rect 24500 8204 25564 8260
rect 25620 8204 25630 8260
rect 28354 8204 28364 8260
rect 28420 8204 30268 8260
rect 30324 8204 30334 8260
rect 30594 8204 30604 8260
rect 30660 8204 31388 8260
rect 31444 8204 31454 8260
rect 33730 8204 33740 8260
rect 33796 8204 35756 8260
rect 35812 8204 37772 8260
rect 37828 8204 37838 8260
rect 40002 8204 40012 8260
rect 40068 8204 41132 8260
rect 41188 8204 41198 8260
rect 42578 8204 42588 8260
rect 42644 8204 43484 8260
rect 43540 8204 45276 8260
rect 45332 8204 45342 8260
rect 47282 8204 47292 8260
rect 47348 8204 50876 8260
rect 50932 8204 50942 8260
rect 51762 8204 51772 8260
rect 51828 8204 53900 8260
rect 53956 8204 53966 8260
rect 8306 8092 8316 8148
rect 8372 8092 9660 8148
rect 9716 8092 9726 8148
rect 15474 8092 15484 8148
rect 15540 8092 16268 8148
rect 16324 8092 17836 8148
rect 17892 8092 17902 8148
rect 26786 8092 26796 8148
rect 26852 8092 29148 8148
rect 29204 8092 29214 8148
rect 42018 8092 42028 8148
rect 42084 8092 43708 8148
rect 43764 8092 45052 8148
rect 45108 8092 45724 8148
rect 45780 8092 45790 8148
rect 52994 8092 53004 8148
rect 53060 8092 54236 8148
rect 54292 8092 54302 8148
rect 9202 7980 9212 8036
rect 9268 7980 12684 8036
rect 12740 7980 12750 8036
rect 13010 7980 13020 8036
rect 13076 7980 14140 8036
rect 14196 7980 14206 8036
rect 18274 7980 18284 8036
rect 18340 7980 20524 8036
rect 20580 7980 20590 8036
rect 34850 7980 34860 8036
rect 34916 7980 35532 8036
rect 35588 7980 36316 8036
rect 36372 7980 36382 8036
rect 41794 7980 41804 8036
rect 41860 7980 42700 8036
rect 42756 7980 43820 8036
rect 43876 7980 44716 8036
rect 44772 7980 44782 8036
rect 48962 7980 48972 8036
rect 49028 7980 49756 8036
rect 49812 7980 52892 8036
rect 52948 7980 53228 8036
rect 53284 7980 53788 8036
rect 53844 7980 53854 8036
rect 8978 7868 8988 7924
rect 9044 7868 11900 7924
rect 11956 7868 12796 7924
rect 12852 7868 14924 7924
rect 14980 7868 14990 7924
rect 48290 7868 48300 7924
rect 48356 7868 48860 7924
rect 48916 7868 48926 7924
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 50546 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50830 7868
rect 15372 7756 15596 7812
rect 15652 7756 15662 7812
rect 39778 7756 39788 7812
rect 39844 7756 40460 7812
rect 40516 7756 40526 7812
rect 15372 7700 15428 7756
rect 8754 7644 8764 7700
rect 8820 7644 9548 7700
rect 9604 7644 9614 7700
rect 15362 7644 15372 7700
rect 15428 7644 15438 7700
rect 23548 7644 28028 7700
rect 28084 7644 28094 7700
rect 41122 7644 41132 7700
rect 41188 7644 43372 7700
rect 43428 7644 44380 7700
rect 44436 7644 44446 7700
rect 45714 7644 45724 7700
rect 45780 7644 47068 7700
rect 47124 7644 47134 7700
rect 47618 7644 47628 7700
rect 47684 7644 48748 7700
rect 48804 7644 48814 7700
rect 50754 7644 50764 7700
rect 50820 7644 51100 7700
rect 51156 7644 51166 7700
rect 9314 7532 9324 7588
rect 9380 7532 11788 7588
rect 11844 7532 12348 7588
rect 12404 7532 12414 7588
rect 12674 7532 12684 7588
rect 12740 7532 19404 7588
rect 19460 7532 20300 7588
rect 20356 7532 20366 7588
rect 23548 7476 23604 7644
rect 26562 7532 26572 7588
rect 26628 7532 27804 7588
rect 27860 7532 27870 7588
rect 31378 7532 31388 7588
rect 31444 7532 33068 7588
rect 33124 7532 34300 7588
rect 34356 7532 34366 7588
rect 40226 7532 40236 7588
rect 40292 7532 42252 7588
rect 42308 7532 42318 7588
rect 50194 7532 50204 7588
rect 50260 7532 52444 7588
rect 52500 7532 52510 7588
rect 15092 7420 16044 7476
rect 16100 7420 16110 7476
rect 16594 7420 16604 7476
rect 16660 7420 18172 7476
rect 18228 7420 18238 7476
rect 19954 7420 19964 7476
rect 20020 7420 23548 7476
rect 23604 7420 23614 7476
rect 25442 7420 25452 7476
rect 25508 7420 27244 7476
rect 27300 7420 27310 7476
rect 28130 7420 28140 7476
rect 28196 7420 29148 7476
rect 29204 7420 30604 7476
rect 30660 7420 30670 7476
rect 31938 7420 31948 7476
rect 32004 7420 33292 7476
rect 33348 7420 34076 7476
rect 34132 7420 34142 7476
rect 36418 7420 36428 7476
rect 36484 7420 36988 7476
rect 37044 7420 37548 7476
rect 37604 7420 37614 7476
rect 38994 7420 39004 7476
rect 39060 7420 39452 7476
rect 39508 7420 39518 7476
rect 39890 7420 39900 7476
rect 39956 7420 43932 7476
rect 43988 7420 43998 7476
rect 46834 7420 46844 7476
rect 46900 7420 48076 7476
rect 48132 7420 48142 7476
rect 49410 7420 49420 7476
rect 49476 7420 51436 7476
rect 51492 7420 51502 7476
rect 15092 7364 15148 7420
rect 39452 7364 39508 7420
rect 14242 7308 14252 7364
rect 14308 7308 15148 7364
rect 26002 7308 26012 7364
rect 26068 7308 27020 7364
rect 27076 7308 27692 7364
rect 27748 7308 27758 7364
rect 28914 7308 28924 7364
rect 28980 7308 30268 7364
rect 30324 7308 30334 7364
rect 39452 7308 41468 7364
rect 41524 7308 41534 7364
rect 42130 7308 42140 7364
rect 42196 7308 43820 7364
rect 43876 7308 43886 7364
rect 46050 7308 46060 7364
rect 46116 7308 47964 7364
rect 48020 7308 48030 7364
rect 9090 7196 9100 7252
rect 9156 7196 9772 7252
rect 9828 7196 9838 7252
rect 10994 7196 11004 7252
rect 11060 7196 12236 7252
rect 12292 7196 12302 7252
rect 33506 7196 33516 7252
rect 33572 7196 34636 7252
rect 34692 7196 35308 7252
rect 35364 7196 36540 7252
rect 36596 7196 36606 7252
rect 38434 7196 38444 7252
rect 38500 7196 40684 7252
rect 40740 7196 40750 7252
rect 42242 7196 42252 7252
rect 42308 7196 42924 7252
rect 42980 7196 42990 7252
rect 38210 7084 38220 7140
rect 38276 7084 40516 7140
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 38546 6972 38556 7028
rect 38612 6972 40236 7028
rect 40292 6972 40302 7028
rect 40460 6916 40516 7084
rect 37426 6860 37436 6916
rect 37492 6860 38668 6916
rect 38724 6860 38734 6916
rect 40460 6860 43932 6916
rect 43988 6860 43998 6916
rect 50866 6860 50876 6916
rect 50932 6860 53004 6916
rect 53060 6860 53452 6916
rect 53508 6860 53518 6916
rect 11666 6748 11676 6804
rect 11732 6748 13132 6804
rect 13188 6748 13580 6804
rect 13636 6748 13646 6804
rect 18050 6748 18060 6804
rect 18116 6748 22204 6804
rect 22260 6748 22270 6804
rect 23986 6748 23996 6804
rect 24052 6748 26348 6804
rect 26404 6748 28924 6804
rect 28980 6748 28990 6804
rect 35858 6748 35868 6804
rect 35924 6748 37212 6804
rect 37268 6748 37278 6804
rect 42690 6748 42700 6804
rect 42756 6748 44940 6804
rect 44996 6748 45006 6804
rect 12450 6636 12460 6692
rect 12516 6636 16492 6692
rect 16548 6636 16558 6692
rect 17266 6636 17276 6692
rect 17332 6636 18732 6692
rect 18788 6636 19404 6692
rect 19460 6636 19470 6692
rect 20514 6636 20524 6692
rect 20580 6636 22092 6692
rect 22148 6636 22158 6692
rect 22530 6636 22540 6692
rect 22596 6636 24108 6692
rect 24164 6636 24174 6692
rect 30930 6636 30940 6692
rect 30996 6636 32396 6692
rect 32452 6636 32462 6692
rect 34290 6636 34300 6692
rect 34356 6636 35084 6692
rect 35140 6636 35150 6692
rect 39106 6636 39116 6692
rect 39172 6636 39452 6692
rect 39508 6636 39518 6692
rect 43138 6636 43148 6692
rect 43204 6636 44156 6692
rect 44212 6636 45388 6692
rect 45444 6636 45454 6692
rect 47282 6636 47292 6692
rect 47348 6636 49308 6692
rect 49364 6636 49374 6692
rect 50418 6636 50428 6692
rect 50484 6636 51436 6692
rect 51492 6636 51502 6692
rect 16156 6580 16212 6636
rect 11330 6524 11340 6580
rect 11396 6524 12348 6580
rect 12404 6524 12414 6580
rect 16146 6524 16156 6580
rect 16212 6524 16222 6580
rect 22418 6524 22428 6580
rect 22484 6524 23660 6580
rect 23716 6524 24780 6580
rect 24836 6524 24846 6580
rect 30482 6524 30492 6580
rect 30548 6524 32732 6580
rect 32788 6524 35644 6580
rect 35700 6524 41020 6580
rect 41076 6524 41086 6580
rect 47506 6524 47516 6580
rect 47572 6524 49532 6580
rect 49588 6524 50316 6580
rect 50372 6524 50382 6580
rect 11778 6412 11788 6468
rect 11844 6412 12572 6468
rect 12628 6412 15148 6468
rect 15204 6412 15214 6468
rect 16482 6412 16492 6468
rect 16548 6412 17724 6468
rect 17780 6412 17790 6468
rect 17948 6412 20188 6468
rect 20244 6412 25340 6468
rect 25396 6412 25406 6468
rect 33842 6412 33852 6468
rect 33908 6412 34636 6468
rect 34692 6412 36428 6468
rect 36484 6412 36494 6468
rect 42130 6412 42140 6468
rect 42196 6412 45612 6468
rect 45668 6412 45678 6468
rect 46050 6412 46060 6468
rect 46116 6412 47068 6468
rect 47124 6412 47134 6468
rect 50372 6412 50540 6468
rect 50596 6412 50606 6468
rect 17948 6356 18004 6412
rect 15250 6300 15260 6356
rect 15316 6300 18004 6356
rect 31042 6300 31052 6356
rect 31108 6300 32060 6356
rect 32116 6300 36204 6356
rect 36260 6300 42924 6356
rect 42980 6300 42990 6356
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 37090 6188 37100 6244
rect 37156 6188 41356 6244
rect 41412 6188 41422 6244
rect 50372 6132 50428 6412
rect 50546 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50830 6300
rect 33506 6076 33516 6132
rect 33572 6076 36316 6132
rect 36372 6076 36382 6132
rect 39218 6076 39228 6132
rect 39284 6076 40908 6132
rect 40964 6076 40974 6132
rect 49858 6076 49868 6132
rect 49924 6076 52220 6132
rect 52276 6076 52668 6132
rect 52724 6076 52734 6132
rect 11554 5964 11564 6020
rect 11620 5964 12348 6020
rect 12404 5964 12414 6020
rect 34178 5964 34188 6020
rect 34244 5964 39788 6020
rect 39844 5964 39854 6020
rect 42578 5964 42588 6020
rect 42644 5964 43596 6020
rect 43652 5964 44604 6020
rect 44660 5964 44670 6020
rect 20738 5852 20748 5908
rect 20804 5852 21644 5908
rect 21700 5852 21710 5908
rect 30930 5852 30940 5908
rect 30996 5852 33740 5908
rect 33796 5852 33806 5908
rect 34402 5852 34412 5908
rect 34468 5852 38668 5908
rect 41906 5852 41916 5908
rect 41972 5852 44044 5908
rect 44100 5852 44110 5908
rect 48962 5852 48972 5908
rect 49028 5852 50204 5908
rect 50260 5852 51324 5908
rect 51380 5852 51390 5908
rect 38612 5796 38668 5852
rect 18386 5740 18396 5796
rect 18452 5740 20860 5796
rect 20916 5740 20926 5796
rect 32162 5740 32172 5796
rect 32228 5740 35868 5796
rect 35924 5740 35934 5796
rect 38612 5740 39564 5796
rect 39620 5740 39630 5796
rect 41122 5740 41132 5796
rect 41188 5740 42476 5796
rect 42532 5740 42542 5796
rect 45154 5740 45164 5796
rect 45220 5740 46396 5796
rect 46452 5740 46462 5796
rect 46620 5740 49868 5796
rect 49924 5740 49934 5796
rect 46620 5684 46676 5740
rect 31826 5628 31836 5684
rect 31892 5628 34524 5684
rect 34580 5628 34590 5684
rect 43810 5628 43820 5684
rect 43876 5628 44380 5684
rect 44436 5628 45948 5684
rect 46004 5628 46620 5684
rect 46676 5628 46686 5684
rect 48850 5628 48860 5684
rect 48916 5628 49980 5684
rect 50036 5628 50046 5684
rect 50306 5628 50316 5684
rect 50372 5628 52108 5684
rect 52164 5628 52174 5684
rect 20514 5516 20524 5572
rect 20580 5516 21868 5572
rect 21924 5516 21934 5572
rect 30930 5516 30940 5572
rect 30996 5516 34300 5572
rect 34356 5516 34366 5572
rect 43698 5516 43708 5572
rect 43764 5516 45836 5572
rect 45892 5516 45902 5572
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 30034 5404 30044 5460
rect 30100 5404 32172 5460
rect 32228 5404 32238 5460
rect 39330 5404 39340 5460
rect 39396 5404 43932 5460
rect 43988 5404 43998 5460
rect 31948 5292 33068 5348
rect 33124 5292 33134 5348
rect 35746 5292 35756 5348
rect 35812 5292 39004 5348
rect 39060 5292 40236 5348
rect 40292 5292 40302 5348
rect 43474 5292 43484 5348
rect 43540 5292 45164 5348
rect 45220 5292 47964 5348
rect 48020 5292 49084 5348
rect 49140 5292 49150 5348
rect 31948 5236 32004 5292
rect 28578 5180 28588 5236
rect 28644 5180 31500 5236
rect 31556 5180 31948 5236
rect 32004 5180 32014 5236
rect 32274 5180 32284 5236
rect 32340 5180 33516 5236
rect 33572 5180 33582 5236
rect 36418 5180 36428 5236
rect 36484 5180 36764 5236
rect 36820 5180 38668 5236
rect 39218 5180 39228 5236
rect 39284 5180 44156 5236
rect 44212 5180 44222 5236
rect 38612 5124 38668 5180
rect 28354 5068 28364 5124
rect 28420 5068 29260 5124
rect 29316 5068 29326 5124
rect 29698 5068 29708 5124
rect 29764 5068 29876 5124
rect 30034 5068 30044 5124
rect 30100 5068 31612 5124
rect 31668 5068 32060 5124
rect 32116 5068 32126 5124
rect 35746 5068 35756 5124
rect 35812 5068 36652 5124
rect 36708 5068 36718 5124
rect 38612 5068 38892 5124
rect 38948 5068 38958 5124
rect 39442 5068 39452 5124
rect 39508 5068 40348 5124
rect 40404 5068 40414 5124
rect 40562 5068 40572 5124
rect 40628 5068 41468 5124
rect 41524 5068 41534 5124
rect 43810 5068 43820 5124
rect 43876 5068 44828 5124
rect 44884 5068 44894 5124
rect 45938 5068 45948 5124
rect 46004 5068 47180 5124
rect 47236 5068 47246 5124
rect 48066 5068 48076 5124
rect 48132 5068 48412 5124
rect 48468 5068 49980 5124
rect 50036 5068 50046 5124
rect 29820 5012 29876 5068
rect 29820 4956 30492 5012
rect 30548 4956 35084 5012
rect 35140 4956 35150 5012
rect 44258 4956 44268 5012
rect 44324 4956 45612 5012
rect 45668 4956 45678 5012
rect 28690 4844 28700 4900
rect 28756 4844 30380 4900
rect 30436 4844 31724 4900
rect 31780 4844 31790 4900
rect 34514 4844 34524 4900
rect 34580 4844 35980 4900
rect 36036 4844 36046 4900
rect 36194 4844 36204 4900
rect 36260 4844 43260 4900
rect 43316 4844 43820 4900
rect 43876 4844 43886 4900
rect 29250 4732 29260 4788
rect 29316 4732 32956 4788
rect 33012 4732 33022 4788
rect 34402 4732 34412 4788
rect 34468 4732 39116 4788
rect 39172 4732 39182 4788
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 32162 4508 32172 4564
rect 32228 4508 32238 4564
rect 36306 4508 36316 4564
rect 36372 4508 39228 4564
rect 39284 4508 39294 4564
rect 32172 4452 32228 4508
rect 32172 4396 34860 4452
rect 34916 4396 40908 4452
rect 40964 4396 40974 4452
rect 42252 4340 42308 4844
rect 43026 4732 43036 4788
rect 43092 4732 45388 4788
rect 45444 4732 45454 4788
rect 50546 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50830 4732
rect 42914 4508 42924 4564
rect 42980 4508 43596 4564
rect 43652 4508 43662 4564
rect 43148 4396 46396 4452
rect 46452 4396 47404 4452
rect 47460 4396 47470 4452
rect 43148 4340 43204 4396
rect 33954 4284 33964 4340
rect 34020 4284 36988 4340
rect 37044 4284 37054 4340
rect 42252 4284 42700 4340
rect 42756 4284 42766 4340
rect 43138 4284 43148 4340
rect 43204 4284 43214 4340
rect 45602 4284 45612 4340
rect 45668 4284 46284 4340
rect 46340 4284 46350 4340
rect 42018 4172 42028 4228
rect 42084 4172 43372 4228
rect 43428 4172 43438 4228
rect 45938 4172 45948 4228
rect 46004 4172 48188 4228
rect 48244 4172 48254 4228
rect 28466 4060 28476 4116
rect 28532 4060 29484 4116
rect 29540 4060 29550 4116
rect 33618 4060 33628 4116
rect 33684 4060 41132 4116
rect 41188 4060 41198 4116
rect 37650 3948 37660 4004
rect 37716 3948 44940 4004
rect 44996 3948 47292 4004
rect 47348 3948 47358 4004
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 36306 3836 36316 3892
rect 36372 3836 44492 3892
rect 44548 3836 47740 3892
rect 47796 3836 47806 3892
rect 34962 3724 34972 3780
rect 35028 3724 42140 3780
rect 42196 3724 42206 3780
rect 43922 3724 43932 3780
rect 43988 3724 46844 3780
rect 46900 3724 46910 3780
rect 30258 3612 30268 3668
rect 30324 3612 32396 3668
rect 32452 3612 32462 3668
rect 35634 3612 35644 3668
rect 35700 3612 36988 3668
rect 37044 3612 37054 3668
rect 38994 3612 39004 3668
rect 39060 3612 41804 3668
rect 41860 3612 41870 3668
rect 43138 3612 43148 3668
rect 43204 3612 47628 3668
rect 47684 3612 49308 3668
rect 49364 3612 49374 3668
rect 31602 3500 31612 3556
rect 31668 3500 32620 3556
rect 32676 3500 35308 3556
rect 35364 3500 35374 3556
rect 38322 3500 38332 3556
rect 38388 3500 45164 3556
rect 45220 3500 45230 3556
rect 47282 3500 47292 3556
rect 47348 3500 48188 3556
rect 48244 3500 48860 3556
rect 48916 3500 48926 3556
rect 45164 3444 45220 3500
rect 28354 3388 28364 3444
rect 28420 3388 30940 3444
rect 30996 3388 31006 3444
rect 38994 3388 39004 3444
rect 39060 3388 45108 3444
rect 45164 3388 48748 3444
rect 48804 3388 48814 3444
rect 45052 3332 45108 3388
rect 35970 3276 35980 3332
rect 36036 3276 43484 3332
rect 43540 3276 43550 3332
rect 45052 3276 45948 3332
rect 46004 3276 46014 3332
rect 32162 3164 32172 3220
rect 32228 3164 35532 3220
rect 35588 3164 42700 3220
rect 42756 3164 42766 3220
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 50546 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50830 3164
rect 39666 2604 39676 2660
rect 39732 2604 46508 2660
rect 46564 2604 46574 2660
rect 34290 2492 34300 2548
rect 34356 2492 43932 2548
rect 43988 2492 43998 2548
<< via3 >>
rect 19836 56420 19892 56476
rect 19940 56420 19996 56476
rect 20044 56420 20100 56476
rect 50556 56420 50612 56476
rect 50660 56420 50716 56476
rect 50764 56420 50820 56476
rect 4476 55636 4532 55692
rect 4580 55636 4636 55692
rect 4684 55636 4740 55692
rect 35196 55636 35252 55692
rect 35300 55636 35356 55692
rect 35404 55636 35460 55692
rect 19836 54852 19892 54908
rect 19940 54852 19996 54908
rect 20044 54852 20100 54908
rect 50556 54852 50612 54908
rect 50660 54852 50716 54908
rect 50764 54852 50820 54908
rect 32508 54460 32564 54516
rect 4476 54068 4532 54124
rect 4580 54068 4636 54124
rect 4684 54068 4740 54124
rect 35196 54068 35252 54124
rect 35300 54068 35356 54124
rect 35404 54068 35460 54124
rect 19836 53284 19892 53340
rect 19940 53284 19996 53340
rect 20044 53284 20100 53340
rect 50556 53284 50612 53340
rect 50660 53284 50716 53340
rect 50764 53284 50820 53340
rect 4476 52500 4532 52556
rect 4580 52500 4636 52556
rect 4684 52500 4740 52556
rect 35196 52500 35252 52556
rect 35300 52500 35356 52556
rect 35404 52500 35460 52556
rect 19836 51716 19892 51772
rect 19940 51716 19996 51772
rect 20044 51716 20100 51772
rect 50556 51716 50612 51772
rect 50660 51716 50716 51772
rect 50764 51716 50820 51772
rect 4476 50932 4532 50988
rect 4580 50932 4636 50988
rect 4684 50932 4740 50988
rect 35196 50932 35252 50988
rect 35300 50932 35356 50988
rect 35404 50932 35460 50988
rect 19836 50148 19892 50204
rect 19940 50148 19996 50204
rect 20044 50148 20100 50204
rect 50556 50148 50612 50204
rect 50660 50148 50716 50204
rect 50764 50148 50820 50204
rect 2828 49644 2884 49700
rect 4476 49364 4532 49420
rect 4580 49364 4636 49420
rect 4684 49364 4740 49420
rect 35196 49364 35252 49420
rect 35300 49364 35356 49420
rect 35404 49364 35460 49420
rect 3388 49196 3444 49252
rect 3500 48860 3556 48916
rect 3836 48860 3892 48916
rect 19836 48580 19892 48636
rect 19940 48580 19996 48636
rect 20044 48580 20100 48636
rect 50556 48580 50612 48636
rect 50660 48580 50716 48636
rect 50764 48580 50820 48636
rect 3500 48076 3556 48132
rect 4476 47796 4532 47852
rect 4580 47796 4636 47852
rect 4684 47796 4740 47852
rect 35196 47796 35252 47852
rect 35300 47796 35356 47852
rect 35404 47796 35460 47852
rect 3388 47404 3444 47460
rect 3836 47068 3892 47124
rect 19836 47012 19892 47068
rect 19940 47012 19996 47068
rect 20044 47012 20100 47068
rect 50556 47012 50612 47068
rect 50660 47012 50716 47068
rect 50764 47012 50820 47068
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 50556 45444 50612 45500
rect 50660 45444 50716 45500
rect 50764 45444 50820 45500
rect 3388 45276 3444 45332
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 26572 44044 26628 44100
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 50556 43876 50612 43932
rect 50660 43876 50716 43932
rect 50764 43876 50820 43932
rect 6860 43708 6916 43764
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 50556 42308 50612 42364
rect 50660 42308 50716 42364
rect 50764 42308 50820 42364
rect 2828 41916 2884 41972
rect 25676 41804 25732 41860
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 50556 40740 50612 40796
rect 50660 40740 50716 40796
rect 50764 40740 50820 40796
rect 32508 40236 32564 40292
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 48860 39788 48916 39844
rect 48860 39228 48916 39284
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 50556 39172 50612 39228
rect 50660 39172 50716 39228
rect 50764 39172 50820 39228
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 6860 38108 6916 38164
rect 25676 37660 25732 37716
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 50556 37604 50612 37660
rect 50660 37604 50716 37660
rect 50764 37604 50820 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 26572 36764 26628 36820
rect 2156 36540 2212 36596
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 50556 36036 50612 36092
rect 50660 36036 50716 36092
rect 50764 36036 50820 36092
rect 3276 35420 3332 35476
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 2156 35196 2212 35252
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 3276 34860 3332 34916
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 50556 34468 50612 34524
rect 50660 34468 50716 34524
rect 50764 34468 50820 34524
rect 3724 34188 3780 34244
rect 32620 34076 32676 34132
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 3724 33516 3780 33572
rect 31948 33068 32004 33124
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 50556 32900 50612 32956
rect 50660 32900 50716 32956
rect 50764 32900 50820 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 50556 31332 50612 31388
rect 50660 31332 50716 31388
rect 50764 31332 50820 31388
rect 33292 31164 33348 31220
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 34972 29708 35028 29764
rect 50556 29764 50612 29820
rect 50660 29764 50716 29820
rect 50764 29764 50820 29820
rect 26460 29260 26516 29316
rect 33740 29260 33796 29316
rect 34860 29148 34916 29204
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 27692 28812 27748 28868
rect 32844 28364 32900 28420
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 50556 28196 50612 28252
rect 50660 28196 50716 28252
rect 50764 28196 50820 28252
rect 34636 27468 34692 27524
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 32172 27132 32228 27188
rect 32844 27132 32900 27188
rect 27692 27020 27748 27076
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 50556 26628 50612 26684
rect 50660 26628 50716 26684
rect 50764 26628 50820 26684
rect 23884 26572 23940 26628
rect 26460 26460 26516 26516
rect 32172 26348 32228 26404
rect 23884 25900 23940 25956
rect 31948 25900 32004 25956
rect 34524 25900 34580 25956
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 2044 25564 2100 25620
rect 32620 25452 32676 25508
rect 34972 25340 35028 25396
rect 34972 25116 35028 25172
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 50556 25060 50612 25116
rect 50660 25060 50716 25116
rect 50764 25060 50820 25116
rect 33740 25004 33796 25060
rect 34860 25004 34916 25060
rect 34636 24556 34692 24612
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 7420 23884 7476 23940
rect 34972 23884 35028 23940
rect 34524 23660 34580 23716
rect 34972 23660 35028 23716
rect 7420 23548 7476 23604
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 50556 23492 50612 23548
rect 50660 23492 50716 23548
rect 50764 23492 50820 23548
rect 34748 23212 34804 23268
rect 23772 22988 23828 23044
rect 34860 22876 34916 22932
rect 2380 22764 2436 22820
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 34748 22316 34804 22372
rect 3612 21980 3668 22036
rect 23772 21980 23828 22036
rect 30156 21980 30212 22036
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 2828 21868 2884 21924
rect 50556 21924 50612 21980
rect 50660 21924 50716 21980
rect 50764 21924 50820 21980
rect 3276 21644 3332 21700
rect 3276 21196 3332 21252
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 1820 20860 1876 20916
rect 6300 20860 6356 20916
rect 2828 20524 2884 20580
rect 4844 20524 4900 20580
rect 4060 20412 4116 20468
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 50556 20356 50612 20412
rect 50660 20356 50716 20412
rect 50764 20356 50820 20412
rect 3836 20076 3892 20132
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 1708 19516 1764 19572
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 50556 18788 50612 18844
rect 50660 18788 50716 18844
rect 50764 18788 50820 18844
rect 4060 18620 4116 18676
rect 33292 18620 33348 18676
rect 1820 18284 1876 18340
rect 3836 18284 3892 18340
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 2044 17500 2100 17556
rect 3612 17500 3668 17556
rect 4844 17500 4900 17556
rect 1708 17388 1764 17444
rect 34972 17388 35028 17444
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 50556 17220 50612 17276
rect 50660 17220 50716 17276
rect 50764 17220 50820 17276
rect 2380 17164 2436 17220
rect 28028 16828 28084 16884
rect 30156 16716 30212 16772
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 28588 16268 28644 16324
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 50556 15652 50612 15708
rect 50660 15652 50716 15708
rect 50764 15652 50820 15708
rect 34860 15036 34916 15092
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 50556 14084 50612 14140
rect 50660 14084 50716 14140
rect 50764 14084 50820 14140
rect 2828 13692 2884 13748
rect 28028 13468 28084 13524
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 6300 13020 6356 13076
rect 28588 13020 28644 13076
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 50556 12516 50612 12572
rect 50660 12516 50716 12572
rect 50764 12516 50820 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 50556 10948 50612 11004
rect 50660 10948 50716 11004
rect 50764 10948 50820 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 50556 9380 50612 9436
rect 50660 9380 50716 9436
rect 50764 9380 50820 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 50556 7812 50612 7868
rect 50660 7812 50716 7868
rect 50764 7812 50820 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 50556 6244 50612 6300
rect 50660 6244 50716 6300
rect 50764 6244 50820 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 50556 4676 50612 4732
rect 50660 4676 50716 4732
rect 50764 4676 50820 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
rect 50556 3108 50612 3164
rect 50660 3108 50716 3164
rect 50764 3108 50820 3164
<< metal4 >>
rect 4448 55692 4768 56508
rect 4448 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4768 55692
rect 4448 54124 4768 55636
rect 4448 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4768 54124
rect 4448 52556 4768 54068
rect 4448 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4768 52556
rect 4448 50988 4768 52500
rect 4448 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4768 50988
rect 2828 49700 2884 49710
rect 2828 41972 2884 49644
rect 4448 49420 4768 50932
rect 4448 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4768 49420
rect 3388 49252 3444 49262
rect 3388 47460 3444 49196
rect 3500 48916 3556 48926
rect 3500 48132 3556 48860
rect 3500 48066 3556 48076
rect 3836 48916 3892 48926
rect 3388 45332 3444 47404
rect 3836 47124 3892 48860
rect 3836 47058 3892 47068
rect 4448 47852 4768 49364
rect 4448 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4768 47852
rect 3388 45266 3444 45276
rect 4448 46284 4768 47796
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 2828 41906 2884 41916
rect 4448 44716 4768 46228
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 19808 56476 20128 56508
rect 19808 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20128 56476
rect 19808 54908 20128 56420
rect 19808 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20128 54908
rect 19808 53340 20128 54852
rect 35168 55692 35488 56508
rect 35168 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35488 55692
rect 19808 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20128 53340
rect 19808 51772 20128 53284
rect 19808 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20128 51772
rect 19808 50204 20128 51716
rect 19808 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20128 50204
rect 19808 48636 20128 50148
rect 19808 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20128 48636
rect 19808 47068 20128 48580
rect 19808 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20128 47068
rect 19808 45500 20128 47012
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 19808 43932 20128 45444
rect 32508 54516 32564 54526
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 6860 43764 6916 43774
rect 6860 38164 6916 43708
rect 6860 38098 6916 38108
rect 19808 42364 20128 43876
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 26572 44100 26628 44110
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 2156 36596 2212 36606
rect 2156 35252 2212 36540
rect 2156 35186 2212 35196
rect 3276 35476 3332 35486
rect 3276 34916 3332 35420
rect 3276 34850 3332 34860
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 3724 34244 3780 34254
rect 3724 33572 3780 34188
rect 3724 33506 3780 33516
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 2044 25620 2100 25630
rect 1820 20916 1876 20926
rect 1708 19572 1764 19582
rect 1708 17444 1764 19516
rect 1820 18340 1876 20860
rect 1820 18274 1876 18284
rect 2044 17556 2100 25564
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 2044 17490 2100 17500
rect 2380 22820 2436 22830
rect 1708 17378 1764 17388
rect 2380 17220 2436 22764
rect 4448 22764 4768 24276
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 25676 41860 25732 41870
rect 25676 37716 25732 41804
rect 25676 37650 25732 37660
rect 19808 36092 20128 37604
rect 26572 36820 26628 44044
rect 32508 40292 32564 54460
rect 32508 40226 32564 40236
rect 35168 54124 35488 55636
rect 35168 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35488 54124
rect 35168 52556 35488 54068
rect 35168 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35488 52556
rect 35168 50988 35488 52500
rect 35168 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35488 50988
rect 35168 49420 35488 50932
rect 35168 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35488 49420
rect 35168 47852 35488 49364
rect 35168 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35488 47852
rect 35168 46284 35488 47796
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 26572 36754 26628 36764
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 50528 56476 50848 56508
rect 50528 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50848 56476
rect 50528 54908 50848 56420
rect 50528 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50848 54908
rect 50528 53340 50848 54852
rect 50528 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50848 53340
rect 50528 51772 50848 53284
rect 50528 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50848 51772
rect 50528 50204 50848 51716
rect 50528 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50848 50204
rect 50528 48636 50848 50148
rect 50528 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50848 48636
rect 50528 47068 50848 48580
rect 50528 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50848 47068
rect 50528 45500 50848 47012
rect 50528 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50848 45500
rect 50528 43932 50848 45444
rect 50528 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50848 43932
rect 50528 42364 50848 43876
rect 50528 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50848 42364
rect 50528 40796 50848 42308
rect 50528 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50848 40796
rect 48860 39844 48916 39854
rect 48860 39284 48916 39788
rect 48860 39218 48916 39228
rect 50528 39228 50848 40740
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 32620 34132 32676 34142
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 31948 33124 32004 33134
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 26460 29316 26516 29326
rect 19808 25116 20128 26628
rect 23884 26628 23940 26638
rect 23884 25956 23940 26572
rect 26460 26516 26516 29260
rect 27692 28868 27748 28878
rect 27692 27076 27748 28812
rect 27692 27010 27748 27020
rect 26460 26450 26516 26460
rect 23884 25890 23940 25900
rect 31948 25956 32004 33068
rect 32172 27188 32228 27198
rect 32172 26404 32228 27132
rect 32172 26338 32228 26348
rect 31948 25890 32004 25900
rect 32620 25508 32676 34076
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 33292 31220 33348 31230
rect 32844 28420 32900 28430
rect 32844 27188 32900 28364
rect 32844 27122 32900 27132
rect 32620 25442 32676 25452
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 7420 23940 7476 23950
rect 7420 23604 7476 23884
rect 7420 23538 7476 23548
rect 19808 23548 20128 25060
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 3612 22036 3668 22046
rect 2380 17154 2436 17164
rect 2828 21924 2884 21934
rect 2828 20580 2884 21868
rect 3276 21700 3332 21710
rect 3276 21252 3332 21644
rect 3276 21186 3332 21196
rect 2828 13748 2884 20524
rect 3612 17556 3668 21980
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4060 20468 4116 20478
rect 3836 20132 3892 20142
rect 3836 18340 3892 20076
rect 4060 18676 4116 20412
rect 4060 18610 4116 18620
rect 4448 19628 4768 21140
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 23772 23044 23828 23054
rect 23772 22036 23828 22988
rect 23772 21970 23828 21980
rect 30156 22036 30212 22046
rect 6300 20916 6356 20926
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 3836 18274 3892 18284
rect 3612 17490 3668 17500
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 2828 13682 2884 13692
rect 4448 16492 4768 18004
rect 4844 20580 4900 20590
rect 4844 17556 4900 20524
rect 4844 17490 4900 17500
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 6300 13076 6356 20860
rect 6300 13010 6356 13020
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 12572 20128 14084
rect 28028 16884 28084 16894
rect 28028 13524 28084 16828
rect 30156 16772 30212 21980
rect 33292 18676 33348 31164
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 34972 29764 35028 29774
rect 33740 29316 33796 29326
rect 33740 25060 33796 29260
rect 34860 29204 34916 29214
rect 34636 27524 34692 27534
rect 33740 24994 33796 25004
rect 34524 25956 34580 25966
rect 34524 23716 34580 25900
rect 34636 24612 34692 27468
rect 34860 25060 34916 29148
rect 34972 25396 35028 29708
rect 34972 25330 35028 25340
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 34860 24994 34916 25004
rect 34972 25172 35028 25182
rect 34636 24546 34692 24556
rect 34972 23940 35028 25116
rect 34972 23874 35028 23884
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 34524 23650 34580 23660
rect 34972 23716 35028 23726
rect 34748 23268 34804 23278
rect 34748 22372 34804 23212
rect 34748 22306 34804 22316
rect 34860 22932 34916 22942
rect 33292 18610 33348 18620
rect 30156 16706 30212 16716
rect 28028 13458 28084 13468
rect 28588 16324 28644 16334
rect 28588 13076 28644 16268
rect 34860 15092 34916 22876
rect 34972 17444 35028 23660
rect 34972 17378 35028 17388
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 34860 15026 34916 15036
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 28588 13010 28644 13020
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
rect 50528 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50848 39228
rect 50528 37660 50848 39172
rect 50528 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50848 37660
rect 50528 36092 50848 37604
rect 50528 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50848 36092
rect 50528 34524 50848 36036
rect 50528 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50848 34524
rect 50528 32956 50848 34468
rect 50528 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50848 32956
rect 50528 31388 50848 32900
rect 50528 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50848 31388
rect 50528 29820 50848 31332
rect 50528 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50848 29820
rect 50528 28252 50848 29764
rect 50528 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50848 28252
rect 50528 26684 50848 28196
rect 50528 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50848 26684
rect 50528 25116 50848 26628
rect 50528 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50848 25116
rect 50528 23548 50848 25060
rect 50528 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50848 23548
rect 50528 21980 50848 23492
rect 50528 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50848 21980
rect 50528 20412 50848 21924
rect 50528 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50848 20412
rect 50528 18844 50848 20356
rect 50528 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50848 18844
rect 50528 17276 50848 18788
rect 50528 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50848 17276
rect 50528 15708 50848 17220
rect 50528 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50848 15708
rect 50528 14140 50848 15652
rect 50528 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50848 14140
rect 50528 12572 50848 14084
rect 50528 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50848 12572
rect 50528 11004 50848 12516
rect 50528 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50848 11004
rect 50528 9436 50848 10948
rect 50528 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50848 9436
rect 50528 7868 50848 9380
rect 50528 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50848 7868
rect 50528 6300 50848 7812
rect 50528 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50848 6300
rect 50528 4732 50848 6244
rect 50528 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50848 4732
rect 50528 3164 50848 4676
rect 50528 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50848 3164
rect 50528 3076 50848 3108
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1767_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 19712 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1768_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18256 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1769_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19152 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1770_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18816 0 -1 28224
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1771_
timestamp 1698431365
transform 1 0 21168 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1772_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 22064 0 -1 28224
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1773_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21168 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1774_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 37520 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1775_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 39088 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1776_
timestamp 1698431365
transform 1 0 4480 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1777_
timestamp 1698431365
transform 1 0 14784 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1778_
timestamp 1698431365
transform 1 0 21168 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1779_
timestamp 1698431365
transform 1 0 17248 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1780_
timestamp 1698431365
transform 1 0 19824 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1781_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13664 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1782_
timestamp 1698431365
transform 1 0 10192 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1783_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11312 0 1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1784_
timestamp 1698431365
transform 1 0 5712 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1785_
timestamp 1698431365
transform 1 0 5712 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1786_
timestamp 1698431365
transform 1 0 2240 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1787_
timestamp 1698431365
transform 1 0 7616 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1788_
timestamp 1698431365
transform -1 0 2912 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1789_
timestamp 1698431365
transform 1 0 1568 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1790_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 7840 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1791_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 7616 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1792_
timestamp 1698431365
transform 1 0 5712 0 -1 32928
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1793_
timestamp 1698431365
transform 1 0 9408 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or3_2  _1794_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 8288 0 1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1795_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9968 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1796_
timestamp 1698431365
transform 1 0 7056 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1797_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 8960 0 -1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1798_
timestamp 1698431365
transform 1 0 1568 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1799_
timestamp 1698431365
transform -1 0 7056 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1800_
timestamp 1698431365
transform 1 0 2128 0 -1 31360
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1801_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 5152 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1802_
timestamp 1698431365
transform 1 0 5488 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1803_
timestamp 1698431365
transform -1 0 7616 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1804_
timestamp 1698431365
transform 1 0 4480 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1805_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3360 0 -1 31360
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1806_
timestamp 1698431365
transform 1 0 6608 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1807_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5712 0 1 29792
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1808_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10640 0 1 29792
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1809_
timestamp 1698431365
transform -1 0 15120 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1810_
timestamp 1698431365
transform 1 0 9520 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1811_
timestamp 1698431365
transform 1 0 10416 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _1812_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5264 0 -1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _1813_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 7168 0 -1 29792
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1814_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 8064 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1815_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7504 0 -1 31360
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1816_
timestamp 1698431365
transform 1 0 8960 0 1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1817_
timestamp 1698431365
transform 1 0 6608 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1818_
timestamp 1698431365
transform -1 0 7840 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1819_
timestamp 1698431365
transform 1 0 1568 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1820_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2240 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1821_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3136 0 1 32928
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1822_
timestamp 1698431365
transform -1 0 5712 0 -1 34496
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1823_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2240 0 -1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1824_
timestamp 1698431365
transform 1 0 4480 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1825_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3248 0 -1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1826_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6608 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _1827_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9744 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1828_
timestamp 1698431365
transform 1 0 14000 0 1 32928
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1829_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 16912 0 1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1830_
timestamp 1698431365
transform 1 0 12768 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1831_
timestamp 1698431365
transform 1 0 10416 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1832_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 12208 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1833_
timestamp 1698431365
transform -1 0 9184 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1834_
timestamp 1698431365
transform 1 0 8064 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1835_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9408 0 -1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1836_
timestamp 1698431365
transform 1 0 10864 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai33_4  _1837_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 16912 0 -1 32928
box -86 -86 5798 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1838_
timestamp 1698431365
transform -1 0 7952 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1839_
timestamp 1698431365
transform -1 0 9184 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1840_
timestamp 1698431365
transform 1 0 7952 0 1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1841_
timestamp 1698431365
transform -1 0 5488 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1842_
timestamp 1698431365
transform -1 0 5040 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1843_
timestamp 1698431365
transform -1 0 2800 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1844_
timestamp 1698431365
transform 1 0 1568 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1845_
timestamp 1698431365
transform 1 0 1904 0 -1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1846_
timestamp 1698431365
transform -1 0 4480 0 1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1847_
timestamp 1698431365
transform -1 0 3472 0 1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1848_
timestamp 1698431365
transform 1 0 3696 0 1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _1849_
timestamp 1698431365
transform 1 0 5936 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1850_
timestamp 1698431365
transform 1 0 13328 0 1 34496
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1851_
timestamp 1698431365
transform 1 0 16688 0 1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1852_
timestamp 1698431365
transform 1 0 18816 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1853_
timestamp 1698431365
transform 1 0 17920 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1854_
timestamp 1698431365
transform -1 0 15904 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1855_
timestamp 1698431365
transform 1 0 13104 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1856_
timestamp 1698431365
transform 1 0 13328 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1857_
timestamp 1698431365
transform 1 0 15344 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1858_
timestamp 1698431365
transform 1 0 9408 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1859_
timestamp 1698431365
transform 1 0 13776 0 -1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1860_
timestamp 1698431365
transform 1 0 8064 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1861_
timestamp 1698431365
transform 1 0 9408 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1862_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7616 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1863_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 8848 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1864_
timestamp 1698431365
transform 1 0 7616 0 1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1865_
timestamp 1698431365
transform 1 0 8960 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1866_
timestamp 1698431365
transform -1 0 11536 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1867_
timestamp 1698431365
transform -1 0 11200 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1868_
timestamp 1698431365
transform 1 0 3696 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1869_
timestamp 1698431365
transform -1 0 7168 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1870_
timestamp 1698431365
transform 1 0 4368 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1871_
timestamp 1698431365
transform -1 0 5936 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1872_
timestamp 1698431365
transform 1 0 4480 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1873_
timestamp 1698431365
transform -1 0 6608 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1874_
timestamp 1698431365
transform 1 0 2240 0 1 43904
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1875_
timestamp 1698431365
transform 1 0 1680 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1876_
timestamp 1698431365
transform 1 0 6160 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1877_
timestamp 1698431365
transform -1 0 3584 0 -1 45472
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1878_
timestamp 1698431365
transform 1 0 5488 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1879_
timestamp 1698431365
transform 1 0 4032 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1880_
timestamp 1698431365
transform -1 0 3920 0 1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1881_
timestamp 1698431365
transform 1 0 1904 0 -1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1882_
timestamp 1698431365
transform 1 0 2800 0 -1 42336
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _1883_
timestamp 1698431365
transform 1 0 5488 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1884_
timestamp 1698431365
transform 1 0 10528 0 1 37632
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1885_
timestamp 1698431365
transform 1 0 17248 0 -1 37632
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1886_
timestamp 1698431365
transform 1 0 19488 0 1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1887_
timestamp 1698431365
transform 1 0 21056 0 -1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1888_
timestamp 1698431365
transform 1 0 19600 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1889_
timestamp 1698431365
transform 1 0 20272 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1890_
timestamp 1698431365
transform 1 0 15904 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1891_
timestamp 1698431365
transform -1 0 15344 0 -1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1892_
timestamp 1698431365
transform -1 0 3024 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1893_
timestamp 1698431365
transform 1 0 6384 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1894_
timestamp 1698431365
transform -1 0 7168 0 1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1895_
timestamp 1698431365
transform 1 0 5712 0 1 39200
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1896_
timestamp 1698431365
transform 1 0 11200 0 -1 37632
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1897_
timestamp 1698431365
transform 1 0 14896 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1898_
timestamp 1698431365
transform -1 0 19264 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai33_1  _1899_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 19376 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1900_
timestamp 1698431365
transform -1 0 16576 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1901_
timestamp 1698431365
transform 1 0 8400 0 1 39200
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1902_
timestamp 1698431365
transform 1 0 10080 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1903_
timestamp 1698431365
transform 1 0 10864 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1904_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 11312 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1905_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 12432 0 -1 39200
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1906_
timestamp 1698431365
transform 1 0 13664 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1907_
timestamp 1698431365
transform 1 0 14896 0 -1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1908_
timestamp 1698431365
transform 1 0 9968 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1909_
timestamp 1698431365
transform -1 0 14448 0 1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1910_
timestamp 1698431365
transform -1 0 9184 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1911_
timestamp 1698431365
transform 1 0 6944 0 1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1912_
timestamp 1698431365
transform 1 0 9184 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1913_
timestamp 1698431365
transform 1 0 12096 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1914_
timestamp 1698431365
transform -1 0 7728 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1915_
timestamp 1698431365
transform 1 0 5712 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1916_
timestamp 1698431365
transform 1 0 5488 0 1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1917_
timestamp 1698431365
transform -1 0 7392 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1918_
timestamp 1698431365
transform 1 0 3360 0 -1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1919_
timestamp 1698431365
transform 1 0 4816 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1920_
timestamp 1698431365
transform -1 0 3472 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1921_
timestamp 1698431365
transform -1 0 2912 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1922_
timestamp 1698431365
transform 1 0 1904 0 -1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1923_
timestamp 1698431365
transform 1 0 2352 0 1 45472
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1924_
timestamp 1698431365
transform 1 0 3808 0 1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _1925_
timestamp 1698431365
transform 1 0 5600 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _1926_
timestamp 1698431365
transform 1 0 11536 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1927_
timestamp 1698431365
transform 1 0 15120 0 1 39200
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1928_
timestamp 1698431365
transform 1 0 18816 0 -1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1929_
timestamp 1698431365
transform 1 0 21840 0 1 37632
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1930_
timestamp 1698431365
transform 1 0 21168 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1931_
timestamp 1698431365
transform 1 0 24080 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1932_
timestamp 1698431365
transform 1 0 24416 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1933_
timestamp 1698431365
transform 1 0 24752 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1934_
timestamp 1698431365
transform 1 0 25536 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1935_
timestamp 1698431365
transform 1 0 25872 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1936_
timestamp 1698431365
transform 1 0 26656 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1937_
timestamp 1698431365
transform 1 0 21168 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1938_
timestamp 1698431365
transform 1 0 22064 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1939_
timestamp 1698431365
transform -1 0 23744 0 -1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1940_
timestamp 1698431365
transform 1 0 17696 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1941_
timestamp 1698431365
transform 1 0 21168 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1942_
timestamp 1698431365
transform 1 0 17584 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  _1943_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 18592 0 1 37632
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1944_
timestamp 1698431365
transform 1 0 15120 0 -1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1945_
timestamp 1698431365
transform 1 0 18368 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1946_
timestamp 1698431365
transform 1 0 18816 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1947_
timestamp 1698431365
transform -1 0 16912 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1948_
timestamp 1698431365
transform 1 0 9184 0 1 42336
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1949_
timestamp 1698431365
transform -1 0 10864 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1950_
timestamp 1698431365
transform 1 0 4480 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1951_
timestamp 1698431365
transform 1 0 3920 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1952_
timestamp 1698431365
transform -1 0 5712 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1953_
timestamp 1698431365
transform 1 0 5936 0 -1 42336
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1954_
timestamp 1698431365
transform -1 0 10864 0 -1 42336
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1955_
timestamp 1698431365
transform 1 0 10640 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1956_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 12768 0 1 42336
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1957_
timestamp 1698431365
transform -1 0 15120 0 1 42336
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1958_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 17136 0 1 40768
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1959_
timestamp 1698431365
transform 1 0 9408 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1960_
timestamp 1698431365
transform -1 0 16128 0 -1 45472
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1961_
timestamp 1698431365
transform 1 0 6384 0 -1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1962_
timestamp 1698431365
transform 1 0 9072 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1963_
timestamp 1698431365
transform -1 0 10192 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1964_
timestamp 1698431365
transform -1 0 6160 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1965_
timestamp 1698431365
transform 1 0 6160 0 1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1966_
timestamp 1698431365
transform -1 0 5264 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1967_
timestamp 1698431365
transform -1 0 5152 0 -1 45472
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1968_
timestamp 1698431365
transform -1 0 5936 0 -1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1969_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 -1 45472
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1970_
timestamp 1698431365
transform 1 0 6160 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1971_
timestamp 1698431365
transform -1 0 6048 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1972_
timestamp 1698431365
transform 1 0 2688 0 1 47040
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1973_
timestamp 1698431365
transform -1 0 4144 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1974_
timestamp 1698431365
transform -1 0 4144 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1975_
timestamp 1698431365
transform 1 0 2912 0 -1 48608
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1976_
timestamp 1698431365
transform 1 0 4256 0 -1 48608
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_2  _1977_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6720 0 1 45472
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _1978_
timestamp 1698431365
transform 1 0 11872 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1979_
timestamp 1698431365
transform 1 0 17248 0 -1 42336
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1980_
timestamp 1698431365
transform -1 0 20384 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1981_
timestamp 1698431365
transform 1 0 21168 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1982_
timestamp 1698431365
transform 1 0 17584 0 1 40768
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1983_
timestamp 1698431365
transform 1 0 18368 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1984_
timestamp 1698431365
transform 1 0 11088 0 -1 42336
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _1985_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13664 0 -1 42336
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1986_
timestamp 1698431365
transform 1 0 15456 0 1 42336
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1987_
timestamp 1698431365
transform 1 0 19824 0 -1 40768
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1988_
timestamp 1698431365
transform 1 0 21392 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1989_
timestamp 1698431365
transform 1 0 22064 0 -1 40768
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1990_
timestamp 1698431365
transform -1 0 28000 0 1 39200
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1991_
timestamp 1698431365
transform -1 0 29680 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1992_
timestamp 1698431365
transform 1 0 27216 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1993_
timestamp 1698431365
transform 1 0 30576 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1994_
timestamp 1698431365
transform 1 0 30688 0 1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1995_
timestamp 1698431365
transform 1 0 21168 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1996_
timestamp 1698431365
transform 1 0 27888 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1997_
timestamp 1698431365
transform 1 0 28560 0 -1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1998_
timestamp 1698431365
transform 1 0 28112 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1999_
timestamp 1698431365
transform 1 0 29008 0 1 31360
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2000_
timestamp 1698431365
transform -1 0 30128 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2001_
timestamp 1698431365
transform -1 0 21952 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2002_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 -1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2003_
timestamp 1698431365
transform 1 0 22064 0 -1 28224
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2004_
timestamp 1698431365
transform -1 0 22736 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2005_
timestamp 1698431365
transform -1 0 21056 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2006_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15456 0 1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2007_
timestamp 1698431365
transform 1 0 14224 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2008_
timestamp 1698431365
transform 1 0 24976 0 1 40768
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2009_
timestamp 1698431365
transform -1 0 26208 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2010_
timestamp 1698431365
transform 1 0 25760 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2011_
timestamp 1698431365
transform 1 0 23856 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2012_
timestamp 1698431365
transform -1 0 22736 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2013_
timestamp 1698431365
transform -1 0 23520 0 -1 42336
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2014_
timestamp 1698431365
transform -1 0 23968 0 1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2015_
timestamp 1698431365
transform -1 0 22400 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2016_
timestamp 1698431365
transform 1 0 17472 0 -1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2017_
timestamp 1698431365
transform 1 0 19040 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2018_
timestamp 1698431365
transform 1 0 20384 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2019_
timestamp 1698431365
transform -1 0 16912 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2020_
timestamp 1698431365
transform 1 0 8176 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2021_
timestamp 1698431365
transform -1 0 11312 0 -1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2022_
timestamp 1698431365
transform 1 0 10416 0 1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2023_
timestamp 1698431365
transform 1 0 5936 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2024_
timestamp 1698431365
transform 1 0 10416 0 1 43904
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _2025_
timestamp 1698431365
transform -1 0 13104 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2026_
timestamp 1698431365
transform 1 0 11760 0 -1 43904
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  _2027_
timestamp 1698431365
transform 1 0 13440 0 1 43904
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2028_
timestamp 1698431365
transform -1 0 15456 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2029_
timestamp 1698431365
transform 1 0 8288 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2030_
timestamp 1698431365
transform -1 0 14336 0 -1 50176
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2031_
timestamp 1698431365
transform 1 0 7168 0 1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2032_
timestamp 1698431365
transform 1 0 9296 0 1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2033_
timestamp 1698431365
transform -1 0 11760 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2034_
timestamp 1698431365
transform 1 0 6608 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2035_
timestamp 1698431365
transform 1 0 3920 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2036_
timestamp 1698431365
transform 1 0 4704 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2037_
timestamp 1698431365
transform 1 0 6048 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2038_
timestamp 1698431365
transform 1 0 6384 0 1 50176
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2039_
timestamp 1698431365
transform 1 0 5488 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2040_
timestamp 1698431365
transform -1 0 8960 0 -1 48608
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2041_
timestamp 1698431365
transform 1 0 6608 0 -1 50176
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2042_
timestamp 1698431365
transform 1 0 11088 0 -1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2043_
timestamp 1698431365
transform 1 0 17248 0 -1 45472
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2044_
timestamp 1698431365
transform 1 0 20832 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2045_
timestamp 1698431365
transform 1 0 23520 0 1 42336
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2046_
timestamp 1698431365
transform -1 0 26880 0 -1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2047_
timestamp 1698431365
transform 1 0 11536 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2048_
timestamp 1698431365
transform 1 0 11200 0 -1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2049_
timestamp 1698431365
transform 1 0 17360 0 1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2050_
timestamp 1698431365
transform 1 0 16800 0 1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2051_
timestamp 1698431365
transform 1 0 16128 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2052_
timestamp 1698431365
transform 1 0 26096 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2053_
timestamp 1698431365
transform 1 0 23520 0 -1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2054_
timestamp 1698431365
transform 1 0 25088 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2055_
timestamp 1698431365
transform -1 0 27104 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2056_
timestamp 1698431365
transform 1 0 27104 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2057_
timestamp 1698431365
transform -1 0 20832 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2058_
timestamp 1698431365
transform -1 0 19600 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2059_
timestamp 1698431365
transform -1 0 19824 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2060_
timestamp 1698431365
transform 1 0 13552 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2061_
timestamp 1698431365
transform 1 0 14448 0 -1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2062_
timestamp 1698431365
transform 1 0 15456 0 1 45472
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2063_
timestamp 1698431365
transform 1 0 19264 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2064_
timestamp 1698431365
transform 1 0 21168 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2065_
timestamp 1698431365
transform 1 0 22960 0 1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2066_
timestamp 1698431365
transform 1 0 21280 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2067_
timestamp 1698431365
transform 1 0 18592 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2068_
timestamp 1698431365
transform 1 0 21952 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2069_
timestamp 1698431365
transform 1 0 18368 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2070_
timestamp 1698431365
transform 1 0 17472 0 1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2071_
timestamp 1698431365
transform 1 0 19376 0 1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2072_
timestamp 1698431365
transform -1 0 16576 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2073_
timestamp 1698431365
transform -1 0 11088 0 -1 48608
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2074_
timestamp 1698431365
transform -1 0 11872 0 -1 45472
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_2  _2075_
timestamp 1698431365
transform 1 0 7504 0 1 48608
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2076_
timestamp 1698431365
transform 1 0 10416 0 1 47040
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2077_
timestamp 1698431365
transform -1 0 12992 0 -1 47040
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2078_
timestamp 1698431365
transform 1 0 13104 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2079_
timestamp 1698431365
transform 1 0 13440 0 1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2080_
timestamp 1698431365
transform -1 0 14896 0 1 51744
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2081_
timestamp 1698431365
transform 1 0 6944 0 1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2082_
timestamp 1698431365
transform 1 0 8064 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2083_
timestamp 1698431365
transform 1 0 11648 0 1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2084_
timestamp 1698431365
transform 1 0 5488 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2085_
timestamp 1698431365
transform 1 0 9968 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2086_
timestamp 1698431365
transform 1 0 6944 0 -1 51744
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2087_
timestamp 1698431365
transform 1 0 9968 0 -1 53312
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2088_
timestamp 1698431365
transform 1 0 12768 0 -1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2089_
timestamp 1698431365
transform 1 0 14896 0 1 47040
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2090_
timestamp 1698431365
transform -1 0 22064 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2091_
timestamp 1698431365
transform 1 0 21504 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2092_
timestamp 1698431365
transform 1 0 19264 0 -1 48608
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2093_
timestamp 1698431365
transform 1 0 19824 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2094_
timestamp 1698431365
transform 1 0 10528 0 -1 50176
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _2095_
timestamp 1698431365
transform 1 0 13328 0 1 48608
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2096_
timestamp 1698431365
transform 1 0 14448 0 -1 48608
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2097_
timestamp 1698431365
transform 1 0 20160 0 -1 47040
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2098_
timestamp 1698431365
transform 1 0 22960 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2099_
timestamp 1698431365
transform 1 0 22848 0 1 45472
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2100_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 30016 0 -1 42336
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2101_
timestamp 1698431365
transform -1 0 30912 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2102_
timestamp 1698431365
transform 1 0 30576 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2103_
timestamp 1698431365
transform 1 0 29904 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2104_
timestamp 1698431365
transform -1 0 29904 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2105_
timestamp 1698431365
transform -1 0 10528 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2106_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 21616 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2107_
timestamp 1698431365
transform -1 0 22512 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2108_
timestamp 1698431365
transform 1 0 18816 0 1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2109_
timestamp 1698431365
transform 1 0 18032 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2110_
timestamp 1698431365
transform 1 0 13552 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2111_
timestamp 1698431365
transform 1 0 26992 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2112_
timestamp 1698431365
transform 1 0 28448 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2113_
timestamp 1698431365
transform 1 0 27552 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2114_
timestamp 1698431365
transform 1 0 26096 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2115_
timestamp 1698431365
transform 1 0 22064 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2116_
timestamp 1698431365
transform 1 0 22736 0 1 47040
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2117_
timestamp 1698431365
transform 1 0 22960 0 -1 47040
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2118_
timestamp 1698431365
transform 1 0 18256 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2119_
timestamp 1698431365
transform -1 0 22176 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2120_
timestamp 1698431365
transform 1 0 20384 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2121_
timestamp 1698431365
transform 1 0 15904 0 1 48608
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2122_
timestamp 1698431365
transform 1 0 20160 0 1 48608
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2123_
timestamp 1698431365
transform -1 0 21504 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2124_
timestamp 1698431365
transform 1 0 15232 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2125_
timestamp 1698431365
transform -1 0 18704 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2126_
timestamp 1698431365
transform 1 0 9968 0 1 51744
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2127_
timestamp 1698431365
transform 1 0 13328 0 1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2128_
timestamp 1698431365
transform -1 0 12768 0 -1 51744
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2129_
timestamp 1698431365
transform 1 0 11760 0 -1 53312
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  _2130_
timestamp 1698431365
transform 1 0 13328 0 1 50176
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2131_
timestamp 1698431365
transform 1 0 15344 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2132_
timestamp 1698431365
transform 1 0 10640 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2133_
timestamp 1698431365
transform -1 0 12656 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _2134_
timestamp 1698431365
transform 1 0 14896 0 1 51744
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2135_
timestamp 1698431365
transform 1 0 16912 0 1 51744
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2136_
timestamp 1698431365
transform 1 0 21168 0 -1 50176
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2137_
timestamp 1698431365
transform 1 0 23632 0 1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2138_
timestamp 1698431365
transform -1 0 28784 0 1 43904
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _2139_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 16016 0 1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2140_
timestamp 1698431365
transform 1 0 15344 0 -1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2141_
timestamp 1698431365
transform 1 0 14112 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2142_
timestamp 1698431365
transform 1 0 24304 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2143_
timestamp 1698431365
transform 1 0 26096 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2144_
timestamp 1698431365
transform -1 0 30576 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2145_
timestamp 1698431365
transform -1 0 28672 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2146_
timestamp 1698431365
transform 1 0 26656 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2147_
timestamp 1698431365
transform 1 0 27328 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2148_
timestamp 1698431365
transform 1 0 26880 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2149_
timestamp 1698431365
transform 1 0 22176 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2150_
timestamp 1698431365
transform 1 0 25536 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2151_
timestamp 1698431365
transform 1 0 21392 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2152_
timestamp 1698431365
transform 1 0 19040 0 1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2153_
timestamp 1698431365
transform -1 0 20160 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2154_
timestamp 1698431365
transform 1 0 17248 0 -1 51744
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2155_
timestamp 1698431365
transform 1 0 18704 0 -1 50176
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2156_
timestamp 1698431365
transform -1 0 22176 0 1 48608
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _2157_
timestamp 1698431365
transform 1 0 22176 0 1 48608
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2158_
timestamp 1698431365
transform 1 0 23408 0 1 48608
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2159_
timestamp 1698431365
transform -1 0 22848 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2160_
timestamp 1698431365
transform -1 0 20832 0 1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2161_
timestamp 1698431365
transform 1 0 19936 0 -1 51744
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2162_
timestamp 1698431365
transform 1 0 21392 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2163_
timestamp 1698431365
transform 1 0 19936 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2164_
timestamp 1698431365
transform 1 0 16016 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2165_
timestamp 1698431365
transform 1 0 17248 0 -1 53312
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2166_
timestamp 1698431365
transform 1 0 20272 0 -1 53312
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2167_
timestamp 1698431365
transform 1 0 21728 0 -1 53312
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2168_
timestamp 1698431365
transform 1 0 23632 0 1 50176
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2169_
timestamp 1698431365
transform -1 0 28112 0 1 47040
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2170_
timestamp 1698431365
transform -1 0 18144 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2171_
timestamp 1698431365
transform 1 0 23296 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2172_
timestamp 1698431365
transform 1 0 23856 0 1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2173_
timestamp 1698431365
transform 1 0 22736 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2174_
timestamp 1698431365
transform 1 0 26880 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2175_
timestamp 1698431365
transform -1 0 28672 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2176_
timestamp 1698431365
transform 1 0 25872 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2177_
timestamp 1698431365
transform 1 0 18704 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2178_
timestamp 1698431365
transform 1 0 25424 0 -1 47040
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2179_
timestamp 1698431365
transform 1 0 26096 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2180_
timestamp 1698431365
transform 1 0 26208 0 -1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2181_
timestamp 1698431365
transform 1 0 25536 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2182_
timestamp 1698431365
transform 1 0 18928 0 -1 53312
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2183_
timestamp 1698431365
transform 1 0 21168 0 1 51744
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2184_
timestamp 1698431365
transform -1 0 22848 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _2185_
timestamp 1698431365
transform 1 0 22736 0 1 51744
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2186_
timestamp 1698431365
transform 1 0 20720 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2187_
timestamp 1698431365
transform 1 0 24304 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2188_
timestamp 1698431365
transform -1 0 22064 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2189_
timestamp 1698431365
transform -1 0 22736 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2190_
timestamp 1698431365
transform 1 0 24640 0 1 53312
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2191_
timestamp 1698431365
transform 1 0 25536 0 1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2192_
timestamp 1698431365
transform 1 0 26208 0 -1 50176
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _2193_
timestamp 1698431365
transform 1 0 19600 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2194_
timestamp 1698431365
transform -1 0 21616 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2195_
timestamp 1698431365
transform 1 0 19264 0 1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2196_
timestamp 1698431365
transform -1 0 21392 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2197_
timestamp 1698431365
transform -1 0 26208 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2198_
timestamp 1698431365
transform -1 0 28784 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2199_
timestamp 1698431365
transform -1 0 28224 0 1 48608
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2200_
timestamp 1698431365
transform 1 0 24304 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2201_
timestamp 1698431365
transform -1 0 24640 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2202_
timestamp 1698431365
transform 1 0 25536 0 -1 53312
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2203_
timestamp 1698431365
transform -1 0 28448 0 -1 51744
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2204_
timestamp 1698431365
transform -1 0 24640 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2205_
timestamp 1698431365
transform -1 0 23408 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2206_
timestamp 1698431365
transform -1 0 28448 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2207_
timestamp 1698431365
transform 1 0 29680 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2208_
timestamp 1698431365
transform 1 0 29008 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2209_
timestamp 1698431365
transform -1 0 25872 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2210_
timestamp 1698431365
transform 1 0 26880 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2211_
timestamp 1698431365
transform 1 0 26320 0 1 50176
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2212_
timestamp 1698431365
transform 1 0 24640 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2213_
timestamp 1698431365
transform 1 0 25312 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2214_
timestamp 1698431365
transform -1 0 26544 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2215_
timestamp 1698431365
transform -1 0 28112 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2216_
timestamp 1698431365
transform 1 0 26544 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2217_
timestamp 1698431365
transform 1 0 23184 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2218_
timestamp 1698431365
transform 1 0 24976 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2219_
timestamp 1698431365
transform 1 0 30352 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2220_
timestamp 1698431365
transform -1 0 37520 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2221_
timestamp 1698431365
transform -1 0 30240 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2222_
timestamp 1698431365
transform 1 0 33936 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2223_
timestamp 1698431365
transform 1 0 34832 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2224_
timestamp 1698431365
transform -1 0 40208 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2225_
timestamp 1698431365
transform -1 0 40432 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2226_
timestamp 1698431365
transform -1 0 40208 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2227_
timestamp 1698431365
transform 1 0 38640 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2228_
timestamp 1698431365
transform -1 0 36176 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2229_
timestamp 1698431365
transform -1 0 37296 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2230_
timestamp 1698431365
transform 1 0 29568 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _2231_
timestamp 1698431365
transform -1 0 32368 0 1 4704
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _2232_
timestamp 1698431365
transform 1 0 31472 0 -1 4704
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2233_
timestamp 1698431365
transform -1 0 32368 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2234_
timestamp 1698431365
transform 1 0 31136 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2235_
timestamp 1698431365
transform -1 0 31248 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2236_
timestamp 1698431365
transform 1 0 42560 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2237_
timestamp 1698431365
transform 1 0 30240 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2238_
timestamp 1698431365
transform -1 0 39424 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2239_
timestamp 1698431365
transform -1 0 36624 0 1 4704
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2240_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 31584 0 -1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2241_
timestamp 1698431365
transform -1 0 32144 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2242_
timestamp 1698431365
transform 1 0 30352 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2243_
timestamp 1698431365
transform -1 0 37744 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2244_
timestamp 1698431365
transform 1 0 34048 0 1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2245_
timestamp 1698431365
transform 1 0 32704 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2246_
timestamp 1698431365
transform -1 0 31584 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2247_
timestamp 1698431365
transform -1 0 35840 0 -1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2248_
timestamp 1698431365
transform 1 0 32928 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_2  _2249_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 36512 0 -1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2250_
timestamp 1698431365
transform 1 0 30240 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _2251_
timestamp 1698431365
transform 1 0 36512 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2252_
timestamp 1698431365
transform -1 0 33600 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_2  _2253_
timestamp 1698431365
transform 1 0 30688 0 1 7840
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2254_
timestamp 1698431365
transform -1 0 33712 0 1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2255_
timestamp 1698431365
transform 1 0 32368 0 1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2256_
timestamp 1698431365
transform -1 0 36624 0 -1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2257_
timestamp 1698431365
transform 1 0 31808 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2258_
timestamp 1698431365
transform 1 0 34384 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _2259_
timestamp 1698431365
transform -1 0 35952 0 1 7840
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _2260_
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2261_
timestamp 1698431365
transform 1 0 33600 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  _2262_
timestamp 1698431365
transform 1 0 33152 0 -1 10976
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2263_
timestamp 1698431365
transform -1 0 41216 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2264_
timestamp 1698431365
transform -1 0 38640 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _2265_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 32928 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _2266_
timestamp 1698431365
transform 1 0 32592 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _2267_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 34496 0 -1 6272
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2268_
timestamp 1698431365
transform 1 0 35952 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2269_
timestamp 1698431365
transform -1 0 44464 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2270_
timestamp 1698431365
transform -1 0 40544 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2271_
timestamp 1698431365
transform 1 0 33936 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2272_
timestamp 1698431365
transform -1 0 39872 0 -1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_2  _2273_
timestamp 1698431365
transform 1 0 36848 0 1 7840
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2274_
timestamp 1698431365
transform -1 0 35952 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2275_
timestamp 1698431365
transform 1 0 33264 0 -1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2276_
timestamp 1698431365
transform 1 0 35504 0 1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2277_
timestamp 1698431365
transform 1 0 36064 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2278_
timestamp 1698431365
transform 1 0 34384 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2279_
timestamp 1698431365
transform 1 0 35280 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2280_
timestamp 1698431365
transform 1 0 33152 0 1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2281_
timestamp 1698431365
transform 1 0 32256 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai33_4  _2282_
timestamp 1698431365
transform 1 0 33712 0 -1 14112
box -86 -86 5798 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2283_
timestamp 1698431365
transform 1 0 36064 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2284_
timestamp 1698431365
transform -1 0 38640 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2285_
timestamp 1698431365
transform 1 0 36736 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2286_
timestamp 1698431365
transform 1 0 36848 0 1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2287_
timestamp 1698431365
transform 1 0 37408 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2288_
timestamp 1698431365
transform -1 0 39424 0 -1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2289_
timestamp 1698431365
transform -1 0 40992 0 1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2290_
timestamp 1698431365
transform -1 0 45920 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _2291_
timestamp 1698431365
transform -1 0 43680 0 -1 4704
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2292_
timestamp 1698431365
transform 1 0 44688 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2293_
timestamp 1698431365
transform -1 0 46592 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2294_
timestamp 1698431365
transform 1 0 42896 0 1 4704
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2295_
timestamp 1698431365
transform -1 0 42448 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2296_
timestamp 1698431365
transform 1 0 39648 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2297_
timestamp 1698431365
transform 1 0 40768 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2298_
timestamp 1698431365
transform -1 0 42672 0 1 4704
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2299_
timestamp 1698431365
transform 1 0 36848 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2300_
timestamp 1698431365
transform -1 0 39424 0 1 14112
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2301_
timestamp 1698431365
transform 1 0 36848 0 1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2302_
timestamp 1698431365
transform -1 0 37632 0 -1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2303_
timestamp 1698431365
transform 1 0 35504 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2304_
timestamp 1698431365
transform 1 0 39536 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2305_
timestamp 1698431365
transform 1 0 34384 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2306_
timestamp 1698431365
transform 1 0 36176 0 -1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2307_
timestamp 1698431365
transform 1 0 37184 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2308_
timestamp 1698431365
transform 1 0 37520 0 -1 15680
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2309_
timestamp 1698431365
transform 1 0 38640 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2310_
timestamp 1698431365
transform 1 0 39088 0 -1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2311_
timestamp 1698431365
transform -1 0 43232 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2312_
timestamp 1698431365
transform -1 0 32704 0 1 9408
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2313_
timestamp 1698431365
transform 1 0 35840 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2314_
timestamp 1698431365
transform 1 0 35056 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2315_
timestamp 1698431365
transform 1 0 38528 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2316_
timestamp 1698431365
transform -1 0 40208 0 -1 10976
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2317_
timestamp 1698431365
transform 1 0 38640 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2318_
timestamp 1698431365
transform -1 0 41440 0 1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2319_
timestamp 1698431365
transform 1 0 37968 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2320_
timestamp 1698431365
transform 1 0 39424 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2321_
timestamp 1698431365
transform 1 0 42224 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2322_
timestamp 1698431365
transform 1 0 37408 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2323_
timestamp 1698431365
transform -1 0 42224 0 -1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2324_
timestamp 1698431365
transform -1 0 41888 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2325_
timestamp 1698431365
transform 1 0 38976 0 -1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2326_
timestamp 1698431365
transform 1 0 37968 0 1 6272
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  _2327_
timestamp 1698431365
transform -1 0 45584 0 -1 7840
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2328_
timestamp 1698431365
transform -1 0 43344 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2329_
timestamp 1698431365
transform 1 0 43680 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2330_
timestamp 1698431365
transform 1 0 45808 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2331_
timestamp 1698431365
transform -1 0 48272 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2332_
timestamp 1698431365
transform -1 0 46816 0 1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2333_
timestamp 1698431365
transform 1 0 44688 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_2  _2334_
timestamp 1698431365
transform -1 0 44464 0 1 6272
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2335_
timestamp 1698431365
transform -1 0 43344 0 -1 10976
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2336_
timestamp 1698431365
transform -1 0 42896 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2337_
timestamp 1698431365
transform -1 0 41552 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2338_
timestamp 1698431365
transform -1 0 39536 0 1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2339_
timestamp 1698431365
transform 1 0 38976 0 -1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2340_
timestamp 1698431365
transform 1 0 38416 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2341_
timestamp 1698431365
transform 1 0 40768 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2342_
timestamp 1698431365
transform -1 0 39088 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2343_
timestamp 1698431365
transform 1 0 37632 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2344_
timestamp 1698431365
transform 1 0 37296 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai33_4  _2345_
timestamp 1698431365
transform 1 0 38416 0 1 17248
box -86 -86 5798 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2346_
timestamp 1698431365
transform -1 0 42112 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2347_
timestamp 1698431365
transform -1 0 40544 0 -1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2348_
timestamp 1698431365
transform 1 0 38080 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2349_
timestamp 1698431365
transform 1 0 39536 0 1 12544
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2350_
timestamp 1698431365
transform 1 0 39648 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2351_
timestamp 1698431365
transform 1 0 40768 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2352_
timestamp 1698431365
transform 1 0 39760 0 1 9408
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2353_
timestamp 1698431365
transform -1 0 42336 0 -1 12544
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  _2354_
timestamp 1698431365
transform -1 0 45584 0 -1 15680
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2355_
timestamp 1698431365
transform 1 0 43232 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2356_
timestamp 1698431365
transform 1 0 43232 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2357_
timestamp 1698431365
transform 1 0 47712 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2358_
timestamp 1698431365
transform 1 0 42784 0 1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2359_
timestamp 1698431365
transform -1 0 44464 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2360_
timestamp 1698431365
transform 1 0 42896 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2361_
timestamp 1698431365
transform -1 0 45584 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2362_
timestamp 1698431365
transform 1 0 43680 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2363_
timestamp 1698431365
transform -1 0 45472 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2364_
timestamp 1698431365
transform -1 0 46256 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2365_
timestamp 1698431365
transform -1 0 43792 0 -1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2366_
timestamp 1698431365
transform 1 0 43344 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2367_
timestamp 1698431365
transform -1 0 45136 0 -1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2368_
timestamp 1698431365
transform 1 0 45584 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2369_
timestamp 1698431365
transform -1 0 47376 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2370_
timestamp 1698431365
transform 1 0 46816 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2371_
timestamp 1698431365
transform 1 0 47824 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2372_
timestamp 1698431365
transform 1 0 49840 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2373_
timestamp 1698431365
transform -1 0 52416 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2374_
timestamp 1698431365
transform -1 0 49168 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _2375_
timestamp 1698431365
transform -1 0 51184 0 -1 6272
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2376_
timestamp 1698431365
transform -1 0 49168 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2377_
timestamp 1698431365
transform -1 0 47264 0 1 10976
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2378_
timestamp 1698431365
transform 1 0 42784 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_2  _2379_
timestamp 1698431365
transform 1 0 40992 0 -1 17248
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2380_
timestamp 1698431365
transform 1 0 38976 0 1 20384
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2381_
timestamp 1698431365
transform -1 0 40768 0 1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2382_
timestamp 1698431365
transform 1 0 39984 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2383_
timestamp 1698431365
transform 1 0 40768 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2384_
timestamp 1698431365
transform -1 0 41776 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2385_
timestamp 1698431365
transform 1 0 40096 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2386_
timestamp 1698431365
transform -1 0 42112 0 -1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2387_
timestamp 1698431365
transform -1 0 41440 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2388_
timestamp 1698431365
transform -1 0 42224 0 -1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2389_
timestamp 1698431365
transform 1 0 41888 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2390_
timestamp 1698431365
transform 1 0 42672 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2391_
timestamp 1698431365
transform -1 0 49952 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2392_
timestamp 1698431365
transform -1 0 43904 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2393_
timestamp 1698431365
transform 1 0 43344 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2394_
timestamp 1698431365
transform 1 0 42448 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2395_
timestamp 1698431365
transform 1 0 43792 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2396_
timestamp 1698431365
transform -1 0 44464 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2397_
timestamp 1698431365
transform -1 0 45360 0 -1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2398_
timestamp 1698431365
transform 1 0 40768 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2399_
timestamp 1698431365
transform 1 0 44688 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2400_
timestamp 1698431365
transform 1 0 41664 0 -1 9408
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2401_
timestamp 1698431365
transform -1 0 43680 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2402_
timestamp 1698431365
transform 1 0 43904 0 -1 10976
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2403_
timestamp 1698431365
transform 1 0 44688 0 1 12544
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2404_
timestamp 1698431365
transform -1 0 44464 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2405_
timestamp 1698431365
transform -1 0 46256 0 1 14112
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2406_
timestamp 1698431365
transform 1 0 45584 0 -1 15680
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2407_
timestamp 1698431365
transform 1 0 44688 0 1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2408_
timestamp 1698431365
transform 1 0 46368 0 -1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2409_
timestamp 1698431365
transform 1 0 47264 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2410_
timestamp 1698431365
transform -1 0 49728 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2411_
timestamp 1698431365
transform 1 0 46816 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2412_
timestamp 1698431365
transform 1 0 47376 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2413_
timestamp 1698431365
transform -1 0 47712 0 1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2414_
timestamp 1698431365
transform 1 0 46704 0 -1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2415_
timestamp 1698431365
transform 1 0 48608 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2416_
timestamp 1698431365
transform 1 0 47488 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2417_
timestamp 1698431365
transform -1 0 52192 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2418_
timestamp 1698431365
transform 1 0 48944 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2419_
timestamp 1698431365
transform 1 0 51184 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2420_
timestamp 1698431365
transform -1 0 51632 0 1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2421_
timestamp 1698431365
transform 1 0 50288 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2422_
timestamp 1698431365
transform -1 0 50736 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_2  _2423_
timestamp 1698431365
transform 1 0 50736 0 -1 7840
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2424_
timestamp 1698431365
transform -1 0 51744 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2425_
timestamp 1698431365
transform 1 0 45808 0 -1 17248
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2426_
timestamp 1698431365
transform -1 0 47040 0 -1 18816
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2427_
timestamp 1698431365
transform -1 0 45584 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2428_
timestamp 1698431365
transform -1 0 45584 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2429_
timestamp 1698431365
transform 1 0 41664 0 1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2430_
timestamp 1698431365
transform 1 0 42224 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2431_
timestamp 1698431365
transform -1 0 50400 0 -1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2432_
timestamp 1698431365
transform -1 0 50064 0 -1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2433_
timestamp 1698431365
transform -1 0 49616 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2434_
timestamp 1698431365
transform -1 0 47600 0 1 17248
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2435_
timestamp 1698431365
transform -1 0 43568 0 -1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2436_
timestamp 1698431365
transform -1 0 45584 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2437_
timestamp 1698431365
transform -1 0 44464 0 1 21952
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2438_
timestamp 1698431365
transform -1 0 42224 0 1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2439_
timestamp 1698431365
transform -1 0 41440 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2440_
timestamp 1698431365
transform -1 0 35616 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2441_
timestamp 1698431365
transform 1 0 32928 0 -1 25088
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2442_
timestamp 1698431365
transform 1 0 31136 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2443_
timestamp 1698431365
transform 1 0 32368 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2444_
timestamp 1698431365
transform -1 0 32704 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2445_
timestamp 1698431365
transform -1 0 33600 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2446_
timestamp 1698431365
transform 1 0 31696 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2447_
timestamp 1698431365
transform -1 0 31808 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2448_
timestamp 1698431365
transform 1 0 30912 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2449_
timestamp 1698431365
transform 1 0 31584 0 1 32928
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2450_
timestamp 1698431365
transform -1 0 25648 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2451_
timestamp 1698431365
transform -1 0 31808 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2452_
timestamp 1698431365
transform 1 0 35616 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2453_
timestamp 1698431365
transform 1 0 41440 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2454_
timestamp 1698431365
transform -1 0 41440 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2455_
timestamp 1698431365
transform -1 0 42896 0 -1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2456_
timestamp 1698431365
transform 1 0 43792 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2457_
timestamp 1698431365
transform -1 0 44464 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2458_
timestamp 1698431365
transform 1 0 43344 0 1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2459_
timestamp 1698431365
transform -1 0 44912 0 -1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2460_
timestamp 1698431365
transform 1 0 45808 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2461_
timestamp 1698431365
transform -1 0 48384 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2462_
timestamp 1698431365
transform -1 0 47040 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2463_
timestamp 1698431365
transform 1 0 45808 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2464_
timestamp 1698431365
transform 1 0 48272 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2465_
timestamp 1698431365
transform 1 0 48608 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2466_
timestamp 1698431365
transform -1 0 48384 0 -1 14112
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  _2467_
timestamp 1698431365
transform -1 0 51968 0 1 14112
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2468_
timestamp 1698431365
transform 1 0 34832 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2469_
timestamp 1698431365
transform 1 0 50288 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2470_
timestamp 1698431365
transform 1 0 50064 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2471_
timestamp 1698431365
transform 1 0 47936 0 1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2472_
timestamp 1698431365
transform 1 0 49728 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2473_
timestamp 1698431365
transform 1 0 51408 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2474_
timestamp 1698431365
transform -1 0 50288 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2475_
timestamp 1698431365
transform 1 0 52528 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2476_
timestamp 1698431365
transform -1 0 53760 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2477_
timestamp 1698431365
transform 1 0 53760 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2478_
timestamp 1698431365
transform -1 0 53648 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2479_
timestamp 1698431365
transform 1 0 49168 0 1 7840
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _2480_
timestamp 1698431365
transform 1 0 48608 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2481_
timestamp 1698431365
transform -1 0 53648 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2482_
timestamp 1698431365
transform 1 0 53648 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2483_
timestamp 1698431365
transform -1 0 51856 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2484_
timestamp 1698431365
transform -1 0 53312 0 -1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2485_
timestamp 1698431365
transform -1 0 54656 0 -1 12544
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2486_
timestamp 1698431365
transform 1 0 49952 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2487_
timestamp 1698431365
transform 1 0 48160 0 1 17248
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2488_
timestamp 1698431365
transform 1 0 45584 0 -1 21952
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2489_
timestamp 1698431365
transform -1 0 47040 0 1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2490_
timestamp 1698431365
transform -1 0 45136 0 -1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2491_
timestamp 1698431365
transform -1 0 44016 0 -1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2492_
timestamp 1698431365
transform 1 0 35168 0 1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2493_
timestamp 1698431365
transform -1 0 33712 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2494_
timestamp 1698431365
transform 1 0 29904 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _2495_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 32928 0 -1 31360
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2496_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25872 0 1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2497_
timestamp 1698431365
transform 1 0 25088 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2498_
timestamp 1698431365
transform -1 0 24192 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2499_
timestamp 1698431365
transform 1 0 44688 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2500_
timestamp 1698431365
transform -1 0 45696 0 -1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2501_
timestamp 1698431365
transform 1 0 45136 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2502_
timestamp 1698431365
transform -1 0 46256 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2503_
timestamp 1698431365
transform 1 0 46592 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2504_
timestamp 1698431365
transform 1 0 47040 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2505_
timestamp 1698431365
transform 1 0 43568 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2506_
timestamp 1698431365
transform 1 0 48608 0 -1 18816
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2507_
timestamp 1698431365
transform -1 0 49504 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2508_
timestamp 1698431365
transform -1 0 48160 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2509_
timestamp 1698431365
transform -1 0 48384 0 -1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2510_
timestamp 1698431365
transform 1 0 46256 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2511_
timestamp 1698431365
transform 1 0 49168 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2512_
timestamp 1698431365
transform -1 0 49840 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2513_
timestamp 1698431365
transform -1 0 53424 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2514_
timestamp 1698431365
transform 1 0 50064 0 1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2515_
timestamp 1698431365
transform 1 0 50736 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2516_
timestamp 1698431365
transform 1 0 50736 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2517_
timestamp 1698431365
transform -1 0 52304 0 1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2518_
timestamp 1698431365
transform 1 0 50624 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2519_
timestamp 1698431365
transform 1 0 52528 0 1 14112
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2520_
timestamp 1698431365
transform 1 0 50848 0 -1 15680
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2521_
timestamp 1698431365
transform 1 0 52528 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2522_
timestamp 1698431365
transform 1 0 53424 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2523_
timestamp 1698431365
transform 1 0 52528 0 1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2524_
timestamp 1698431365
transform 1 0 53200 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2525_
timestamp 1698431365
transform 1 0 53200 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2526_
timestamp 1698431365
transform 1 0 54544 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2527_
timestamp 1698431365
transform 1 0 54656 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2528_
timestamp 1698431365
transform 1 0 53872 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2529_
timestamp 1698431365
transform 1 0 53648 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2530_
timestamp 1698431365
transform 1 0 54320 0 1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2531_
timestamp 1698431365
transform 1 0 53536 0 -1 15680
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2532_
timestamp 1698431365
transform 1 0 51296 0 -1 17248
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2533_
timestamp 1698431365
transform 1 0 51744 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2534_
timestamp 1698431365
transform 1 0 52528 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2535_
timestamp 1698431365
transform -1 0 51408 0 -1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2536_
timestamp 1698431365
transform 1 0 48272 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2537_
timestamp 1698431365
transform -1 0 53984 0 -1 18816
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2538_
timestamp 1698431365
transform 1 0 49952 0 1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2539_
timestamp 1698431365
transform -1 0 50736 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2540_
timestamp 1698431365
transform -1 0 50848 0 1 23520
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2541_
timestamp 1698431365
transform -1 0 46704 0 1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2542_
timestamp 1698431365
transform -1 0 45696 0 -1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2543_
timestamp 1698431365
transform 1 0 33712 0 1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _2544_
timestamp 1698431365
transform 1 0 33040 0 1 29792
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2545_
timestamp 1698431365
transform 1 0 25088 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2546_
timestamp 1698431365
transform 1 0 23856 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2547_
timestamp 1698431365
transform 1 0 23408 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2548_
timestamp 1698431365
transform 1 0 26432 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2549_
timestamp 1698431365
transform -1 0 33488 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2550_
timestamp 1698431365
transform -1 0 28672 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2551_
timestamp 1698431365
transform 1 0 25088 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2552_
timestamp 1698431365
transform -1 0 35168 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2553_
timestamp 1698431365
transform -1 0 33600 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2554_
timestamp 1698431365
transform 1 0 33824 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2555_
timestamp 1698431365
transform 1 0 46704 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2556_
timestamp 1698431365
transform -1 0 46816 0 1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2557_
timestamp 1698431365
transform 1 0 48384 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2558_
timestamp 1698431365
transform -1 0 50624 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2559_
timestamp 1698431365
transform -1 0 50736 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2560_
timestamp 1698431365
transform -1 0 51632 0 1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2561_
timestamp 1698431365
transform -1 0 51408 0 -1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2562_
timestamp 1698431365
transform 1 0 49280 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2563_
timestamp 1698431365
transform 1 0 51744 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2564_
timestamp 1698431365
transform -1 0 55328 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2565_
timestamp 1698431365
transform -1 0 53760 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2566_
timestamp 1698431365
transform 1 0 51184 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2567_
timestamp 1698431365
transform 1 0 53760 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2568_
timestamp 1698431365
transform 1 0 54208 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2569_
timestamp 1698431365
transform 1 0 54096 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2570_
timestamp 1698431365
transform 1 0 54096 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2571_
timestamp 1698431365
transform 1 0 55216 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2572_
timestamp 1698431365
transform -1 0 57232 0 -1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2573_
timestamp 1698431365
transform -1 0 56224 0 1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2574_
timestamp 1698431365
transform 1 0 54768 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2575_
timestamp 1698431365
transform 1 0 55104 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2576_
timestamp 1698431365
transform -1 0 56672 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _2577_
timestamp 1698431365
transform 1 0 56224 0 1 15680
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2578_
timestamp 1698431365
transform -1 0 58240 0 1 18816
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2579_
timestamp 1698431365
transform 1 0 51856 0 -1 23520
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2580_
timestamp 1698431365
transform -1 0 53312 0 -1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2581_
timestamp 1698431365
transform -1 0 48384 0 -1 28224
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2582_
timestamp 1698431365
transform -1 0 35280 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2583_
timestamp 1698431365
transform -1 0 33488 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2584_
timestamp 1698431365
transform 1 0 30352 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2585_
timestamp 1698431365
transform 1 0 31920 0 1 34496
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2586_
timestamp 1698431365
transform -1 0 32704 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2587_
timestamp 1698431365
transform 1 0 47264 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2588_
timestamp 1698431365
transform -1 0 48160 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2589_
timestamp 1698431365
transform 1 0 47264 0 1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2590_
timestamp 1698431365
transform -1 0 50848 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2591_
timestamp 1698431365
transform 1 0 47264 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2592_
timestamp 1698431365
transform 1 0 54656 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2593_
timestamp 1698431365
transform 1 0 50848 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2594_
timestamp 1698431365
transform -1 0 58016 0 1 17248
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2595_
timestamp 1698431365
transform -1 0 55104 0 -1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2596_
timestamp 1698431365
transform -1 0 53648 0 -1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _2597_
timestamp 1698431365
transform -1 0 55664 0 -1 23520
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2598_
timestamp 1698431365
transform -1 0 54656 0 1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2599_
timestamp 1698431365
transform -1 0 52304 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2600_
timestamp 1698431365
transform -1 0 57792 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2601_
timestamp 1698431365
transform -1 0 57008 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2602_
timestamp 1698431365
transform 1 0 55664 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2603_
timestamp 1698431365
transform 1 0 55552 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2604_
timestamp 1698431365
transform 1 0 55328 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2605_
timestamp 1698431365
transform 1 0 56560 0 -1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2606_
timestamp 1698431365
transform -1 0 57904 0 -1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2607_
timestamp 1698431365
transform 1 0 52864 0 1 23520
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2608_
timestamp 1698431365
transform -1 0 57904 0 -1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2609_
timestamp 1698431365
transform -1 0 50064 0 -1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2610_
timestamp 1698431365
transform -1 0 49952 0 -1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2611_
timestamp 1698431365
transform -1 0 36176 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2612_
timestamp 1698431365
transform 1 0 33712 0 1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2613_
timestamp 1698431365
transform 1 0 30800 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2614_
timestamp 1698431365
transform 1 0 31472 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _2615_
timestamp 1698431365
transform 1 0 33824 0 -1 28224
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2616_
timestamp 1698431365
transform 1 0 32032 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2617_
timestamp 1698431365
transform -1 0 27552 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2618_
timestamp 1698431365
transform 1 0 25536 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2619_
timestamp 1698431365
transform 1 0 27328 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2620_
timestamp 1698431365
transform 1 0 27216 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2621_
timestamp 1698431365
transform -1 0 25872 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2622_
timestamp 1698431365
transform -1 0 26880 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2623_
timestamp 1698431365
transform -1 0 50288 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2624_
timestamp 1698431365
transform -1 0 50400 0 1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2625_
timestamp 1698431365
transform -1 0 53088 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2626_
timestamp 1698431365
transform 1 0 56112 0 1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2627_
timestamp 1698431365
transform -1 0 57904 0 -1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2628_
timestamp 1698431365
transform -1 0 57120 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _2629_
timestamp 1698431365
transform 1 0 55664 0 1 21952
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2630_
timestamp 1698431365
transform -1 0 55216 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2631_
timestamp 1698431365
transform 1 0 53424 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2632_
timestamp 1698431365
transform 1 0 54768 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2633_
timestamp 1698431365
transform -1 0 56112 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2634_
timestamp 1698431365
transform -1 0 55440 0 1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2635_
timestamp 1698431365
transform -1 0 55328 0 -1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2636_
timestamp 1698431365
transform -1 0 52304 0 1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2637_
timestamp 1698431365
transform -1 0 50960 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2638_
timestamp 1698431365
transform -1 0 38192 0 1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2639_
timestamp 1698431365
transform -1 0 31136 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _2640_
timestamp 1698431365
transform 1 0 33264 0 -1 29792
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2641_
timestamp 1698431365
transform 1 0 30688 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2642_
timestamp 1698431365
transform 1 0 29568 0 1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2643_
timestamp 1698431365
transform -1 0 29680 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2644_
timestamp 1698431365
transform -1 0 53424 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2645_
timestamp 1698431365
transform 1 0 55328 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2646_
timestamp 1698431365
transform 1 0 54208 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2647_
timestamp 1698431365
transform -1 0 53872 0 1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2648_
timestamp 1698431365
transform -1 0 52192 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2649_
timestamp 1698431365
transform -1 0 52416 0 -1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2650_
timestamp 1698431365
transform -1 0 52304 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2651_
timestamp 1698431365
transform 1 0 36064 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2652_
timestamp 1698431365
transform -1 0 38304 0 1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _2653_
timestamp 1698431365
transform 1 0 33824 0 1 26656
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2654_
timestamp 1698431365
transform -1 0 28000 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2655_
timestamp 1698431365
transform 1 0 28224 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2656_
timestamp 1698431365
transform 1 0 27440 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2657_
timestamp 1698431365
transform -1 0 52864 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2658_
timestamp 1698431365
transform 1 0 52416 0 -1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2659_
timestamp 1698431365
transform -1 0 40544 0 1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _2660_
timestamp 1698431365
transform 1 0 33936 0 1 25088
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2661_
timestamp 1698431365
transform 1 0 26208 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2662_
timestamp 1698431365
transform 1 0 26768 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2663_
timestamp 1698431365
transform 1 0 26320 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2664_
timestamp 1698431365
transform 1 0 3920 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2665_
timestamp 1698431365
transform 1 0 13440 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2666_
timestamp 1698431365
transform 1 0 22400 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2667_
timestamp 1698431365
transform 1 0 25088 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2668_
timestamp 1698431365
transform -1 0 22848 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2669_
timestamp 1698431365
transform 1 0 18256 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2670_
timestamp 1698431365
transform 1 0 19264 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2671_
timestamp 1698431365
transform 1 0 16016 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2672_
timestamp 1698431365
transform 1 0 18368 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2673_
timestamp 1698431365
transform 1 0 11200 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2674_
timestamp 1698431365
transform -1 0 14672 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2675_
timestamp 1698431365
transform 1 0 2240 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _2676_
timestamp 1698431365
transform 1 0 2688 0 1 23520
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2677_
timestamp 1698431365
transform 1 0 1792 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _2678_
timestamp 1698431365
transform 1 0 2688 0 -1 25088
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2679_
timestamp 1698431365
transform 1 0 1792 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2680_
timestamp 1698431365
transform 1 0 4368 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2681_
timestamp 1698431365
transform 1 0 2688 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2682_
timestamp 1698431365
transform 1 0 3584 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2683_
timestamp 1698431365
transform 1 0 2912 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2684_
timestamp 1698431365
transform 1 0 2128 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2685_
timestamp 1698431365
transform 1 0 4144 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2686_
timestamp 1698431365
transform 1 0 4368 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2687_
timestamp 1698431365
transform 1 0 4928 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2688_
timestamp 1698431365
transform 1 0 7392 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2689_
timestamp 1698431365
transform -1 0 8512 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2690_
timestamp 1698431365
transform 1 0 8400 0 1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2691_
timestamp 1698431365
transform -1 0 9632 0 1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2692_
timestamp 1698431365
transform 1 0 5488 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2693_
timestamp 1698431365
transform 1 0 6608 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_2  _2694_
timestamp 1698431365
transform 1 0 2128 0 -1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2695_
timestamp 1698431365
transform 1 0 1904 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _2696_
timestamp 1698431365
transform 1 0 2800 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2697_
timestamp 1698431365
transform 1 0 6272 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_2  _2698_
timestamp 1698431365
transform 1 0 6048 0 1 26656
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2699_
timestamp 1698431365
transform 1 0 10416 0 -1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2700_
timestamp 1698431365
transform 1 0 12768 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2701_
timestamp 1698431365
transform 1 0 11088 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2702_
timestamp 1698431365
transform -1 0 12320 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _2703_
timestamp 1698431365
transform 1 0 3024 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _2704_
timestamp 1698431365
transform 1 0 1680 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _2705_
timestamp 1698431365
transform 1 0 3584 0 -1 21952
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2706_
timestamp 1698431365
transform 1 0 4592 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2707_
timestamp 1698431365
transform -1 0 9184 0 -1 25088
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2708_
timestamp 1698431365
transform 1 0 9632 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai33_4  _2709_
timestamp 1698431365
transform -1 0 15120 0 -1 25088
box -86 -86 5798 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2710_
timestamp 1698431365
transform 1 0 8512 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2711_
timestamp 1698431365
transform -1 0 7056 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2712_
timestamp 1698431365
transform 1 0 3584 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2713_
timestamp 1698431365
transform 1 0 3584 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2714_
timestamp 1698431365
transform 1 0 2912 0 1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2715_
timestamp 1698431365
transform 1 0 5936 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2716_
timestamp 1698431365
transform 1 0 10528 0 1 23520
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2717_
timestamp 1698431365
transform 1 0 13440 0 1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2718_
timestamp 1698431365
transform 1 0 18368 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2719_
timestamp 1698431365
transform -1 0 16016 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2720_
timestamp 1698431365
transform 1 0 11312 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2721_
timestamp 1698431365
transform 1 0 12208 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _2722_
timestamp 1698431365
transform 1 0 12096 0 -1 23520
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2723_
timestamp 1698431365
transform 1 0 10192 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2724_
timestamp 1698431365
transform -1 0 11424 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2725_
timestamp 1698431365
transform 1 0 7840 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2726_
timestamp 1698431365
transform 1 0 5712 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2727_
timestamp 1698431365
transform -1 0 6608 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2728_
timestamp 1698431365
transform 1 0 7056 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2729_
timestamp 1698431365
transform 1 0 6832 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _2730_
timestamp 1698431365
transform 1 0 7952 0 -1 21952
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2731_
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2732_
timestamp 1698431365
transform 1 0 3696 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2733_
timestamp 1698431365
transform -1 0 8288 0 -1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _2734_
timestamp 1698431365
transform 1 0 3360 0 1 15680
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2735_
timestamp 1698431365
transform 1 0 4592 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2736_
timestamp 1698431365
transform 1 0 2688 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2737_
timestamp 1698431365
transform 1 0 4144 0 -1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2738_
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2739_
timestamp 1698431365
transform 1 0 4256 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2740_
timestamp 1698431365
transform 1 0 5152 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_2  _2741_
timestamp 1698431365
transform 1 0 6048 0 -1 18816
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2742_
timestamp 1698431365
transform 1 0 9856 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2743_
timestamp 1698431365
transform 1 0 14784 0 1 23520
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2744_
timestamp 1698431365
transform 1 0 18928 0 -1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  _2745_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19824 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2746_
timestamp 1698431365
transform 1 0 18816 0 -1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2747_
timestamp 1698431365
transform 1 0 16352 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2748_
timestamp 1698431365
transform 1 0 15120 0 -1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2749_
timestamp 1698431365
transform 1 0 16464 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2750_
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2751_
timestamp 1698431365
transform 1 0 11536 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2752_
timestamp 1698431365
transform 1 0 16240 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2753_
timestamp 1698431365
transform 1 0 11648 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2754_
timestamp 1698431365
transform 1 0 5824 0 -1 26656
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2755_
timestamp 1698431365
transform 1 0 6384 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _2756_
timestamp 1698431365
transform 1 0 5936 0 -1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2757_
timestamp 1698431365
transform 1 0 7504 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2758_
timestamp 1698431365
transform -1 0 10304 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2759_
timestamp 1698431365
transform 1 0 9184 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _2760_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 8176 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2761_
timestamp 1698431365
transform 1 0 9408 0 -1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2762_
timestamp 1698431365
transform 1 0 10864 0 -1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2763_
timestamp 1698431365
transform 1 0 13328 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2764_
timestamp 1698431365
transform -1 0 14224 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2765_
timestamp 1698431365
transform -1 0 13104 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2766_
timestamp 1698431365
transform -1 0 12768 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2767_
timestamp 1698431365
transform -1 0 5152 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2768_
timestamp 1698431365
transform 1 0 4816 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2769_
timestamp 1698431365
transform 1 0 5936 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2770_
timestamp 1698431365
transform 1 0 8848 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2771_
timestamp 1698431365
transform 1 0 9408 0 -1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2772_
timestamp 1698431365
transform -1 0 7728 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2773_
timestamp 1698431365
transform 1 0 5152 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2774_
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2775_
timestamp 1698431365
transform 1 0 4704 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2776_
timestamp 1698431365
transform 1 0 5264 0 -1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2777_
timestamp 1698431365
transform -1 0 7168 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2778_
timestamp 1698431365
transform 1 0 5712 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2779_
timestamp 1698431365
transform 1 0 10080 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2780_
timestamp 1698431365
transform 1 0 13776 0 -1 21952
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2781_
timestamp 1698431365
transform 1 0 17360 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2782_
timestamp 1698431365
transform 1 0 20048 0 -1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2783_
timestamp 1698431365
transform 1 0 21616 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2784_
timestamp 1698431365
transform 1 0 19936 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2785_
timestamp 1698431365
transform -1 0 22288 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2786_
timestamp 1698431365
transform 1 0 17696 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2787_
timestamp 1698431365
transform 1 0 15680 0 1 25088
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2788_
timestamp 1698431365
transform 1 0 6272 0 1 17248
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  _2789_
timestamp 1698431365
transform 1 0 7952 0 1 18816
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2790_
timestamp 1698431365
transform 1 0 10192 0 1 17248
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2791_
timestamp 1698431365
transform 1 0 13664 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2792_
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2793_
timestamp 1698431365
transform 1 0 17696 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  _2794_
timestamp 1698431365
transform 1 0 18368 0 -1 21952
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2795_
timestamp 1698431365
transform 1 0 17360 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2796_
timestamp 1698431365
transform 1 0 15568 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2797_
timestamp 1698431365
transform -1 0 14784 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2798_
timestamp 1698431365
transform 1 0 13328 0 1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2799_
timestamp 1698431365
transform 1 0 14672 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2800_
timestamp 1698431365
transform -1 0 15344 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2801_
timestamp 1698431365
transform -1 0 15792 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _2802_
timestamp 1698431365
transform -1 0 16240 0 1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2803_
timestamp 1698431365
transform 1 0 16128 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2804_
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2805_
timestamp 1698431365
transform 1 0 12320 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2806_
timestamp 1698431365
transform -1 0 17808 0 1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2807_
timestamp 1698431365
transform 1 0 10528 0 1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2808_
timestamp 1698431365
transform 1 0 13552 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2809_
timestamp 1698431365
transform 1 0 15792 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2810_
timestamp 1698431365
transform 1 0 8848 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2811_
timestamp 1698431365
transform -1 0 11984 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2812_
timestamp 1698431365
transform 1 0 8512 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2813_
timestamp 1698431365
transform 1 0 9520 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2814_
timestamp 1698431365
transform 1 0 5824 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2815_
timestamp 1698431365
transform 1 0 6608 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2816_
timestamp 1698431365
transform 1 0 6272 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _2817_
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2818_
timestamp 1698431365
transform 1 0 9856 0 -1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2819_
timestamp 1698431365
transform 1 0 8176 0 -1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2820_
timestamp 1698431365
transform 1 0 6608 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2821_
timestamp 1698431365
transform 1 0 6160 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2822_
timestamp 1698431365
transform 1 0 5936 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2823_
timestamp 1698431365
transform 1 0 5600 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2824_
timestamp 1698431365
transform -1 0 7280 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2825_
timestamp 1698431365
transform 1 0 5936 0 1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_2  _2826_
timestamp 1698431365
transform 1 0 8400 0 1 10976
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2827_
timestamp 1698431365
transform 1 0 10864 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2828_
timestamp 1698431365
transform 1 0 15232 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2829_
timestamp 1698431365
transform 1 0 17584 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2830_
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2831_
timestamp 1698431365
transform 1 0 23184 0 -1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2832_
timestamp 1698431365
transform -1 0 26768 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2833_
timestamp 1698431365
transform 1 0 26880 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2834_
timestamp 1698431365
transform -1 0 24752 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2835_
timestamp 1698431365
transform -1 0 22512 0 1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2836_
timestamp 1698431365
transform 1 0 24192 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2837_
timestamp 1698431365
transform 1 0 20608 0 -1 20384
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2838_
timestamp 1698431365
transform 1 0 19936 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2839_
timestamp 1698431365
transform 1 0 20272 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  _2840_
timestamp 1698431365
transform 1 0 16128 0 1 20384
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2841_
timestamp 1698431365
transform 1 0 18144 0 1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2842_
timestamp 1698431365
transform -1 0 20944 0 1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2843_
timestamp 1698431365
transform -1 0 19936 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2844_
timestamp 1698431365
transform 1 0 21168 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2845_
timestamp 1698431365
transform -1 0 20608 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2846_
timestamp 1698431365
transform -1 0 14000 0 -1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2847_
timestamp 1698431365
transform 1 0 12768 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2848_
timestamp 1698431365
transform 1 0 8176 0 -1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _2849_
timestamp 1698431365
transform 1 0 7840 0 1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2850_
timestamp 1698431365
transform 1 0 8848 0 1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2851_
timestamp 1698431365
transform 1 0 10528 0 1 14112
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2852_
timestamp 1698431365
transform 1 0 12992 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2853_
timestamp 1698431365
transform 1 0 15008 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2854_
timestamp 1698431365
transform -1 0 16352 0 -1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2855_
timestamp 1698431365
transform 1 0 18480 0 1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2856_
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2857_
timestamp 1698431365
transform 1 0 17472 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2858_
timestamp 1698431365
transform 1 0 12432 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2859_
timestamp 1698431365
transform -1 0 18592 0 1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2860_
timestamp 1698431365
transform 1 0 13552 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2861_
timestamp 1698431365
transform 1 0 11760 0 1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2862_
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2863_
timestamp 1698431365
transform 1 0 15120 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2864_
timestamp 1698431365
transform 1 0 10304 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2865_
timestamp 1698431365
transform -1 0 12992 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2866_
timestamp 1698431365
transform 1 0 6496 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2867_
timestamp 1698431365
transform 1 0 7280 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2868_
timestamp 1698431365
transform 1 0 7056 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2869_
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2870_
timestamp 1698431365
transform -1 0 11872 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2871_
timestamp 1698431365
transform 1 0 5712 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2872_
timestamp 1698431365
transform 1 0 9184 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2873_
timestamp 1698431365
transform -1 0 7280 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2874_
timestamp 1698431365
transform 1 0 7280 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2875_
timestamp 1698431365
transform 1 0 7504 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_2  _2876_
timestamp 1698431365
transform 1 0 7952 0 1 7840
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2877_
timestamp 1698431365
transform 1 0 11872 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2878_
timestamp 1698431365
transform 1 0 15680 0 1 12544
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2879_
timestamp 1698431365
transform 1 0 18928 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2880_
timestamp 1698431365
transform 1 0 21168 0 1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2881_
timestamp 1698431365
transform 1 0 21280 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2882_
timestamp 1698431365
transform 1 0 23520 0 1 20384
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2883_
timestamp 1698431365
transform -1 0 26880 0 -1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2884_
timestamp 1698431365
transform 1 0 23408 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2885_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25088 0 -1 26656
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2886_
timestamp 1698431365
transform -1 0 34272 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2887_
timestamp 1698431365
transform 1 0 23184 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2888_
timestamp 1698431365
transform -1 0 24416 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2889_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 23968 0 1 25088
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2890_
timestamp 1698431365
transform 1 0 26432 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2891_
timestamp 1698431365
transform 1 0 23968 0 1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2892_
timestamp 1698431365
transform -1 0 26320 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2893_
timestamp 1698431365
transform 1 0 27552 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2894_
timestamp 1698431365
transform 1 0 24304 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2895_
timestamp 1698431365
transform -1 0 17024 0 -1 15680
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _2896_
timestamp 1698431365
transform 1 0 16016 0 1 14112
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2897_
timestamp 1698431365
transform 1 0 18592 0 -1 15680
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2898_
timestamp 1698431365
transform 1 0 20832 0 -1 18816
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2899_
timestamp 1698431365
transform -1 0 22512 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  _2900_
timestamp 1698431365
transform 1 0 22512 0 1 17248
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2901_
timestamp 1698431365
transform -1 0 24192 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2902_
timestamp 1698431365
transform 1 0 23184 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2903_
timestamp 1698431365
transform -1 0 24416 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2904_
timestamp 1698431365
transform 1 0 21168 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2905_
timestamp 1698431365
transform -1 0 23184 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2906_
timestamp 1698431365
transform 1 0 18592 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2907_
timestamp 1698431365
transform -1 0 20272 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2908_
timestamp 1698431365
transform 1 0 14112 0 1 9408
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2909_
timestamp 1698431365
transform -1 0 14784 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2910_
timestamp 1698431365
transform 1 0 8064 0 1 9408
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  _2911_
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2912_
timestamp 1698431365
transform 1 0 12096 0 -1 9408
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2913_
timestamp 1698431365
transform -1 0 15680 0 1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _2914_
timestamp 1698431365
transform -1 0 17360 0 1 10976
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2915_
timestamp 1698431365
transform 1 0 17472 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2916_
timestamp 1698431365
transform -1 0 19488 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2917_
timestamp 1698431365
transform 1 0 17696 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2918_
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2919_
timestamp 1698431365
transform -1 0 16128 0 -1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2920_
timestamp 1698431365
transform -1 0 16800 0 -1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2921_
timestamp 1698431365
transform -1 0 17248 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2922_
timestamp 1698431365
transform 1 0 12544 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2923_
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2924_
timestamp 1698431365
transform 1 0 8512 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2925_
timestamp 1698431365
transform -1 0 12096 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2926_
timestamp 1698431365
transform 1 0 10640 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2927_
timestamp 1698431365
transform -1 0 12544 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2928_
timestamp 1698431365
transform 1 0 10528 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2929_
timestamp 1698431365
transform 1 0 11200 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2930_
timestamp 1698431365
transform -1 0 9184 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2931_
timestamp 1698431365
transform -1 0 10304 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2932_
timestamp 1698431365
transform 1 0 11088 0 1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2933_
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2934_
timestamp 1698431365
transform 1 0 16128 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2935_
timestamp 1698431365
transform 1 0 18368 0 -1 12544
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2936_
timestamp 1698431365
transform 1 0 21616 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2937_
timestamp 1698431365
transform 1 0 25088 0 -1 17248
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2938_
timestamp 1698431365
transform 1 0 27328 0 -1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2939_
timestamp 1698431365
transform 1 0 27440 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2940_
timestamp 1698431365
transform 1 0 28224 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2941_
timestamp 1698431365
transform 1 0 22960 0 1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2942_
timestamp 1698431365
transform 1 0 23856 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2943_
timestamp 1698431365
transform -1 0 29904 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2944_
timestamp 1698431365
transform -1 0 28784 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2945_
timestamp 1698431365
transform -1 0 28896 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2946_
timestamp 1698431365
transform 1 0 27552 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2947_
timestamp 1698431365
transform 1 0 27216 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2948_
timestamp 1698431365
transform -1 0 37744 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2949_
timestamp 1698431365
transform -1 0 36176 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2950_
timestamp 1698431365
transform 1 0 25088 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2951_
timestamp 1698431365
transform 1 0 26544 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2952_
timestamp 1698431365
transform 1 0 24976 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2953_
timestamp 1698431365
transform 1 0 23184 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2954_
timestamp 1698431365
transform -1 0 23968 0 1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2955_
timestamp 1698431365
transform 1 0 22288 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _2956_
timestamp 1698431365
transform 1 0 23408 0 -1 14112
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2957_
timestamp 1698431365
transform -1 0 27552 0 1 14112
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2958_
timestamp 1698431365
transform 1 0 21280 0 1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2959_
timestamp 1698431365
transform 1 0 22288 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2960_
timestamp 1698431365
transform -1 0 17024 0 -1 12544
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  _2961_
timestamp 1698431365
transform 1 0 17472 0 -1 10976
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2962_
timestamp 1698431365
transform 1 0 19600 0 1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2963_
timestamp 1698431365
transform -1 0 22848 0 1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2964_
timestamp 1698431365
transform 1 0 22512 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2965_
timestamp 1698431365
transform 1 0 19040 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2966_
timestamp 1698431365
transform -1 0 21728 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2967_
timestamp 1698431365
transform -1 0 16688 0 1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2968_
timestamp 1698431365
transform 1 0 15008 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2969_
timestamp 1698431365
transform -1 0 18816 0 -1 9408
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2970_
timestamp 1698431365
transform -1 0 20944 0 1 9408
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2971_
timestamp 1698431365
transform 1 0 20160 0 -1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2972_
timestamp 1698431365
transform 1 0 12656 0 -1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2973_
timestamp 1698431365
transform 1 0 13776 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2974_
timestamp 1698431365
transform 1 0 15680 0 -1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2975_
timestamp 1698431365
transform 1 0 15120 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2976_
timestamp 1698431365
transform -1 0 12544 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2977_
timestamp 1698431365
transform -1 0 12768 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2978_
timestamp 1698431365
transform 1 0 16016 0 1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2979_
timestamp 1698431365
transform 1 0 17696 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2980_
timestamp 1698431365
transform 1 0 19824 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2981_
timestamp 1698431365
transform 1 0 23632 0 1 10976
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2982_
timestamp 1698431365
transform 1 0 25536 0 -1 15680
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2983_
timestamp 1698431365
transform -1 0 30464 0 1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2984_
timestamp 1698431365
transform 1 0 31808 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2985_
timestamp 1698431365
transform 1 0 28224 0 -1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2986_
timestamp 1698431365
transform 1 0 29568 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2987_
timestamp 1698431365
transform 1 0 10528 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2988_
timestamp 1698431365
transform 1 0 13664 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2989_
timestamp 1698431365
transform 1 0 14896 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2990_
timestamp 1698431365
transform -1 0 36512 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2991_
timestamp 1698431365
transform 1 0 29680 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2992_
timestamp 1698431365
transform 1 0 33152 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2993_
timestamp 1698431365
transform -1 0 35056 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2994_
timestamp 1698431365
transform 1 0 36848 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2995_
timestamp 1698431365
transform 1 0 27216 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2996_
timestamp 1698431365
transform 1 0 25536 0 1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2997_
timestamp 1698431365
transform 1 0 26880 0 1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2998_
timestamp 1698431365
transform 1 0 26096 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2999_
timestamp 1698431365
transform 1 0 20944 0 -1 12544
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _3000_
timestamp 1698431365
transform 1 0 23632 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _3001_
timestamp 1698431365
transform 1 0 22288 0 1 12544
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  _3002_
timestamp 1698431365
transform 1 0 25088 0 -1 12544
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3003_
timestamp 1698431365
transform -1 0 25088 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _3004_
timestamp 1698431365
transform 1 0 19488 0 1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _3005_
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3006_
timestamp 1698431365
transform 1 0 23856 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _3007_
timestamp 1698431365
transform 1 0 19264 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3008_
timestamp 1698431365
transform -1 0 23744 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _3009_
timestamp 1698431365
transform 1 0 17808 0 -1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _3010_
timestamp 1698431365
transform 1 0 18368 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  _3011_
timestamp 1698431365
transform 1 0 18368 0 -1 6272
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3012_
timestamp 1698431365
transform 1 0 20048 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3013_
timestamp 1698431365
transform 1 0 16016 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3014_
timestamp 1698431365
transform -1 0 18368 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3015_
timestamp 1698431365
transform 1 0 21392 0 1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _3016_
timestamp 1698431365
transform 1 0 22064 0 -1 7840
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _3017_
timestamp 1698431365
transform 1 0 23856 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _3018_
timestamp 1698431365
transform 1 0 26208 0 1 12544
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _3019_
timestamp 1698431365
transform 1 0 29120 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _3020_
timestamp 1698431365
transform 1 0 29008 0 1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3021_
timestamp 1698431365
transform 1 0 29120 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3022_
timestamp 1698431365
transform 1 0 12208 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _3023_
timestamp 1698431365
transform 1 0 14336 0 -1 26656
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3024_
timestamp 1698431365
transform 1 0 29904 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3025_
timestamp 1698431365
transform -1 0 32032 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3026_
timestamp 1698431365
transform -1 0 30912 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3027_
timestamp 1698431365
transform 1 0 27664 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3028_
timestamp 1698431365
transform -1 0 31472 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3029_
timestamp 1698431365
transform -1 0 30352 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3030_
timestamp 1698431365
transform -1 0 37968 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3031_
timestamp 1698431365
transform 1 0 26656 0 -1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3032_
timestamp 1698431365
transform 1 0 28000 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3033_
timestamp 1698431365
transform 1 0 25648 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _3034_
timestamp 1698431365
transform -1 0 24864 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _3035_
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _3036_
timestamp 1698431365
transform 1 0 25760 0 1 9408
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _3037_
timestamp 1698431365
transform 1 0 26880 0 1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3038_
timestamp 1698431365
transform 1 0 27888 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3039_
timestamp 1698431365
transform 1 0 24304 0 1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _3040_
timestamp 1698431365
transform 1 0 27104 0 -1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3041_
timestamp 1698431365
transform 1 0 27216 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3042_
timestamp 1698431365
transform 1 0 25536 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3043_
timestamp 1698431365
transform 1 0 27664 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _3044_
timestamp 1698431365
transform 1 0 21728 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _3045_
timestamp 1698431365
transform 1 0 22848 0 1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3046_
timestamp 1698431365
transform -1 0 31360 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _3047_
timestamp 1698431365
transform 1 0 29008 0 1 9408
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _3048_
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _3049_
timestamp 1698431365
transform -1 0 31584 0 1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _3050_
timestamp 1698431365
transform -1 0 30128 0 1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3051_
timestamp 1698431365
transform 1 0 30576 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3052_
timestamp 1698431365
transform 1 0 18144 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _3053_
timestamp 1698431365
transform 1 0 19488 0 1 25088
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3054_
timestamp 1698431365
transform 1 0 30800 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3055_
timestamp 1698431365
transform 1 0 35056 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3056_
timestamp 1698431365
transform 1 0 35728 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _3057_
timestamp 1698431365
transform -1 0 30016 0 -1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _3058_
timestamp 1698431365
transform 1 0 27776 0 -1 9408
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3059_
timestamp 1698431365
transform 1 0 29904 0 -1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _3060_
timestamp 1698431365
transform -1 0 31584 0 -1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3061_
timestamp 1698431365
transform 1 0 27888 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _3062_
timestamp 1698431365
transform -1 0 28784 0 1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3063_
timestamp 1698431365
transform -1 0 28784 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _3064_
timestamp 1698431365
transform 1 0 28784 0 -1 10976
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3065_
timestamp 1698431365
transform 1 0 28224 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3066_
timestamp 1698431365
transform -1 0 27104 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _3067_
timestamp 1698431365
transform 1 0 29008 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3068_
timestamp 1698431365
transform 1 0 28560 0 -1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3069_
timestamp 1698431365
transform 1 0 29904 0 -1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _3070_
timestamp 1698431365
transform 1 0 30688 0 1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3071_
timestamp 1698431365
transform 1 0 29568 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3072_
timestamp 1698431365
transform -1 0 31920 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3073_
timestamp 1698431365
transform -1 0 30128 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _3074_
timestamp 1698431365
transform -1 0 29904 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3075_
timestamp 1698431365
transform -1 0 21952 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3076_
timestamp 1698431365
transform 1 0 20496 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _3077_
timestamp 1698431365
transform 1 0 30128 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3078_
timestamp 1698431365
transform -1 0 34944 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3079_
timestamp 1698431365
transform 1 0 33152 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3080_
timestamp 1698431365
transform -1 0 34832 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3081_
timestamp 1698431365
transform -1 0 32256 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3082_
timestamp 1698431365
transform 1 0 30800 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3083_
timestamp 1698431365
transform -1 0 30800 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3084_
timestamp 1698431365
transform -1 0 31696 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3085_
timestamp 1698431365
transform 1 0 28448 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _3086_
timestamp 1698431365
transform 1 0 29680 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3087_
timestamp 1698431365
transform 1 0 31248 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3088_
timestamp 1698431365
transform 1 0 30688 0 -1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _3089_
timestamp 1698431365
transform -1 0 32368 0 1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _3090_
timestamp 1698431365
transform 1 0 32368 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3091_
timestamp 1698431365
transform -1 0 23632 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3092_
timestamp 1698431365
transform 1 0 22512 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _3093_
timestamp 1698431365
transform 1 0 32928 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3094_
timestamp 1698431365
transform -1 0 34496 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3095_
timestamp 1698431365
transform 1 0 35952 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3096_
timestamp 1698431365
transform 1 0 33600 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _3097_
timestamp 1698431365
transform 1 0 31696 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _3098_
timestamp 1698431365
transform 1 0 26768 0 1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _3099_
timestamp 1698431365
transform 1 0 27328 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _3100_
timestamp 1698431365
transform 1 0 30128 0 1 20384
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3101_
timestamp 1698431365
transform -1 0 35392 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3102_
timestamp 1698431365
transform -1 0 36176 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3103_
timestamp 1698431365
transform 1 0 34720 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _3104_
timestamp 1698431365
transform 1 0 29904 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3105_
timestamp 1698431365
transform 1 0 32928 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _3106_
timestamp 1698431365
transform 1 0 37072 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _3107_
timestamp 1698431365
transform 1 0 40880 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3108_
timestamp 1698431365
transform 1 0 37296 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3109_
timestamp 1698431365
transform -1 0 39648 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3110_
timestamp 1698431365
transform -1 0 37408 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _3111_
timestamp 1698431365
transform -1 0 34048 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3112_
timestamp 1698431365
transform -1 0 34944 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3113_
timestamp 1698431365
transform 1 0 35056 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3114_
timestamp 1698431365
transform -1 0 32480 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _3115_
timestamp 1698431365
transform -1 0 30464 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _3116_
timestamp 1698431365
transform 1 0 29568 0 1 51744
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _3117_
timestamp 1698431365
transform 1 0 29008 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _3118_
timestamp 1698431365
transform -1 0 30912 0 -1 51744
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _3119_
timestamp 1698431365
transform 1 0 30912 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3120_
timestamp 1698431365
transform -1 0 36624 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _3121_
timestamp 1698431365
transform 1 0 30800 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _3122_
timestamp 1698431365
transform -1 0 33600 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _3123_
timestamp 1698431365
transform 1 0 34944 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _3124_
timestamp 1698431365
transform 1 0 30352 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _3125_
timestamp 1698431365
transform 1 0 34048 0 -1 51744
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _3126_
timestamp 1698431365
transform 1 0 30016 0 -1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3127_
timestamp 1698431365
transform 1 0 29680 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3128_
timestamp 1698431365
transform 1 0 30240 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _3129_
timestamp 1698431365
transform -1 0 30016 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _3130_
timestamp 1698431365
transform 1 0 31360 0 1 48608
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _3131_
timestamp 1698431365
transform -1 0 32256 0 1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3132_
timestamp 1698431365
transform 1 0 29568 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _3133_
timestamp 1698431365
transform 1 0 30352 0 1 48608
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_2  _3134_
timestamp 1698431365
transform 1 0 31248 0 -1 53312
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _3135_
timestamp 1698431365
transform 1 0 30464 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _3136_
timestamp 1698431365
transform 1 0 32928 0 -1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _3137_
timestamp 1698431365
transform -1 0 32704 0 -1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_2  _3138_
timestamp 1698431365
transform 1 0 28784 0 -1 47040
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3139_
timestamp 1698431365
transform -1 0 31920 0 -1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  _3140_
timestamp 1698431365
transform 1 0 31472 0 -1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3141_
timestamp 1698431365
transform 1 0 34160 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _3142_
timestamp 1698431365
transform -1 0 35168 0 -1 45472
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _3143_
timestamp 1698431365
transform -1 0 34944 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _3144_
timestamp 1698431365
transform 1 0 31360 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _3145_
timestamp 1698431365
transform 1 0 32032 0 1 51744
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3146_
timestamp 1698431365
transform 1 0 30688 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _3147_
timestamp 1698431365
transform -1 0 34048 0 1 45472
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _3148_
timestamp 1698431365
transform 1 0 31584 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai33_4  _3149_
timestamp 1698431365
transform 1 0 32928 0 -1 47040
box -86 -86 5798 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3150_
timestamp 1698431365
transform 1 0 32144 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3151_
timestamp 1698431365
transform -1 0 33040 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3152_
timestamp 1698431365
transform -1 0 36624 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3153_
timestamp 1698431365
transform 1 0 32144 0 -1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3154_
timestamp 1698431365
transform -1 0 36288 0 1 53312
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _3155_
timestamp 1698431365
transform 1 0 32928 0 -1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _3156_
timestamp 1698431365
transform -1 0 35280 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _3157_
timestamp 1698431365
transform 1 0 32928 0 1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _3158_
timestamp 1698431365
transform 1 0 33712 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3159_
timestamp 1698431365
transform -1 0 36288 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _3160_
timestamp 1698431365
transform -1 0 33936 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3161_
timestamp 1698431365
transform -1 0 35952 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  _3162_
timestamp 1698431365
transform -1 0 35728 0 1 42336
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3163_
timestamp 1698431365
transform 1 0 35616 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3164_
timestamp 1698431365
transform -1 0 36512 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3165_
timestamp 1698431365
transform -1 0 38528 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _3166_
timestamp 1698431365
transform 1 0 32032 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3167_
timestamp 1698431365
transform -1 0 35952 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3168_
timestamp 1698431365
transform -1 0 36624 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _3169_
timestamp 1698431365
transform 1 0 34160 0 1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _3170_
timestamp 1698431365
transform 1 0 35392 0 1 48608
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _3171_
timestamp 1698431365
transform 1 0 33824 0 1 47040
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3172_
timestamp 1698431365
transform 1 0 36624 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _3173_
timestamp 1698431365
transform -1 0 38080 0 1 50176
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _3174_
timestamp 1698431365
transform 1 0 36848 0 1 51744
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3175_
timestamp 1698431365
transform -1 0 39648 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3176_
timestamp 1698431365
transform -1 0 37968 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _3177_
timestamp 1698431365
transform 1 0 38080 0 1 51744
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _3178_
timestamp 1698431365
transform 1 0 38640 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _3179_
timestamp 1698431365
transform 1 0 35280 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _3180_
timestamp 1698431365
transform 1 0 39760 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_2  _3181_
timestamp 1698431365
transform 1 0 36624 0 -1 54880
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _3182_
timestamp 1698431365
transform 1 0 35392 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _3183_
timestamp 1698431365
transform 1 0 34048 0 -1 42336
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _3184_
timestamp 1698431365
transform 1 0 35168 0 1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _3185_
timestamp 1698431365
transform -1 0 37296 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3186_
timestamp 1698431365
transform -1 0 37968 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _3187_
timestamp 1698431365
transform 1 0 36848 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3188_
timestamp 1698431365
transform 1 0 35728 0 -1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3189_
timestamp 1698431365
transform -1 0 38080 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _3190_
timestamp 1698431365
transform -1 0 36624 0 1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3191_
timestamp 1698431365
transform 1 0 36960 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _3192_
timestamp 1698431365
transform 1 0 38192 0 1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3193_
timestamp 1698431365
transform -1 0 41664 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _3194_
timestamp 1698431365
transform 1 0 29008 0 1 45472
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _3195_
timestamp 1698431365
transform 1 0 32704 0 1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _3196_
timestamp 1698431365
transform 1 0 32928 0 -1 48608
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3197_
timestamp 1698431365
transform -1 0 33936 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3198_
timestamp 1698431365
transform -1 0 35168 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _3199_
timestamp 1698431365
transform 1 0 36848 0 1 48608
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _3200_
timestamp 1698431365
transform -1 0 37968 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _3201_
timestamp 1698431365
transform 1 0 36288 0 -1 48608
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3202_
timestamp 1698431365
transform 1 0 37856 0 1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _3203_
timestamp 1698431365
transform -1 0 40544 0 -1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _3204_
timestamp 1698431365
transform 1 0 35728 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3205_
timestamp 1698431365
transform -1 0 39312 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3206_
timestamp 1698431365
transform -1 0 39760 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3207_
timestamp 1698431365
transform -1 0 40320 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _3208_
timestamp 1698431365
transform -1 0 40432 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _3209_
timestamp 1698431365
transform 1 0 36624 0 -1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _3210_
timestamp 1698431365
transform -1 0 38976 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _3211_
timestamp 1698431365
transform 1 0 38080 0 -1 50176
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3212_
timestamp 1698431365
transform 1 0 36064 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _3213_
timestamp 1698431365
transform 1 0 37744 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3214_
timestamp 1698431365
transform 1 0 42448 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3215_
timestamp 1698431365
transform -1 0 43568 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3216_
timestamp 1698431365
transform -1 0 43232 0 -1 53312
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3217_
timestamp 1698431365
transform 1 0 42336 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _3218_
timestamp 1698431365
transform 1 0 39088 0 1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _3219_
timestamp 1698431365
transform 1 0 38640 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _3220_
timestamp 1698431365
transform 1 0 37632 0 1 43904
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _3221_
timestamp 1698431365
transform -1 0 40208 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _3222_
timestamp 1698431365
transform 1 0 37296 0 -1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _3223_
timestamp 1698431365
transform 1 0 38752 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3224_
timestamp 1698431365
transform 1 0 37744 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _3225_
timestamp 1698431365
transform 1 0 39648 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3226_
timestamp 1698431365
transform -1 0 35728 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _3227_
timestamp 1698431365
transform 1 0 36624 0 -1 42336
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _3228_
timestamp 1698431365
transform 1 0 36848 0 1 53312
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  _3229_
timestamp 1698431365
transform -1 0 42896 0 1 50176
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _3230_
timestamp 1698431365
transform 1 0 37968 0 -1 48608
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _3231_
timestamp 1698431365
transform 1 0 40208 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3232_
timestamp 1698431365
transform -1 0 40320 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3233_
timestamp 1698431365
transform 1 0 38416 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  _3234_
timestamp 1698431365
transform -1 0 40544 0 -1 40768
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _3235_
timestamp 1698431365
transform 1 0 40768 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3236_
timestamp 1698431365
transform 1 0 40768 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _3237_
timestamp 1698431365
transform 1 0 40768 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _3238_
timestamp 1698431365
transform 1 0 41440 0 -1 47040
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3239_
timestamp 1698431365
transform 1 0 36848 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3240_
timestamp 1698431365
transform 1 0 41440 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _3241_
timestamp 1698431365
transform 1 0 41552 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _3242_
timestamp 1698431365
transform -1 0 40544 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _3243_
timestamp 1698431365
transform 1 0 39424 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _3244_
timestamp 1698431365
transform -1 0 40544 0 -1 42336
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3245_
timestamp 1698431365
transform 1 0 43008 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _3246_
timestamp 1698431365
transform -1 0 44464 0 1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3247_
timestamp 1698431365
transform 1 0 41664 0 1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _3248_
timestamp 1698431365
transform -1 0 44016 0 1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3249_
timestamp 1698431365
transform 1 0 41328 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3250_
timestamp 1698431365
transform 1 0 42112 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3251_
timestamp 1698431365
transform 1 0 43680 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3252_
timestamp 1698431365
transform 1 0 41328 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3253_
timestamp 1698431365
transform 1 0 44464 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3254_
timestamp 1698431365
transform 1 0 40768 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3255_
timestamp 1698431365
transform -1 0 44800 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _3256_
timestamp 1698431365
transform 1 0 40768 0 -1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _3257_
timestamp 1698431365
transform -1 0 44128 0 1 50176
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _3258_
timestamp 1698431365
transform 1 0 41328 0 -1 48608
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _3259_
timestamp 1698431365
transform 1 0 44800 0 1 50176
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _3260_
timestamp 1698431365
transform 1 0 43232 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3261_
timestamp 1698431365
transform 1 0 44688 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3262_
timestamp 1698431365
transform 1 0 47936 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _3263_
timestamp 1698431365
transform 1 0 43008 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3264_
timestamp 1698431365
transform -1 0 49392 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3265_
timestamp 1698431365
transform -1 0 49840 0 1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _3266_
timestamp 1698431365
transform 1 0 44912 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _3267_
timestamp 1698431365
transform 1 0 43344 0 -1 47040
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _3268_
timestamp 1698431365
transform 1 0 42000 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _3269_
timestamp 1698431365
transform 1 0 40544 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _3270_
timestamp 1698431365
transform 1 0 39648 0 1 37632
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _3271_
timestamp 1698431365
transform -1 0 42224 0 1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3272_
timestamp 1698431365
transform -1 0 41664 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _3273_
timestamp 1698431365
transform -1 0 41328 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3274_
timestamp 1698431365
transform 1 0 39536 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3275_
timestamp 1698431365
transform 1 0 40768 0 -1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3276_
timestamp 1698431365
transform -1 0 40768 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _3277_
timestamp 1698431365
transform 1 0 40768 0 1 39200
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _3278_
timestamp 1698431365
transform -1 0 43792 0 1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3279_
timestamp 1698431365
transform 1 0 48608 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  _3280_
timestamp 1698431365
transform 1 0 39424 0 1 42336
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3281_
timestamp 1698431365
transform -1 0 46032 0 1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _3282_
timestamp 1698431365
transform -1 0 43456 0 -1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _3283_
timestamp 1698431365
transform 1 0 43456 0 1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3284_
timestamp 1698431365
transform -1 0 44352 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3285_
timestamp 1698431365
transform 1 0 45360 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _3286_
timestamp 1698431365
transform 1 0 42560 0 -1 47040
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3287_
timestamp 1698431365
transform 1 0 40544 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _3288_
timestamp 1698431365
transform -1 0 43344 0 -1 51744
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _3289_
timestamp 1698431365
transform -1 0 45136 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _3290_
timestamp 1698431365
transform -1 0 44464 0 -1 50176
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _3291_
timestamp 1698431365
transform 1 0 44016 0 -1 48608
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3292_
timestamp 1698431365
transform 1 0 44688 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _3293_
timestamp 1698431365
transform 1 0 45696 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _3294_
timestamp 1698431365
transform 1 0 44688 0 1 43904
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _3295_
timestamp 1698431365
transform -1 0 44464 0 -1 45472
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _3296_
timestamp 1698431365
transform -1 0 46592 0 -1 42336
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _3297_
timestamp 1698431365
transform 1 0 46592 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3298_
timestamp 1698431365
transform 1 0 45920 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _3299_
timestamp 1698431365
transform 1 0 46928 0 -1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3300_
timestamp 1698431365
transform 1 0 45696 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3301_
timestamp 1698431365
transform 1 0 46592 0 -1 48608
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _3302_
timestamp 1698431365
transform -1 0 47936 0 1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3303_
timestamp 1698431365
transform 1 0 46592 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3304_
timestamp 1698431365
transform 1 0 47264 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3305_
timestamp 1698431365
transform 1 0 47712 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3306_
timestamp 1698431365
transform 1 0 46256 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _3307_
timestamp 1698431365
transform -1 0 48048 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _3308_
timestamp 1698431365
transform 1 0 45136 0 -1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _3309_
timestamp 1698431365
transform 1 0 46368 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3310_
timestamp 1698431365
transform -1 0 47376 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3311_
timestamp 1698431365
transform 1 0 49952 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3312_
timestamp 1698431365
transform -1 0 51184 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3313_
timestamp 1698431365
transform -1 0 51408 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3314_
timestamp 1698431365
transform 1 0 48608 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3315_
timestamp 1698431365
transform 1 0 49280 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_2  _3316_
timestamp 1698431365
transform 1 0 48608 0 -1 50176
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _3317_
timestamp 1698431365
transform 1 0 47264 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _3318_
timestamp 1698431365
transform 1 0 46704 0 1 40768
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3319_
timestamp 1698431365
transform -1 0 47488 0 -1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3320_
timestamp 1698431365
transform -1 0 47488 0 -1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _3321_
timestamp 1698431365
transform -1 0 45360 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _3322_
timestamp 1698431365
transform 1 0 40768 0 -1 36064
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3323_
timestamp 1698431365
transform -1 0 40432 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _3324_
timestamp 1698431365
transform -1 0 38416 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _3325_
timestamp 1698431365
transform -1 0 34160 0 -1 34496
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3326_
timestamp 1698431365
transform -1 0 32704 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3327_
timestamp 1698431365
transform 1 0 31360 0 1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _3328_
timestamp 1698431365
transform -1 0 31360 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3329_
timestamp 1698431365
transform -1 0 37408 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3330_
timestamp 1698431365
transform 1 0 45136 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _3331_
timestamp 1698431365
transform 1 0 42224 0 1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3332_
timestamp 1698431365
transform 1 0 42560 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3333_
timestamp 1698431365
transform -1 0 42336 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3334_
timestamp 1698431365
transform 1 0 43680 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _3335_
timestamp 1698431365
transform 1 0 41328 0 -1 42336
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _3336_
timestamp 1698431365
transform -1 0 47264 0 1 42336
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _3337_
timestamp 1698431365
transform -1 0 47712 0 1 39200
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _3338_
timestamp 1698431365
transform 1 0 43456 0 -1 40768
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3339_
timestamp 1698431365
transform 1 0 43568 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  _3340_
timestamp 1698431365
transform -1 0 45920 0 -1 37632
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3341_
timestamp 1698431365
transform 1 0 45472 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3342_
timestamp 1698431365
transform 1 0 45136 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3343_
timestamp 1698431365
transform 1 0 46592 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _3344_
timestamp 1698431365
transform 1 0 46256 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3345_
timestamp 1698431365
transform -1 0 48160 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _3346_
timestamp 1698431365
transform 1 0 47488 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3347_
timestamp 1698431365
transform 1 0 48608 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _3348_
timestamp 1698431365
transform 1 0 47600 0 -1 45472
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3349_
timestamp 1698431365
transform -1 0 45360 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _3350_
timestamp 1698431365
transform 1 0 45136 0 1 51744
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  _3351_
timestamp 1698431365
transform -1 0 51184 0 1 50176
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _3352_
timestamp 1698431365
transform -1 0 51184 0 -1 47040
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _3353_
timestamp 1698431365
transform -1 0 50064 0 1 45472
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _3354_
timestamp 1698431365
transform -1 0 50176 0 1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _3355_
timestamp 1698431365
transform 1 0 48608 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3356_
timestamp 1698431365
transform 1 0 48832 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3357_
timestamp 1698431365
transform 1 0 50176 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3358_
timestamp 1698431365
transform 1 0 50512 0 1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _3359_
timestamp 1698431365
transform 1 0 50624 0 1 45472
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _3360_
timestamp 1698431365
transform -1 0 50400 0 -1 45472
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3361_
timestamp 1698431365
transform 1 0 50512 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3362_
timestamp 1698431365
transform 1 0 51184 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _3363_
timestamp 1698431365
transform 1 0 49392 0 -1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3364_
timestamp 1698431365
transform 1 0 51408 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3365_
timestamp 1698431365
transform 1 0 52528 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _3366_
timestamp 1698431365
transform 1 0 52640 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _3367_
timestamp 1698431365
transform 1 0 53088 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3368_
timestamp 1698431365
transform 1 0 53536 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3369_
timestamp 1698431365
transform -1 0 53312 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3370_
timestamp 1698431365
transform -1 0 52080 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3371_
timestamp 1698431365
transform 1 0 51744 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _3372_
timestamp 1698431365
transform -1 0 51744 0 1 48608
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _3373_
timestamp 1698431365
transform -1 0 55216 0 1 47040
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _3374_
timestamp 1698431365
transform 1 0 50512 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _3375_
timestamp 1698431365
transform 1 0 48608 0 -1 40768
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _3376_
timestamp 1698431365
transform 1 0 46368 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _3377_
timestamp 1698431365
transform -1 0 46144 0 -1 36064
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _3378_
timestamp 1698431365
transform 1 0 41552 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _3379_
timestamp 1698431365
transform -1 0 44128 0 1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3380_
timestamp 1698431365
transform -1 0 43120 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3381_
timestamp 1698431365
transform -1 0 42560 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _3382_
timestamp 1698431365
transform -1 0 38864 0 -1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _3383_
timestamp 1698431365
transform 1 0 33712 0 1 34496
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _3384_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 34832 0 1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3385_
timestamp 1698431365
transform 1 0 35728 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3386_
timestamp 1698431365
transform 1 0 36848 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3387_
timestamp 1698431365
transform -1 0 46032 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3388_
timestamp 1698431365
transform -1 0 44800 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3389_
timestamp 1698431365
transform 1 0 46032 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3390_
timestamp 1698431365
transform 1 0 49392 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _3391_
timestamp 1698431365
transform -1 0 49168 0 1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _3392_
timestamp 1698431365
transform 1 0 47712 0 1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _3393_
timestamp 1698431365
transform 1 0 47152 0 -1 37632
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _3394_
timestamp 1698431365
transform 1 0 46928 0 1 34496
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _3395_
timestamp 1698431365
transform 1 0 49168 0 -1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _3396_
timestamp 1698431365
transform -1 0 52640 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _3397_
timestamp 1698431365
transform 1 0 47264 0 1 43904
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  _3398_
timestamp 1698431365
transform -1 0 54096 0 -1 42336
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3399_
timestamp 1698431365
transform -1 0 52528 0 -1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _3400_
timestamp 1698431365
transform 1 0 50176 0 -1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _3401_
timestamp 1698431365
transform 1 0 49840 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3402_
timestamp 1698431365
transform 1 0 52528 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3403_
timestamp 1698431365
transform 1 0 51744 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _3404_
timestamp 1698431365
transform -1 0 52864 0 -1 45472
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _3405_
timestamp 1698431365
transform -1 0 52192 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _3406_
timestamp 1698431365
transform -1 0 52304 0 1 42336
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _3407_
timestamp 1698431365
transform 1 0 49616 0 1 40768
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _3408_
timestamp 1698431365
transform 1 0 54096 0 -1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3409_
timestamp 1698431365
transform 1 0 51968 0 -1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3410_
timestamp 1698431365
transform 1 0 53312 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _3411_
timestamp 1698431365
transform 1 0 52864 0 -1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3412_
timestamp 1698431365
transform 1 0 52528 0 1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _3413_
timestamp 1698431365
transform -1 0 53984 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3414_
timestamp 1698431365
transform 1 0 52976 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _3415_
timestamp 1698431365
transform 1 0 53648 0 1 45472
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _3416_
timestamp 1698431365
transform -1 0 56672 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _3417_
timestamp 1698431365
transform -1 0 56224 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _3418_
timestamp 1698431365
transform -1 0 52304 0 1 36064
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _3419_
timestamp 1698431365
transform -1 0 48384 0 -1 34496
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _3420_
timestamp 1698431365
transform -1 0 44240 0 -1 34496
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _3421_
timestamp 1698431365
transform -1 0 44912 0 -1 32928
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3422_
timestamp 1698431365
transform -1 0 37520 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3423_
timestamp 1698431365
transform 1 0 31920 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3424_
timestamp 1698431365
transform 1 0 33040 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _3425_
timestamp 1698431365
transform 1 0 34832 0 -1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3426_
timestamp 1698431365
transform -1 0 36848 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3427_
timestamp 1698431365
transform 1 0 35392 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _3428_
timestamp 1698431365
transform 1 0 33712 0 -1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _3429_
timestamp 1698431365
transform -1 0 33824 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3430_
timestamp 1698431365
transform 1 0 29120 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3431_
timestamp 1698431365
transform -1 0 45360 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3432_
timestamp 1698431365
transform -1 0 48720 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _3433_
timestamp 1698431365
transform -1 0 47376 0 1 32928
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3434_
timestamp 1698431365
transform 1 0 49056 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _3435_
timestamp 1698431365
transform 1 0 49504 0 1 37632
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _3436_
timestamp 1698431365
transform -1 0 53424 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _3437_
timestamp 1698431365
transform -1 0 52640 0 -1 36064
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  _3438_
timestamp 1698431365
transform -1 0 53424 0 -1 37632
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3439_
timestamp 1698431365
transform 1 0 51744 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _3440_
timestamp 1698431365
transform -1 0 55328 0 -1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _3441_
timestamp 1698431365
transform 1 0 52752 0 -1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3442_
timestamp 1698431365
transform 1 0 55104 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _3443_
timestamp 1698431365
transform -1 0 51744 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3444_
timestamp 1698431365
transform 1 0 53312 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3445_
timestamp 1698431365
transform 1 0 54880 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _3446_
timestamp 1698431365
transform 1 0 53984 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  _3447_
timestamp 1698431365
transform -1 0 58352 0 1 42336
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3448_
timestamp 1698431365
transform 1 0 52528 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3449_
timestamp 1698431365
transform 1 0 53984 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3450_
timestamp 1698431365
transform -1 0 54992 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3451_
timestamp 1698431365
transform 1 0 53648 0 1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _3452_
timestamp 1698431365
transform 1 0 53424 0 1 37632
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _3453_
timestamp 1698431365
transform -1 0 56224 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _3454_
timestamp 1698431365
transform -1 0 51632 0 1 32928
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _3455_
timestamp 1698431365
transform -1 0 45696 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _3456_
timestamp 1698431365
transform -1 0 46704 0 -1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3457_
timestamp 1698431365
transform -1 0 33712 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3458_
timestamp 1698431365
transform 1 0 30352 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _3459_
timestamp 1698431365
transform 1 0 31920 0 1 40768
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3460_
timestamp 1698431365
transform 1 0 33712 0 1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _3461_
timestamp 1698431365
transform -1 0 35392 0 1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3462_
timestamp 1698431365
transform -1 0 30240 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _3463_
timestamp 1698431365
transform -1 0 39424 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3464_
timestamp 1698431365
transform -1 0 50960 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3465_
timestamp 1698431365
transform -1 0 49952 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3466_
timestamp 1698431365
transform -1 0 50176 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _3467_
timestamp 1698431365
transform -1 0 55440 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _3468_
timestamp 1698431365
transform -1 0 54992 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _3469_
timestamp 1698431365
transform 1 0 52528 0 1 34496
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _3470_
timestamp 1698431365
transform -1 0 53200 0 -1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3471_
timestamp 1698431365
transform 1 0 51968 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3472_
timestamp 1698431365
transform -1 0 55104 0 -1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _3473_
timestamp 1698431365
transform 1 0 52528 0 1 32928
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3474_
timestamp 1698431365
transform 1 0 51408 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3475_
timestamp 1698431365
transform 1 0 52640 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3476_
timestamp 1698431365
transform 1 0 53200 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _3477_
timestamp 1698431365
transform 1 0 54992 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _3478_
timestamp 1698431365
transform -1 0 55664 0 -1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3479_
timestamp 1698431365
transform -1 0 55328 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _3480_
timestamp 1698431365
transform -1 0 55216 0 1 31360
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _3481_
timestamp 1698431365
transform -1 0 51968 0 -1 31360
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _3482_
timestamp 1698431365
transform 1 0 48608 0 -1 31360
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _3483_
timestamp 1698431365
transform 1 0 48384 0 1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3484_
timestamp 1698431365
transform -1 0 37856 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3485_
timestamp 1698431365
transform 1 0 33152 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _3486_
timestamp 1698431365
transform 1 0 33824 0 1 39200
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3487_
timestamp 1698431365
transform 1 0 34944 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3488_
timestamp 1698431365
transform 1 0 37856 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3489_
timestamp 1698431365
transform 1 0 37744 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _3490_
timestamp 1698431365
transform 1 0 37856 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _3491_
timestamp 1698431365
transform 1 0 53648 0 -1 32928
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _3492_
timestamp 1698431365
transform -1 0 55104 0 1 29792
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3493_
timestamp 1698431365
transform -1 0 51520 0 1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _3494_
timestamp 1698431365
transform 1 0 48720 0 1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3495_
timestamp 1698431365
transform -1 0 46816 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _3496_
timestamp 1698431365
transform 1 0 56448 0 -1 32928
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3497_
timestamp 1698431365
transform -1 0 55216 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _3498_
timestamp 1698431365
transform -1 0 54544 0 -1 31360
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3499_
timestamp 1698431365
transform 1 0 46928 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3500_
timestamp 1698431365
transform 1 0 52528 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _3501_
timestamp 1698431365
transform -1 0 52304 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3502_
timestamp 1698431365
transform -1 0 48384 0 -1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3503_
timestamp 1698431365
transform -1 0 48272 0 1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _3504_
timestamp 1698431365
transform -1 0 46144 0 1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3505_
timestamp 1698431365
transform 1 0 46144 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3506_
timestamp 1698431365
transform -1 0 44464 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3507_
timestamp 1698431365
transform -1 0 38192 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3508_
timestamp 1698431365
transform -1 0 36624 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3509_
timestamp 1698431365
transform 1 0 36848 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _3510_
timestamp 1698431365
transform -1 0 37744 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3511_
timestamp 1698431365
transform -1 0 36176 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3512_
timestamp 1698431365
transform -1 0 38752 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3513_
timestamp 1698431365
transform 1 0 36960 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3514_
timestamp 1698431365
transform -1 0 46368 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3515_
timestamp 1698431365
transform 1 0 44240 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3516_
timestamp 1698431365
transform -1 0 46256 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _3517_
timestamp 1698431365
transform -1 0 48384 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3518_
timestamp 1698431365
transform 1 0 46144 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3519_
timestamp 1698431365
transform -1 0 45808 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _3520_
timestamp 1698431365
transform -1 0 43792 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _3521_
timestamp 1698431365
transform 1 0 41216 0 -1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3522_
timestamp 1698431365
transform -1 0 38416 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3523_
timestamp 1698431365
transform -1 0 38752 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _3524_
timestamp 1698431365
transform -1 0 42000 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3525_
timestamp 1698431365
transform -1 0 39536 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3526_
timestamp 1698431365
transform -1 0 43456 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3527_
timestamp 1698431365
transform 1 0 42000 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _3528_
timestamp 1698431365
transform -1 0 46032 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _3529_
timestamp 1698431365
transform -1 0 40880 0 1 34496
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _3530_
timestamp 1698431365
transform 1 0 39984 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _3531_
timestamp 1698431365
transform 1 0 40768 0 -1 29792
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3532_
timestamp 1698431365
transform -1 0 39648 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3533_
timestamp 1698431365
transform -1 0 42112 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3534_
timestamp 1698431365
transform 1 0 39648 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3535_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 16352 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3536_
timestamp 1698431365
transform -1 0 18256 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3537_
timestamp 1698431365
transform -1 0 20496 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3538_
timestamp 1698431365
transform -1 0 16576 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3539_
timestamp 1698431365
transform 1 0 24864 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3540_
timestamp 1698431365
transform -1 0 20720 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3541_
timestamp 1698431365
transform 1 0 28112 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3542_
timestamp 1698431365
transform 1 0 25536 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3543_
timestamp 1698431365
transform -1 0 24864 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3544_
timestamp 1698431365
transform -1 0 24864 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _3545_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 24864 0 1 29792
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _3546_
timestamp 1698431365
transform 1 0 30688 0 1 36064
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3547_
timestamp 1698431365
transform -1 0 25984 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3548_
timestamp 1698431365
transform 1 0 26208 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3549_
timestamp 1698431365
transform 1 0 25872 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3550_
timestamp 1698431365
transform 1 0 23968 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _3551_
timestamp 1698431365
transform -1 0 23968 0 -1 26656
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3552_
timestamp 1698431365
transform 1 0 25312 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3553_
timestamp 1698431365
transform 1 0 36176 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _3554_
timestamp 1698431365
transform 1 0 29008 0 1 25088
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3555_
timestamp 1698431365
transform 1 0 35056 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3556_
timestamp 1698431365
transform 1 0 29344 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3557_
timestamp 1698431365
transform 1 0 32704 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3558_
timestamp 1698431365
transform 1 0 34272 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3559_
timestamp 1698431365
transform 1 0 29456 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3560_
timestamp 1698431365
transform 1 0 34608 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _3561_
timestamp 1698431365
transform 1 0 32144 0 1 37632
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _3562_
timestamp 1698431365
transform -1 0 31024 0 -1 34496
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3563_
timestamp 1698431365
transform 1 0 36848 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3564_
timestamp 1698431365
transform 1 0 36848 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3565_
timestamp 1698431365
transform 1 0 40768 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3566_
timestamp 1698431365
transform 1 0 40096 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3567_
timestamp 1698431365
transform 1 0 39648 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3569_
timestamp 1698431365
transform 1 0 42672 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1767__A2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18928 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1767__A3
timestamp 1698431365
transform 1 0 19376 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1768__A1
timestamp 1698431365
transform -1 0 18256 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1769__A1
timestamp 1698431365
transform -1 0 19152 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1770__A1
timestamp 1698431365
transform 1 0 18592 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1770__A2
timestamp 1698431365
transform 1 0 17584 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1771__A1
timestamp 1698431365
transform 1 0 20720 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1771__A2
timestamp 1698431365
transform -1 0 20160 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1771__A3
timestamp 1698431365
transform -1 0 19712 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1772__A1
timestamp 1698431365
transform -1 0 20272 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1772__A2
timestamp 1698431365
transform -1 0 20160 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1772__A3
timestamp 1698431365
transform 1 0 18032 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1772__A4
timestamp 1698431365
transform -1 0 20608 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1779__I
timestamp 1698431365
transform -1 0 16016 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1781__I
timestamp 1698431365
transform 1 0 12880 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1790__A2
timestamp 1698431365
transform 1 0 5488 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1791__A1
timestamp 1698431365
transform 1 0 8400 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1797__A2
timestamp 1698431365
transform -1 0 8064 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1830__A2
timestamp 1698431365
transform -1 0 12768 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1853__A2
timestamp 1698431365
transform -1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1859__A2
timestamp 1698431365
transform 1 0 13552 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1874__A1
timestamp 1698431365
transform 1 0 3696 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1874__A4
timestamp 1698431365
transform 1 0 5040 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1877__A1
timestamp 1698431365
transform 1 0 2464 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1877__B1
timestamp 1698431365
transform -1 0 2576 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1900__A2
timestamp 1698431365
transform 1 0 14896 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1909__A1
timestamp 1698431365
transform -1 0 13776 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1919__I
timestamp 1698431365
transform 1 0 7616 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1920__A2
timestamp 1698431365
transform -1 0 3696 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1921__A1
timestamp 1698431365
transform -1 0 3472 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1931__A2
timestamp 1698431365
transform -1 0 24080 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1933__I
timestamp 1698431365
transform -1 0 23856 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1947__A1
timestamp 1698431365
transform 1 0 16576 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1947__A2
timestamp 1698431365
transform -1 0 16352 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1972__A2
timestamp 1698431365
transform 1 0 4144 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1974__A1
timestamp 1698431365
transform 1 0 4592 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1991__I
timestamp 1698431365
transform -1 0 29008 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1992__A1
timestamp 1698431365
transform 1 0 27776 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1992__A2
timestamp 1698431365
transform -1 0 23744 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1995__I
timestamp 1698431365
transform 1 0 20720 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1996__A1
timestamp 1698431365
transform 1 0 29232 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1996__A2
timestamp 1698431365
transform -1 0 26880 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1997__A1
timestamp 1698431365
transform 1 0 27888 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1998__I
timestamp 1698431365
transform 1 0 26992 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1999__A1
timestamp 1698431365
transform 1 0 31472 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1999__A3
timestamp 1698431365
transform 1 0 27440 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2002__A1
timestamp 1698431365
transform -1 0 18816 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2006__I1
timestamp 1698431365
transform -1 0 15456 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2011__A1
timestamp 1698431365
transform 1 0 25312 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2015__A2
timestamp 1698431365
transform 1 0 22624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2030__A1
timestamp 1698431365
transform 1 0 14560 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2038__A1
timestamp 1698431365
transform 1 0 9184 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2047__A2
timestamp 1698431365
transform 1 0 12320 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2049__A2
timestamp 1698431365
transform 1 0 18704 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2056__A2
timestamp 1698431365
transform 1 0 27104 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2080__A1
timestamp 1698431365
transform 1 0 14896 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2106__A2
timestamp 1698431365
transform 1 0 20720 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2131__A1
timestamp 1698431365
transform 1 0 16128 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2139__B1
timestamp 1698431365
transform 1 0 19152 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2157__A1
timestamp 1698431365
transform 1 0 22288 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2170__A2
timestamp 1698431365
transform 1 0 17136 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2172__A2
timestamp 1698431365
transform 1 0 25760 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2175__A1
timestamp 1698431365
transform 1 0 27328 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2187__A1
timestamp 1698431365
transform 1 0 25312 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2193__B1
timestamp 1698431365
transform 1 0 21840 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2193__B2
timestamp 1698431365
transform -1 0 21168 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2195__I1
timestamp 1698431365
transform -1 0 19264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2195__S
timestamp 1698431365
transform 1 0 20496 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2201__A1
timestamp 1698431365
transform -1 0 23744 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2204__A2
timestamp 1698431365
transform -1 0 23856 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2206__A2
timestamp 1698431365
transform 1 0 29344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2207__A1
timestamp 1698431365
transform 1 0 30464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2214__A2
timestamp 1698431365
transform 1 0 26544 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2215__A1
timestamp 1698431365
transform 1 0 28112 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2218__A1
timestamp 1698431365
transform 1 0 22176 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2224__A2
timestamp 1698431365
transform 1 0 42112 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2225__I
timestamp 1698431365
transform 1 0 42448 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2226__I
timestamp 1698431365
transform -1 0 40656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2228__I
timestamp 1698431365
transform -1 0 36848 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2277__A2
timestamp 1698431365
transform 1 0 37072 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2304__A2
timestamp 1698431365
transform -1 0 41104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2310__A2
timestamp 1698431365
transform -1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2330__A2
timestamp 1698431365
transform 1 0 46592 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2340__A2
timestamp 1698431365
transform -1 0 38416 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2373__A2
timestamp 1698431365
transform 1 0 52640 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2383__A1
timestamp 1698431365
transform -1 0 42224 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2420__A1
timestamp 1698431365
transform 1 0 49504 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2422__A1
timestamp 1698431365
transform 1 0 49952 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2441__A2
timestamp 1698431365
transform 1 0 33264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2441__A3
timestamp 1698431365
transform -1 0 32256 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2445__A1
timestamp 1698431365
transform 1 0 33152 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2448__A1
timestamp 1698431365
transform 1 0 30128 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2456__A1
timestamp 1698431365
transform 1 0 44912 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2469__A1
timestamp 1698431365
transform 1 0 50064 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2492__A1
timestamp 1698431365
transform 1 0 37072 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2492__B1
timestamp 1698431365
transform -1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2495__B1
timestamp 1698431365
transform 1 0 36400 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2495__B2
timestamp 1698431365
transform 1 0 32816 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2496__A1
timestamp 1698431365
transform -1 0 26432 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2496__A2
timestamp 1698431365
transform 1 0 23072 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2497__A1
timestamp 1698431365
transform -1 0 22848 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2501__I
timestamp 1698431365
transform 1 0 46032 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2522__A1
timestamp 1698431365
transform 1 0 53200 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2544__B1
timestamp 1698431365
transform 1 0 36400 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2544__B2
timestamp 1698431365
transform 1 0 33152 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2546__A1
timestamp 1698431365
transform -1 0 24304 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2549__A1
timestamp 1698431365
transform 1 0 34384 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2549__A2
timestamp 1698431365
transform 1 0 31920 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2550__A1
timestamp 1698431365
transform -1 0 30128 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2574__A1
timestamp 1698431365
transform 1 0 54544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2583__A1
timestamp 1698431365
transform 1 0 32144 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2584__A2
timestamp 1698431365
transform 1 0 29680 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2597__A1
timestamp 1698431365
transform -1 0 54432 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2611__A2
timestamp 1698431365
transform 1 0 36400 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2619__A2
timestamp 1698431365
transform 1 0 28112 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2621__A1
timestamp 1698431365
transform 1 0 24640 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2631__A1
timestamp 1698431365
transform 1 0 52080 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2640__B2
timestamp 1698431365
transform 1 0 32480 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2641__A2
timestamp 1698431365
transform 1 0 30464 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2642__I1
timestamp 1698431365
transform -1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2642__S
timestamp 1698431365
transform -1 0 29568 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2645__A1
timestamp 1698431365
transform 1 0 53760 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2651__A2
timestamp 1698431365
transform -1 0 36064 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2654__A2
timestamp 1698431365
transform -1 0 25536 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2655__A1
timestamp 1698431365
transform 1 0 29232 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2660__A2
timestamp 1698431365
transform 1 0 37968 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2660__C
timestamp 1698431365
transform 1 0 33712 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2661__A2
timestamp 1698431365
transform 1 0 27104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2662__A1
timestamp 1698431365
transform 1 0 27440 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2668__A2
timestamp 1698431365
transform 1 0 22848 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2669__I
timestamp 1698431365
transform 1 0 15904 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2673__I
timestamp 1698431365
transform -1 0 10528 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2702__A2
timestamp 1698431365
transform 1 0 12544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2707__A1
timestamp 1698431365
transform 1 0 5712 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2724__A2
timestamp 1698431365
transform 1 0 13552 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2746__A2
timestamp 1698431365
transform -1 0 18816 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2755__A1
timestamp 1698431365
transform -1 0 5936 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2756__A1
timestamp 1698431365
transform -1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2774__A2
timestamp 1698431365
transform -1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2785__A2
timestamp 1698431365
transform 1 0 25536 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2796__A2
timestamp 1698431365
transform 1 0 15344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2822__A2
timestamp 1698431365
transform 1 0 5712 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2824__A1
timestamp 1698431365
transform 1 0 6496 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2838__A1
timestamp 1698431365
transform 1 0 20944 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2873__A1
timestamp 1698431365
transform -1 0 5712 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2875__A1
timestamp 1698431365
transform 1 0 7616 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2884__A2
timestamp 1698431365
transform -1 0 24752 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2885__B2
timestamp 1698431365
transform -1 0 26544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2886__A2
timestamp 1698431365
transform 1 0 34496 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2888__A1
timestamp 1698431365
transform 1 0 24192 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2888__A2
timestamp 1698431365
transform -1 0 22736 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2901__I
timestamp 1698431365
transform 1 0 23520 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2925__A2
timestamp 1698431365
transform 1 0 12768 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2940__A1
timestamp 1698431365
transform 1 0 29120 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2941__A1
timestamp 1698431365
transform 1 0 25088 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2941__B1
timestamp 1698431365
transform 1 0 23296 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2942__A1
timestamp 1698431365
transform -1 0 25200 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2942__A2
timestamp 1698431365
transform 1 0 23632 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2944__C
timestamp 1698431365
transform 1 0 29232 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2945__A2
timestamp 1698431365
transform 1 0 28560 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2946__A1
timestamp 1698431365
transform 1 0 28336 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2948__A1
timestamp 1698431365
transform -1 0 39088 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2948__A2
timestamp 1698431365
transform 1 0 38416 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2975__A2
timestamp 1698431365
transform 1 0 14896 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2993__A2
timestamp 1698431365
transform 1 0 35168 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3012__A2
timestamp 1698431365
transform 1 0 19824 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3023__A1
timestamp 1698431365
transform -1 0 15568 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3028__A1
timestamp 1698431365
transform -1 0 31696 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3030__A2
timestamp 1698431365
transform 1 0 38192 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3042__I
timestamp 1698431365
transform 1 0 25312 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3053__A1
timestamp 1698431365
transform 1 0 20496 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3073__A1
timestamp 1698431365
transform 1 0 29232 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3075__A1
timestamp 1698431365
transform 1 0 22176 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3077__C
timestamp 1698431365
transform 1 0 29344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3089__B
timestamp 1698431365
transform -1 0 33376 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3091__A1
timestamp 1698431365
transform 1 0 24080 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3093__C
timestamp 1698431365
transform -1 0 33712 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3100__C
timestamp 1698431365
transform -1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3102__A1
timestamp 1698431365
transform 1 0 36400 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3107__I
timestamp 1698431365
transform 1 0 41776 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3108__A2
timestamp 1698431365
transform -1 0 37296 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3109__I
timestamp 1698431365
transform 1 0 40544 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3111__I
timestamp 1698431365
transform 1 0 34048 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3159__A2
timestamp 1698431365
transform 1 0 37296 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3186__A2
timestamp 1698431365
transform 1 0 38192 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3214__A2
timestamp 1698431365
transform -1 0 42448 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3225__A2
timestamp 1698431365
transform 1 0 39872 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3236__A2
timestamp 1698431365
transform 1 0 41104 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3262__A2
timestamp 1698431365
transform -1 0 47936 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3264__A1
timestamp 1698431365
transform 1 0 49616 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3274__A1
timestamp 1698431365
transform -1 0 39536 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3278__A1
timestamp 1698431365
transform 1 0 44016 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3313__A1
timestamp 1698431365
transform 1 0 50848 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3315__A1
timestamp 1698431365
transform 1 0 49056 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3324__A2
timestamp 1698431365
transform -1 0 38864 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3325__B2
timestamp 1698431365
transform 1 0 32704 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3327__S
timestamp 1698431365
transform 1 0 31136 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3329__A1
timestamp 1698431365
transform -1 0 37632 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3329__A2
timestamp 1698431365
transform 1 0 36624 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3341__I
timestamp 1698431365
transform 1 0 46144 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3382__A1
timestamp 1698431365
transform 1 0 39984 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3382__B1
timestamp 1698431365
transform -1 0 39760 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3383__A1
timestamp 1698431365
transform 1 0 34160 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3424__A1
timestamp 1698431365
transform -1 0 33936 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3428__I1
timestamp 1698431365
transform 1 0 35616 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3428__S
timestamp 1698431365
transform 1 0 33488 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3430__A1
timestamp 1698431365
transform 1 0 28896 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3459__A1
timestamp 1698431365
transform -1 0 31920 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3484__A1
timestamp 1698431365
transform 1 0 39648 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3486__A1
timestamp 1698431365
transform 1 0 34048 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3508__A1
timestamp 1698431365
transform -1 0 36064 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3510__C
timestamp 1698431365
transform 1 0 36624 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3512__A1
timestamp 1698431365
transform -1 0 39984 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3512__A2
timestamp 1698431365
transform -1 0 38640 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3521__B
timestamp 1698431365
transform 1 0 40992 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3522__A1
timestamp 1698431365
transform 1 0 38640 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3526__A2
timestamp 1698431365
transform 1 0 43680 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3531__B2
timestamp 1698431365
transform 1 0 39872 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3531__C
timestamp 1698431365
transform 1 0 40320 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3532__A2
timestamp 1698431365
transform -1 0 40432 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3533__A2
timestamp 1698431365
transform -1 0 42560 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3535__CLK
timestamp 1698431365
transform 1 0 16576 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3537__CLK
timestamp 1698431365
transform 1 0 20272 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3539__CLK
timestamp 1698431365
transform 1 0 24640 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3540__CLK
timestamp 1698431365
transform 1 0 21392 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3541__CLK
timestamp 1698431365
transform 1 0 31584 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3542__CLK
timestamp 1698431365
transform 1 0 25312 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3543__CLK
timestamp 1698431365
transform 1 0 25312 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3544__CLK
timestamp 1698431365
transform 1 0 22960 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3546__CLK
timestamp 1698431365
transform 1 0 34832 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3548__CLK
timestamp 1698431365
transform 1 0 25984 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3553__CLK
timestamp 1698431365
transform 1 0 39424 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3554__CLK
timestamp 1698431365
transform 1 0 32480 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3555__CLK
timestamp 1698431365
transform 1 0 38528 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3556__CLK
timestamp 1698431365
transform 1 0 33152 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3557__CLK
timestamp 1698431365
transform 1 0 37072 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3558__CLK
timestamp 1698431365
transform 1 0 37744 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3559__CLK
timestamp 1698431365
transform 1 0 33264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3560__CLK
timestamp 1698431365
transform 1 0 39088 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3561__CLK
timestamp 1698431365
transform 1 0 35840 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3562__CLK
timestamp 1698431365
transform 1 0 30464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3563__CLK
timestamp 1698431365
transform 1 0 40320 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3564__CLK
timestamp 1698431365
transform 1 0 40992 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3565__CLK
timestamp 1698431365
transform -1 0 40880 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3566__CLK
timestamp 1698431365
transform 1 0 39872 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3567__CLK
timestamp 1698431365
transform -1 0 39648 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698431365
transform -1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform 1 0 2464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform -1 0 24304 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform -1 0 26320 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform 1 0 28560 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform 1 0 4704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform -1 0 2016 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform 1 0 3584 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698431365
transform 1 0 3136 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698431365
transform 1 0 3920 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698431365
transform 1 0 3136 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698431365
transform 1 0 2912 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698431365
transform 1 0 1792 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698431365
transform 1 0 3808 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1698431365
transform 1 0 2464 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1698431365
transform 1 0 3136 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1698431365
transform 1 0 4256 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1698431365
transform 1 0 6272 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1698431365
transform 1 0 1792 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1698431365
transform 1 0 46816 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1698431365
transform 1 0 45584 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1698431365
transform 1 0 47040 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input22_I
timestamp 1698431365
transform 1 0 49280 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input23_I
timestamp 1698431365
transform 1 0 48832 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input24_I
timestamp 1698431365
transform -1 0 49840 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input25_I
timestamp 1698431365
transform 1 0 3360 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input26_I
timestamp 1698431365
transform 1 0 3808 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input27_I
timestamp 1698431365
transform 1 0 3584 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input28_I
timestamp 1698431365
transform 1 0 3584 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input29_I
timestamp 1698431365
transform 1 0 8512 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input30_I
timestamp 1698431365
transform 1 0 4032 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input31_I
timestamp 1698431365
transform 1 0 4928 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input32_I
timestamp 1698431365
transform 1 0 2464 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input33_I
timestamp 1698431365
transform 1 0 2464 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input34_I
timestamp 1698431365
transform -1 0 28560 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input35_I
timestamp 1698431365
transform -1 0 29008 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input36_I
timestamp 1698431365
transform -1 0 30352 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input37_I
timestamp 1698431365
transform 1 0 42000 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input38_I
timestamp 1698431365
transform 1 0 43680 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input39_I
timestamp 1698431365
transform 1 0 40992 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input40_I
timestamp 1698431365
transform 1 0 8848 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input41_I
timestamp 1698431365
transform -1 0 49840 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input42_I
timestamp 1698431365
transform -1 0 51072 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input43_I
timestamp 1698431365
transform -1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input44_I
timestamp 1698431365
transform 1 0 1792 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input45_I
timestamp 1698431365
transform -1 0 2128 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input46_I
timestamp 1698431365
transform 1 0 2464 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input47_I
timestamp 1698431365
transform 1 0 2912 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input48_I
timestamp 1698431365
transform 1 0 42448 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input49_I
timestamp 1698431365
transform -1 0 28336 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input50_I
timestamp 1698431365
transform 1 0 9632 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input51_I
timestamp 1698431365
transform 1 0 47712 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input52_I
timestamp 1698431365
transform 1 0 47264 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input53_I
timestamp 1698431365
transform 1 0 48160 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input54_I
timestamp 1698431365
transform 1 0 48832 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input55_I
timestamp 1698431365
transform -1 0 58352 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input56_I
timestamp 1698431365
transform -1 0 57680 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input57_I
timestamp 1698431365
transform 1 0 1792 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input58_I
timestamp 1698431365
transform 1 0 6720 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input59_I
timestamp 1698431365
transform 1 0 2464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input60_I
timestamp 1698431365
transform 1 0 3136 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input61_I
timestamp 1698431365
transform 1 0 3584 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input62_I
timestamp 1698431365
transform 1 0 2464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input63_I
timestamp 1698431365
transform 1 0 5712 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input64_I
timestamp 1698431365
transform -1 0 22288 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input65_I
timestamp 1698431365
transform 1 0 25312 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input66_I
timestamp 1698431365
transform 1 0 28112 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input67_I
timestamp 1698431365
transform 1 0 31248 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input68_I
timestamp 1698431365
transform 1 0 36400 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input69_I
timestamp 1698431365
transform 1 0 43008 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input70_I
timestamp 1698431365
transform 1 0 42560 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input71_I
timestamp 1698431365
transform 1 0 42448 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input72_I
timestamp 1698431365
transform 1 0 2800 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input73_I
timestamp 1698431365
transform -1 0 57680 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input74_I
timestamp 1698431365
transform -1 0 57680 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input75_I
timestamp 1698431365
transform 1 0 8176 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input76_I
timestamp 1698431365
transform 1 0 3696 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input77_I
timestamp 1698431365
transform 1 0 4480 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input78_I
timestamp 1698431365
transform 1 0 9408 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input79_I
timestamp 1698431365
transform -1 0 23520 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input80_I
timestamp 1698431365
transform -1 0 29344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input81_I
timestamp 1698431365
transform -1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input82_I
timestamp 1698431365
transform 1 0 5712 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output83_I
timestamp 1698431365
transform 1 0 8960 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output84_I
timestamp 1698431365
transform -1 0 8176 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output85_I
timestamp 1698431365
transform 1 0 42112 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output86_I
timestamp 1698431365
transform -1 0 4368 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output87_I
timestamp 1698431365
transform 1 0 32144 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output88_I
timestamp 1698431365
transform 1 0 32368 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output89_I
timestamp 1698431365
transform 1 0 27664 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output90_I
timestamp 1698431365
transform -1 0 4704 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output91_I
timestamp 1698431365
transform 1 0 29344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output92_I
timestamp 1698431365
transform 1 0 58128 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output93_I
timestamp 1698431365
transform 1 0 36400 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output98_I
timestamp 1698431365
transform 1 0 40320 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output100_I
timestamp 1698431365
transform 1 0 56000 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output101_I
timestamp 1698431365
transform 1 0 41552 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output102_I
timestamp 1698431365
transform 1 0 27440 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output104_I
timestamp 1698431365
transform 1 0 57344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output109_I
timestamp 1698431365
transform 1 0 27888 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output110_I
timestamp 1698431365
transform -1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output111_I
timestamp 1698431365
transform 1 0 31808 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output112_I
timestamp 1698431365
transform 1 0 31696 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output113_I
timestamp 1698431365
transform -1 0 5488 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output114_I
timestamp 1698431365
transform 1 0 9296 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 27104 0 -1 31360
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1698431365
transform -1 0 27328 0 1 28224
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1698431365
transform -1 0 27552 0 1 32928
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1698431365
transform 1 0 34832 0 -1 26656
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1698431365
transform 1 0 33600 0 -1 32928
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698431365
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 16800 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_154 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18592 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_162 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19488 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_167 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 20048 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_169
timestamp 1698431365
transform 1 0 20272 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_172
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_180 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21504 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_184
timestamp 1698431365
transform 1 0 21952 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_193
timestamp 1698431365
transform 1 0 22960 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_201
timestamp 1698431365
transform 1 0 23856 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_203
timestamp 1698431365
transform 1 0 24080 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_350
timestamp 1698431365
transform 1 0 40544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_406
timestamp 1698431365
transform 1 0 46816 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_422
timestamp 1698431365
transform 1 0 48608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_426
timestamp 1698431365
transform 1 0 49056 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_430
timestamp 1698431365
transform 1 0 49504 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_432
timestamp 1698431365
transform 1 0 49728 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_439
timestamp 1698431365
transform 1 0 50512 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_441
timestamp 1698431365
transform 1 0 50736 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_444
timestamp 1698431365
transform 1 0 51072 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_478
timestamp 1698431365
transform 1 0 54880 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_494
timestamp 1698431365
transform 1 0 56672 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_502
timestamp 1698431365
transform 1 0 57568 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_506
timestamp 1698431365
transform 1 0 58016 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_508
timestamp 1698431365
transform 1 0 58240 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698431365
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698431365
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_142
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_206
timestamp 1698431365
transform 1 0 24416 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_212
timestamp 1698431365
transform 1 0 25088 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_216
timestamp 1698431365
transform 1 0 25536 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_232
timestamp 1698431365
transform 1 0 27328 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_234
timestamp 1698431365
transform 1 0 27552 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_237
timestamp 1698431365
transform 1 0 27888 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_267
timestamp 1698431365
transform 1 0 31248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698431365
transform 1 0 40096 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_358
timestamp 1698431365
transform 1 0 41440 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_404
timestamp 1698431365
transform 1 0 46592 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_408
timestamp 1698431365
transform 1 0 47040 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_412
timestamp 1698431365
transform 1 0 47488 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_416
timestamp 1698431365
transform 1 0 47936 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_422
timestamp 1698431365
transform 1 0 48608 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_426
timestamp 1698431365
transform 1 0 49056 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_430
timestamp 1698431365
transform 1 0 49504 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_433
timestamp 1698431365
transform 1 0 49840 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_465
timestamp 1698431365
transform 1 0 53424 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_481
timestamp 1698431365
transform 1 0 55216 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_489
timestamp 1698431365
transform 1 0 56112 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_492
timestamp 1698431365
transform 1 0 56448 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_508
timestamp 1698431365
transform 1 0 58240 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698431365
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698431365
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_107
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_139
timestamp 1698431365
transform 1 0 16912 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_143
timestamp 1698431365
transform 1 0 17360 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_145
timestamp 1698431365
transform 1 0 17584 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_177
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_181
timestamp 1698431365
transform 1 0 21616 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_190
timestamp 1698431365
transform 1 0 22624 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_222
timestamp 1698431365
transform 1 0 26208 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_238
timestamp 1698431365
transform 1 0 28000 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_247
timestamp 1698431365
transform 1 0 29008 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_249
timestamp 1698431365
transform 1 0 29232 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_303
timestamp 1698431365
transform 1 0 35280 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_305
timestamp 1698431365
transform 1 0 35504 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_317
timestamp 1698431365
transform 1 0 36848 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_369
timestamp 1698431365
transform 1 0 42672 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_393
timestamp 1698431365
transform 1 0 45360 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_419
timestamp 1698431365
transform 1 0 48272 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_423
timestamp 1698431365
transform 1 0 48720 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_439
timestamp 1698431365
transform 1 0 50512 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_457
timestamp 1698431365
transform 1 0 52528 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_489
timestamp 1698431365
transform 1 0 56112 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_505
timestamp 1698431365
transform 1 0 57904 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698431365
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_88
timestamp 1698431365
transform 1 0 11200 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_100
timestamp 1698431365
transform 1 0 12544 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_113
timestamp 1698431365
transform 1 0 14000 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_129
timestamp 1698431365
transform 1 0 15792 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698431365
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_142
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_150
timestamp 1698431365
transform 1 0 18144 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_195
timestamp 1698431365
transform 1 0 23184 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_203
timestamp 1698431365
transform 1 0 24080 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_207
timestamp 1698431365
transform 1 0 24528 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_209
timestamp 1698431365
transform 1 0 24752 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_212
timestamp 1698431365
transform 1 0 25088 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_244
timestamp 1698431365
transform 1 0 28672 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_274
timestamp 1698431365
transform 1 0 32032 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_290
timestamp 1698431365
transform 1 0 33824 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_365
timestamp 1698431365
transform 1 0 42224 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_394
timestamp 1698431365
transform 1 0 45472 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_396
timestamp 1698431365
transform 1 0 45696 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_402
timestamp 1698431365
transform 1 0 46368 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_406
timestamp 1698431365
transform 1 0 46816 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_410
timestamp 1698431365
transform 1 0 47264 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_418
timestamp 1698431365
transform 1 0 48160 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_456
timestamp 1698431365
transform 1 0 52416 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_460
timestamp 1698431365
transform 1 0 52864 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_476
timestamp 1698431365
transform 1 0 54656 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_484
timestamp 1698431365
transform 1 0 55552 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_488
timestamp 1698431365
transform 1 0 56000 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_492
timestamp 1698431365
transform 1 0 56448 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_508
timestamp 1698431365
transform 1 0 58240 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_69
timestamp 1698431365
transform 1 0 9072 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_75
timestamp 1698431365
transform 1 0 9744 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_79
timestamp 1698431365
transform 1 0 10192 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_81
timestamp 1698431365
transform 1 0 10416 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_102
timestamp 1698431365
transform 1 0 12768 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_104
timestamp 1698431365
transform 1 0 12992 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_160
timestamp 1698431365
transform 1 0 19264 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_164
timestamp 1698431365
transform 1 0 19712 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_172
timestamp 1698431365
transform 1 0 20608 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_174
timestamp 1698431365
transform 1 0 20832 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_177
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_191
timestamp 1698431365
transform 1 0 22736 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_217
timestamp 1698431365
transform 1 0 25648 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_233
timestamp 1698431365
transform 1 0 27440 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_240
timestamp 1698431365
transform 1 0 28224 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_244
timestamp 1698431365
transform 1 0 28672 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_247
timestamp 1698431365
transform 1 0 29008 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_255
timestamp 1698431365
transform 1 0 29904 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_275
timestamp 1698431365
transform 1 0 32144 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_311
timestamp 1698431365
transform 1 0 36176 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_356
timestamp 1698431365
transform 1 0 41216 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_393
timestamp 1698431365
transform 1 0 45360 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_397
timestamp 1698431365
transform 1 0 45808 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_414
timestamp 1698431365
transform 1 0 47712 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_432
timestamp 1698431365
transform 1 0 49728 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_449
timestamp 1698431365
transform 1 0 51632 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_453
timestamp 1698431365
transform 1 0 52080 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_465
timestamp 1698431365
transform 1 0 53424 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_497
timestamp 1698431365
transform 1 0 57008 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_505
timestamp 1698431365
transform 1 0 57904 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_34
timestamp 1698431365
transform 1 0 5152 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_50
timestamp 1698431365
transform 1 0 6944 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_58
timestamp 1698431365
transform 1 0 7840 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_82
timestamp 1698431365
transform 1 0 10528 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_100
timestamp 1698431365
transform 1 0 12544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_104
timestamp 1698431365
transform 1 0 12992 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_108
timestamp 1698431365
transform 1 0 13440 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_110
timestamp 1698431365
transform 1 0 13664 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_117
timestamp 1698431365
transform 1 0 14448 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_138
timestamp 1698431365
transform 1 0 16800 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_142
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_146
timestamp 1698431365
transform 1 0 17696 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_157
timestamp 1698431365
transform 1 0 18928 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_159
timestamp 1698431365
transform 1 0 19152 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_177
timestamp 1698431365
transform 1 0 21168 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_209
timestamp 1698431365
transform 1 0 24752 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_212
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_268
timestamp 1698431365
transform 1 0 31360 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_294
timestamp 1698431365
transform 1 0 34272 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_314
timestamp 1698431365
transform 1 0 36512 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_333
timestamp 1698431365
transform 1 0 38640 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_335
timestamp 1698431365
transform 1 0 38864 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_346
timestamp 1698431365
transform 1 0 40096 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_401
timestamp 1698431365
transform 1 0 46256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_434
timestamp 1698431365
transform 1 0 49952 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_469
timestamp 1698431365
transform 1 0 53872 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_485
timestamp 1698431365
transform 1 0 55664 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_489
timestamp 1698431365
transform 1 0 56112 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_492
timestamp 1698431365
transform 1 0 56448 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_508
timestamp 1698431365
transform 1 0 58240 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_45
timestamp 1698431365
transform 1 0 6384 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_119
timestamp 1698431365
transform 1 0 14672 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_121
timestamp 1698431365
transform 1 0 14896 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_161
timestamp 1698431365
transform 1 0 19376 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_200
timestamp 1698431365
transform 1 0 23744 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_230
timestamp 1698431365
transform 1 0 27104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_255
timestamp 1698431365
transform 1 0 29904 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_259
timestamp 1698431365
transform 1 0 30352 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_261
timestamp 1698431365
transform 1 0 30576 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_362
timestamp 1698431365
transform 1 0 41888 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_366
timestamp 1698431365
transform 1 0 42336 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_395
timestamp 1698431365
transform 1 0 45584 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_397
timestamp 1698431365
transform 1 0 45808 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_451
timestamp 1698431365
transform 1 0 51856 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_475
timestamp 1698431365
transform 1 0 54544 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_507
timestamp 1698431365
transform 1 0 58128 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_8
timestamp 1698431365
transform 1 0 2240 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_12
timestamp 1698431365
transform 1 0 2688 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_28
timestamp 1698431365
transform 1 0 4480 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_36
timestamp 1698431365
transform 1 0 5376 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_61
timestamp 1698431365
transform 1 0 8176 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_63
timestamp 1698431365
transform 1 0 8400 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_80
timestamp 1698431365
transform 1 0 10304 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_132
timestamp 1698431365
transform 1 0 16128 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_156
timestamp 1698431365
transform 1 0 18816 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_164
timestamp 1698431365
transform 1 0 19712 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_194
timestamp 1698431365
transform 1 0 23072 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_222
timestamp 1698431365
transform 1 0 26208 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_230
timestamp 1698431365
transform 1 0 27104 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_270
timestamp 1698431365
transform 1 0 31584 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_277
timestamp 1698431365
transform 1 0 32368 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_279
timestamp 1698431365
transform 1 0 32592 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_296
timestamp 1698431365
transform 1 0 34496 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_298
timestamp 1698431365
transform 1 0 34720 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_340
timestamp 1698431365
transform 1 0 39424 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_367
timestamp 1698431365
transform 1 0 42448 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_369
timestamp 1698431365
transform 1 0 42672 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_391
timestamp 1698431365
transform 1 0 45136 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_401
timestamp 1698431365
transform 1 0 46256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_405
timestamp 1698431365
transform 1 0 46704 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_411
timestamp 1698431365
transform 1 0 47376 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_419
timestamp 1698431365
transform 1 0 48272 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_430
timestamp 1698431365
transform 1 0 49504 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_464
timestamp 1698431365
transform 1 0 53312 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_480
timestamp 1698431365
transform 1 0 55104 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_488
timestamp 1698431365
transform 1 0 56000 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_492
timestamp 1698431365
transform 1 0 56448 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_508
timestamp 1698431365
transform 1 0 58240 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_53
timestamp 1698431365
transform 1 0 7280 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_83
timestamp 1698431365
transform 1 0 10640 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_104
timestamp 1698431365
transform 1 0 12992 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_111
timestamp 1698431365
transform 1 0 13776 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_113
timestamp 1698431365
transform 1 0 14000 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_121
timestamp 1698431365
transform 1 0 14896 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_123
timestamp 1698431365
transform 1 0 15120 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_142
timestamp 1698431365
transform 1 0 17248 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_182
timestamp 1698431365
transform 1 0 21728 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_190
timestamp 1698431365
transform 1 0 22624 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_194
timestamp 1698431365
transform 1 0 23072 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_212
timestamp 1698431365
transform 1 0 25088 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_216
timestamp 1698431365
transform 1 0 25536 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_229
timestamp 1698431365
transform 1 0 26992 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_237
timestamp 1698431365
transform 1 0 27888 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_270
timestamp 1698431365
transform 1 0 31584 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_272
timestamp 1698431365
transform 1 0 31808 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_288
timestamp 1698431365
transform 1 0 33600 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_309
timestamp 1698431365
transform 1 0 35952 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_313
timestamp 1698431365
transform 1 0 36400 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_341
timestamp 1698431365
transform 1 0 39536 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_366
timestamp 1698431365
transform 1 0 42336 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_382
timestamp 1698431365
transform 1 0 44128 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_384
timestamp 1698431365
transform 1 0 44352 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_395
timestamp 1698431365
transform 1 0 45584 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_427
timestamp 1698431365
transform 1 0 49168 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_443
timestamp 1698431365
transform 1 0 50960 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_447
timestamp 1698431365
transform 1 0 51408 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_454
timestamp 1698431365
transform 1 0 52192 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_457
timestamp 1698431365
transform 1 0 52528 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_459
timestamp 1698431365
transform 1 0 52752 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_476
timestamp 1698431365
transform 1 0 54656 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_508
timestamp 1698431365
transform 1 0 58240 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_8
timestamp 1698431365
transform 1 0 2240 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_12
timestamp 1698431365
transform 1 0 2688 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_28
timestamp 1698431365
transform 1 0 4480 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_36
timestamp 1698431365
transform 1 0 5376 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_38
timestamp 1698431365
transform 1 0 5600 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_54
timestamp 1698431365
transform 1 0 7392 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_58
timestamp 1698431365
transform 1 0 7840 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698431365
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_138
timestamp 1698431365
transform 1 0 16800 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_187
timestamp 1698431365
transform 1 0 22288 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_197
timestamp 1698431365
transform 1 0 23408 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_205
timestamp 1698431365
transform 1 0 24304 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_209
timestamp 1698431365
transform 1 0 24752 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_212
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_228
timestamp 1698431365
transform 1 0 26880 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_236
timestamp 1698431365
transform 1 0 27776 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_242
timestamp 1698431365
transform 1 0 28448 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_244
timestamp 1698431365
transform 1 0 28672 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_268
timestamp 1698431365
transform 1 0 31360 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_282
timestamp 1698431365
transform 1 0 32928 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_347
timestamp 1698431365
transform 1 0 40208 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_349
timestamp 1698431365
transform 1 0 40432 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_375
timestamp 1698431365
transform 1 0 43344 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_379
timestamp 1698431365
transform 1 0 43792 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_403
timestamp 1698431365
transform 1 0 46480 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_405
timestamp 1698431365
transform 1 0 46704 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_422
timestamp 1698431365
transform 1 0 48608 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_438
timestamp 1698431365
transform 1 0 50400 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_454
timestamp 1698431365
transform 1 0 52192 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_458
timestamp 1698431365
transform 1 0 52640 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_460
timestamp 1698431365
transform 1 0 52864 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_481
timestamp 1698431365
transform 1 0 55216 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_489
timestamp 1698431365
transform 1 0 56112 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_492
timestamp 1698431365
transform 1 0 56448 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_508
timestamp 1698431365
transform 1 0 58240 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_8
timestamp 1698431365
transform 1 0 2240 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_12
timestamp 1698431365
transform 1 0 2688 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_28
timestamp 1698431365
transform 1 0 4480 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_32
timestamp 1698431365
transform 1 0 4928 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_42
timestamp 1698431365
transform 1 0 6048 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_61
timestamp 1698431365
transform 1 0 8176 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_91
timestamp 1698431365
transform 1 0 11536 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_143
timestamp 1698431365
transform 1 0 17360 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_162
timestamp 1698431365
transform 1 0 19488 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_177
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_192
timestamp 1698431365
transform 1 0 22848 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_196
timestamp 1698431365
transform 1 0 23296 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_198
timestamp 1698431365
transform 1 0 23520 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_223
timestamp 1698431365
transform 1 0 26320 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_227
timestamp 1698431365
transform 1 0 26768 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698431365
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_247
timestamp 1698431365
transform 1 0 29008 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_263
timestamp 1698431365
transform 1 0 30800 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_271
timestamp 1698431365
transform 1 0 31696 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_275
timestamp 1698431365
transform 1 0 32144 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_301
timestamp 1698431365
transform 1 0 35056 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_309
timestamp 1698431365
transform 1 0 35952 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_358
timestamp 1698431365
transform 1 0 41440 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_374
timestamp 1698431365
transform 1 0 43232 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_383
timestamp 1698431365
transform 1 0 44240 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_420
timestamp 1698431365
transform 1 0 48384 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_450
timestamp 1698431365
transform 1 0 51744 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_454
timestamp 1698431365
transform 1 0 52192 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_473
timestamp 1698431365
transform 1 0 54320 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_505
timestamp 1698431365
transform 1 0 57904 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_8
timestamp 1698431365
transform 1 0 2240 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_12
timestamp 1698431365
transform 1 0 2688 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_16
timestamp 1698431365
transform 1 0 3136 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_24
timestamp 1698431365
transform 1 0 4032 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_28
timestamp 1698431365
transform 1 0 4480 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_55
timestamp 1698431365
transform 1 0 7504 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_59
timestamp 1698431365
transform 1 0 7952 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_115
timestamp 1698431365
transform 1 0 14224 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_207
timestamp 1698431365
transform 1 0 24528 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_209
timestamp 1698431365
transform 1 0 24752 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_267
timestamp 1698431365
transform 1 0 31248 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_275
timestamp 1698431365
transform 1 0 32144 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_279
timestamp 1698431365
transform 1 0 32592 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_282
timestamp 1698431365
transform 1 0 32928 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_298
timestamp 1698431365
transform 1 0 34720 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_321
timestamp 1698431365
transform 1 0 37296 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_366
timestamp 1698431365
transform 1 0 42336 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_393
timestamp 1698431365
transform 1 0 45360 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_401
timestamp 1698431365
transform 1 0 46256 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_443
timestamp 1698431365
transform 1 0 50960 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_481
timestamp 1698431365
transform 1 0 55216 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_489
timestamp 1698431365
transform 1 0 56112 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_492
timestamp 1698431365
transform 1 0 56448 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_508
timestamp 1698431365
transform 1 0 58240 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_14
timestamp 1698431365
transform 1 0 2912 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_18
timestamp 1698431365
transform 1 0 3360 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_22
timestamp 1698431365
transform 1 0 3808 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_30
timestamp 1698431365
transform 1 0 4704 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698431365
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_37
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_46
timestamp 1698431365
transform 1 0 6496 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_53
timestamp 1698431365
transform 1 0 7280 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_61
timestamp 1698431365
transform 1 0 8176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_65
timestamp 1698431365
transform 1 0 8624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_79
timestamp 1698431365
transform 1 0 10192 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_95
timestamp 1698431365
transform 1 0 11984 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_107
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_151
timestamp 1698431365
transform 1 0 18256 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_153
timestamp 1698431365
transform 1 0 18480 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_162
timestamp 1698431365
transform 1 0 19488 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_177
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_210
timestamp 1698431365
transform 1 0 24864 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_214
timestamp 1698431365
transform 1 0 25312 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_216
timestamp 1698431365
transform 1 0 25536 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_270
timestamp 1698431365
transform 1 0 31584 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_278
timestamp 1698431365
transform 1 0 32480 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_309
timestamp 1698431365
transform 1 0 35952 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_313
timestamp 1698431365
transform 1 0 36400 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_317
timestamp 1698431365
transform 1 0 36848 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_321
timestamp 1698431365
transform 1 0 37296 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_325
timestamp 1698431365
transform 1 0 37744 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_327
timestamp 1698431365
transform 1 0 37968 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_371
timestamp 1698431365
transform 1 0 42896 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_431
timestamp 1698431365
transform 1 0 49616 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_439
timestamp 1698431365
transform 1 0 50512 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_441
timestamp 1698431365
transform 1 0 50736 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_469
timestamp 1698431365
transform 1 0 53872 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_485
timestamp 1698431365
transform 1 0 55664 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_501
timestamp 1698431365
transform 1 0 57456 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_14
timestamp 1698431365
transform 1 0 2912 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_18
timestamp 1698431365
transform 1 0 3360 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_22
timestamp 1698431365
transform 1 0 3808 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_26
timestamp 1698431365
transform 1 0 4256 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_34
timestamp 1698431365
transform 1 0 5152 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_38
timestamp 1698431365
transform 1 0 5600 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_48
timestamp 1698431365
transform 1 0 6720 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_56
timestamp 1698431365
transform 1 0 7616 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_60
timestamp 1698431365
transform 1 0 8064 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_83
timestamp 1698431365
transform 1 0 10640 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_114
timestamp 1698431365
transform 1 0 14112 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_122
timestamp 1698431365
transform 1 0 15008 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_129
timestamp 1698431365
transform 1 0 15792 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_137
timestamp 1698431365
transform 1 0 16688 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_139
timestamp 1698431365
transform 1 0 16912 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_142
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_152
timestamp 1698431365
transform 1 0 18368 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_184
timestamp 1698431365
transform 1 0 21952 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_186
timestamp 1698431365
transform 1 0 22176 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_208
timestamp 1698431365
transform 1 0 24640 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_212
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_220
timestamp 1698431365
transform 1 0 25984 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_243
timestamp 1698431365
transform 1 0 28560 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_251
timestamp 1698431365
transform 1 0 29456 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_255
timestamp 1698431365
transform 1 0 29904 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_270
timestamp 1698431365
transform 1 0 31584 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_274
timestamp 1698431365
transform 1 0 32032 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_282
timestamp 1698431365
transform 1 0 32928 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_286
timestamp 1698431365
transform 1 0 33376 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_288
timestamp 1698431365
transform 1 0 33600 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_348
timestamp 1698431365
transform 1 0 40320 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_367
timestamp 1698431365
transform 1 0 42448 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_369
timestamp 1698431365
transform 1 0 42672 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_399
timestamp 1698431365
transform 1 0 46032 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_403
timestamp 1698431365
transform 1 0 46480 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_405
timestamp 1698431365
transform 1 0 46704 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_432
timestamp 1698431365
transform 1 0 49728 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_469
timestamp 1698431365
transform 1 0 53872 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_471
timestamp 1698431365
transform 1 0 54096 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_485
timestamp 1698431365
transform 1 0 55664 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_489
timestamp 1698431365
transform 1 0 56112 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_492
timestamp 1698431365
transform 1 0 56448 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_508
timestamp 1698431365
transform 1 0 58240 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_16
timestamp 1698431365
transform 1 0 3136 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_20
timestamp 1698431365
transform 1 0 3584 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_24
timestamp 1698431365
transform 1 0 4032 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_30
timestamp 1698431365
transform 1 0 4704 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698431365
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_41
timestamp 1698431365
transform 1 0 5936 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_43
timestamp 1698431365
transform 1 0 6160 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_54
timestamp 1698431365
transform 1 0 7392 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_107
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_115
timestamp 1698431365
transform 1 0 14224 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_119
timestamp 1698431365
transform 1 0 14672 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_121
timestamp 1698431365
transform 1 0 14896 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_130
timestamp 1698431365
transform 1 0 15904 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_154
timestamp 1698431365
transform 1 0 18592 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_156
timestamp 1698431365
transform 1 0 18816 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_169
timestamp 1698431365
transform 1 0 20272 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_173
timestamp 1698431365
transform 1 0 20720 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_183
timestamp 1698431365
transform 1 0 21840 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_202
timestamp 1698431365
transform 1 0 23968 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_234
timestamp 1698431365
transform 1 0 27552 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_238
timestamp 1698431365
transform 1 0 28000 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_247
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_249
timestamp 1698431365
transform 1 0 29232 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_270
timestamp 1698431365
transform 1 0 31584 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_274
timestamp 1698431365
transform 1 0 32032 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_276
timestamp 1698431365
transform 1 0 32256 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_293
timestamp 1698431365
transform 1 0 34160 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_309
timestamp 1698431365
transform 1 0 35952 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_340
timestamp 1698431365
transform 1 0 39424 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_401
timestamp 1698431365
transform 1 0 46256 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_452
timestamp 1698431365
transform 1 0 51968 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_454
timestamp 1698431365
transform 1 0 52192 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_494
timestamp 1698431365
transform 1 0 56672 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_502
timestamp 1698431365
transform 1 0 57568 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_506
timestamp 1698431365
transform 1 0 58016 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_508
timestamp 1698431365
transform 1 0 58240 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_28
timestamp 1698431365
transform 1 0 4480 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_30
timestamp 1698431365
transform 1 0 4704 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_68
timestamp 1698431365
transform 1 0 8960 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_72
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_89
timestamp 1698431365
transform 1 0 11312 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_95
timestamp 1698431365
transform 1 0 11984 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_103
timestamp 1698431365
transform 1 0 12880 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_105
timestamp 1698431365
transform 1 0 13104 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_113
timestamp 1698431365
transform 1 0 14000 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_142
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_150
timestamp 1698431365
transform 1 0 18144 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_177
timestamp 1698431365
transform 1 0 21168 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_212
timestamp 1698431365
transform 1 0 25088 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_239
timestamp 1698431365
transform 1 0 28112 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_275
timestamp 1698431365
transform 1 0 32144 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_279
timestamp 1698431365
transform 1 0 32592 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_282
timestamp 1698431365
transform 1 0 32928 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_284
timestamp 1698431365
transform 1 0 33152 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_302
timestamp 1698431365
transform 1 0 35168 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_304
timestamp 1698431365
transform 1 0 35392 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_347
timestamp 1698431365
transform 1 0 40208 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_349
timestamp 1698431365
transform 1 0 40432 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_419
timestamp 1698431365
transform 1 0 48272 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_489
timestamp 1698431365
transform 1 0 56112 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_499
timestamp 1698431365
transform 1 0 57232 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_507
timestamp 1698431365
transform 1 0 58128 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_8
timestamp 1698431365
transform 1 0 2240 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_45
timestamp 1698431365
transform 1 0 6384 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_57
timestamp 1698431365
transform 1 0 7728 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_70
timestamp 1698431365
transform 1 0 9184 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_78
timestamp 1698431365
transform 1 0 10080 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_94
timestamp 1698431365
transform 1 0 11872 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_102
timestamp 1698431365
transform 1 0 12768 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_104
timestamp 1698431365
transform 1 0 12992 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_107
timestamp 1698431365
transform 1 0 13328 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_119
timestamp 1698431365
transform 1 0 14672 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_123
timestamp 1698431365
transform 1 0 15120 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_172
timestamp 1698431365
transform 1 0 20608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1698431365
transform 1 0 20832 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_206
timestamp 1698431365
transform 1 0 24416 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_210
timestamp 1698431365
transform 1 0 24864 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_241
timestamp 1698431365
transform 1 0 28336 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_247
timestamp 1698431365
transform 1 0 29008 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_251
timestamp 1698431365
transform 1 0 29456 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_261
timestamp 1698431365
transform 1 0 30576 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_277
timestamp 1698431365
transform 1 0 32368 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_281
timestamp 1698431365
transform 1 0 32816 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_288
timestamp 1698431365
transform 1 0 33600 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_290
timestamp 1698431365
transform 1 0 33824 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_297
timestamp 1698431365
transform 1 0 34608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_312
timestamp 1698431365
transform 1 0 36288 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_314
timestamp 1698431365
transform 1 0 36512 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_329
timestamp 1698431365
transform 1 0 38192 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_364
timestamp 1698431365
transform 1 0 42112 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_372
timestamp 1698431365
transform 1 0 43008 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_396
timestamp 1698431365
transform 1 0 45696 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_400
timestamp 1698431365
transform 1 0 46144 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_431
timestamp 1698431365
transform 1 0 49616 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_437
timestamp 1698431365
transform 1 0 50288 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_439
timestamp 1698431365
transform 1 0 50512 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_450
timestamp 1698431365
transform 1 0 51744 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_454
timestamp 1698431365
transform 1 0 52192 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_457
timestamp 1698431365
transform 1 0 52528 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_461
timestamp 1698431365
transform 1 0 52976 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_470
timestamp 1698431365
transform 1 0 53984 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_508
timestamp 1698431365
transform 1 0 58240 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_42
timestamp 1698431365
transform 1 0 6048 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_46
timestamp 1698431365
transform 1 0 6496 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_50
timestamp 1698431365
transform 1 0 6944 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_52
timestamp 1698431365
transform 1 0 7168 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_62
timestamp 1698431365
transform 1 0 8288 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_72
timestamp 1698431365
transform 1 0 9408 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_88
timestamp 1698431365
transform 1 0 11200 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_134
timestamp 1698431365
transform 1 0 16352 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_138
timestamp 1698431365
transform 1 0 16800 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_166
timestamp 1698431365
transform 1 0 19936 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_174
timestamp 1698431365
transform 1 0 20832 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_177
timestamp 1698431365
transform 1 0 21168 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_207
timestamp 1698431365
transform 1 0 24528 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1698431365
transform 1 0 24752 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_235
timestamp 1698431365
transform 1 0 27664 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_247
timestamp 1698431365
transform 1 0 29008 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_256
timestamp 1698431365
transform 1 0 30016 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_260
timestamp 1698431365
transform 1 0 30464 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_274
timestamp 1698431365
transform 1 0 32032 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_278
timestamp 1698431365
transform 1 0 32480 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_282
timestamp 1698431365
transform 1 0 32928 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_290
timestamp 1698431365
transform 1 0 33824 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_294
timestamp 1698431365
transform 1 0 34272 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_313
timestamp 1698431365
transform 1 0 36400 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_317
timestamp 1698431365
transform 1 0 36848 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_319
timestamp 1698431365
transform 1 0 37072 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_326
timestamp 1698431365
transform 1 0 37856 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_328
timestamp 1698431365
transform 1 0 38080 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_346
timestamp 1698431365
transform 1 0 40096 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_352
timestamp 1698431365
transform 1 0 40768 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_382
timestamp 1698431365
transform 1 0 44128 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_390
timestamp 1698431365
transform 1 0 45024 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_394
timestamp 1698431365
transform 1 0 45472 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_396
timestamp 1698431365
transform 1 0 45696 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_422
timestamp 1698431365
transform 1 0 48608 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_438
timestamp 1698431365
transform 1 0 50400 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_469
timestamp 1698431365
transform 1 0 53872 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_473
timestamp 1698431365
transform 1 0 54320 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_492
timestamp 1698431365
transform 1 0 56448 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_506
timestamp 1698431365
transform 1 0 58016 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_508
timestamp 1698431365
transform 1 0 58240 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_20
timestamp 1698431365
transform 1 0 3584 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_33
timestamp 1698431365
transform 1 0 5040 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_37
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_41
timestamp 1698431365
transform 1 0 5936 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_43
timestamp 1698431365
transform 1 0 6160 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_75
timestamp 1698431365
transform 1 0 9744 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_102
timestamp 1698431365
transform 1 0 12768 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_104
timestamp 1698431365
transform 1 0 12992 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_120
timestamp 1698431365
transform 1 0 14784 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_135
timestamp 1698431365
transform 1 0 16464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_137
timestamp 1698431365
transform 1 0 16688 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_147
timestamp 1698431365
transform 1 0 17808 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_149
timestamp 1698431365
transform 1 0 18032 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_182
timestamp 1698431365
transform 1 0 21728 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_232
timestamp 1698431365
transform 1 0 27328 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_240
timestamp 1698431365
transform 1 0 28224 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_244
timestamp 1698431365
transform 1 0 28672 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_275
timestamp 1698431365
transform 1 0 32144 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_311
timestamp 1698431365
transform 1 0 36176 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_317
timestamp 1698431365
transform 1 0 36848 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_325
timestamp 1698431365
transform 1 0 37744 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_329
timestamp 1698431365
transform 1 0 38192 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_382
timestamp 1698431365
transform 1 0 44128 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_384
timestamp 1698431365
transform 1 0 44352 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_387
timestamp 1698431365
transform 1 0 44688 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_389
timestamp 1698431365
transform 1 0 44912 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_413
timestamp 1698431365
transform 1 0 47600 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_417
timestamp 1698431365
transform 1 0 48048 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_446
timestamp 1698431365
transform 1 0 51296 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_454
timestamp 1698431365
transform 1 0 52192 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_457
timestamp 1698431365
transform 1 0 52528 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_473
timestamp 1698431365
transform 1 0 54320 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_481
timestamp 1698431365
transform 1 0 55216 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_506
timestamp 1698431365
transform 1 0 58016 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_508
timestamp 1698431365
transform 1 0 58240 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_72
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_76
timestamp 1698431365
transform 1 0 9856 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_125
timestamp 1698431365
transform 1 0 15344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_142
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_144
timestamp 1698431365
transform 1 0 17472 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_204
timestamp 1698431365
transform 1 0 24192 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_230
timestamp 1698431365
transform 1 0 27104 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_237
timestamp 1698431365
transform 1 0 27888 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_239
timestamp 1698431365
transform 1 0 28112 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_247
timestamp 1698431365
transform 1 0 29008 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_255
timestamp 1698431365
transform 1 0 29904 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_257
timestamp 1698431365
transform 1 0 30128 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_279
timestamp 1698431365
transform 1 0 32592 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_282
timestamp 1698431365
transform 1 0 32928 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_286
timestamp 1698431365
transform 1 0 33376 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_294
timestamp 1698431365
transform 1 0 34272 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_298
timestamp 1698431365
transform 1 0 34720 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_311
timestamp 1698431365
transform 1 0 36176 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_315
timestamp 1698431365
transform 1 0 36624 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_339
timestamp 1698431365
transform 1 0 39312 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_482
timestamp 1698431365
transform 1 0 55328 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_504
timestamp 1698431365
transform 1 0 57792 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_508
timestamp 1698431365
transform 1 0 58240 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698431365
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_37
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_51
timestamp 1698431365
transform 1 0 7056 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_102
timestamp 1698431365
transform 1 0 12768 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_104
timestamp 1698431365
transform 1 0 12992 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_142
timestamp 1698431365
transform 1 0 17248 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_201
timestamp 1698431365
transform 1 0 23856 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_223
timestamp 1698431365
transform 1 0 26320 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_230
timestamp 1698431365
transform 1 0 27104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_232
timestamp 1698431365
transform 1 0 27328 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_241
timestamp 1698431365
transform 1 0 28336 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_260
timestamp 1698431365
transform 1 0 30464 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_285
timestamp 1698431365
transform 1 0 33264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_289
timestamp 1698431365
transform 1 0 33712 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_305
timestamp 1698431365
transform 1 0 35504 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_313
timestamp 1698431365
transform 1 0 36400 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_347
timestamp 1698431365
transform 1 0 40208 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_351
timestamp 1698431365
transform 1 0 40656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_355
timestamp 1698431365
transform 1 0 41104 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_359
timestamp 1698431365
transform 1 0 41552 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_395
timestamp 1698431365
transform 1 0 45584 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_399
timestamp 1698431365
transform 1 0 46032 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_414
timestamp 1698431365
transform 1 0 47712 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_418
timestamp 1698431365
transform 1 0 48160 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_424
timestamp 1698431365
transform 1 0 48832 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_434
timestamp 1698431365
transform 1 0 49952 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_447
timestamp 1698431365
transform 1 0 51408 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_457
timestamp 1698431365
transform 1 0 52528 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_459
timestamp 1698431365
transform 1 0 52752 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_482
timestamp 1698431365
transform 1 0 55328 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_508
timestamp 1698431365
transform 1 0 58240 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_2
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_4
timestamp 1698431365
transform 1 0 1792 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_57
timestamp 1698431365
transform 1 0 7728 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_65
timestamp 1698431365
transform 1 0 8624 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_69
timestamp 1698431365
transform 1 0 9072 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_139
timestamp 1698431365
transform 1 0 16912 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_155
timestamp 1698431365
transform 1 0 18704 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_165
timestamp 1698431365
transform 1 0 19824 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_196
timestamp 1698431365
transform 1 0 23296 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_200
timestamp 1698431365
transform 1 0 23744 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_209
timestamp 1698431365
transform 1 0 24752 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_218
timestamp 1698431365
transform 1 0 25760 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_226
timestamp 1698431365
transform 1 0 26656 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_230
timestamp 1698431365
transform 1 0 27104 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_247
timestamp 1698431365
transform 1 0 29008 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_249
timestamp 1698431365
transform 1 0 29232 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_273
timestamp 1698431365
transform 1 0 31920 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_277
timestamp 1698431365
transform 1 0 32368 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_292
timestamp 1698431365
transform 1 0 34048 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_323
timestamp 1698431365
transform 1 0 37520 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_327
timestamp 1698431365
transform 1 0 37968 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_343
timestamp 1698431365
transform 1 0 39760 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_345
timestamp 1698431365
transform 1 0 39984 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_364
timestamp 1698431365
transform 1 0 42112 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_385
timestamp 1698431365
transform 1 0 44464 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_417
timestamp 1698431365
transform 1 0 48048 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_419
timestamp 1698431365
transform 1 0 48272 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_430
timestamp 1698431365
transform 1 0 49504 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_438
timestamp 1698431365
transform 1 0 50400 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_450
timestamp 1698431365
transform 1 0 51744 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_458
timestamp 1698431365
transform 1 0 52640 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_480
timestamp 1698431365
transform 1 0 55104 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_488
timestamp 1698431365
transform 1 0 56000 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_497
timestamp 1698431365
transform 1 0 57008 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_505
timestamp 1698431365
transform 1 0 57904 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_8
timestamp 1698431365
transform 1 0 2240 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698431365
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_47
timestamp 1698431365
transform 1 0 6608 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_59
timestamp 1698431365
transform 1 0 7952 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_90
timestamp 1698431365
transform 1 0 11424 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_97
timestamp 1698431365
transform 1 0 12208 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_107
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_111
timestamp 1698431365
transform 1 0 13776 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_119
timestamp 1698431365
transform 1 0 14672 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_123
timestamp 1698431365
transform 1 0 15120 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_127
timestamp 1698431365
transform 1 0 15568 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_129
timestamp 1698431365
transform 1 0 15792 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_189
timestamp 1698431365
transform 1 0 22512 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_191
timestamp 1698431365
transform 1 0 22736 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_194
timestamp 1698431365
transform 1 0 23072 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_222
timestamp 1698431365
transform 1 0 26208 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_226
timestamp 1698431365
transform 1 0 26656 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_240
timestamp 1698431365
transform 1 0 28224 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_244
timestamp 1698431365
transform 1 0 28672 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_247
timestamp 1698431365
transform 1 0 29008 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_314
timestamp 1698431365
transform 1 0 36512 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_317
timestamp 1698431365
transform 1 0 36848 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_321
timestamp 1698431365
transform 1 0 37296 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_329
timestamp 1698431365
transform 1 0 38192 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_333
timestamp 1698431365
transform 1 0 38640 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_335
timestamp 1698431365
transform 1 0 38864 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_359
timestamp 1698431365
transform 1 0 41552 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_382
timestamp 1698431365
transform 1 0 44128 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_384
timestamp 1698431365
transform 1 0 44352 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_387
timestamp 1698431365
transform 1 0 44688 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_395
timestamp 1698431365
transform 1 0 45584 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_402
timestamp 1698431365
transform 1 0 46368 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_412
timestamp 1698431365
transform 1 0 47488 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_416
timestamp 1698431365
transform 1 0 47936 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_418
timestamp 1698431365
transform 1 0 48160 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_433
timestamp 1698431365
transform 1 0 49840 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_451
timestamp 1698431365
transform 1 0 51856 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_457
timestamp 1698431365
transform 1 0 52528 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_473
timestamp 1698431365
transform 1 0 54320 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_481
timestamp 1698431365
transform 1 0 55216 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_483
timestamp 1698431365
transform 1 0 55440 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_501
timestamp 1698431365
transform 1 0 57456 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_2
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_6
timestamp 1698431365
transform 1 0 2016 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_56
timestamp 1698431365
transform 1 0 7616 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_58
timestamp 1698431365
transform 1 0 7840 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_98
timestamp 1698431365
transform 1 0 12320 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_102
timestamp 1698431365
transform 1 0 12768 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_110
timestamp 1698431365
transform 1 0 13664 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_134
timestamp 1698431365
transform 1 0 16352 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_138
timestamp 1698431365
transform 1 0 16800 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_208
timestamp 1698431365
transform 1 0 24640 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_212
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_246
timestamp 1698431365
transform 1 0 28896 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_279
timestamp 1698431365
transform 1 0 32592 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_282
timestamp 1698431365
transform 1 0 32928 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_286
timestamp 1698431365
transform 1 0 33376 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_296
timestamp 1698431365
transform 1 0 34496 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_311
timestamp 1698431365
transform 1 0 36176 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_315
timestamp 1698431365
transform 1 0 36624 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_323
timestamp 1698431365
transform 1 0 37520 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_327
timestamp 1698431365
transform 1 0 37968 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_349
timestamp 1698431365
transform 1 0 40432 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_365
timestamp 1698431365
transform 1 0 42224 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_369
timestamp 1698431365
transform 1 0 42672 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_373
timestamp 1698431365
transform 1 0 43120 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_418
timestamp 1698431365
transform 1 0 48160 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_422
timestamp 1698431365
transform 1 0 48608 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_426
timestamp 1698431365
transform 1 0 49056 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_434
timestamp 1698431365
transform 1 0 49952 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_438
timestamp 1698431365
transform 1 0 50400 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_447
timestamp 1698431365
transform 1 0 51408 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_449
timestamp 1698431365
transform 1 0 51632 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_458
timestamp 1698431365
transform 1 0 52640 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_467
timestamp 1698431365
transform 1 0 53648 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_471
timestamp 1698431365
transform 1 0 54096 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_474
timestamp 1698431365
transform 1 0 54432 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_481
timestamp 1698431365
transform 1 0 55216 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_489
timestamp 1698431365
transform 1 0 56112 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_505
timestamp 1698431365
transform 1 0 57904 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_2
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_37
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_70
timestamp 1698431365
transform 1 0 9184 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_74
timestamp 1698431365
transform 1 0 9632 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_115
timestamp 1698431365
transform 1 0 14224 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_131
timestamp 1698431365
transform 1 0 16016 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_139
timestamp 1698431365
transform 1 0 16912 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_172
timestamp 1698431365
transform 1 0 20608 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_174
timestamp 1698431365
transform 1 0 20832 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_177
timestamp 1698431365
transform 1 0 21168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_192
timestamp 1698431365
transform 1 0 22848 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_202
timestamp 1698431365
transform 1 0 23968 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_210
timestamp 1698431365
transform 1 0 24864 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_214
timestamp 1698431365
transform 1 0 25312 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_218
timestamp 1698431365
transform 1 0 25760 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_227
timestamp 1698431365
transform 1 0 26768 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_247
timestamp 1698431365
transform 1 0 29008 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_251
timestamp 1698431365
transform 1 0 29456 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_259
timestamp 1698431365
transform 1 0 30352 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_276
timestamp 1698431365
transform 1 0 32256 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_284
timestamp 1698431365
transform 1 0 33152 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_304
timestamp 1698431365
transform 1 0 35392 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_330
timestamp 1698431365
transform 1 0 38304 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_338
timestamp 1698431365
transform 1 0 39200 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_358
timestamp 1698431365
transform 1 0 41440 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_395
timestamp 1698431365
transform 1 0 45584 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_402
timestamp 1698431365
transform 1 0 46368 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_418
timestamp 1698431365
transform 1 0 48160 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_426
timestamp 1698431365
transform 1 0 49056 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_430
timestamp 1698431365
transform 1 0 49504 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_432
timestamp 1698431365
transform 1 0 49728 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_441
timestamp 1698431365
transform 1 0 50736 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_476
timestamp 1698431365
transform 1 0 54656 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_508
timestamp 1698431365
transform 1 0 58240 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_2
timestamp 1698431365
transform 1 0 1568 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_6
timestamp 1698431365
transform 1 0 2016 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_69
timestamp 1698431365
transform 1 0 9072 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_85
timestamp 1698431365
transform 1 0 10864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_87
timestamp 1698431365
transform 1 0 11088 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_94
timestamp 1698431365
transform 1 0 11872 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_124
timestamp 1698431365
transform 1 0 15232 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_139
timestamp 1698431365
transform 1 0 16912 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_142
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_152
timestamp 1698431365
transform 1 0 18368 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_156
timestamp 1698431365
transform 1 0 18816 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_164
timestamp 1698431365
transform 1 0 19712 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_166
timestamp 1698431365
transform 1 0 19936 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_180
timestamp 1698431365
transform 1 0 21504 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_205
timestamp 1698431365
transform 1 0 24304 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698431365
transform 1 0 24752 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_212
timestamp 1698431365
transform 1 0 25088 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_228
timestamp 1698431365
transform 1 0 26880 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_230
timestamp 1698431365
transform 1 0 27104 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_239
timestamp 1698431365
transform 1 0 28112 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_247
timestamp 1698431365
transform 1 0 29008 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_251
timestamp 1698431365
transform 1 0 29456 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_257
timestamp 1698431365
transform 1 0 30128 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_266
timestamp 1698431365
transform 1 0 31136 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_274
timestamp 1698431365
transform 1 0 32032 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_278
timestamp 1698431365
transform 1 0 32480 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_282
timestamp 1698431365
transform 1 0 32928 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_290
timestamp 1698431365
transform 1 0 33824 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_299
timestamp 1698431365
transform 1 0 34832 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_330
timestamp 1698431365
transform 1 0 38304 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_334
timestamp 1698431365
transform 1 0 38752 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_342
timestamp 1698431365
transform 1 0 39648 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_344
timestamp 1698431365
transform 1 0 39872 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_361
timestamp 1698431365
transform 1 0 41776 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_365
timestamp 1698431365
transform 1 0 42224 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_385
timestamp 1698431365
transform 1 0 44464 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_422
timestamp 1698431365
transform 1 0 48608 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_430
timestamp 1698431365
transform 1 0 49504 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_447
timestamp 1698431365
transform 1 0 51408 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_505
timestamp 1698431365
transform 1 0 57904 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_2
timestamp 1698431365
transform 1 0 1568 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_31
timestamp 1698431365
transform 1 0 4816 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_37
timestamp 1698431365
transform 1 0 5488 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_72
timestamp 1698431365
transform 1 0 9408 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_107
timestamp 1698431365
transform 1 0 13328 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_119
timestamp 1698431365
transform 1 0 14672 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_143
timestamp 1698431365
transform 1 0 17360 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_145
timestamp 1698431365
transform 1 0 17584 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_157
timestamp 1698431365
transform 1 0 18928 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_159
timestamp 1698431365
transform 1 0 19152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_177
timestamp 1698431365
transform 1 0 21168 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_185
timestamp 1698431365
transform 1 0 22064 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_187
timestamp 1698431365
transform 1 0 22288 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_199
timestamp 1698431365
transform 1 0 23632 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_209
timestamp 1698431365
transform 1 0 24752 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_213
timestamp 1698431365
transform 1 0 25200 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_243
timestamp 1698431365
transform 1 0 28560 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_247
timestamp 1698431365
transform 1 0 29008 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_273
timestamp 1698431365
transform 1 0 31920 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_281
timestamp 1698431365
transform 1 0 32816 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_287
timestamp 1698431365
transform 1 0 33488 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_291
timestamp 1698431365
transform 1 0 33936 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_293
timestamp 1698431365
transform 1 0 34160 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_300
timestamp 1698431365
transform 1 0 34944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_304
timestamp 1698431365
transform 1 0 35392 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_306
timestamp 1698431365
transform 1 0 35616 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_312
timestamp 1698431365
transform 1 0 36288 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_314
timestamp 1698431365
transform 1 0 36512 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_327
timestamp 1698431365
transform 1 0 37968 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_331
timestamp 1698431365
transform 1 0 38416 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_335
timestamp 1698431365
transform 1 0 38864 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_337
timestamp 1698431365
transform 1 0 39088 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_350
timestamp 1698431365
transform 1 0 40544 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_352
timestamp 1698431365
transform 1 0 40768 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_365
timestamp 1698431365
transform 1 0 42224 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_373
timestamp 1698431365
transform 1 0 43120 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_377
timestamp 1698431365
transform 1 0 43568 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_384
timestamp 1698431365
transform 1 0 44352 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_387
timestamp 1698431365
transform 1 0 44688 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_391
timestamp 1698431365
transform 1 0 45136 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_395
timestamp 1698431365
transform 1 0 45584 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_408
timestamp 1698431365
transform 1 0 47040 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_416
timestamp 1698431365
transform 1 0 47936 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_418
timestamp 1698431365
transform 1 0 48160 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_449
timestamp 1698431365
transform 1 0 51632 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_457
timestamp 1698431365
transform 1 0 52528 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_459
timestamp 1698431365
transform 1 0 52752 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_2
timestamp 1698431365
transform 1 0 1568 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_23
timestamp 1698431365
transform 1 0 3920 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_37
timestamp 1698431365
transform 1 0 5488 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_53
timestamp 1698431365
transform 1 0 7280 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_55
timestamp 1698431365
transform 1 0 7504 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_170
timestamp 1698431365
transform 1 0 20384 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_184
timestamp 1698431365
transform 1 0 21952 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_188
timestamp 1698431365
transform 1 0 22400 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_196
timestamp 1698431365
transform 1 0 23296 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_198
timestamp 1698431365
transform 1 0 23520 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_201
timestamp 1698431365
transform 1 0 23856 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_205
timestamp 1698431365
transform 1 0 24304 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_209
timestamp 1698431365
transform 1 0 24752 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_212
timestamp 1698431365
transform 1 0 25088 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_220
timestamp 1698431365
transform 1 0 25984 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_222
timestamp 1698431365
transform 1 0 26208 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_225
timestamp 1698431365
transform 1 0 26544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_232
timestamp 1698431365
transform 1 0 27328 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_239
timestamp 1698431365
transform 1 0 28112 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_243
timestamp 1698431365
transform 1 0 28560 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_251
timestamp 1698431365
transform 1 0 29456 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_265
timestamp 1698431365
transform 1 0 31024 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_273
timestamp 1698431365
transform 1 0 31920 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_276
timestamp 1698431365
transform 1 0 32256 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_289
timestamp 1698431365
transform 1 0 33712 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_340
timestamp 1698431365
transform 1 0 39424 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_347
timestamp 1698431365
transform 1 0 40208 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_349
timestamp 1698431365
transform 1 0 40432 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_371
timestamp 1698431365
transform 1 0 42896 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_375
timestamp 1698431365
transform 1 0 43344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_377
timestamp 1698431365
transform 1 0 43568 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_397
timestamp 1698431365
transform 1 0 45808 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_401
timestamp 1698431365
transform 1 0 46256 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_417
timestamp 1698431365
transform 1 0 48048 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_419
timestamp 1698431365
transform 1 0 48272 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_422
timestamp 1698431365
transform 1 0 48608 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_424
timestamp 1698431365
transform 1 0 48832 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_441
timestamp 1698431365
transform 1 0 50736 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_449
timestamp 1698431365
transform 1 0 51632 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_451
timestamp 1698431365
transform 1 0 51856 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_505
timestamp 1698431365
transform 1 0 57904 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_28
timestamp 1698431365
transform 1 0 4480 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_43
timestamp 1698431365
transform 1 0 6160 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_59
timestamp 1698431365
transform 1 0 7952 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_87
timestamp 1698431365
transform 1 0 11088 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_103
timestamp 1698431365
transform 1 0 12880 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_107
timestamp 1698431365
transform 1 0 13328 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_126
timestamp 1698431365
transform 1 0 15456 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_160
timestamp 1698431365
transform 1 0 19264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_169
timestamp 1698431365
transform 1 0 20272 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_173
timestamp 1698431365
transform 1 0 20720 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_177
timestamp 1698431365
transform 1 0 21168 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_185
timestamp 1698431365
transform 1 0 22064 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_189
timestamp 1698431365
transform 1 0 22512 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_231
timestamp 1698431365
transform 1 0 27216 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_241
timestamp 1698431365
transform 1 0 28336 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_288
timestamp 1698431365
transform 1 0 33600 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_290
timestamp 1698431365
transform 1 0 33824 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_314
timestamp 1698431365
transform 1 0 36512 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_317
timestamp 1698431365
transform 1 0 36848 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_319
timestamp 1698431365
transform 1 0 37072 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_325
timestamp 1698431365
transform 1 0 37744 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_329
timestamp 1698431365
transform 1 0 38192 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_333
timestamp 1698431365
transform 1 0 38640 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_337
timestamp 1698431365
transform 1 0 39088 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_339
timestamp 1698431365
transform 1 0 39312 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_342
timestamp 1698431365
transform 1 0 39648 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_362
timestamp 1698431365
transform 1 0 41888 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_366
timestamp 1698431365
transform 1 0 42336 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_382
timestamp 1698431365
transform 1 0 44128 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_384
timestamp 1698431365
transform 1 0 44352 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_418
timestamp 1698431365
transform 1 0 48160 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_426
timestamp 1698431365
transform 1 0 49056 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_428
timestamp 1698431365
transform 1 0 49280 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_442
timestamp 1698431365
transform 1 0 50848 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_450
timestamp 1698431365
transform 1 0 51744 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_452
timestamp 1698431365
transform 1 0 51968 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_462
timestamp 1698431365
transform 1 0 53088 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_464
timestamp 1698431365
transform 1 0 53312 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_20
timestamp 1698431365
transform 1 0 3584 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_24
timestamp 1698431365
transform 1 0 4032 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_28
timestamp 1698431365
transform 1 0 4480 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_38
timestamp 1698431365
transform 1 0 5600 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_63
timestamp 1698431365
transform 1 0 8400 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_67
timestamp 1698431365
transform 1 0 8848 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_69
timestamp 1698431365
transform 1 0 9072 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_80
timestamp 1698431365
transform 1 0 10304 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_93
timestamp 1698431365
transform 1 0 11760 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_123
timestamp 1698431365
transform 1 0 15120 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_127
timestamp 1698431365
transform 1 0 15568 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_131
timestamp 1698431365
transform 1 0 16016 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_133
timestamp 1698431365
transform 1 0 16240 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_138
timestamp 1698431365
transform 1 0 16800 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_142
timestamp 1698431365
transform 1 0 17248 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_155
timestamp 1698431365
transform 1 0 18704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_159
timestamp 1698431365
transform 1 0 19152 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_163
timestamp 1698431365
transform 1 0 19600 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_202
timestamp 1698431365
transform 1 0 23968 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_206
timestamp 1698431365
transform 1 0 24416 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_237
timestamp 1698431365
transform 1 0 27888 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_241
timestamp 1698431365
transform 1 0 28336 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_247
timestamp 1698431365
transform 1 0 29008 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_282
timestamp 1698431365
transform 1 0 32928 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_294
timestamp 1698431365
transform 1 0 34272 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_298
timestamp 1698431365
transform 1 0 34720 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_349
timestamp 1698431365
transform 1 0 40432 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_352
timestamp 1698431365
transform 1 0 40768 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_356
timestamp 1698431365
transform 1 0 41216 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_358
timestamp 1698431365
transform 1 0 41440 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_364
timestamp 1698431365
transform 1 0 42112 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_368
timestamp 1698431365
transform 1 0 42560 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_401
timestamp 1698431365
transform 1 0 46256 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_409
timestamp 1698431365
transform 1 0 47152 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_416
timestamp 1698431365
transform 1 0 47936 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_440
timestamp 1698431365
transform 1 0 50624 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_448
timestamp 1698431365
transform 1 0 51520 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_465
timestamp 1698431365
transform 1 0 53424 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_467
timestamp 1698431365
transform 1 0 53648 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_498
timestamp 1698431365
transform 1 0 57120 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_502
timestamp 1698431365
transform 1 0 57568 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_14
timestamp 1698431365
transform 1 0 2912 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_18
timestamp 1698431365
transform 1 0 3360 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_22
timestamp 1698431365
transform 1 0 3808 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_30
timestamp 1698431365
transform 1 0 4704 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698431365
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_37
timestamp 1698431365
transform 1 0 5488 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_41
timestamp 1698431365
transform 1 0 5936 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_70
timestamp 1698431365
transform 1 0 9184 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_102
timestamp 1698431365
transform 1 0 12768 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_104
timestamp 1698431365
transform 1 0 12992 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_107
timestamp 1698431365
transform 1 0 13328 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_115
timestamp 1698431365
transform 1 0 14224 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_119
timestamp 1698431365
transform 1 0 14672 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_121
timestamp 1698431365
transform 1 0 14896 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_151
timestamp 1698431365
transform 1 0 18256 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_153
timestamp 1698431365
transform 1 0 18480 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_164
timestamp 1698431365
transform 1 0 19712 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_168
timestamp 1698431365
transform 1 0 20160 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_172
timestamp 1698431365
transform 1 0 20608 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_174
timestamp 1698431365
transform 1 0 20832 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_187
timestamp 1698431365
transform 1 0 22288 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_228
timestamp 1698431365
transform 1 0 26880 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_232
timestamp 1698431365
transform 1 0 27328 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_241
timestamp 1698431365
transform 1 0 28336 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_255
timestamp 1698431365
transform 1 0 29904 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_257
timestamp 1698431365
transform 1 0 30128 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_266
timestamp 1698431365
transform 1 0 31136 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_268
timestamp 1698431365
transform 1 0 31360 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_271
timestamp 1698431365
transform 1 0 31696 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_287
timestamp 1698431365
transform 1 0 33488 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_289
timestamp 1698431365
transform 1 0 33712 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_313
timestamp 1698431365
transform 1 0 36400 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_375
timestamp 1698431365
transform 1 0 43344 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_383
timestamp 1698431365
transform 1 0 44240 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_387
timestamp 1698431365
transform 1 0 44688 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_391
timestamp 1698431365
transform 1 0 45136 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_406
timestamp 1698431365
transform 1 0 46816 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_438
timestamp 1698431365
transform 1 0 50400 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_469
timestamp 1698431365
transform 1 0 53872 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_471
timestamp 1698431365
transform 1 0 54096 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_480
timestamp 1698431365
transform 1 0 55104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_482
timestamp 1698431365
transform 1 0 55328 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_14
timestamp 1698431365
transform 1 0 2912 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_18
timestamp 1698431365
transform 1 0 3360 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_22
timestamp 1698431365
transform 1 0 3808 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_54
timestamp 1698431365
transform 1 0 7392 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_72
timestamp 1698431365
transform 1 0 9408 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_104
timestamp 1698431365
transform 1 0 12992 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_120
timestamp 1698431365
transform 1 0 14784 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_128
timestamp 1698431365
transform 1 0 15680 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_138
timestamp 1698431365
transform 1 0 16800 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_142
timestamp 1698431365
transform 1 0 17248 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_144
timestamp 1698431365
transform 1 0 17472 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_147
timestamp 1698431365
transform 1 0 17808 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_192
timestamp 1698431365
transform 1 0 22848 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_194
timestamp 1698431365
transform 1 0 23072 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_206
timestamp 1698431365
transform 1 0 24416 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_212
timestamp 1698431365
transform 1 0 25088 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_248
timestamp 1698431365
transform 1 0 29120 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_271
timestamp 1698431365
transform 1 0 31696 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_275
timestamp 1698431365
transform 1 0 32144 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_277
timestamp 1698431365
transform 1 0 32368 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_282
timestamp 1698431365
transform 1 0 32928 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_313
timestamp 1698431365
transform 1 0 36400 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_317
timestamp 1698431365
transform 1 0 36848 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_326
timestamp 1698431365
transform 1 0 37856 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_328
timestamp 1698431365
transform 1 0 38080 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_381
timestamp 1698431365
transform 1 0 44016 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_383
timestamp 1698431365
transform 1 0 44240 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_434
timestamp 1698431365
transform 1 0 49952 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_438
timestamp 1698431365
transform 1 0 50400 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_440
timestamp 1698431365
transform 1 0 50624 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_469
timestamp 1698431365
transform 1 0 53872 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_485
timestamp 1698431365
transform 1 0 55664 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_489
timestamp 1698431365
transform 1 0 56112 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_492
timestamp 1698431365
transform 1 0 56448 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_500
timestamp 1698431365
transform 1 0 57344 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_503
timestamp 1698431365
transform 1 0 57680 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_507
timestamp 1698431365
transform 1 0 58128 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_2
timestamp 1698431365
transform 1 0 1568 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_20
timestamp 1698431365
transform 1 0 3584 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_28
timestamp 1698431365
transform 1 0 4480 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_32
timestamp 1698431365
transform 1 0 4928 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698431365
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_43
timestamp 1698431365
transform 1 0 6160 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_75
timestamp 1698431365
transform 1 0 9744 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_91
timestamp 1698431365
transform 1 0 11536 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_99
timestamp 1698431365
transform 1 0 12432 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_103
timestamp 1698431365
transform 1 0 12880 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_136
timestamp 1698431365
transform 1 0 16576 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_153
timestamp 1698431365
transform 1 0 18480 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_165
timestamp 1698431365
transform 1 0 19824 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_169
timestamp 1698431365
transform 1 0 20272 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_177
timestamp 1698431365
transform 1 0 21168 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_181
timestamp 1698431365
transform 1 0 21616 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_283
timestamp 1698431365
transform 1 0 33040 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_311
timestamp 1698431365
transform 1 0 36176 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_329
timestamp 1698431365
transform 1 0 38192 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_341
timestamp 1698431365
transform 1 0 39536 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_345
timestamp 1698431365
transform 1 0 39984 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_349
timestamp 1698431365
transform 1 0 40432 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_376
timestamp 1698431365
transform 1 0 43456 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_380
timestamp 1698431365
transform 1 0 43904 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_384
timestamp 1698431365
transform 1 0 44352 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_387
timestamp 1698431365
transform 1 0 44688 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_419
timestamp 1698431365
transform 1 0 48272 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_427
timestamp 1698431365
transform 1 0 49168 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_457
timestamp 1698431365
transform 1 0 52528 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_473
timestamp 1698431365
transform 1 0 54320 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_481
timestamp 1698431365
transform 1 0 55216 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_28
timestamp 1698431365
transform 1 0 4480 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_32
timestamp 1698431365
transform 1 0 4928 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_72
timestamp 1698431365
transform 1 0 9408 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_104
timestamp 1698431365
transform 1 0 12992 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_112
timestamp 1698431365
transform 1 0 13888 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_120
timestamp 1698431365
transform 1 0 14784 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_124
timestamp 1698431365
transform 1 0 15232 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_142
timestamp 1698431365
transform 1 0 17248 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_146
timestamp 1698431365
transform 1 0 17696 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_148
timestamp 1698431365
transform 1 0 17920 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_151
timestamp 1698431365
transform 1 0 18256 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_159
timestamp 1698431365
transform 1 0 19152 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_161
timestamp 1698431365
transform 1 0 19376 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_164
timestamp 1698431365
transform 1 0 19712 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_176
timestamp 1698431365
transform 1 0 21056 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_201
timestamp 1698431365
transform 1 0 23856 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_205
timestamp 1698431365
transform 1 0 24304 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_207
timestamp 1698431365
transform 1 0 24528 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_212
timestamp 1698431365
transform 1 0 25088 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_246
timestamp 1698431365
transform 1 0 28896 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_253
timestamp 1698431365
transform 1 0 29680 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_257
timestamp 1698431365
transform 1 0 30128 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_278
timestamp 1698431365
transform 1 0 32480 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_282
timestamp 1698431365
transform 1 0 32928 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_284
timestamp 1698431365
transform 1 0 33152 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_314
timestamp 1698431365
transform 1 0 36512 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_333
timestamp 1698431365
transform 1 0 38640 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_341
timestamp 1698431365
transform 1 0 39536 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_343
timestamp 1698431365
transform 1 0 39760 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698431365
transform 1 0 40096 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_375
timestamp 1698431365
transform 1 0 43344 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_383
timestamp 1698431365
transform 1 0 44240 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_402
timestamp 1698431365
transform 1 0 46368 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_418
timestamp 1698431365
transform 1 0 48160 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_422
timestamp 1698431365
transform 1 0 48608 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_486
timestamp 1698431365
transform 1 0 55776 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_492
timestamp 1698431365
transform 1 0 56448 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_508
timestamp 1698431365
transform 1 0 58240 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698431365
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_37
timestamp 1698431365
transform 1 0 5488 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_62
timestamp 1698431365
transform 1 0 8288 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_66
timestamp 1698431365
transform 1 0 8736 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698431365
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_107
timestamp 1698431365
transform 1 0 13328 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_121
timestamp 1698431365
transform 1 0 14896 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_123
timestamp 1698431365
transform 1 0 15120 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_141
timestamp 1698431365
transform 1 0 17136 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_155
timestamp 1698431365
transform 1 0 18704 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_171
timestamp 1698431365
transform 1 0 20496 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_177
timestamp 1698431365
transform 1 0 21168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_210
timestamp 1698431365
transform 1 0 24864 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_218
timestamp 1698431365
transform 1 0 25760 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_224
timestamp 1698431365
transform 1 0 26432 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_244
timestamp 1698431365
transform 1 0 28672 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_257
timestamp 1698431365
transform 1 0 30128 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_265
timestamp 1698431365
transform 1 0 31024 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_280
timestamp 1698431365
transform 1 0 32704 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_282
timestamp 1698431365
transform 1 0 32928 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_314
timestamp 1698431365
transform 1 0 36512 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_329
timestamp 1698431365
transform 1 0 38192 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_337
timestamp 1698431365
transform 1 0 39088 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_339
timestamp 1698431365
transform 1 0 39312 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_405
timestamp 1698431365
transform 1 0 46704 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_419
timestamp 1698431365
transform 1 0 48272 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_448
timestamp 1698431365
transform 1 0 51520 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_452
timestamp 1698431365
transform 1 0 51968 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_454
timestamp 1698431365
transform 1 0 52192 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_480
timestamp 1698431365
transform 1 0 55104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_482
timestamp 1698431365
transform 1 0 55328 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_2
timestamp 1698431365
transform 1 0 1568 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_6
timestamp 1698431365
transform 1 0 2016 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_33
timestamp 1698431365
transform 1 0 5040 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_53
timestamp 1698431365
transform 1 0 7280 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_85
timestamp 1698431365
transform 1 0 10864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_87
timestamp 1698431365
transform 1 0 11088 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_101
timestamp 1698431365
transform 1 0 12656 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_134
timestamp 1698431365
transform 1 0 16352 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_138
timestamp 1698431365
transform 1 0 16800 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_189
timestamp 1698431365
transform 1 0 22512 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_209
timestamp 1698431365
transform 1 0 24752 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_222
timestamp 1698431365
transform 1 0 26208 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_317
timestamp 1698431365
transform 1 0 36848 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_319
timestamp 1698431365
transform 1 0 37072 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_340
timestamp 1698431365
transform 1 0 39424 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_344
timestamp 1698431365
transform 1 0 39872 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_348
timestamp 1698431365
transform 1 0 40320 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_352
timestamp 1698431365
transform 1 0 40768 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_375
timestamp 1698431365
transform 1 0 43344 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_399
timestamp 1698431365
transform 1 0 46032 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_481
timestamp 1698431365
transform 1 0 55216 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_489
timestamp 1698431365
transform 1 0 56112 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_492
timestamp 1698431365
transform 1 0 56448 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_508
timestamp 1698431365
transform 1 0 58240 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698431365
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_56
timestamp 1698431365
transform 1 0 7616 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_60
timestamp 1698431365
transform 1 0 8064 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_82
timestamp 1698431365
transform 1 0 10528 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_86
timestamp 1698431365
transform 1 0 10976 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_88
timestamp 1698431365
transform 1 0 11200 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_98
timestamp 1698431365
transform 1 0 12320 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_102
timestamp 1698431365
transform 1 0 12768 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_104
timestamp 1698431365
transform 1 0 12992 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_107
timestamp 1698431365
transform 1 0 13328 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_123
timestamp 1698431365
transform 1 0 15120 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_153
timestamp 1698431365
transform 1 0 18480 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_157
timestamp 1698431365
transform 1 0 18928 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_161
timestamp 1698431365
transform 1 0 19376 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_171
timestamp 1698431365
transform 1 0 20496 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_183
timestamp 1698431365
transform 1 0 21840 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_185
timestamp 1698431365
transform 1 0 22064 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_188
timestamp 1698431365
transform 1 0 22400 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_192
timestamp 1698431365
transform 1 0 22848 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_196
timestamp 1698431365
transform 1 0 23296 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_204
timestamp 1698431365
transform 1 0 24192 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_216
timestamp 1698431365
transform 1 0 25536 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_218
timestamp 1698431365
transform 1 0 25760 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_229
timestamp 1698431365
transform 1 0 26992 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_261
timestamp 1698431365
transform 1 0 30576 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_279
timestamp 1698431365
transform 1 0 32592 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_283
timestamp 1698431365
transform 1 0 33040 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_311
timestamp 1698431365
transform 1 0 36176 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_346
timestamp 1698431365
transform 1 0 40096 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_350
timestamp 1698431365
transform 1 0 40544 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_382
timestamp 1698431365
transform 1 0 44128 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_384
timestamp 1698431365
transform 1 0 44352 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_387
timestamp 1698431365
transform 1 0 44688 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_406
timestamp 1698431365
transform 1 0 46816 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_433
timestamp 1698431365
transform 1 0 49840 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_441
timestamp 1698431365
transform 1 0 50736 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_445
timestamp 1698431365
transform 1 0 51184 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_457
timestamp 1698431365
transform 1 0 52528 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_481
timestamp 1698431365
transform 1 0 55216 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_34
timestamp 1698431365
transform 1 0 5152 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_36
timestamp 1698431365
transform 1 0 5376 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_68
timestamp 1698431365
transform 1 0 8960 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_81
timestamp 1698431365
transform 1 0 10416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_85
timestamp 1698431365
transform 1 0 10864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_87
timestamp 1698431365
transform 1 0 11088 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_139
timestamp 1698431365
transform 1 0 16912 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_152
timestamp 1698431365
transform 1 0 18368 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_156
timestamp 1698431365
transform 1 0 18816 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_164
timestamp 1698431365
transform 1 0 19712 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_168
timestamp 1698431365
transform 1 0 20160 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_170
timestamp 1698431365
transform 1 0 20384 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_220
timestamp 1698431365
transform 1 0 25984 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_227
timestamp 1698431365
transform 1 0 26768 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_231
timestamp 1698431365
transform 1 0 27216 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_235
timestamp 1698431365
transform 1 0 27664 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_267
timestamp 1698431365
transform 1 0 31248 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_271
timestamp 1698431365
transform 1 0 31696 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_279
timestamp 1698431365
transform 1 0 32592 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_282
timestamp 1698431365
transform 1 0 32928 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_286
timestamp 1698431365
transform 1 0 33376 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_338
timestamp 1698431365
transform 1 0 39200 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_346
timestamp 1698431365
transform 1 0 40096 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_352
timestamp 1698431365
transform 1 0 40768 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_360
timestamp 1698431365
transform 1 0 41664 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_373
timestamp 1698431365
transform 1 0 43120 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_375
timestamp 1698431365
transform 1 0 43344 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_389
timestamp 1698431365
transform 1 0 44912 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_405
timestamp 1698431365
transform 1 0 46704 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_413
timestamp 1698431365
transform 1 0 47600 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_417
timestamp 1698431365
transform 1 0 48048 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_419
timestamp 1698431365
transform 1 0 48272 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_422
timestamp 1698431365
transform 1 0 48608 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_426
timestamp 1698431365
transform 1 0 49056 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_428
timestamp 1698431365
transform 1 0 49280 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_434
timestamp 1698431365
transform 1 0 49952 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_442
timestamp 1698431365
transform 1 0 50848 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_446
timestamp 1698431365
transform 1 0 51296 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_465
timestamp 1698431365
transform 1 0 53424 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_480
timestamp 1698431365
transform 1 0 55104 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_488
timestamp 1698431365
transform 1 0 56000 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_505
timestamp 1698431365
transform 1 0 57904 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_14
timestamp 1698431365
transform 1 0 2912 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_37
timestamp 1698431365
transform 1 0 5488 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_39
timestamp 1698431365
transform 1 0 5712 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_61
timestamp 1698431365
transform 1 0 8176 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_65
timestamp 1698431365
transform 1 0 8624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_69
timestamp 1698431365
transform 1 0 9072 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_73
timestamp 1698431365
transform 1 0 9520 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_104
timestamp 1698431365
transform 1 0 12992 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_107
timestamp 1698431365
transform 1 0 13328 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_111
timestamp 1698431365
transform 1 0 13776 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_126
timestamp 1698431365
transform 1 0 15456 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_177
timestamp 1698431365
transform 1 0 21168 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_234
timestamp 1698431365
transform 1 0 27552 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_244
timestamp 1698431365
transform 1 0 28672 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_247
timestamp 1698431365
transform 1 0 29008 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_251
timestamp 1698431365
transform 1 0 29456 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_255
timestamp 1698431365
transform 1 0 29904 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_269
timestamp 1698431365
transform 1 0 31472 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_277
timestamp 1698431365
transform 1 0 32368 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_279
timestamp 1698431365
transform 1 0 32592 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_282
timestamp 1698431365
transform 1 0 32928 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_290
timestamp 1698431365
transform 1 0 33824 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_312
timestamp 1698431365
transform 1 0 36288 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_314
timestamp 1698431365
transform 1 0 36512 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_323
timestamp 1698431365
transform 1 0 37520 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_325
timestamp 1698431365
transform 1 0 37744 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_334
timestamp 1698431365
transform 1 0 38752 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_342
timestamp 1698431365
transform 1 0 39648 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_344
timestamp 1698431365
transform 1 0 39872 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_357
timestamp 1698431365
transform 1 0 41328 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_382
timestamp 1698431365
transform 1 0 44128 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_384
timestamp 1698431365
transform 1 0 44352 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_393
timestamp 1698431365
transform 1 0 45360 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_397
timestamp 1698431365
transform 1 0 45808 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_423
timestamp 1698431365
transform 1 0 48720 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_425
timestamp 1698431365
transform 1 0 48944 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_449
timestamp 1698431365
transform 1 0 51632 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_453
timestamp 1698431365
transform 1 0 52080 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_482
timestamp 1698431365
transform 1 0 55328 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_58
timestamp 1698431365
transform 1 0 7840 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_67
timestamp 1698431365
transform 1 0 8848 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_69
timestamp 1698431365
transform 1 0 9072 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_72
timestamp 1698431365
transform 1 0 9408 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_101
timestamp 1698431365
transform 1 0 12656 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_117
timestamp 1698431365
transform 1 0 14448 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_119
timestamp 1698431365
transform 1 0 14672 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_130
timestamp 1698431365
transform 1 0 15904 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_138
timestamp 1698431365
transform 1 0 16800 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_142
timestamp 1698431365
transform 1 0 17248 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_179
timestamp 1698431365
transform 1 0 21392 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_217
timestamp 1698431365
transform 1 0 25648 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_227
timestamp 1698431365
transform 1 0 26768 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_265
timestamp 1698431365
transform 1 0 31024 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_293
timestamp 1698431365
transform 1 0 34160 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_297
timestamp 1698431365
transform 1 0 34608 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_308
timestamp 1698431365
transform 1 0 35840 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_312
timestamp 1698431365
transform 1 0 36288 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_314
timestamp 1698431365
transform 1 0 36512 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_317
timestamp 1698431365
transform 1 0 36848 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_321
timestamp 1698431365
transform 1 0 37296 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_324
timestamp 1698431365
transform 1 0 37632 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_332
timestamp 1698431365
transform 1 0 38528 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_336
timestamp 1698431365
transform 1 0 38976 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_349
timestamp 1698431365
transform 1 0 40432 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_366
timestamp 1698431365
transform 1 0 42336 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_388
timestamp 1698431365
transform 1 0 44800 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_390
timestamp 1698431365
transform 1 0 45024 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_422
timestamp 1698431365
transform 1 0 48608 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_443
timestamp 1698431365
transform 1 0 50960 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_447
timestamp 1698431365
transform 1 0 51408 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_449
timestamp 1698431365
transform 1 0 51632 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_468
timestamp 1698431365
transform 1 0 53760 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_484
timestamp 1698431365
transform 1 0 55552 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_488
timestamp 1698431365
transform 1 0 56000 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_492
timestamp 1698431365
transform 1 0 56448 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_508
timestamp 1698431365
transform 1 0 58240 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_32
timestamp 1698431365
transform 1 0 4928 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698431365
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_37
timestamp 1698431365
transform 1 0 5488 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_45
timestamp 1698431365
transform 1 0 6384 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_80
timestamp 1698431365
transform 1 0 10304 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_86
timestamp 1698431365
transform 1 0 10976 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_102
timestamp 1698431365
transform 1 0 12768 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_104
timestamp 1698431365
transform 1 0 12992 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_136
timestamp 1698431365
transform 1 0 16576 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_150
timestamp 1698431365
transform 1 0 18144 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_154
timestamp 1698431365
transform 1 0 18592 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_177
timestamp 1698431365
transform 1 0 21168 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_181
timestamp 1698431365
transform 1 0 21616 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_185
timestamp 1698431365
transform 1 0 22064 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_244
timestamp 1698431365
transform 1 0 28672 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_247
timestamp 1698431365
transform 1 0 29008 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_258
timestamp 1698431365
transform 1 0 30240 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_270
timestamp 1698431365
transform 1 0 31584 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_272
timestamp 1698431365
transform 1 0 31808 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_280
timestamp 1698431365
transform 1 0 32704 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_282
timestamp 1698431365
transform 1 0 32928 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_305
timestamp 1698431365
transform 1 0 35504 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_312
timestamp 1698431365
transform 1 0 36288 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_314
timestamp 1698431365
transform 1 0 36512 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_322
timestamp 1698431365
transform 1 0 37408 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_331
timestamp 1698431365
transform 1 0 38416 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_335
timestamp 1698431365
transform 1 0 38864 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_359
timestamp 1698431365
transform 1 0 41552 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_363
timestamp 1698431365
transform 1 0 42000 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_383
timestamp 1698431365
transform 1 0 44240 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_404
timestamp 1698431365
transform 1 0 46592 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_406
timestamp 1698431365
transform 1 0 46816 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_436
timestamp 1698431365
transform 1 0 50176 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_444
timestamp 1698431365
transform 1 0 51072 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_448
timestamp 1698431365
transform 1 0 51520 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_468
timestamp 1698431365
transform 1 0 53760 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_479
timestamp 1698431365
transform 1 0 54992 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_495
timestamp 1698431365
transform 1 0 56784 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_503
timestamp 1698431365
transform 1 0 57680 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_507
timestamp 1698431365
transform 1 0 58128 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_30
timestamp 1698431365
transform 1 0 4704 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_55
timestamp 1698431365
transform 1 0 7504 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_72
timestamp 1698431365
transform 1 0 9408 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_76
timestamp 1698431365
transform 1 0 9856 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_80
timestamp 1698431365
transform 1 0 10304 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_87
timestamp 1698431365
transform 1 0 11088 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_95
timestamp 1698431365
transform 1 0 11984 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_99
timestamp 1698431365
transform 1 0 12432 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_150
timestamp 1698431365
transform 1 0 18144 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_154
timestamp 1698431365
transform 1 0 18592 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_162
timestamp 1698431365
transform 1 0 19488 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_170
timestamp 1698431365
transform 1 0 20384 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_174
timestamp 1698431365
transform 1 0 20832 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_177
timestamp 1698431365
transform 1 0 21168 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_193
timestamp 1698431365
transform 1 0 22960 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_195
timestamp 1698431365
transform 1 0 23184 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_202
timestamp 1698431365
transform 1 0 23968 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_206
timestamp 1698431365
transform 1 0 24416 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_212
timestamp 1698431365
transform 1 0 25088 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_216
timestamp 1698431365
transform 1 0 25536 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_220
timestamp 1698431365
transform 1 0 25984 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_228
timestamp 1698431365
transform 1 0 26880 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_242
timestamp 1698431365
transform 1 0 28448 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_248
timestamp 1698431365
transform 1 0 29120 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_252
timestamp 1698431365
transform 1 0 29568 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_262
timestamp 1698431365
transform 1 0 30688 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_270
timestamp 1698431365
transform 1 0 31584 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_272
timestamp 1698431365
transform 1 0 31808 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_287
timestamp 1698431365
transform 1 0 33488 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_291
timestamp 1698431365
transform 1 0 33936 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_295
timestamp 1698431365
transform 1 0 34384 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_335
timestamp 1698431365
transform 1 0 38864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_339
timestamp 1698431365
transform 1 0 39312 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_343
timestamp 1698431365
transform 1 0 39760 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_347
timestamp 1698431365
transform 1 0 40208 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_349
timestamp 1698431365
transform 1 0 40432 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_376
timestamp 1698431365
transform 1 0 43456 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_400
timestamp 1698431365
transform 1 0 46144 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_416
timestamp 1698431365
transform 1 0 47936 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_422
timestamp 1698431365
transform 1 0 48608 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_426
timestamp 1698431365
transform 1 0 49056 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_428
timestamp 1698431365
transform 1 0 49280 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_458
timestamp 1698431365
transform 1 0 52640 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_460
timestamp 1698431365
transform 1 0 52864 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_492
timestamp 1698431365
transform 1 0 56448 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_500
timestamp 1698431365
transform 1 0 57344 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698431365
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_53
timestamp 1698431365
transform 1 0 7280 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_59
timestamp 1698431365
transform 1 0 7952 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_63
timestamp 1698431365
transform 1 0 8400 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_71
timestamp 1698431365
transform 1 0 9296 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_75
timestamp 1698431365
transform 1 0 9744 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_77
timestamp 1698431365
transform 1 0 9968 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_96
timestamp 1698431365
transform 1 0 12096 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_100
timestamp 1698431365
transform 1 0 12544 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_102
timestamp 1698431365
transform 1 0 12768 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_107
timestamp 1698431365
transform 1 0 13328 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_109
timestamp 1698431365
transform 1 0 13552 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_139
timestamp 1698431365
transform 1 0 16912 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_143
timestamp 1698431365
transform 1 0 17360 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_145
timestamp 1698431365
transform 1 0 17584 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_161
timestamp 1698431365
transform 1 0 19376 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_183
timestamp 1698431365
transform 1 0 21840 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_187
timestamp 1698431365
transform 1 0 22288 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_197
timestamp 1698431365
transform 1 0 23408 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_201
timestamp 1698431365
transform 1 0 23856 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_205
timestamp 1698431365
transform 1 0 24304 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_207
timestamp 1698431365
transform 1 0 24528 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_214
timestamp 1698431365
transform 1 0 25312 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_255
timestamp 1698431365
transform 1 0 29904 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_259
timestamp 1698431365
transform 1 0 30352 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_261
timestamp 1698431365
transform 1 0 30576 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_293
timestamp 1698431365
transform 1 0 34160 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_297
timestamp 1698431365
transform 1 0 34608 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_301
timestamp 1698431365
transform 1 0 35056 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_309
timestamp 1698431365
transform 1 0 35952 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_313
timestamp 1698431365
transform 1 0 36400 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_317
timestamp 1698431365
transform 1 0 36848 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_325
timestamp 1698431365
transform 1 0 37744 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_331
timestamp 1698431365
transform 1 0 38416 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_335
timestamp 1698431365
transform 1 0 38864 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_343
timestamp 1698431365
transform 1 0 39760 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_365
timestamp 1698431365
transform 1 0 42224 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_369
timestamp 1698431365
transform 1 0 42672 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_379
timestamp 1698431365
transform 1 0 43792 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_383
timestamp 1698431365
transform 1 0 44240 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_387
timestamp 1698431365
transform 1 0 44688 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_391
timestamp 1698431365
transform 1 0 45136 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_393
timestamp 1698431365
transform 1 0 45360 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_400
timestamp 1698431365
transform 1 0 46144 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_465
timestamp 1698431365
transform 1 0 53424 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_467
timestamp 1698431365
transform 1 0 53648 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_78
timestamp 1698431365
transform 1 0 10080 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_120
timestamp 1698431365
transform 1 0 14784 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_134
timestamp 1698431365
transform 1 0 16352 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_138
timestamp 1698431365
transform 1 0 16800 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_170
timestamp 1698431365
transform 1 0 20384 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_174
timestamp 1698431365
transform 1 0 20832 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_186
timestamp 1698431365
transform 1 0 22176 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_208
timestamp 1698431365
transform 1 0 24640 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_212
timestamp 1698431365
transform 1 0 25088 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_216
timestamp 1698431365
transform 1 0 25536 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_233
timestamp 1698431365
transform 1 0 27440 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_268
timestamp 1698431365
transform 1 0 31360 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_272
timestamp 1698431365
transform 1 0 31808 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_282
timestamp 1698431365
transform 1 0 32928 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_286
timestamp 1698431365
transform 1 0 33376 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_304
timestamp 1698431365
transform 1 0 35392 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_308
timestamp 1698431365
transform 1 0 35840 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_316
timestamp 1698431365
transform 1 0 36736 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_318
timestamp 1698431365
transform 1 0 36960 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_352
timestamp 1698431365
transform 1 0 40768 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_354
timestamp 1698431365
transform 1 0 40992 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_398
timestamp 1698431365
transform 1 0 45920 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_402
timestamp 1698431365
transform 1 0 46368 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_465
timestamp 1698431365
transform 1 0 53424 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_467
timestamp 1698431365
transform 1 0 53648 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_486
timestamp 1698431365
transform 1 0 55776 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_492
timestamp 1698431365
transform 1 0 56448 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_500
timestamp 1698431365
transform 1 0 57344 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_2
timestamp 1698431365
transform 1 0 1568 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_19
timestamp 1698431365
transform 1 0 3472 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_33
timestamp 1698431365
transform 1 0 5040 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_52
timestamp 1698431365
transform 1 0 7168 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_78
timestamp 1698431365
transform 1 0 10080 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_107
timestamp 1698431365
transform 1 0 13328 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_160
timestamp 1698431365
transform 1 0 19264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_162
timestamp 1698431365
transform 1 0 19488 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_169
timestamp 1698431365
transform 1 0 20272 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_173
timestamp 1698431365
transform 1 0 20720 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_222
timestamp 1698431365
transform 1 0 26208 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_224
timestamp 1698431365
transform 1 0 26432 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_227
timestamp 1698431365
transform 1 0 26768 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_235
timestamp 1698431365
transform 1 0 27664 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_241
timestamp 1698431365
transform 1 0 28336 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_247
timestamp 1698431365
transform 1 0 29008 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_251
timestamp 1698431365
transform 1 0 29456 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_258
timestamp 1698431365
transform 1 0 30240 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_262
timestamp 1698431365
transform 1 0 30688 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_270
timestamp 1698431365
transform 1 0 31584 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_274
timestamp 1698431365
transform 1 0 32032 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_306
timestamp 1698431365
transform 1 0 35616 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_331
timestamp 1698431365
transform 1 0 38416 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_339
timestamp 1698431365
transform 1 0 39312 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_341
timestamp 1698431365
transform 1 0 39536 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_366
timestamp 1698431365
transform 1 0 42336 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_374
timestamp 1698431365
transform 1 0 43232 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_376
timestamp 1698431365
transform 1 0 43456 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_383
timestamp 1698431365
transform 1 0 44240 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_387
timestamp 1698431365
transform 1 0 44688 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_397
timestamp 1698431365
transform 1 0 45808 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_411
timestamp 1698431365
transform 1 0 47376 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_427
timestamp 1698431365
transform 1 0 49168 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_429
timestamp 1698431365
transform 1 0 49392 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_454
timestamp 1698431365
transform 1 0 52192 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_457
timestamp 1698431365
transform 1 0 52528 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_489
timestamp 1698431365
transform 1 0 56112 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_505
timestamp 1698431365
transform 1 0 57904 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_2
timestamp 1698431365
transform 1 0 1568 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_4
timestamp 1698431365
transform 1 0 1792 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_18
timestamp 1698431365
transform 1 0 3360 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_20
timestamp 1698431365
transform 1 0 3584 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_33
timestamp 1698431365
transform 1 0 5040 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_66
timestamp 1698431365
transform 1 0 8736 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_72
timestamp 1698431365
transform 1 0 9408 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_99
timestamp 1698431365
transform 1 0 12432 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_107
timestamp 1698431365
transform 1 0 13328 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_109
timestamp 1698431365
transform 1 0 13552 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_118
timestamp 1698431365
transform 1 0 14560 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_120
timestamp 1698431365
transform 1 0 14784 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_127
timestamp 1698431365
transform 1 0 15568 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_136
timestamp 1698431365
transform 1 0 16576 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_153
timestamp 1698431365
transform 1 0 18480 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_155
timestamp 1698431365
transform 1 0 18704 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_168
timestamp 1698431365
transform 1 0 20160 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_193
timestamp 1698431365
transform 1 0 22960 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_208
timestamp 1698431365
transform 1 0 24640 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_212
timestamp 1698431365
transform 1 0 25088 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_216
timestamp 1698431365
transform 1 0 25536 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_222
timestamp 1698431365
transform 1 0 26208 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_254
timestamp 1698431365
transform 1 0 29792 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_262
timestamp 1698431365
transform 1 0 30688 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_268
timestamp 1698431365
transform 1 0 31360 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_276
timestamp 1698431365
transform 1 0 32256 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_282
timestamp 1698431365
transform 1 0 32928 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_290
timestamp 1698431365
transform 1 0 33824 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_294
timestamp 1698431365
transform 1 0 34272 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_302
timestamp 1698431365
transform 1 0 35168 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_306
timestamp 1698431365
transform 1 0 35616 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_310
timestamp 1698431365
transform 1 0 36064 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_312
timestamp 1698431365
transform 1 0 36288 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_334
timestamp 1698431365
transform 1 0 38752 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_398
timestamp 1698431365
transform 1 0 45920 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_418
timestamp 1698431365
transform 1 0 48160 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_449
timestamp 1698431365
transform 1 0 51632 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_469
timestamp 1698431365
transform 1 0 53872 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_471
timestamp 1698431365
transform 1 0 54096 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_485
timestamp 1698431365
transform 1 0 55664 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_489
timestamp 1698431365
transform 1 0 56112 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_492
timestamp 1698431365
transform 1 0 56448 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_508
timestamp 1698431365
transform 1 0 58240 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_31
timestamp 1698431365
transform 1 0 4816 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_37
timestamp 1698431365
transform 1 0 5488 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_62
timestamp 1698431365
transform 1 0 8288 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_70
timestamp 1698431365
transform 1 0 9184 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_74
timestamp 1698431365
transform 1 0 9632 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_76
timestamp 1698431365
transform 1 0 9856 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_93
timestamp 1698431365
transform 1 0 11760 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_101
timestamp 1698431365
transform 1 0 12656 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_107
timestamp 1698431365
transform 1 0 13328 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_111
timestamp 1698431365
transform 1 0 13776 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_119
timestamp 1698431365
transform 1 0 14672 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_152
timestamp 1698431365
transform 1 0 18368 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_170
timestamp 1698431365
transform 1 0 20384 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_174
timestamp 1698431365
transform 1 0 20832 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_183
timestamp 1698431365
transform 1 0 21840 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_206
timestamp 1698431365
transform 1 0 24416 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_208
timestamp 1698431365
transform 1 0 24640 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_238
timestamp 1698431365
transform 1 0 28000 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_242
timestamp 1698431365
transform 1 0 28448 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_247
timestamp 1698431365
transform 1 0 29008 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_249
timestamp 1698431365
transform 1 0 29232 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_267
timestamp 1698431365
transform 1 0 31248 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_283
timestamp 1698431365
transform 1 0 33040 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_287
timestamp 1698431365
transform 1 0 33488 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_289
timestamp 1698431365
transform 1 0 33712 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_297
timestamp 1698431365
transform 1 0 34608 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_301
timestamp 1698431365
transform 1 0 35056 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_327
timestamp 1698431365
transform 1 0 37968 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_331
timestamp 1698431365
transform 1 0 38416 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_335
timestamp 1698431365
transform 1 0 38864 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_348
timestamp 1698431365
transform 1 0 40320 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_387
timestamp 1698431365
transform 1 0 44688 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_432
timestamp 1698431365
transform 1 0 49728 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_441
timestamp 1698431365
transform 1 0 50736 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_463
timestamp 1698431365
transform 1 0 53200 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_487
timestamp 1698431365
transform 1 0 55888 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_503
timestamp 1698431365
transform 1 0 57680 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_507
timestamp 1698431365
transform 1 0 58128 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_57
timestamp 1698431365
transform 1 0 7728 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_59
timestamp 1698431365
transform 1 0 7952 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_66
timestamp 1698431365
transform 1 0 8736 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_72
timestamp 1698431365
transform 1 0 9408 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_80
timestamp 1698431365
transform 1 0 10304 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_89
timestamp 1698431365
transform 1 0 11312 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_120
timestamp 1698431365
transform 1 0 14784 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_122
timestamp 1698431365
transform 1 0 15008 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_135
timestamp 1698431365
transform 1 0 16464 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_139
timestamp 1698431365
transform 1 0 16912 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_142
timestamp 1698431365
transform 1 0 17248 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_150
timestamp 1698431365
transform 1 0 18144 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_172
timestamp 1698431365
transform 1 0 20608 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_176
timestamp 1698431365
transform 1 0 21056 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_208
timestamp 1698431365
transform 1 0 24640 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_212
timestamp 1698431365
transform 1 0 25088 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_282
timestamp 1698431365
transform 1 0 32928 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_297
timestamp 1698431365
transform 1 0 34608 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_360
timestamp 1698431365
transform 1 0 41664 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_362
timestamp 1698431365
transform 1 0 41888 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_457
timestamp 1698431365
transform 1 0 52528 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_482
timestamp 1698431365
transform 1 0 55328 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_492
timestamp 1698431365
transform 1 0 56448 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_508
timestamp 1698431365
transform 1 0 58240 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_34
timestamp 1698431365
transform 1 0 5152 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_62
timestamp 1698431365
transform 1 0 8288 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_66
timestamp 1698431365
transform 1 0 8736 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_80
timestamp 1698431365
transform 1 0 10304 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_102
timestamp 1698431365
transform 1 0 12768 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_104
timestamp 1698431365
transform 1 0 12992 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_107
timestamp 1698431365
transform 1 0 13328 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_141
timestamp 1698431365
transform 1 0 17136 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_170
timestamp 1698431365
transform 1 0 20384 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_174
timestamp 1698431365
transform 1 0 20832 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_177
timestamp 1698431365
transform 1 0 21168 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_202
timestamp 1698431365
transform 1 0 23968 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_210
timestamp 1698431365
transform 1 0 24864 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_231
timestamp 1698431365
transform 1 0 27216 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_239
timestamp 1698431365
transform 1 0 28112 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_243
timestamp 1698431365
transform 1 0 28560 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_253
timestamp 1698431365
transform 1 0 29680 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_261
timestamp 1698431365
transform 1 0 30576 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_268
timestamp 1698431365
transform 1 0 31360 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_270
timestamp 1698431365
transform 1 0 31584 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_280
timestamp 1698431365
transform 1 0 32704 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_317
timestamp 1698431365
transform 1 0 36848 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_347
timestamp 1698431365
transform 1 0 40208 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_349
timestamp 1698431365
transform 1 0 40432 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_384
timestamp 1698431365
transform 1 0 44352 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_399
timestamp 1698431365
transform 1 0 46032 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_403
timestamp 1698431365
transform 1 0 46480 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_428
timestamp 1698431365
transform 1 0 49280 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_430
timestamp 1698431365
transform 1 0 49504 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_457
timestamp 1698431365
transform 1 0 52528 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_490
timestamp 1698431365
transform 1 0 56224 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_506
timestamp 1698431365
transform 1 0 58016 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_508
timestamp 1698431365
transform 1 0 58240 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_39
timestamp 1698431365
transform 1 0 5712 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_85
timestamp 1698431365
transform 1 0 10864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_133
timestamp 1698431365
transform 1 0 16240 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_139
timestamp 1698431365
transform 1 0 16912 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_165
timestamp 1698431365
transform 1 0 19824 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_181
timestamp 1698431365
transform 1 0 21616 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_212
timestamp 1698431365
transform 1 0 25088 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_228
timestamp 1698431365
transform 1 0 26880 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_256
timestamp 1698431365
transform 1 0 30016 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_264
timestamp 1698431365
transform 1 0 30912 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_268
timestamp 1698431365
transform 1 0 31360 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_279
timestamp 1698431365
transform 1 0 32592 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_282
timestamp 1698431365
transform 1 0 32928 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_328
timestamp 1698431365
transform 1 0 38080 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_330
timestamp 1698431365
transform 1 0 38304 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_404
timestamp 1698431365
transform 1 0 46592 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_406
timestamp 1698431365
transform 1 0 46816 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_416
timestamp 1698431365
transform 1 0 47936 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_480
timestamp 1698431365
transform 1 0 55104 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_488
timestamp 1698431365
transform 1 0 56000 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_492
timestamp 1698431365
transform 1 0 56448 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_508
timestamp 1698431365
transform 1 0 58240 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_34
timestamp 1698431365
transform 1 0 5152 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_37
timestamp 1698431365
transform 1 0 5488 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_67
timestamp 1698431365
transform 1 0 8848 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_69
timestamp 1698431365
transform 1 0 9072 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_83
timestamp 1698431365
transform 1 0 10640 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_87
timestamp 1698431365
transform 1 0 11088 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_102
timestamp 1698431365
transform 1 0 12768 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_104
timestamp 1698431365
transform 1 0 12992 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_107
timestamp 1698431365
transform 1 0 13328 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_123
timestamp 1698431365
transform 1 0 15120 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_125
timestamp 1698431365
transform 1 0 15344 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_149
timestamp 1698431365
transform 1 0 18032 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_163
timestamp 1698431365
transform 1 0 19600 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_167
timestamp 1698431365
transform 1 0 20048 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_169
timestamp 1698431365
transform 1 0 20272 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_188
timestamp 1698431365
transform 1 0 22400 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_192
timestamp 1698431365
transform 1 0 22848 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_196
timestamp 1698431365
transform 1 0 23296 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_221
timestamp 1698431365
transform 1 0 26096 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_238
timestamp 1698431365
transform 1 0 28000 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_242
timestamp 1698431365
transform 1 0 28448 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_244
timestamp 1698431365
transform 1 0 28672 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_247
timestamp 1698431365
transform 1 0 29008 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_255
timestamp 1698431365
transform 1 0 29904 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_312
timestamp 1698431365
transform 1 0 36288 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_314
timestamp 1698431365
transform 1 0 36512 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_321
timestamp 1698431365
transform 1 0 37296 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_328
timestamp 1698431365
transform 1 0 38080 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_338
timestamp 1698431365
transform 1 0 39200 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_383
timestamp 1698431365
transform 1 0 44240 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_462
timestamp 1698431365
transform 1 0 53088 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_2
timestamp 1698431365
transform 1 0 1568 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_4
timestamp 1698431365
transform 1 0 1792 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_57
timestamp 1698431365
transform 1 0 7728 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_61
timestamp 1698431365
transform 1 0 8176 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_69
timestamp 1698431365
transform 1 0 9072 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_80
timestamp 1698431365
transform 1 0 10304 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_82
timestamp 1698431365
transform 1 0 10528 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_91
timestamp 1698431365
transform 1 0 11536 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_116
timestamp 1698431365
transform 1 0 14336 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_130
timestamp 1698431365
transform 1 0 15904 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_134
timestamp 1698431365
transform 1 0 16352 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_138
timestamp 1698431365
transform 1 0 16800 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_142
timestamp 1698431365
transform 1 0 17248 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_156
timestamp 1698431365
transform 1 0 18816 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_203
timestamp 1698431365
transform 1 0 24080 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_207
timestamp 1698431365
transform 1 0 24528 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_209
timestamp 1698431365
transform 1 0 24752 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_217
timestamp 1698431365
transform 1 0 25648 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_225
timestamp 1698431365
transform 1 0 26544 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_248
timestamp 1698431365
transform 1 0 29120 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_256
timestamp 1698431365
transform 1 0 30016 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_260
timestamp 1698431365
transform 1 0 30464 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_278
timestamp 1698431365
transform 1 0 32480 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_288
timestamp 1698431365
transform 1 0 33600 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_294
timestamp 1698431365
transform 1 0 34272 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_302
timestamp 1698431365
transform 1 0 35168 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_306
timestamp 1698431365
transform 1 0 35616 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_319
timestamp 1698431365
transform 1 0 37072 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_323
timestamp 1698431365
transform 1 0 37520 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_339
timestamp 1698431365
transform 1 0 39312 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_348
timestamp 1698431365
transform 1 0 40320 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_352
timestamp 1698431365
transform 1 0 40768 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_354
timestamp 1698431365
transform 1 0 40992 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_392
timestamp 1698431365
transform 1 0 45248 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_400
timestamp 1698431365
transform 1 0 46144 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_412
timestamp 1698431365
transform 1 0 47488 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_430
timestamp 1698431365
transform 1 0 49504 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_438
timestamp 1698431365
transform 1 0 50400 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_468
timestamp 1698431365
transform 1 0 53760 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_484
timestamp 1698431365
transform 1 0 55552 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_488
timestamp 1698431365
transform 1 0 56000 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_492
timestamp 1698431365
transform 1 0 56448 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_508
timestamp 1698431365
transform 1 0 58240 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_19
timestamp 1698431365
transform 1 0 3472 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_21
timestamp 1698431365
transform 1 0 3696 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_54
timestamp 1698431365
transform 1 0 7392 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_58
timestamp 1698431365
transform 1 0 7840 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_60
timestamp 1698431365
transform 1 0 8064 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_79
timestamp 1698431365
transform 1 0 10192 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_107
timestamp 1698431365
transform 1 0 13328 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_151
timestamp 1698431365
transform 1 0 18256 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_159
timestamp 1698431365
transform 1 0 19152 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_168
timestamp 1698431365
transform 1 0 20160 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_172
timestamp 1698431365
transform 1 0 20608 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_174
timestamp 1698431365
transform 1 0 20832 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_185
timestamp 1698431365
transform 1 0 22064 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_206
timestamp 1698431365
transform 1 0 24416 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_214
timestamp 1698431365
transform 1 0 25312 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_247
timestamp 1698431365
transform 1 0 29008 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_263
timestamp 1698431365
transform 1 0 30800 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_271
timestamp 1698431365
transform 1 0 31696 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_273
timestamp 1698431365
transform 1 0 31920 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_314
timestamp 1698431365
transform 1 0 36512 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_322
timestamp 1698431365
transform 1 0 37408 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_401
timestamp 1698431365
transform 1 0 46256 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_403
timestamp 1698431365
transform 1 0 46480 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_433
timestamp 1698431365
transform 1 0 49840 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_437
timestamp 1698431365
transform 1 0 50288 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_454
timestamp 1698431365
transform 1 0 52192 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_457
timestamp 1698431365
transform 1 0 52528 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_494
timestamp 1698431365
transform 1 0 56672 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_502
timestamp 1698431365
transform 1 0 57568 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_506
timestamp 1698431365
transform 1 0 58016 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_508
timestamp 1698431365
transform 1 0 58240 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_8
timestamp 1698431365
transform 1 0 2240 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_10
timestamp 1698431365
transform 1 0 2464 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_20
timestamp 1698431365
transform 1 0 3584 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_61
timestamp 1698431365
transform 1 0 8176 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_72
timestamp 1698431365
transform 1 0 9408 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_132
timestamp 1698431365
transform 1 0 16128 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_139
timestamp 1698431365
transform 1 0 16912 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_173
timestamp 1698431365
transform 1 0 20720 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_189
timestamp 1698431365
transform 1 0 22512 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_201
timestamp 1698431365
transform 1 0 23856 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_209
timestamp 1698431365
transform 1 0 24752 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_212
timestamp 1698431365
transform 1 0 25088 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_220
timestamp 1698431365
transform 1 0 25984 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_53_237
timestamp 1698431365
transform 1 0 27888 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_269
timestamp 1698431365
transform 1 0 31472 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_278
timestamp 1698431365
transform 1 0 32480 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_282
timestamp 1698431365
transform 1 0 32928 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_291
timestamp 1698431365
transform 1 0 33936 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_302
timestamp 1698431365
transform 1 0 35168 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_339
timestamp 1698431365
transform 1 0 39312 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_347
timestamp 1698431365
transform 1 0 40208 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_349
timestamp 1698431365
transform 1 0 40432 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_352
timestamp 1698431365
transform 1 0 40768 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_356
timestamp 1698431365
transform 1 0 41216 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_358
timestamp 1698431365
transform 1 0 41440 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_367
timestamp 1698431365
transform 1 0 42448 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_393
timestamp 1698431365
transform 1 0 45360 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_395
timestamp 1698431365
transform 1 0 45584 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_404
timestamp 1698431365
transform 1 0 46592 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_412
timestamp 1698431365
transform 1 0 47488 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_422
timestamp 1698431365
transform 1 0 48608 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_438
timestamp 1698431365
transform 1 0 50400 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_446
timestamp 1698431365
transform 1 0 51296 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_470
timestamp 1698431365
transform 1 0 53984 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_479
timestamp 1698431365
transform 1 0 54992 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_487
timestamp 1698431365
transform 1 0 55888 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_489
timestamp 1698431365
transform 1 0 56112 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_492
timestamp 1698431365
transform 1 0 56448 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_508
timestamp 1698431365
transform 1 0 58240 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_2
timestamp 1698431365
transform 1 0 1568 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_76
timestamp 1698431365
transform 1 0 9856 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_78
timestamp 1698431365
transform 1 0 10080 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_107
timestamp 1698431365
transform 1 0 13328 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_117
timestamp 1698431365
transform 1 0 14448 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_125
timestamp 1698431365
transform 1 0 15344 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_149
timestamp 1698431365
transform 1 0 18032 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_153
timestamp 1698431365
transform 1 0 18480 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_160
timestamp 1698431365
transform 1 0 19264 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_168
timestamp 1698431365
transform 1 0 20160 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_172
timestamp 1698431365
transform 1 0 20608 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_174
timestamp 1698431365
transform 1 0 20832 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_177
timestamp 1698431365
transform 1 0 21168 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_215
timestamp 1698431365
transform 1 0 25424 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_225
timestamp 1698431365
transform 1 0 26544 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_227
timestamp 1698431365
transform 1 0 26768 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_236
timestamp 1698431365
transform 1 0 27776 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_244
timestamp 1698431365
transform 1 0 28672 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_292
timestamp 1698431365
transform 1 0 34048 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_299
timestamp 1698431365
transform 1 0 34832 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_317
timestamp 1698431365
transform 1 0 36848 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_366
timestamp 1698431365
transform 1 0 42336 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_370
timestamp 1698431365
transform 1 0 42784 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_381
timestamp 1698431365
transform 1 0 44016 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_395
timestamp 1698431365
transform 1 0 45584 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_402
timestamp 1698431365
transform 1 0 46368 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_416
timestamp 1698431365
transform 1 0 47936 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_420
timestamp 1698431365
transform 1 0 48384 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_435
timestamp 1698431365
transform 1 0 50064 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_439
timestamp 1698431365
transform 1 0 50512 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_453
timestamp 1698431365
transform 1 0 52080 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_462
timestamp 1698431365
transform 1 0 53088 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_466
timestamp 1698431365
transform 1 0 53536 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_480
timestamp 1698431365
transform 1 0 55104 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_496
timestamp 1698431365
transform 1 0 56896 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_504
timestamp 1698431365
transform 1 0 57792 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_508
timestamp 1698431365
transform 1 0 58240 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_2
timestamp 1698431365
transform 1 0 1568 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_4
timestamp 1698431365
transform 1 0 1792 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_25
timestamp 1698431365
transform 1 0 4144 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_27
timestamp 1698431365
transform 1 0 4368 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_72
timestamp 1698431365
transform 1 0 9408 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_89
timestamp 1698431365
transform 1 0 11312 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_104
timestamp 1698431365
transform 1 0 12992 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_113
timestamp 1698431365
transform 1 0 14000 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_129
timestamp 1698431365
transform 1 0 15792 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_136
timestamp 1698431365
transform 1 0 16576 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_142
timestamp 1698431365
transform 1 0 17248 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_144
timestamp 1698431365
transform 1 0 17472 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_151
timestamp 1698431365
transform 1 0 18256 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_159
timestamp 1698431365
transform 1 0 19152 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_175
timestamp 1698431365
transform 1 0 20944 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_208
timestamp 1698431365
transform 1 0 24640 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_212
timestamp 1698431365
transform 1 0 25088 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_214
timestamp 1698431365
transform 1 0 25312 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_235
timestamp 1698431365
transform 1 0 27664 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_243
timestamp 1698431365
transform 1 0 28560 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_273
timestamp 1698431365
transform 1 0 31920 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_277
timestamp 1698431365
transform 1 0 32368 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_279
timestamp 1698431365
transform 1 0 32592 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_333
timestamp 1698431365
transform 1 0 38640 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_337
timestamp 1698431365
transform 1 0 39088 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_339
timestamp 1698431365
transform 1 0 39312 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_365
timestamp 1698431365
transform 1 0 42224 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_367
timestamp 1698431365
transform 1 0 42448 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_404
timestamp 1698431365
transform 1 0 46592 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_412
timestamp 1698431365
transform 1 0 47488 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_419
timestamp 1698431365
transform 1 0 48272 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_450
timestamp 1698431365
transform 1 0 51744 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_475
timestamp 1698431365
transform 1 0 54544 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_483
timestamp 1698431365
transform 1 0 55440 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_487
timestamp 1698431365
transform 1 0 55888 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_489
timestamp 1698431365
transform 1 0 56112 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_492
timestamp 1698431365
transform 1 0 56448 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_508
timestamp 1698431365
transform 1 0 58240 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_8
timestamp 1698431365
transform 1 0 2240 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_19
timestamp 1698431365
transform 1 0 3472 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_31
timestamp 1698431365
transform 1 0 4816 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_49
timestamp 1698431365
transform 1 0 6832 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_51
timestamp 1698431365
transform 1 0 7056 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_64
timestamp 1698431365
transform 1 0 8512 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_68
timestamp 1698431365
transform 1 0 8960 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_70
timestamp 1698431365
transform 1 0 9184 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_107
timestamp 1698431365
transform 1 0 13328 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_156
timestamp 1698431365
transform 1 0 18816 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_160
timestamp 1698431365
transform 1 0 19264 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_171
timestamp 1698431365
transform 1 0 20496 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_185
timestamp 1698431365
transform 1 0 22064 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_189
timestamp 1698431365
transform 1 0 22512 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_198
timestamp 1698431365
transform 1 0 23520 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_211
timestamp 1698431365
transform 1 0 24976 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_239
timestamp 1698431365
transform 1 0 28112 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_243
timestamp 1698431365
transform 1 0 28560 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_247
timestamp 1698431365
transform 1 0 29008 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_255
timestamp 1698431365
transform 1 0 29904 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_257
timestamp 1698431365
transform 1 0 30128 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_276
timestamp 1698431365
transform 1 0 32256 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_314
timestamp 1698431365
transform 1 0 36512 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_317
timestamp 1698431365
transform 1 0 36848 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_325
timestamp 1698431365
transform 1 0 37744 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_343
timestamp 1698431365
transform 1 0 39760 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_351
timestamp 1698431365
transform 1 0 40656 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_353
timestamp 1698431365
transform 1 0 40880 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_383
timestamp 1698431365
transform 1 0 44240 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_387
timestamp 1698431365
transform 1 0 44688 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_403
timestamp 1698431365
transform 1 0 46480 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_407
timestamp 1698431365
transform 1 0 46928 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_409
timestamp 1698431365
transform 1 0 47152 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_451
timestamp 1698431365
transform 1 0 51856 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_481
timestamp 1698431365
transform 1 0 55216 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_497
timestamp 1698431365
transform 1 0 57008 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_505
timestamp 1698431365
transform 1 0 57904 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_2
timestamp 1698431365
transform 1 0 1568 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_68
timestamp 1698431365
transform 1 0 8960 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_72
timestamp 1698431365
transform 1 0 9408 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_116
timestamp 1698431365
transform 1 0 14336 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_142
timestamp 1698431365
transform 1 0 17248 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_150
timestamp 1698431365
transform 1 0 18144 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_157
timestamp 1698431365
transform 1 0 18928 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_159
timestamp 1698431365
transform 1 0 19152 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_167
timestamp 1698431365
transform 1 0 20048 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_192
timestamp 1698431365
transform 1 0 22848 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_208
timestamp 1698431365
transform 1 0 24640 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_212
timestamp 1698431365
transform 1 0 25088 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_229
timestamp 1698431365
transform 1 0 26992 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_245
timestamp 1698431365
transform 1 0 28784 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_249
timestamp 1698431365
transform 1 0 29232 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_251
timestamp 1698431365
transform 1 0 29456 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_258
timestamp 1698431365
transform 1 0 30240 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_268
timestamp 1698431365
transform 1 0 31360 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_272
timestamp 1698431365
transform 1 0 31808 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_274
timestamp 1698431365
transform 1 0 32032 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_302
timestamp 1698431365
transform 1 0 35168 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_352
timestamp 1698431365
transform 1 0 40768 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_356
timestamp 1698431365
transform 1 0 41216 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_416
timestamp 1698431365
transform 1 0 47936 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_422
timestamp 1698431365
transform 1 0 48608 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_438
timestamp 1698431365
transform 1 0 50400 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_445
timestamp 1698431365
transform 1 0 51184 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_469
timestamp 1698431365
transform 1 0 53872 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_485
timestamp 1698431365
transform 1 0 55664 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_489
timestamp 1698431365
transform 1 0 56112 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_492
timestamp 1698431365
transform 1 0 56448 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_508
timestamp 1698431365
transform 1 0 58240 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_19
timestamp 1698431365
transform 1 0 3472 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_25
timestamp 1698431365
transform 1 0 4144 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_27
timestamp 1698431365
transform 1 0 4368 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_83
timestamp 1698431365
transform 1 0 10640 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_93
timestamp 1698431365
transform 1 0 11760 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_101
timestamp 1698431365
transform 1 0 12656 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_142
timestamp 1698431365
transform 1 0 17248 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_150
timestamp 1698431365
transform 1 0 18144 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_177
timestamp 1698431365
transform 1 0 21168 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_210
timestamp 1698431365
transform 1 0 24864 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_218
timestamp 1698431365
transform 1 0 25760 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_222
timestamp 1698431365
transform 1 0 26208 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_224
timestamp 1698431365
transform 1 0 26432 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_247
timestamp 1698431365
transform 1 0 29008 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_251
timestamp 1698431365
transform 1 0 29456 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_291
timestamp 1698431365
transform 1 0 33936 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_303
timestamp 1698431365
transform 1 0 35280 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_332
timestamp 1698431365
transform 1 0 38528 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_362
timestamp 1698431365
transform 1 0 41888 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_378
timestamp 1698431365
transform 1 0 43680 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_382
timestamp 1698431365
transform 1 0 44128 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_384
timestamp 1698431365
transform 1 0 44352 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_387
timestamp 1698431365
transform 1 0 44688 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_411
timestamp 1698431365
transform 1 0 47376 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_419
timestamp 1698431365
transform 1 0 48272 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_423
timestamp 1698431365
transform 1 0 48720 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_425
timestamp 1698431365
transform 1 0 48944 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_433
timestamp 1698431365
transform 1 0 49840 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_450
timestamp 1698431365
transform 1 0 51744 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_454
timestamp 1698431365
transform 1 0 52192 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_457
timestamp 1698431365
transform 1 0 52528 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_464
timestamp 1698431365
transform 1 0 53312 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_58_470
timestamp 1698431365
transform 1 0 53984 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_502
timestamp 1698431365
transform 1 0 57568 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_506
timestamp 1698431365
transform 1 0 58016 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_508
timestamp 1698431365
transform 1 0 58240 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_2
timestamp 1698431365
transform 1 0 1568 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_4
timestamp 1698431365
transform 1 0 1792 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_7
timestamp 1698431365
transform 1 0 2128 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_11
timestamp 1698431365
transform 1 0 2576 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_15
timestamp 1698431365
transform 1 0 3024 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_19
timestamp 1698431365
transform 1 0 3472 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_23
timestamp 1698431365
transform 1 0 3920 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_27
timestamp 1698431365
transform 1 0 4368 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_31
timestamp 1698431365
transform 1 0 4816 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_72
timestamp 1698431365
transform 1 0 9408 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_80
timestamp 1698431365
transform 1 0 10304 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_105
timestamp 1698431365
transform 1 0 13104 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_116
timestamp 1698431365
transform 1 0 14336 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_120
timestamp 1698431365
transform 1 0 14784 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_130
timestamp 1698431365
transform 1 0 15904 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_138
timestamp 1698431365
transform 1 0 16800 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_142
timestamp 1698431365
transform 1 0 17248 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_150
timestamp 1698431365
transform 1 0 18144 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_154
timestamp 1698431365
transform 1 0 18592 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_176
timestamp 1698431365
transform 1 0 21056 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_200
timestamp 1698431365
transform 1 0 23744 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_208
timestamp 1698431365
transform 1 0 24640 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_212
timestamp 1698431365
transform 1 0 25088 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_245
timestamp 1698431365
transform 1 0 28784 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_247
timestamp 1698431365
transform 1 0 29008 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_266
timestamp 1698431365
transform 1 0 31136 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_327
timestamp 1698431365
transform 1 0 37968 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_341
timestamp 1698431365
transform 1 0 39536 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_349
timestamp 1698431365
transform 1 0 40432 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_352
timestamp 1698431365
transform 1 0 40768 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_356
timestamp 1698431365
transform 1 0 41216 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_363
timestamp 1698431365
transform 1 0 42000 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_391
timestamp 1698431365
transform 1 0 45136 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_399
timestamp 1698431365
transform 1 0 46032 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_401
timestamp 1698431365
transform 1 0 46256 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_416
timestamp 1698431365
transform 1 0 47936 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_472
timestamp 1698431365
transform 1 0 54208 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_488
timestamp 1698431365
transform 1 0 56000 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_492
timestamp 1698431365
transform 1 0 56448 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_508
timestamp 1698431365
transform 1 0 58240 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_8
timestamp 1698431365
transform 1 0 2240 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_12
timestamp 1698431365
transform 1 0 2688 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_16
timestamp 1698431365
transform 1 0 3136 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_18
timestamp 1698431365
transform 1 0 3360 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_21
timestamp 1698431365
transform 1 0 3696 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_25
timestamp 1698431365
transform 1 0 4144 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_33
timestamp 1698431365
transform 1 0 5040 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_43
timestamp 1698431365
transform 1 0 6160 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_68
timestamp 1698431365
transform 1 0 8960 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_72
timestamp 1698431365
transform 1 0 9408 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_88
timestamp 1698431365
transform 1 0 11200 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_102
timestamp 1698431365
transform 1 0 12768 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_104
timestamp 1698431365
transform 1 0 12992 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_155
timestamp 1698431365
transform 1 0 18704 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_163
timestamp 1698431365
transform 1 0 19600 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_165
timestamp 1698431365
transform 1 0 19824 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_171
timestamp 1698431365
transform 1 0 20496 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_177
timestamp 1698431365
transform 1 0 21168 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_186
timestamp 1698431365
transform 1 0 22176 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_192
timestamp 1698431365
transform 1 0 22848 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_196
timestamp 1698431365
transform 1 0 23296 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_198
timestamp 1698431365
transform 1 0 23520 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_212
timestamp 1698431365
transform 1 0 25088 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_221
timestamp 1698431365
transform 1 0 26096 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_236
timestamp 1698431365
transform 1 0 27776 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_244
timestamp 1698431365
transform 1 0 28672 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_247
timestamp 1698431365
transform 1 0 29008 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_255
timestamp 1698431365
transform 1 0 29904 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_267
timestamp 1698431365
transform 1 0 31248 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_306
timestamp 1698431365
transform 1 0 35616 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_317
timestamp 1698431365
transform 1 0 36848 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_382
timestamp 1698431365
transform 1 0 44128 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_384
timestamp 1698431365
transform 1 0 44352 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_387
timestamp 1698431365
transform 1 0 44688 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_397
timestamp 1698431365
transform 1 0 45808 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_401
timestamp 1698431365
transform 1 0 46256 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_453
timestamp 1698431365
transform 1 0 52080 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_60_466
timestamp 1698431365
transform 1 0 53536 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_498
timestamp 1698431365
transform 1 0 57120 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_506
timestamp 1698431365
transform 1 0 58016 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_508
timestamp 1698431365
transform 1 0 58240 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_2
timestamp 1698431365
transform 1 0 1568 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_6
timestamp 1698431365
transform 1 0 2016 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_38
timestamp 1698431365
transform 1 0 5600 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_46
timestamp 1698431365
transform 1 0 6496 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_65
timestamp 1698431365
transform 1 0 8624 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_69
timestamp 1698431365
transform 1 0 9072 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_72
timestamp 1698431365
transform 1 0 9408 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_76
timestamp 1698431365
transform 1 0 9856 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_82
timestamp 1698431365
transform 1 0 10528 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_139
timestamp 1698431365
transform 1 0 16912 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_184
timestamp 1698431365
transform 1 0 21952 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_191
timestamp 1698431365
transform 1 0 22736 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_199
timestamp 1698431365
transform 1 0 23632 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_203
timestamp 1698431365
transform 1 0 24080 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_212
timestamp 1698431365
transform 1 0 25088 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_242
timestamp 1698431365
transform 1 0 28448 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_250
timestamp 1698431365
transform 1 0 29344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_252
timestamp 1698431365
transform 1 0 29568 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_272
timestamp 1698431365
transform 1 0 31808 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_288
timestamp 1698431365
transform 1 0 33600 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_327
timestamp 1698431365
transform 1 0 37968 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_342
timestamp 1698431365
transform 1 0 39648 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_362
timestamp 1698431365
transform 1 0 41888 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_417
timestamp 1698431365
transform 1 0 48048 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_419
timestamp 1698431365
transform 1 0 48272 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_428
timestamp 1698431365
transform 1 0 49280 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_453
timestamp 1698431365
transform 1 0 52080 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_485
timestamp 1698431365
transform 1 0 55664 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_489
timestamp 1698431365
transform 1 0 56112 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_492
timestamp 1698431365
transform 1 0 56448 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_508
timestamp 1698431365
transform 1 0 58240 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_62_2
timestamp 1698431365
transform 1 0 1568 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_34
timestamp 1698431365
transform 1 0 5152 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_37
timestamp 1698431365
transform 1 0 5488 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_45
timestamp 1698431365
transform 1 0 6384 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_49
timestamp 1698431365
transform 1 0 6832 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_62
timestamp 1698431365
transform 1 0 8288 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_70
timestamp 1698431365
transform 1 0 9184 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_74
timestamp 1698431365
transform 1 0 9632 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_76
timestamp 1698431365
transform 1 0 9856 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_90
timestamp 1698431365
transform 1 0 11424 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_92
timestamp 1698431365
transform 1 0 11648 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_101
timestamp 1698431365
transform 1 0 12656 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_107
timestamp 1698431365
transform 1 0 13328 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_111
timestamp 1698431365
transform 1 0 13776 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_174
timestamp 1698431365
transform 1 0 20832 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_190
timestamp 1698431365
transform 1 0 22624 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_214
timestamp 1698431365
transform 1 0 25312 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_234
timestamp 1698431365
transform 1 0 27552 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_242
timestamp 1698431365
transform 1 0 28448 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_244
timestamp 1698431365
transform 1 0 28672 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_247
timestamp 1698431365
transform 1 0 29008 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_251
timestamp 1698431365
transform 1 0 29456 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_271
timestamp 1698431365
transform 1 0 31696 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_273
timestamp 1698431365
transform 1 0 31920 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_380
timestamp 1698431365
transform 1 0 43904 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_384
timestamp 1698431365
transform 1 0 44352 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_387
timestamp 1698431365
transform 1 0 44688 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_415
timestamp 1698431365
transform 1 0 47824 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_433
timestamp 1698431365
transform 1 0 49840 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_440
timestamp 1698431365
transform 1 0 50624 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_444
timestamp 1698431365
transform 1 0 51072 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_452
timestamp 1698431365
transform 1 0 51968 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_454
timestamp 1698431365
transform 1 0 52192 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_62_457
timestamp 1698431365
transform 1 0 52528 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_489
timestamp 1698431365
transform 1 0 56112 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_505
timestamp 1698431365
transform 1 0 57904 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_2
timestamp 1698431365
transform 1 0 1568 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_66
timestamp 1698431365
transform 1 0 8736 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_72
timestamp 1698431365
transform 1 0 9408 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_76
timestamp 1698431365
transform 1 0 9856 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_89
timestamp 1698431365
transform 1 0 11312 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_116
timestamp 1698431365
transform 1 0 14336 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_120
timestamp 1698431365
transform 1 0 14784 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_123
timestamp 1698431365
transform 1 0 15120 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_130
timestamp 1698431365
transform 1 0 15904 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_134
timestamp 1698431365
transform 1 0 16352 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_138
timestamp 1698431365
transform 1 0 16800 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_155
timestamp 1698431365
transform 1 0 18704 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_212
timestamp 1698431365
transform 1 0 25088 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_229
timestamp 1698431365
transform 1 0 26992 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_245
timestamp 1698431365
transform 1 0 28784 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_263
timestamp 1698431365
transform 1 0 30800 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_314
timestamp 1698431365
transform 1 0 36512 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_349
timestamp 1698431365
transform 1 0 40432 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_360
timestamp 1698431365
transform 1 0 41664 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_388
timestamp 1698431365
transform 1 0 44800 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_418
timestamp 1698431365
transform 1 0 48160 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_422
timestamp 1698431365
transform 1 0 48608 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_429
timestamp 1698431365
transform 1 0 49392 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_63_433
timestamp 1698431365
transform 1 0 49840 0 -1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_465
timestamp 1698431365
transform 1 0 53424 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_481
timestamp 1698431365
transform 1 0 55216 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_489
timestamp 1698431365
transform 1 0 56112 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_492
timestamp 1698431365
transform 1 0 56448 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_508
timestamp 1698431365
transform 1 0 58240 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_64_2
timestamp 1698431365
transform 1 0 1568 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_34
timestamp 1698431365
transform 1 0 5152 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_37
timestamp 1698431365
transform 1 0 5488 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_101
timestamp 1698431365
transform 1 0 12656 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_64_117
timestamp 1698431365
transform 1 0 14448 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_149
timestamp 1698431365
transform 1 0 18032 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_165
timestamp 1698431365
transform 1 0 19824 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_173
timestamp 1698431365
transform 1 0 20720 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_185
timestamp 1698431365
transform 1 0 22064 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_192
timestamp 1698431365
transform 1 0 22848 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_196
timestamp 1698431365
transform 1 0 23296 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_221
timestamp 1698431365
transform 1 0 26096 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_237
timestamp 1698431365
transform 1 0 27888 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_247
timestamp 1698431365
transform 1 0 29008 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_251
timestamp 1698431365
transform 1 0 29456 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_253
timestamp 1698431365
transform 1 0 29680 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_312
timestamp 1698431365
transform 1 0 36288 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_314
timestamp 1698431365
transform 1 0 36512 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_348
timestamp 1698431365
transform 1 0 40320 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_364
timestamp 1698431365
transform 1 0 42112 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_377
timestamp 1698431365
transform 1 0 43568 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_392
timestamp 1698431365
transform 1 0 45248 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_408
timestamp 1698431365
transform 1 0 47040 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_412
timestamp 1698431365
transform 1 0 47488 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_64_416
timestamp 1698431365
transform 1 0 47936 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_448
timestamp 1698431365
transform 1 0 51520 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_452
timestamp 1698431365
transform 1 0 51968 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_454
timestamp 1698431365
transform 1 0 52192 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_64_457
timestamp 1698431365
transform 1 0 52528 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_489
timestamp 1698431365
transform 1 0 56112 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_505
timestamp 1698431365
transform 1 0 57904 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_2
timestamp 1698431365
transform 1 0 1568 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_66
timestamp 1698431365
transform 1 0 8736 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_72
timestamp 1698431365
transform 1 0 9408 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_136
timestamp 1698431365
transform 1 0 16576 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_142
timestamp 1698431365
transform 1 0 17248 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_206
timestamp 1698431365
transform 1 0 24416 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_212
timestamp 1698431365
transform 1 0 25088 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_220
timestamp 1698431365
transform 1 0 25984 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_231
timestamp 1698431365
transform 1 0 27216 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_235
timestamp 1698431365
transform 1 0 27664 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_239
timestamp 1698431365
transform 1 0 28112 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_243
timestamp 1698431365
transform 1 0 28560 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_259
timestamp 1698431365
transform 1 0 30352 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_267
timestamp 1698431365
transform 1 0 31248 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_271
timestamp 1698431365
transform 1 0 31696 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_274
timestamp 1698431365
transform 1 0 32032 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_282
timestamp 1698431365
transform 1 0 32928 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_349
timestamp 1698431365
transform 1 0 40432 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_352
timestamp 1698431365
transform 1 0 40768 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_356
timestamp 1698431365
transform 1 0 41216 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_422
timestamp 1698431365
transform 1 0 48608 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_486
timestamp 1698431365
transform 1 0 55776 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_492
timestamp 1698431365
transform 1 0 56448 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_508
timestamp 1698431365
transform 1 0 58240 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_2
timestamp 1698431365
transform 1 0 1568 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_34
timestamp 1698431365
transform 1 0 5152 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_37
timestamp 1698431365
transform 1 0 5488 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_101
timestamp 1698431365
transform 1 0 12656 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_107
timestamp 1698431365
transform 1 0 13328 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_171
timestamp 1698431365
transform 1 0 20496 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_177
timestamp 1698431365
transform 1 0 21168 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_193
timestamp 1698431365
transform 1 0 22960 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_201
timestamp 1698431365
transform 1 0 23856 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_237
timestamp 1698431365
transform 1 0 27888 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_241
timestamp 1698431365
transform 1 0 28336 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_255
timestamp 1698431365
transform 1 0 29904 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_265
timestamp 1698431365
transform 1 0 31024 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_269
timestamp 1698431365
transform 1 0 31472 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_273
timestamp 1698431365
transform 1 0 31920 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_311
timestamp 1698431365
transform 1 0 36176 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_357
timestamp 1698431365
transform 1 0 41328 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_361
timestamp 1698431365
transform 1 0 41776 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_365
timestamp 1698431365
transform 1 0 42224 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_369
timestamp 1698431365
transform 1 0 42672 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_387
timestamp 1698431365
transform 1 0 44688 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_419
timestamp 1698431365
transform 1 0 48272 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_435
timestamp 1698431365
transform 1 0 50064 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_439
timestamp 1698431365
transform 1 0 50512 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_441
timestamp 1698431365
transform 1 0 50736 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_444
timestamp 1698431365
transform 1 0 51072 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_452
timestamp 1698431365
transform 1 0 51968 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_454
timestamp 1698431365
transform 1 0 52192 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_457
timestamp 1698431365
transform 1 0 52528 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_489
timestamp 1698431365
transform 1 0 56112 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_505
timestamp 1698431365
transform 1 0 57904 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_2
timestamp 1698431365
transform 1 0 1568 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_36
timestamp 1698431365
transform 1 0 5376 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_70
timestamp 1698431365
transform 1 0 9184 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_104
timestamp 1698431365
transform 1 0 12992 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_138
timestamp 1698431365
transform 1 0 16800 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_172
timestamp 1698431365
transform 1 0 20608 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_188
timestamp 1698431365
transform 1 0 22400 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_362
timestamp 1698431365
transform 1 0 41888 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_366
timestamp 1698431365
transform 1 0 42336 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_370
timestamp 1698431365
transform 1 0 42784 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_376
timestamp 1698431365
transform 1 0 43456 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_380
timestamp 1698431365
transform 1 0 43904 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_396
timestamp 1698431365
transform 1 0 45696 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_404
timestamp 1698431365
transform 1 0 46592 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_410
timestamp 1698431365
transform 1 0 47264 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_426
timestamp 1698431365
transform 1 0 49056 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_430
timestamp 1698431365
transform 1 0 49504 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_439
timestamp 1698431365
transform 1 0 50512 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_441
timestamp 1698431365
transform 1 0 50736 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_450
timestamp 1698431365
transform 1 0 51744 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_466
timestamp 1698431365
transform 1 0 53536 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_474
timestamp 1698431365
transform 1 0 54432 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_478
timestamp 1698431365
transform 1 0 54880 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_494
timestamp 1698431365
transform 1 0 56672 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_502
timestamp 1698431365
transform 1 0 57568 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_506
timestamp 1698431365
transform 1 0 58016 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_508
timestamp 1698431365
transform 1 0 58240 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input2
timestamp 1698431365
transform -1 0 25088 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input3
timestamp 1698431365
transform 1 0 26320 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input4
timestamp 1698431365
transform 1 0 29008 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1698431365
transform 1 0 1568 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1698431365
transform 1 0 2912 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1698431365
transform 1 0 1568 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1698431365
transform 1 0 2240 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input9
timestamp 1698431365
transform 1 0 1568 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input10
timestamp 1698431365
transform 1 0 2240 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input11
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input12
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input13
timestamp 1698431365
transform 1 0 2912 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input14
timestamp 1698431365
transform 1 0 2240 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input15
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input16
timestamp 1698431365
transform 1 0 2240 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input17
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input18
timestamp 1698431365
transform 1 0 1568 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input19
timestamp 1698431365
transform -1 0 44128 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input20
timestamp 1698431365
transform -1 0 42560 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input21
timestamp 1698431365
transform -1 0 46816 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input22
timestamp 1698431365
transform -1 0 47936 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input23
timestamp 1698431365
transform 1 0 47936 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input24
timestamp 1698431365
transform 1 0 49840 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input25
timestamp 1698431365
transform -1 0 3584 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input26
timestamp 1698431365
transform -1 0 2912 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input27
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input28
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input29
timestamp 1698431365
transform 1 0 4480 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input30
timestamp 1698431365
transform 1 0 2240 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input31
timestamp 1698431365
transform 1 0 2464 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input32
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input33
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input34
timestamp 1698431365
transform 1 0 29008 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input35
timestamp 1698431365
transform 1 0 29680 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input36
timestamp 1698431365
transform 1 0 30352 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input37
timestamp 1698431365
transform -1 0 40544 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input38
timestamp 1698431365
transform -1 0 41888 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input39
timestamp 1698431365
transform -1 0 40432 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input40
timestamp 1698431365
transform -1 0 6384 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input41
timestamp 1698431365
transform 1 0 49840 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input42
timestamp 1698431365
transform 1 0 51072 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input43
timestamp 1698431365
transform 1 0 5488 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input44
timestamp 1698431365
transform 1 0 1568 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input45
timestamp 1698431365
transform 1 0 2240 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input46
timestamp 1698431365
transform 1 0 1680 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input47
timestamp 1698431365
transform 1 0 1568 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input48
timestamp 1698431365
transform -1 0 41440 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input49
timestamp 1698431365
transform 1 0 28224 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input50
timestamp 1698431365
transform -1 0 6384 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input51
timestamp 1698431365
transform -1 0 44800 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input52
timestamp 1698431365
transform -1 0 45248 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input53
timestamp 1698431365
transform -1 0 46144 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input54
timestamp 1698431365
transform -1 0 45472 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input55
timestamp 1698431365
transform -1 0 58352 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input56
timestamp 1698431365
transform -1 0 58352 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input57
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input58
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input59
timestamp 1698431365
transform 1 0 2240 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input60
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input61
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input62
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input63
timestamp 1698431365
transform 1 0 2912 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input64
timestamp 1698431365
transform 1 0 22288 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input65
timestamp 1698431365
transform -1 0 25088 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input66
timestamp 1698431365
transform 1 0 27216 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input67
timestamp 1698431365
transform -1 0 31808 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input68
timestamp 1698431365
transform -1 0 35616 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input69
timestamp 1698431365
transform -1 0 41216 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input70
timestamp 1698431365
transform -1 0 39424 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input71
timestamp 1698431365
transform -1 0 41328 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input72
timestamp 1698431365
transform 1 0 1568 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input73
timestamp 1698431365
transform -1 0 58352 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input74
timestamp 1698431365
transform -1 0 58352 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input75
timestamp 1698431365
transform 1 0 6384 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input76
timestamp 1698431365
transform 1 0 1568 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input77
timestamp 1698431365
transform 1 0 1568 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input78
timestamp 1698431365
transform 1 0 5376 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input79
timestamp 1698431365
transform 1 0 23520 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input80
timestamp 1698431365
transform 1 0 28112 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input81
timestamp 1698431365
transform -1 0 35616 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input82
timestamp 1698431365
transform 1 0 2240 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  max_cap117
timestamp 1698431365
transform -1 0 21840 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output83 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 4480 0 1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output84
timestamp 1698431365
transform -1 0 4480 0 1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output85
timestamp 1698431365
transform -1 0 38752 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output86
timestamp 1698431365
transform -1 0 4480 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output87
timestamp 1698431365
transform 1 0 32368 0 1 54880
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output88
timestamp 1698431365
transform -1 0 31808 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output89
timestamp 1698431365
transform -1 0 28000 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output90
timestamp 1698431365
transform -1 0 4480 0 -1 15680
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output91
timestamp 1698431365
transform 1 0 28336 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output92
timestamp 1698431365
transform 1 0 55440 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output93
timestamp 1698431365
transform -1 0 34944 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output94
timestamp 1698431365
transform -1 0 4480 0 -1 29792
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output95
timestamp 1698431365
transform 1 0 53312 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output96
timestamp 1698431365
transform 1 0 32368 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output97
timestamp 1698431365
transform 1 0 35840 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output98
timestamp 1698431365
transform -1 0 39984 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output99
timestamp 1698431365
transform 1 0 33040 0 -1 54880
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output100
timestamp 1698431365
transform 1 0 55440 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output101
timestamp 1698431365
transform -1 0 39760 0 1 54880
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output102
timestamp 1698431365
transform -1 0 27216 0 1 54880
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output103
timestamp 1698431365
transform 1 0 55440 0 1 31360
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output104
timestamp 1698431365
transform 1 0 55440 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output105
timestamp 1698431365
transform -1 0 4480 0 1 31360
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output106
timestamp 1698431365
transform 1 0 55440 0 1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output107
timestamp 1698431365
transform 1 0 55440 0 1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output108
timestamp 1698431365
transform -1 0 4480 0 1 29792
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output109
timestamp 1698431365
transform -1 0 28000 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output110
timestamp 1698431365
transform -1 0 4480 0 -1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output111
timestamp 1698431365
transform 1 0 32032 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output112
timestamp 1698431365
transform -1 0 31136 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output113
timestamp 1698431365
transform -1 0 4480 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output114
timestamp 1698431365
transform -1 0 4480 0 -1 34496
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output115
timestamp 1698431365
transform 1 0 55440 0 1 32928
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output116
timestamp 1698431365
transform 1 0 55440 0 1 29792
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  pcpi_exact_mul_118 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20048 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_68 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 58576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_69
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 58576 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_70
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 58576 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_71
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 58576 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_72
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 58576 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_73
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 58576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_74
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 58576 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_75
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 58576 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_76
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 58576 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_77
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 58576 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_78
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 58576 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_79
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 58576 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_80
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 58576 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_81
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 58576 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_82
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 58576 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_83
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 58576 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_84
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 58576 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_85
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 58576 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_86
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 58576 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_87
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 58576 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_88
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 58576 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_89
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 58576 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_90
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 58576 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_91
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 58576 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_92
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 58576 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_93
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 58576 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_94
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 58576 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_95
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 58576 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_96
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 58576 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_97
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 58576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_98
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 58576 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_99
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 58576 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_100
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 58576 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_101
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 58576 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_102
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 58576 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_103
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 58576 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_104
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 58576 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_105
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 58576 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_106
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 58576 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_107
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 58576 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_108
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 58576 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_109
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 58576 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_110
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 58576 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_111
timestamp 1698431365
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698431365
transform -1 0 58576 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_112
timestamp 1698431365
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698431365
transform -1 0 58576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_113
timestamp 1698431365
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698431365
transform -1 0 58576 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_114
timestamp 1698431365
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698431365
transform -1 0 58576 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_115
timestamp 1698431365
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698431365
transform -1 0 58576 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_116
timestamp 1698431365
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698431365
transform -1 0 58576 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_117
timestamp 1698431365
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698431365
transform -1 0 58576 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Left_118
timestamp 1698431365
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1698431365
transform -1 0 58576 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Left_119
timestamp 1698431365
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1698431365
transform -1 0 58576 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Left_120
timestamp 1698431365
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Right_52
timestamp 1698431365
transform -1 0 58576 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Left_121
timestamp 1698431365
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Right_53
timestamp 1698431365
transform -1 0 58576 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Left_122
timestamp 1698431365
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Right_54
timestamp 1698431365
transform -1 0 58576 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Left_123
timestamp 1698431365
transform 1 0 1344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Right_55
timestamp 1698431365
transform -1 0 58576 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Left_124
timestamp 1698431365
transform 1 0 1344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Right_56
timestamp 1698431365
transform -1 0 58576 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Left_125
timestamp 1698431365
transform 1 0 1344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Right_57
timestamp 1698431365
transform -1 0 58576 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Left_126
timestamp 1698431365
transform 1 0 1344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Right_58
timestamp 1698431365
transform -1 0 58576 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Left_127
timestamp 1698431365
transform 1 0 1344 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Right_59
timestamp 1698431365
transform -1 0 58576 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Left_128
timestamp 1698431365
transform 1 0 1344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Right_60
timestamp 1698431365
transform -1 0 58576 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Left_129
timestamp 1698431365
transform 1 0 1344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Right_61
timestamp 1698431365
transform -1 0 58576 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Left_130
timestamp 1698431365
transform 1 0 1344 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Right_62
timestamp 1698431365
transform -1 0 58576 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Left_131
timestamp 1698431365
transform 1 0 1344 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Right_63
timestamp 1698431365
transform -1 0 58576 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Left_132
timestamp 1698431365
transform 1 0 1344 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Right_64
timestamp 1698431365
transform -1 0 58576 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Left_133
timestamp 1698431365
transform 1 0 1344 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Right_65
timestamp 1698431365
transform -1 0 58576 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Left_134
timestamp 1698431365
transform 1 0 1344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Right_66
timestamp 1698431365
transform -1 0 58576 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Left_135
timestamp 1698431365
transform 1 0 1344 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Right_67
timestamp 1698431365
transform -1 0 58576 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_136 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_137
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_138
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_139
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_140
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_141
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_142
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_143
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_144
timestamp 1698431365
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_145
timestamp 1698431365
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_146
timestamp 1698431365
transform 1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_147
timestamp 1698431365
transform 1 0 47040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_148
timestamp 1698431365
transform 1 0 50848 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_149
timestamp 1698431365
transform 1 0 54656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_150
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_151
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_152
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_153
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_154
timestamp 1698431365
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_155
timestamp 1698431365
transform 1 0 48384 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_156
timestamp 1698431365
transform 1 0 56224 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_157
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_158
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_159
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_160
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_161
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_162
timestamp 1698431365
transform 1 0 44464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_163
timestamp 1698431365
transform 1 0 52304 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_164
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_165
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_166
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_167
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_168
timestamp 1698431365
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_169
timestamp 1698431365
transform 1 0 48384 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_170
timestamp 1698431365
transform 1 0 56224 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_171
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_172
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_173
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_174
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_175
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_176
timestamp 1698431365
transform 1 0 44464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_177
timestamp 1698431365
transform 1 0 52304 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_178
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_179
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_180
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_181
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_182
timestamp 1698431365
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_183
timestamp 1698431365
transform 1 0 48384 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_184
timestamp 1698431365
transform 1 0 56224 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_185
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_186
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_187
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_188
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_189
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_190
timestamp 1698431365
transform 1 0 44464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_191
timestamp 1698431365
transform 1 0 52304 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_192
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_193
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_194
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_195
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_196
timestamp 1698431365
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_197
timestamp 1698431365
transform 1 0 48384 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_198
timestamp 1698431365
transform 1 0 56224 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_199
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_200
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_201
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_202
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_203
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_204
timestamp 1698431365
transform 1 0 44464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_205
timestamp 1698431365
transform 1 0 52304 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_206
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_207
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_208
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_209
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_210
timestamp 1698431365
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_211
timestamp 1698431365
transform 1 0 48384 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_212
timestamp 1698431365
transform 1 0 56224 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_213
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_214
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_215
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_216
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_217
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_218
timestamp 1698431365
transform 1 0 44464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_219
timestamp 1698431365
transform 1 0 52304 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_220
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_221
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_222
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_223
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_224
timestamp 1698431365
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_225
timestamp 1698431365
transform 1 0 48384 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_226
timestamp 1698431365
transform 1 0 56224 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_227
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_228
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_229
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_230
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_231
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_232
timestamp 1698431365
transform 1 0 44464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_233
timestamp 1698431365
transform 1 0 52304 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_234
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_235
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_236
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_237
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_238
timestamp 1698431365
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_239
timestamp 1698431365
transform 1 0 48384 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_240
timestamp 1698431365
transform 1 0 56224 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_241
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_242
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_243
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_244
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_245
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_246
timestamp 1698431365
transform 1 0 44464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_247
timestamp 1698431365
transform 1 0 52304 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_248
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_249
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_250
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_251
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_252
timestamp 1698431365
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_253
timestamp 1698431365
transform 1 0 48384 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_254
timestamp 1698431365
transform 1 0 56224 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_255
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_256
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_257
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_258
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_259
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_260
timestamp 1698431365
transform 1 0 44464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_261
timestamp 1698431365
transform 1 0 52304 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_262
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_263
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_264
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_265
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_266
timestamp 1698431365
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_267
timestamp 1698431365
transform 1 0 48384 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_268
timestamp 1698431365
transform 1 0 56224 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_269
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_270
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_271
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_272
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_273
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_274
timestamp 1698431365
transform 1 0 44464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_275
timestamp 1698431365
transform 1 0 52304 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_276
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_277
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_278
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_279
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_280
timestamp 1698431365
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_281
timestamp 1698431365
transform 1 0 48384 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_282
timestamp 1698431365
transform 1 0 56224 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_283
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_284
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_285
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_286
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_287
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_288
timestamp 1698431365
transform 1 0 44464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_289
timestamp 1698431365
transform 1 0 52304 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_290
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_291
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_292
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_293
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_294
timestamp 1698431365
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_295
timestamp 1698431365
transform 1 0 48384 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_296
timestamp 1698431365
transform 1 0 56224 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_297
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_298
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_299
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_300
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_301
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_302
timestamp 1698431365
transform 1 0 44464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_303
timestamp 1698431365
transform 1 0 52304 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_304
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_305
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_306
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_307
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_308
timestamp 1698431365
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_309
timestamp 1698431365
transform 1 0 48384 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_310
timestamp 1698431365
transform 1 0 56224 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_311
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_312
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_313
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_314
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_315
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_316
timestamp 1698431365
transform 1 0 44464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_317
timestamp 1698431365
transform 1 0 52304 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_318
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_319
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_320
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_321
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_322
timestamp 1698431365
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_323
timestamp 1698431365
transform 1 0 48384 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_324
timestamp 1698431365
transform 1 0 56224 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_325
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_326
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_327
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_328
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_329
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_330
timestamp 1698431365
transform 1 0 44464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_331
timestamp 1698431365
transform 1 0 52304 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_332
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_333
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_334
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_335
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_336
timestamp 1698431365
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_337
timestamp 1698431365
transform 1 0 48384 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_338
timestamp 1698431365
transform 1 0 56224 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_339
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_340
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_341
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_342
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_343
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_344
timestamp 1698431365
transform 1 0 44464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_345
timestamp 1698431365
transform 1 0 52304 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_346
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_347
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_348
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_349
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_350
timestamp 1698431365
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_351
timestamp 1698431365
transform 1 0 48384 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_352
timestamp 1698431365
transform 1 0 56224 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_353
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_354
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_355
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_356
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_357
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_358
timestamp 1698431365
transform 1 0 44464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_359
timestamp 1698431365
transform 1 0 52304 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_360
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_361
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_362
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_363
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_364
timestamp 1698431365
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_365
timestamp 1698431365
transform 1 0 48384 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_366
timestamp 1698431365
transform 1 0 56224 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_367
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_368
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_369
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_370
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_371
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_372
timestamp 1698431365
transform 1 0 44464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_373
timestamp 1698431365
transform 1 0 52304 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_374
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_375
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_376
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_377
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_378
timestamp 1698431365
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_379
timestamp 1698431365
transform 1 0 48384 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_380
timestamp 1698431365
transform 1 0 56224 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_381
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_382
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_383
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_384
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_385
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_386
timestamp 1698431365
transform 1 0 44464 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_387
timestamp 1698431365
transform 1 0 52304 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_388
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_389
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_390
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_391
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_392
timestamp 1698431365
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_393
timestamp 1698431365
transform 1 0 48384 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_394
timestamp 1698431365
transform 1 0 56224 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_395
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_396
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_397
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_398
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_399
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_400
timestamp 1698431365
transform 1 0 44464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_401
timestamp 1698431365
transform 1 0 52304 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_402
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_403
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_404
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_405
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_406
timestamp 1698431365
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_407
timestamp 1698431365
transform 1 0 48384 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_408
timestamp 1698431365
transform 1 0 56224 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_409
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_410
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_411
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_412
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_413
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_414
timestamp 1698431365
transform 1 0 44464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_415
timestamp 1698431365
transform 1 0 52304 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_416
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_417
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_418
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_419
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_420
timestamp 1698431365
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_421
timestamp 1698431365
transform 1 0 48384 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_422
timestamp 1698431365
transform 1 0 56224 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_423
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_424
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_425
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_426
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_427
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_428
timestamp 1698431365
transform 1 0 44464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_429
timestamp 1698431365
transform 1 0 52304 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_430
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_431
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_432
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_433
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_434
timestamp 1698431365
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_435
timestamp 1698431365
transform 1 0 48384 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_436
timestamp 1698431365
transform 1 0 56224 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_437
timestamp 1698431365
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_438
timestamp 1698431365
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_439
timestamp 1698431365
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_440
timestamp 1698431365
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_441
timestamp 1698431365
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_442
timestamp 1698431365
transform 1 0 44464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_443
timestamp 1698431365
transform 1 0 52304 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_444
timestamp 1698431365
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_445
timestamp 1698431365
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_446
timestamp 1698431365
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_447
timestamp 1698431365
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_448
timestamp 1698431365
transform 1 0 40544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_449
timestamp 1698431365
transform 1 0 48384 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_450
timestamp 1698431365
transform 1 0 56224 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_451
timestamp 1698431365
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_452
timestamp 1698431365
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_453
timestamp 1698431365
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_454
timestamp 1698431365
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_455
timestamp 1698431365
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_456
timestamp 1698431365
transform 1 0 44464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_457
timestamp 1698431365
transform 1 0 52304 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_458
timestamp 1698431365
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_459
timestamp 1698431365
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_460
timestamp 1698431365
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_461
timestamp 1698431365
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_462
timestamp 1698431365
transform 1 0 40544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_463
timestamp 1698431365
transform 1 0 48384 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_464
timestamp 1698431365
transform 1 0 56224 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_465
timestamp 1698431365
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_466
timestamp 1698431365
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_467
timestamp 1698431365
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_468
timestamp 1698431365
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_469
timestamp 1698431365
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_470
timestamp 1698431365
transform 1 0 44464 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_471
timestamp 1698431365
transform 1 0 52304 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_472
timestamp 1698431365
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_473
timestamp 1698431365
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_474
timestamp 1698431365
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_475
timestamp 1698431365
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_476
timestamp 1698431365
transform 1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_477
timestamp 1698431365
transform 1 0 48384 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_478
timestamp 1698431365
transform 1 0 56224 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_479
timestamp 1698431365
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_480
timestamp 1698431365
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_481
timestamp 1698431365
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_482
timestamp 1698431365
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_483
timestamp 1698431365
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_484
timestamp 1698431365
transform 1 0 44464 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_485
timestamp 1698431365
transform 1 0 52304 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_486
timestamp 1698431365
transform 1 0 9184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_487
timestamp 1698431365
transform 1 0 17024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_488
timestamp 1698431365
transform 1 0 24864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_489
timestamp 1698431365
transform 1 0 32704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_490
timestamp 1698431365
transform 1 0 40544 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_491
timestamp 1698431365
transform 1 0 48384 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_492
timestamp 1698431365
transform 1 0 56224 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_493
timestamp 1698431365
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_494
timestamp 1698431365
transform 1 0 13104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_495
timestamp 1698431365
transform 1 0 20944 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_496
timestamp 1698431365
transform 1 0 28784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_497
timestamp 1698431365
transform 1 0 36624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_498
timestamp 1698431365
transform 1 0 44464 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_499
timestamp 1698431365
transform 1 0 52304 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_500
timestamp 1698431365
transform 1 0 9184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_501
timestamp 1698431365
transform 1 0 17024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_502
timestamp 1698431365
transform 1 0 24864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_503
timestamp 1698431365
transform 1 0 32704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_504
timestamp 1698431365
transform 1 0 40544 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_505
timestamp 1698431365
transform 1 0 48384 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_506
timestamp 1698431365
transform 1 0 56224 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_507
timestamp 1698431365
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_508
timestamp 1698431365
transform 1 0 13104 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_509
timestamp 1698431365
transform 1 0 20944 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_510
timestamp 1698431365
transform 1 0 28784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_511
timestamp 1698431365
transform 1 0 36624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_512
timestamp 1698431365
transform 1 0 44464 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_513
timestamp 1698431365
transform 1 0 52304 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_514
timestamp 1698431365
transform 1 0 9184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_515
timestamp 1698431365
transform 1 0 17024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_516
timestamp 1698431365
transform 1 0 24864 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_517
timestamp 1698431365
transform 1 0 32704 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_518
timestamp 1698431365
transform 1 0 40544 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_519
timestamp 1698431365
transform 1 0 48384 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_520
timestamp 1698431365
transform 1 0 56224 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_521
timestamp 1698431365
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_522
timestamp 1698431365
transform 1 0 13104 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_523
timestamp 1698431365
transform 1 0 20944 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_524
timestamp 1698431365
transform 1 0 28784 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_525
timestamp 1698431365
transform 1 0 36624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_526
timestamp 1698431365
transform 1 0 44464 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_527
timestamp 1698431365
transform 1 0 52304 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_528
timestamp 1698431365
transform 1 0 9184 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_529
timestamp 1698431365
transform 1 0 17024 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_530
timestamp 1698431365
transform 1 0 24864 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_531
timestamp 1698431365
transform 1 0 32704 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_532
timestamp 1698431365
transform 1 0 40544 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_533
timestamp 1698431365
transform 1 0 48384 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_534
timestamp 1698431365
transform 1 0 56224 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_535
timestamp 1698431365
transform 1 0 5264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_536
timestamp 1698431365
transform 1 0 13104 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_537
timestamp 1698431365
transform 1 0 20944 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_538
timestamp 1698431365
transform 1 0 28784 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_539
timestamp 1698431365
transform 1 0 36624 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_540
timestamp 1698431365
transform 1 0 44464 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_541
timestamp 1698431365
transform 1 0 52304 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_542
timestamp 1698431365
transform 1 0 9184 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_543
timestamp 1698431365
transform 1 0 17024 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_544
timestamp 1698431365
transform 1 0 24864 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_545
timestamp 1698431365
transform 1 0 32704 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_546
timestamp 1698431365
transform 1 0 40544 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_547
timestamp 1698431365
transform 1 0 48384 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_548
timestamp 1698431365
transform 1 0 56224 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_549
timestamp 1698431365
transform 1 0 5264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_550
timestamp 1698431365
transform 1 0 13104 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_551
timestamp 1698431365
transform 1 0 20944 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_552
timestamp 1698431365
transform 1 0 28784 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_553
timestamp 1698431365
transform 1 0 36624 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_554
timestamp 1698431365
transform 1 0 44464 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_555
timestamp 1698431365
transform 1 0 52304 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_556
timestamp 1698431365
transform 1 0 9184 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_557
timestamp 1698431365
transform 1 0 17024 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_558
timestamp 1698431365
transform 1 0 24864 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_559
timestamp 1698431365
transform 1 0 32704 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_560
timestamp 1698431365
transform 1 0 40544 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_561
timestamp 1698431365
transform 1 0 48384 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_562
timestamp 1698431365
transform 1 0 56224 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_563
timestamp 1698431365
transform 1 0 5264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_564
timestamp 1698431365
transform 1 0 13104 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_565
timestamp 1698431365
transform 1 0 20944 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_566
timestamp 1698431365
transform 1 0 28784 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_567
timestamp 1698431365
transform 1 0 36624 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_568
timestamp 1698431365
transform 1 0 44464 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_569
timestamp 1698431365
transform 1 0 52304 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_570
timestamp 1698431365
transform 1 0 9184 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_571
timestamp 1698431365
transform 1 0 17024 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_572
timestamp 1698431365
transform 1 0 24864 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_573
timestamp 1698431365
transform 1 0 32704 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_574
timestamp 1698431365
transform 1 0 40544 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_575
timestamp 1698431365
transform 1 0 48384 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_576
timestamp 1698431365
transform 1 0 56224 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_577
timestamp 1698431365
transform 1 0 5264 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_578
timestamp 1698431365
transform 1 0 13104 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_579
timestamp 1698431365
transform 1 0 20944 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_580
timestamp 1698431365
transform 1 0 28784 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_581
timestamp 1698431365
transform 1 0 36624 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_582
timestamp 1698431365
transform 1 0 44464 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_583
timestamp 1698431365
transform 1 0 52304 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_584
timestamp 1698431365
transform 1 0 9184 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_585
timestamp 1698431365
transform 1 0 17024 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_586
timestamp 1698431365
transform 1 0 24864 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_587
timestamp 1698431365
transform 1 0 32704 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_588
timestamp 1698431365
transform 1 0 40544 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_589
timestamp 1698431365
transform 1 0 48384 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_590
timestamp 1698431365
transform 1 0 56224 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_591
timestamp 1698431365
transform 1 0 5264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_592
timestamp 1698431365
transform 1 0 13104 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_593
timestamp 1698431365
transform 1 0 20944 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_594
timestamp 1698431365
transform 1 0 28784 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_595
timestamp 1698431365
transform 1 0 36624 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_596
timestamp 1698431365
transform 1 0 44464 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_597
timestamp 1698431365
transform 1 0 52304 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_598
timestamp 1698431365
transform 1 0 9184 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_599
timestamp 1698431365
transform 1 0 17024 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_600
timestamp 1698431365
transform 1 0 24864 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_601
timestamp 1698431365
transform 1 0 32704 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_602
timestamp 1698431365
transform 1 0 40544 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_603
timestamp 1698431365
transform 1 0 48384 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_604
timestamp 1698431365
transform 1 0 56224 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_605
timestamp 1698431365
transform 1 0 5264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_606
timestamp 1698431365
transform 1 0 13104 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_607
timestamp 1698431365
transform 1 0 20944 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_608
timestamp 1698431365
transform 1 0 28784 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_609
timestamp 1698431365
transform 1 0 36624 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_610
timestamp 1698431365
transform 1 0 44464 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_611
timestamp 1698431365
transform 1 0 52304 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_612
timestamp 1698431365
transform 1 0 5152 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_613
timestamp 1698431365
transform 1 0 8960 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_614
timestamp 1698431365
transform 1 0 12768 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_615
timestamp 1698431365
transform 1 0 16576 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_616
timestamp 1698431365
transform 1 0 20384 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_617
timestamp 1698431365
transform 1 0 24192 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_618
timestamp 1698431365
transform 1 0 28000 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_619
timestamp 1698431365
transform 1 0 31808 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_620
timestamp 1698431365
transform 1 0 35616 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_621
timestamp 1698431365
transform 1 0 39424 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_622
timestamp 1698431365
transform 1 0 43232 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_623
timestamp 1698431365
transform 1 0 47040 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_624
timestamp 1698431365
transform 1 0 50848 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_625
timestamp 1698431365
transform 1 0 54656 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  wire1
timestamp 1698431365
transform 1 0 19712 0 1 39200
box -86 -86 758 870
<< labels >>
flabel metal3 s 0 43008 800 43120 0 FreeSans 448 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 0 10752 800 10864 0 FreeSans 448 0 0 0 pcpi_insn[0]
port 1 nsew signal input
flabel metal2 s 0 0 112 800 0 FreeSans 448 90 0 0 pcpi_insn[10]
port 2 nsew signal input
flabel metal2 s 672 0 784 800 0 FreeSans 448 90 0 0 pcpi_insn[11]
port 3 nsew signal input
flabel metal2 s 24864 59200 24976 60000 0 FreeSans 448 90 0 0 pcpi_insn[12]
port 4 nsew signal input
flabel metal2 s 26208 59200 26320 60000 0 FreeSans 448 90 0 0 pcpi_insn[13]
port 5 nsew signal input
flabel metal2 s 28224 59200 28336 60000 0 FreeSans 448 90 0 0 pcpi_insn[14]
port 6 nsew signal input
flabel metal2 s 1344 0 1456 800 0 FreeSans 448 90 0 0 pcpi_insn[15]
port 7 nsew signal input
flabel metal2 s 2016 0 2128 800 0 FreeSans 448 90 0 0 pcpi_insn[16]
port 8 nsew signal input
flabel metal2 s 2688 0 2800 800 0 FreeSans 448 90 0 0 pcpi_insn[17]
port 9 nsew signal input
flabel metal2 s 3360 0 3472 800 0 FreeSans 448 90 0 0 pcpi_insn[18]
port 10 nsew signal input
flabel metal2 s 4032 0 4144 800 0 FreeSans 448 90 0 0 pcpi_insn[19]
port 11 nsew signal input
flabel metal3 s 0 26880 800 26992 0 FreeSans 448 0 0 0 pcpi_insn[1]
port 12 nsew signal input
flabel metal2 s 4704 0 4816 800 0 FreeSans 448 90 0 0 pcpi_insn[20]
port 13 nsew signal input
flabel metal2 s 5376 0 5488 800 0 FreeSans 448 90 0 0 pcpi_insn[21]
port 14 nsew signal input
flabel metal2 s 6048 0 6160 800 0 FreeSans 448 90 0 0 pcpi_insn[22]
port 15 nsew signal input
flabel metal2 s 6720 0 6832 800 0 FreeSans 448 90 0 0 pcpi_insn[23]
port 16 nsew signal input
flabel metal2 s 7392 0 7504 800 0 FreeSans 448 90 0 0 pcpi_insn[24]
port 17 nsew signal input
flabel metal3 s 0 28224 800 28336 0 FreeSans 448 0 0 0 pcpi_insn[25]
port 18 nsew signal input
flabel metal3 s 0 30240 800 30352 0 FreeSans 448 0 0 0 pcpi_insn[26]
port 19 nsew signal input
flabel metal3 s 0 26208 800 26320 0 FreeSans 448 0 0 0 pcpi_insn[27]
port 20 nsew signal input
flabel metal3 s 0 43680 800 43792 0 FreeSans 448 0 0 0 pcpi_insn[28]
port 21 nsew signal input
flabel metal3 s 0 27552 800 27664 0 FreeSans 448 0 0 0 pcpi_insn[29]
port 22 nsew signal input
flabel metal3 s 0 11424 800 11536 0 FreeSans 448 0 0 0 pcpi_insn[2]
port 23 nsew signal input
flabel metal3 s 0 21504 800 21616 0 FreeSans 448 0 0 0 pcpi_insn[30]
port 24 nsew signal input
flabel metal3 s 0 25536 800 25648 0 FreeSans 448 0 0 0 pcpi_insn[31]
port 25 nsew signal input
flabel metal3 s 0 12096 800 12208 0 FreeSans 448 0 0 0 pcpi_insn[3]
port 26 nsew signal input
flabel metal3 s 0 17472 800 17584 0 FreeSans 448 0 0 0 pcpi_insn[4]
port 27 nsew signal input
flabel metal3 s 0 24192 800 24304 0 FreeSans 448 0 0 0 pcpi_insn[5]
port 28 nsew signal input
flabel metal3 s 0 20160 800 20272 0 FreeSans 448 0 0 0 pcpi_insn[6]
port 29 nsew signal input
flabel metal2 s 8064 0 8176 800 0 FreeSans 448 90 0 0 pcpi_insn[7]
port 30 nsew signal input
flabel metal2 s 8736 0 8848 800 0 FreeSans 448 90 0 0 pcpi_insn[8]
port 31 nsew signal input
flabel metal2 s 9408 0 9520 800 0 FreeSans 448 90 0 0 pcpi_insn[9]
port 32 nsew signal input
flabel metal3 s 0 40320 800 40432 0 FreeSans 448 0 0 0 pcpi_rd[0]
port 33 nsew signal tristate
flabel metal3 s 0 42336 800 42448 0 FreeSans 448 0 0 0 pcpi_rd[10]
port 34 nsew signal tristate
flabel metal2 s 34272 59200 34384 60000 0 FreeSans 448 90 0 0 pcpi_rd[11]
port 35 nsew signal tristate
flabel metal3 s 0 24864 800 24976 0 FreeSans 448 0 0 0 pcpi_rd[12]
port 36 nsew signal tristate
flabel metal2 s 32256 59200 32368 60000 0 FreeSans 448 90 0 0 pcpi_rd[13]
port 37 nsew signal tristate
flabel metal2 s 28896 0 29008 800 0 FreeSans 448 90 0 0 pcpi_rd[14]
port 38 nsew signal tristate
flabel metal2 s 26880 0 26992 800 0 FreeSans 448 90 0 0 pcpi_rd[15]
port 39 nsew signal tristate
flabel metal3 s 0 14784 800 14896 0 FreeSans 448 0 0 0 pcpi_rd[16]
port 40 nsew signal tristate
flabel metal2 s 28224 0 28336 800 0 FreeSans 448 90 0 0 pcpi_rd[17]
port 41 nsew signal tristate
flabel metal3 s 59200 24864 60000 24976 0 FreeSans 448 0 0 0 pcpi_rd[18]
port 42 nsew signal tristate
flabel metal2 s 30240 0 30352 800 0 FreeSans 448 90 0 0 pcpi_rd[19]
port 43 nsew signal tristate
flabel metal3 s 0 28896 800 29008 0 FreeSans 448 0 0 0 pcpi_rd[1]
port 44 nsew signal tristate
flabel metal3 s 59200 24192 60000 24304 0 FreeSans 448 0 0 0 pcpi_rd[20]
port 45 nsew signal tristate
flabel metal2 s 32256 0 32368 800 0 FreeSans 448 90 0 0 pcpi_rd[21]
port 46 nsew signal tristate
flabel metal2 s 35616 0 35728 800 0 FreeSans 448 90 0 0 pcpi_rd[22]
port 47 nsew signal tristate
flabel metal2 s 36960 0 37072 800 0 FreeSans 448 90 0 0 pcpi_rd[23]
port 48 nsew signal tristate
flabel metal2 s 32928 59200 33040 60000 0 FreeSans 448 90 0 0 pcpi_rd[24]
port 49 nsew signal tristate
flabel metal3 s 59200 35616 60000 35728 0 FreeSans 448 0 0 0 pcpi_rd[25]
port 50 nsew signal tristate
flabel metal2 s 35616 59200 35728 60000 0 FreeSans 448 90 0 0 pcpi_rd[26]
port 51 nsew signal tristate
flabel metal2 s 24192 59200 24304 60000 0 FreeSans 448 90 0 0 pcpi_rd[27]
port 52 nsew signal tristate
flabel metal3 s 59200 32256 60000 32368 0 FreeSans 448 0 0 0 pcpi_rd[28]
port 53 nsew signal tristate
flabel metal3 s 59200 26880 60000 26992 0 FreeSans 448 0 0 0 pcpi_rd[29]
port 54 nsew signal tristate
flabel metal3 s 0 30912 800 31024 0 FreeSans 448 0 0 0 pcpi_rd[2]
port 55 nsew signal tristate
flabel metal3 s 59200 28224 60000 28336 0 FreeSans 448 0 0 0 pcpi_rd[30]
port 56 nsew signal tristate
flabel metal3 s 59200 27552 60000 27664 0 FreeSans 448 0 0 0 pcpi_rd[31]
port 57 nsew signal tristate
flabel metal3 s 0 29568 800 29680 0 FreeSans 448 0 0 0 pcpi_rd[3]
port 58 nsew signal tristate
flabel metal2 s 25536 59200 25648 60000 0 FreeSans 448 90 0 0 pcpi_rd[4]
port 59 nsew signal tristate
flabel metal3 s 0 39648 800 39760 0 FreeSans 448 0 0 0 pcpi_rd[5]
port 60 nsew signal tristate
flabel metal2 s 31584 59200 31696 60000 0 FreeSans 448 90 0 0 pcpi_rd[6]
port 61 nsew signal tristate
flabel metal2 s 27552 59200 27664 60000 0 FreeSans 448 90 0 0 pcpi_rd[7]
port 62 nsew signal tristate
flabel metal3 s 0 36960 800 37072 0 FreeSans 448 0 0 0 pcpi_rd[8]
port 63 nsew signal tristate
flabel metal3 s 0 33600 800 33712 0 FreeSans 448 0 0 0 pcpi_rd[9]
port 64 nsew signal tristate
flabel metal3 s 59200 30912 60000 31024 0 FreeSans 448 0 0 0 pcpi_ready
port 65 nsew signal tristate
flabel metal3 s 0 32928 800 33040 0 FreeSans 448 0 0 0 pcpi_rs1[0]
port 66 nsew signal input
flabel metal2 s 34272 0 34384 800 0 FreeSans 448 90 0 0 pcpi_rs1[10]
port 67 nsew signal input
flabel metal2 s 34944 0 35056 800 0 FreeSans 448 90 0 0 pcpi_rs1[11]
port 68 nsew signal input
flabel metal2 s 39648 0 39760 800 0 FreeSans 448 90 0 0 pcpi_rs1[12]
port 69 nsew signal input
flabel metal2 s 43008 0 43120 800 0 FreeSans 448 90 0 0 pcpi_rs1[13]
port 70 nsew signal input
flabel metal2 s 47040 0 47152 800 0 FreeSans 448 90 0 0 pcpi_rs1[14]
port 71 nsew signal input
flabel metal2 s 49728 0 49840 800 0 FreeSans 448 90 0 0 pcpi_rs1[15]
port 72 nsew signal input
flabel metal3 s 0 16800 800 16912 0 FreeSans 448 0 0 0 pcpi_rs1[16]
port 73 nsew signal input
flabel metal3 s 0 18144 800 18256 0 FreeSans 448 0 0 0 pcpi_rs1[17]
port 74 nsew signal input
flabel metal3 s 0 12768 800 12880 0 FreeSans 448 0 0 0 pcpi_rs1[18]
port 75 nsew signal input
flabel metal3 s 0 14112 800 14224 0 FreeSans 448 0 0 0 pcpi_rs1[19]
port 76 nsew signal input
flabel metal3 s 0 37632 800 37744 0 FreeSans 448 0 0 0 pcpi_rs1[1]
port 77 nsew signal input
flabel metal3 s 0 13440 800 13552 0 FreeSans 448 0 0 0 pcpi_rs1[20]
port 78 nsew signal input
flabel metal3 s 0 15456 800 15568 0 FreeSans 448 0 0 0 pcpi_rs1[21]
port 79 nsew signal input
flabel metal3 s 0 10080 800 10192 0 FreeSans 448 0 0 0 pcpi_rs1[22]
port 80 nsew signal input
flabel metal3 s 0 8736 800 8848 0 FreeSans 448 0 0 0 pcpi_rs1[23]
port 81 nsew signal input
flabel metal2 s 28896 59200 29008 60000 0 FreeSans 448 90 0 0 pcpi_rs1[24]
port 82 nsew signal input
flabel metal2 s 29568 59200 29680 60000 0 FreeSans 448 90 0 0 pcpi_rs1[25]
port 83 nsew signal input
flabel metal2 s 30240 59200 30352 60000 0 FreeSans 448 90 0 0 pcpi_rs1[26]
port 84 nsew signal input
flabel metal2 s 38304 59200 38416 60000 0 FreeSans 448 90 0 0 pcpi_rs1[27]
port 85 nsew signal input
flabel metal2 s 36960 59200 37072 60000 0 FreeSans 448 90 0 0 pcpi_rs1[28]
port 86 nsew signal input
flabel metal2 s 37632 59200 37744 60000 0 FreeSans 448 90 0 0 pcpi_rs1[29]
port 87 nsew signal input
flabel metal3 s 0 32256 800 32368 0 FreeSans 448 0 0 0 pcpi_rs1[2]
port 88 nsew signal input
flabel metal2 s 49728 59200 49840 60000 0 FreeSans 448 90 0 0 pcpi_rs1[30]
port 89 nsew signal input
flabel metal2 s 50400 59200 50512 60000 0 FreeSans 448 90 0 0 pcpi_rs1[31]
port 90 nsew signal input
flabel metal3 s 0 35616 800 35728 0 FreeSans 448 0 0 0 pcpi_rs1[3]
port 91 nsew signal input
flabel metal3 s 0 40992 800 41104 0 FreeSans 448 0 0 0 pcpi_rs1[4]
port 92 nsew signal input
flabel metal3 s 0 45024 800 45136 0 FreeSans 448 0 0 0 pcpi_rs1[5]
port 93 nsew signal input
flabel metal3 s 0 44352 800 44464 0 FreeSans 448 0 0 0 pcpi_rs1[6]
port 94 nsew signal input
flabel metal3 s 0 50400 800 50512 0 FreeSans 448 0 0 0 pcpi_rs1[7]
port 95 nsew signal input
flabel metal2 s 33600 0 33712 800 0 FreeSans 448 90 0 0 pcpi_rs1[8]
port 96 nsew signal input
flabel metal2 s 30912 0 31024 800 0 FreeSans 448 90 0 0 pcpi_rs1[9]
port 97 nsew signal input
flabel metal3 s 0 34944 800 35056 0 FreeSans 448 0 0 0 pcpi_rs2[0]
port 98 nsew signal input
flabel metal2 s 36288 0 36400 800 0 FreeSans 448 90 0 0 pcpi_rs2[10]
port 99 nsew signal input
flabel metal2 s 37632 0 37744 800 0 FreeSans 448 90 0 0 pcpi_rs2[11]
port 100 nsew signal input
flabel metal2 s 38976 0 39088 800 0 FreeSans 448 90 0 0 pcpi_rs2[12]
port 101 nsew signal input
flabel metal2 s 38304 0 38416 800 0 FreeSans 448 90 0 0 pcpi_rs2[13]
port 102 nsew signal input
flabel metal3 s 59200 21504 60000 21616 0 FreeSans 448 0 0 0 pcpi_rs2[14]
port 103 nsew signal input
flabel metal3 s 59200 23520 60000 23632 0 FreeSans 448 0 0 0 pcpi_rs2[15]
port 104 nsew signal input
flabel metal3 s 0 22848 800 22960 0 FreeSans 448 0 0 0 pcpi_rs2[16]
port 105 nsew signal input
flabel metal3 s 0 19488 800 19600 0 FreeSans 448 0 0 0 pcpi_rs2[17]
port 106 nsew signal input
flabel metal3 s 0 20832 800 20944 0 FreeSans 448 0 0 0 pcpi_rs2[18]
port 107 nsew signal input
flabel metal3 s 0 16128 800 16240 0 FreeSans 448 0 0 0 pcpi_rs2[19]
port 108 nsew signal input
flabel metal3 s 0 31584 800 31696 0 FreeSans 448 0 0 0 pcpi_rs2[1]
port 109 nsew signal input
flabel metal3 s 0 23520 800 23632 0 FreeSans 448 0 0 0 pcpi_rs2[20]
port 110 nsew signal input
flabel metal3 s 0 18816 800 18928 0 FreeSans 448 0 0 0 pcpi_rs2[21]
port 111 nsew signal input
flabel metal2 s 22176 0 22288 800 0 FreeSans 448 90 0 0 pcpi_rs2[22]
port 112 nsew signal input
flabel metal2 s 24864 0 24976 800 0 FreeSans 448 90 0 0 pcpi_rs2[23]
port 113 nsew signal input
flabel metal2 s 26880 59200 26992 60000 0 FreeSans 448 90 0 0 pcpi_rs2[24]
port 114 nsew signal input
flabel metal2 s 30912 59200 31024 60000 0 FreeSans 448 90 0 0 pcpi_rs2[25]
port 115 nsew signal input
flabel metal2 s 33600 59200 33712 60000 0 FreeSans 448 90 0 0 pcpi_rs2[26]
port 116 nsew signal input
flabel metal2 s 36288 59200 36400 60000 0 FreeSans 448 90 0 0 pcpi_rs2[27]
port 117 nsew signal input
flabel metal2 s 34944 59200 35056 60000 0 FreeSans 448 90 0 0 pcpi_rs2[28]
port 118 nsew signal input
flabel metal2 s 40320 59200 40432 60000 0 FreeSans 448 90 0 0 pcpi_rs2[29]
port 119 nsew signal input
flabel metal3 s 0 36288 800 36400 0 FreeSans 448 0 0 0 pcpi_rs2[2]
port 120 nsew signal input
flabel metal3 s 59200 36960 60000 37072 0 FreeSans 448 0 0 0 pcpi_rs2[30]
port 121 nsew signal input
flabel metal3 s 59200 34944 60000 35056 0 FreeSans 448 0 0 0 pcpi_rs2[31]
port 122 nsew signal input
flabel metal3 s 0 34272 800 34384 0 FreeSans 448 0 0 0 pcpi_rs2[3]
port 123 nsew signal input
flabel metal3 s 0 38304 800 38416 0 FreeSans 448 0 0 0 pcpi_rs2[4]
port 124 nsew signal input
flabel metal3 s 0 41664 800 41776 0 FreeSans 448 0 0 0 pcpi_rs2[5]
port 125 nsew signal input
flabel metal3 s 0 38976 800 39088 0 FreeSans 448 0 0 0 pcpi_rs2[6]
port 126 nsew signal input
flabel metal2 s 23520 59200 23632 60000 0 FreeSans 448 90 0 0 pcpi_rs2[7]
port 127 nsew signal input
flabel metal2 s 32928 0 33040 800 0 FreeSans 448 90 0 0 pcpi_rs2[8]
port 128 nsew signal input
flabel metal2 s 31584 0 31696 800 0 FreeSans 448 90 0 0 pcpi_rs2[9]
port 129 nsew signal input
flabel metal3 s 0 22176 800 22288 0 FreeSans 448 0 0 0 pcpi_valid
port 130 nsew signal input
flabel metal2 s 19488 0 19600 800 0 FreeSans 448 90 0 0 pcpi_wait
port 131 nsew signal tristate
flabel metal3 s 59200 31584 60000 31696 0 FreeSans 448 0 0 0 pcpi_wr
port 132 nsew signal tristate
flabel metal2 s 10080 0 10192 800 0 FreeSans 448 90 0 0 resetn
port 133 nsew signal input
flabel metal4 s 4448 3076 4768 56508 0 FreeSans 1280 90 0 0 vdd
port 134 nsew power bidirectional
flabel metal4 s 35168 3076 35488 56508 0 FreeSans 1280 90 0 0 vdd
port 134 nsew power bidirectional
flabel metal4 s 19808 3076 20128 56508 0 FreeSans 1280 90 0 0 vss
port 135 nsew ground bidirectional
flabel metal4 s 50528 3076 50848 56508 0 FreeSans 1280 90 0 0 vss
port 135 nsew ground bidirectional
rlabel metal1 29960 55664 29960 55664 0 vdd
rlabel metal1 29960 56448 29960 56448 0 vss
rlabel metal2 15400 30576 15400 30576 0 _0000_
rlabel metal3 16968 27160 16968 27160 0 _0001_
rlabel metal2 18536 30464 18536 30464 0 _0002_
rlabel metal2 14616 29120 14616 29120 0 _0003_
rlabel metal2 26152 34440 26152 34440 0 _0004_
rlabel metal3 20328 34216 20328 34216 0 _0005_
rlabel metal2 29288 36848 29288 36848 0 _0006_
rlabel metal2 26488 36904 26488 36904 0 _0007_
rlabel metal2 25144 34048 25144 34048 0 _0008_
rlabel metal2 23912 32200 23912 32200 0 _0009_
rlabel metal2 23688 29848 23688 29848 0 _0010_
rlabel metal2 32200 36120 32200 36120 0 _0011_
rlabel metal3 25816 27160 25816 27160 0 _0012_
rlabel metal3 28168 40488 28168 40488 0 _0013_
rlabel metal2 27720 27440 27720 27440 0 _0014_
rlabel metal2 24920 25872 24920 25872 0 _0015_
rlabel metal2 22960 26152 22960 26152 0 _0016_
rlabel metal2 26264 23576 26264 23576 0 _0017_
rlabel metal2 37128 24360 37128 24360 0 _0018_
rlabel metal2 30016 25592 30016 25592 0 _0019_
rlabel metal2 36064 23240 36064 23240 0 _0020_
rlabel metal2 30296 21896 30296 21896 0 _0021_
rlabel metal2 33656 20944 33656 20944 0 _0022_
rlabel metal2 35112 20104 35112 20104 0 _0023_
rlabel metal2 30408 40712 30408 40712 0 _0024_
rlabel metal2 36008 35336 36008 35336 0 _0025_
rlabel metal2 33096 38192 33096 38192 0 _0026_
rlabel metal2 30072 34272 30072 34272 0 _0027_
rlabel metal2 38472 31192 38472 31192 0 _0028_
rlabel metal2 37800 27216 37800 27216 0 _0029_
rlabel metal2 41720 28000 41720 28000 0 _0030_
rlabel metal2 41048 27440 41048 27440 0 _0031_
rlabel metal2 26768 26824 26768 26824 0 _0032_
rlabel metal2 27720 26320 27720 26320 0 _0033_
rlabel metal2 25984 27048 25984 27048 0 _0034_
rlabel metal2 50064 26488 50064 26488 0 _0035_
rlabel metal2 50344 28224 50344 28224 0 _0036_
rlabel metal2 51912 26040 51912 26040 0 _0037_
rlabel metal2 57288 21224 57288 21224 0 _0038_
rlabel metal2 56840 21896 56840 21896 0 _0039_
rlabel metal2 56616 24248 56616 24248 0 _0040_
rlabel metal2 54824 24920 54824 24920 0 _0041_
rlabel metal2 53592 25872 53592 25872 0 _0042_
rlabel metal2 54600 25592 54600 25592 0 _0043_
rlabel metal2 55608 21672 55608 21672 0 _0044_
rlabel metal2 55048 25536 55048 25536 0 _0045_
rlabel metal2 54656 26152 54656 26152 0 _0046_
rlabel metal3 53088 26376 53088 26376 0 _0047_
rlabel metal2 51016 28224 51016 28224 0 _0048_
rlabel metal2 49784 28784 49784 28784 0 _0049_
rlabel metal3 35896 23128 35896 23128 0 _0050_
rlabel metal2 15176 26656 15176 26656 0 _0051_
rlabel metal2 31416 34272 31416 34272 0 _0052_
rlabel metal2 30968 39060 30968 39060 0 _0053_
rlabel metal2 29848 40432 29848 40432 0 _0054_
rlabel metal2 52472 26264 52472 26264 0 _0055_
rlabel metal3 55272 26488 55272 26488 0 _0056_
rlabel metal2 52696 26488 52696 26488 0 _0057_
rlabel metal2 53256 28056 53256 28056 0 _0058_
rlabel metal2 51800 27832 51800 27832 0 _0059_
rlabel metal2 52136 27776 52136 27776 0 _0060_
rlabel metal3 41104 28504 41104 28504 0 _0061_
rlabel metal3 37016 22344 37016 22344 0 _0062_
rlabel metal3 34216 22120 34216 22120 0 _0063_
rlabel metal3 30856 26824 30856 26824 0 _0064_
rlabel metal3 27664 27048 27664 27048 0 _0065_
rlabel metal2 28280 27944 28280 27944 0 _0066_
rlabel metal2 52584 27160 52584 27160 0 _0067_
rlabel metal2 40376 28280 40376 28280 0 _0068_
rlabel metal3 36456 23856 36456 23856 0 _0069_
rlabel metal2 35784 26040 35784 26040 0 _0070_
rlabel metal4 26488 27888 26488 27888 0 _0071_
rlabel metal2 27216 24920 27216 24920 0 _0072_
rlabel metal2 13720 23856 13720 23856 0 _0073_
rlabel metal3 19096 23688 19096 23688 0 _0074_
rlabel metal2 26376 22288 26376 22288 0 _0075_
rlabel metal3 26096 20104 26096 20104 0 _0076_
rlabel metal2 22624 22568 22624 22568 0 _0077_
rlabel metal2 18760 19152 18760 19152 0 _0078_
rlabel metal3 20440 23912 20440 23912 0 _0079_
rlabel metal2 16744 23464 16744 23464 0 _0080_
rlabel metal2 18592 25368 18592 25368 0 _0081_
rlabel metal3 13104 23352 13104 23352 0 _0082_
rlabel metal2 12936 25648 12936 25648 0 _0083_
rlabel metal2 3416 24304 3416 24304 0 _0084_
rlabel metal2 5992 25424 5992 25424 0 _0085_
rlabel metal2 2296 20832 2296 20832 0 _0086_
rlabel metal2 4760 24752 4760 24752 0 _0087_
rlabel metal2 2632 22288 2632 22288 0 _0088_
rlabel metal4 4872 19040 4872 19040 0 _0089_
rlabel metal2 3304 19376 3304 19376 0 _0090_
rlabel metal2 4872 20496 4872 20496 0 _0091_
rlabel metal2 3416 19600 3416 19600 0 _0092_
rlabel metal2 5096 22064 5096 22064 0 _0093_
rlabel metal2 4928 20888 4928 20888 0 _0094_
rlabel metal3 8176 25368 8176 25368 0 _0095_
rlabel metal2 6328 25088 6328 25088 0 _0096_
rlabel metal3 9464 25480 9464 25480 0 _0097_
rlabel metal2 7784 23352 7784 23352 0 _0098_
rlabel metal3 10696 25200 10696 25200 0 _0099_
rlabel metal2 11144 26320 11144 26320 0 _0100_
rlabel metal2 6328 26040 6328 26040 0 _0101_
rlabel metal3 10024 23912 10024 23912 0 _0102_
rlabel metal4 3304 21448 3304 21448 0 _0103_
rlabel metal2 3752 22736 3752 22736 0 _0104_
rlabel metal2 6888 20888 6888 20888 0 _0105_
rlabel metal2 7224 25032 7224 25032 0 _0106_
rlabel metal2 11480 26096 11480 26096 0 _0107_
rlabel metal3 11984 26264 11984 26264 0 _0108_
rlabel metal2 14056 24248 14056 24248 0 _0109_
rlabel metal3 19712 20104 19712 20104 0 _0110_
rlabel metal3 11984 23128 11984 23128 0 _0111_
rlabel metal2 4312 22344 4312 22344 0 _0112_
rlabel metal2 4536 22008 4536 22008 0 _0113_
rlabel metal2 7224 21280 7224 21280 0 _0114_
rlabel metal2 23688 24528 23688 24528 0 _0115_
rlabel metal3 9464 24696 9464 24696 0 _0116_
rlabel metal2 10808 24920 10808 24920 0 _0117_
rlabel metal2 10752 24024 10752 24024 0 _0118_
rlabel metal2 6664 22568 6664 22568 0 _0119_
rlabel metal2 6776 21280 6776 21280 0 _0120_
rlabel metal2 3640 18760 3640 18760 0 _0121_
rlabel metal2 3976 19880 3976 19880 0 _0122_
rlabel metal2 5992 20440 5992 20440 0 _0123_
rlabel metal2 10136 22848 10136 22848 0 _0124_
rlabel metal3 13440 24024 13440 24024 0 _0125_
rlabel metal2 18312 25872 18312 25872 0 _0126_
rlabel metal2 18088 24248 18088 24248 0 _0127_
rlabel metal2 15512 24360 15512 24360 0 _0128_
rlabel metal2 12040 24024 12040 24024 0 _0129_
rlabel metal2 12488 24696 12488 24696 0 _0130_
rlabel metal2 15624 24304 15624 24304 0 _0131_
rlabel metal3 9408 20664 9408 20664 0 _0132_
rlabel metal2 10920 21056 10920 21056 0 _0133_
rlabel metal2 8120 15848 8120 15848 0 _0134_
rlabel metal3 6608 20776 6608 20776 0 _0135_
rlabel metal2 6328 20328 6328 20328 0 _0136_
rlabel metal2 7560 19992 7560 19992 0 _0137_
rlabel metal2 8512 20776 8512 20776 0 _0138_
rlabel metal2 9128 22456 9128 22456 0 _0139_
rlabel metal3 11088 22344 11088 22344 0 _0140_
rlabel metal2 7784 17192 7784 17192 0 _0141_
rlabel metal2 9464 17920 9464 17920 0 _0142_
rlabel metal3 5096 16072 5096 16072 0 _0143_
rlabel metal2 5040 15960 5040 15960 0 _0144_
rlabel metal2 3192 16072 3192 16072 0 _0145_
rlabel metal2 5824 16296 5824 16296 0 _0146_
rlabel metal3 5432 18312 5432 18312 0 _0147_
rlabel metal2 4984 19264 4984 19264 0 _0148_
rlabel metal3 6832 18424 6832 18424 0 _0149_
rlabel metal2 11592 20384 11592 20384 0 _0150_
rlabel metal2 15400 23856 15400 23856 0 _0151_
rlabel metal3 19152 24584 19152 24584 0 _0152_
rlabel metal2 20384 24696 20384 24696 0 _0153_
rlabel metal2 20888 22456 20888 22456 0 _0154_
rlabel metal2 19656 20160 19656 20160 0 _0155_
rlabel metal2 16632 25760 16632 25760 0 _0156_
rlabel metal2 16296 25088 16296 25088 0 _0157_
rlabel metal2 17136 24696 17136 24696 0 _0158_
rlabel metal2 18256 23128 18256 23128 0 _0159_
rlabel metal2 16632 18928 16632 18928 0 _0160_
rlabel metal2 17080 19376 17080 19376 0 _0161_
rlabel metal2 13720 18144 13720 18144 0 _0162_
rlabel metal3 9184 26264 9184 26264 0 _0163_
rlabel metal2 7784 23912 7784 23912 0 _0164_
rlabel metal2 7560 24192 7560 24192 0 _0165_
rlabel metal2 7952 23688 7952 23688 0 _0166_
rlabel metal2 10360 22680 10360 22680 0 _0167_
rlabel metal2 9912 20944 9912 20944 0 _0168_
rlabel metal2 9128 21224 9128 21224 0 _0169_
rlabel metal2 10472 20720 10472 20720 0 _0170_
rlabel metal3 12936 18424 12936 18424 0 _0171_
rlabel metal3 12936 20104 12936 20104 0 _0172_
rlabel metal2 12936 19600 12936 19600 0 _0173_
rlabel via2 14056 20664 14056 20664 0 _0174_
rlabel metal3 11592 18536 11592 18536 0 _0175_
rlabel metal3 5096 15512 5096 15512 0 _0176_
rlabel metal2 9240 17528 9240 17528 0 _0177_
rlabel metal3 7616 19208 7616 19208 0 _0178_
rlabel metal2 9576 18928 9576 18928 0 _0179_
rlabel metal2 10360 18032 10360 18032 0 _0180_
rlabel metal2 6552 15624 6552 15624 0 _0181_
rlabel metal2 23352 21336 23352 21336 0 _0182_
rlabel metal2 5992 12096 5992 12096 0 _0183_
rlabel metal3 6608 12152 6608 12152 0 _0184_
rlabel metal2 6888 14784 6888 14784 0 _0185_
rlabel metal2 7784 15400 7784 15400 0 _0186_
rlabel metal2 10584 15232 10584 15232 0 _0187_
rlabel metal2 15512 20328 15512 20328 0 _0188_
rlabel metal3 18760 22344 18760 22344 0 _0189_
rlabel metal2 20440 21896 20440 21896 0 _0190_
rlabel metal3 21672 23128 21672 23128 0 _0191_
rlabel metal2 23464 23576 23464 23576 0 _0192_
rlabel metal2 24584 19936 24584 19936 0 _0193_
rlabel metal2 21672 21056 21672 21056 0 _0194_
rlabel metal2 18200 24808 18200 24808 0 _0195_
rlabel metal2 17640 23408 17640 23408 0 _0196_
rlabel metal2 8736 17752 8736 17752 0 _0197_
rlabel metal2 10584 18536 10584 18536 0 _0198_
rlabel metal2 15400 19208 15400 19208 0 _0199_
rlabel metal2 17752 21112 17752 21112 0 _0200_
rlabel metal3 18704 21448 18704 21448 0 _0201_
rlabel metal2 18200 22736 18200 22736 0 _0202_
rlabel metal2 21448 19208 21448 19208 0 _0203_
rlabel metal2 20552 18872 20552 18872 0 _0204_
rlabel metal2 16072 18480 16072 18480 0 _0205_
rlabel metal2 13888 17640 13888 17640 0 _0206_
rlabel metal2 14056 17920 14056 17920 0 _0207_
rlabel metal2 15176 19348 15176 19348 0 _0208_
rlabel metal2 15512 17976 15512 17976 0 _0209_
rlabel metal3 16968 18424 16968 18424 0 _0210_
rlabel metal2 15960 19544 15960 19544 0 _0211_
rlabel metal2 16856 19264 16856 19264 0 _0212_
rlabel metal2 17864 19096 17864 19096 0 _0213_
rlabel metal2 17304 16688 17304 16688 0 _0214_
rlabel metal3 17584 15960 17584 15960 0 _0215_
rlabel metal3 12880 15960 12880 15960 0 _0216_
rlabel metal2 15512 17136 15512 17136 0 _0217_
rlabel metal2 16072 16744 16072 16744 0 _0218_
rlabel metal3 10472 15400 10472 15400 0 _0219_
rlabel metal2 11480 15204 11480 15204 0 _0220_
rlabel metal2 8624 15512 8624 15512 0 _0221_
rlabel metal2 10024 12880 10024 12880 0 _0222_
rlabel metal3 6440 12936 6440 12936 0 _0223_
rlabel metal2 7112 12656 7112 12656 0 _0224_
rlabel metal3 9240 13832 9240 13832 0 _0225_
rlabel metal2 10248 15204 10248 15204 0 _0226_
rlabel metal2 11704 12936 11704 12936 0 _0227_
rlabel metal2 9016 12096 9016 12096 0 _0228_
rlabel metal2 7336 11648 7336 11648 0 _0229_
rlabel metal3 7784 11480 7784 11480 0 _0230_
rlabel metal2 6440 10192 6440 10192 0 _0231_
rlabel metal2 23464 21784 23464 21784 0 _0232_
rlabel metal2 6720 8232 6720 8232 0 _0233_
rlabel metal2 10024 9968 10024 9968 0 _0234_
rlabel metal2 12600 14056 12600 14056 0 _0235_
rlabel metal2 16968 16464 16968 16464 0 _0236_
rlabel metal2 19208 18032 19208 18032 0 _0237_
rlabel metal3 22568 19208 22568 19208 0 _0238_
rlabel metal2 23688 20384 23688 20384 0 _0239_
rlabel metal2 26040 21952 26040 21952 0 _0240_
rlabel metal2 26824 22120 26824 22120 0 _0241_
rlabel metal3 27328 21560 27328 21560 0 _0242_
rlabel metal2 24248 20496 24248 20496 0 _0243_
rlabel metal2 21336 20384 21336 20384 0 _0244_
rlabel metal2 23128 20496 23128 20496 0 _0245_
rlabel metal2 24808 19040 24808 19040 0 _0246_
rlabel metal3 21280 16968 21280 16968 0 _0247_
rlabel metal2 19768 17472 19768 17472 0 _0248_
rlabel metal2 18648 19264 18648 19264 0 _0249_
rlabel metal2 19488 17640 19488 17640 0 _0250_
rlabel metal2 20888 18088 20888 18088 0 _0251_
rlabel metal2 21112 18480 21112 18480 0 _0252_
rlabel metal2 21840 17640 21840 17640 0 _0253_
rlabel metal3 20888 16072 20888 16072 0 _0254_
rlabel metal2 13384 16464 13384 16464 0 _0255_
rlabel metal2 13048 18368 13048 18368 0 _0256_
rlabel metal2 8792 13664 8792 13664 0 _0257_
rlabel metal2 8904 14504 8904 14504 0 _0258_
rlabel metal2 10808 14504 10808 14504 0 _0259_
rlabel metal2 13552 16856 13552 16856 0 _0260_
rlabel metal2 15288 14168 15288 14168 0 _0261_
rlabel metal3 17640 16072 17640 16072 0 _0262_
rlabel metal3 17640 16184 17640 16184 0 _0263_
rlabel metal2 19208 16576 19208 16576 0 _0264_
rlabel metal2 19544 13216 19544 13216 0 _0265_
rlabel metal2 18088 11144 18088 11144 0 _0266_
rlabel metal2 17976 11312 17976 11312 0 _0267_
rlabel metal2 18312 11032 18312 11032 0 _0268_
rlabel metal2 15512 9408 15512 9408 0 _0269_
rlabel metal2 13832 10528 13832 10528 0 _0270_
rlabel metal2 15456 11480 15456 11480 0 _0271_
rlabel metal2 15960 13272 15960 13272 0 _0272_
rlabel metal2 17864 9464 17864 9464 0 _0273_
rlabel metal2 12544 9576 12544 9576 0 _0274_
rlabel metal2 7448 9296 7448 9296 0 _0275_
rlabel metal2 9688 10360 9688 10360 0 _0276_
rlabel metal2 9744 10584 9744 10584 0 _0277_
rlabel metal2 11032 10584 11032 10584 0 _0278_
rlabel metal3 11872 10472 11872 10472 0 _0279_
rlabel metal2 20328 7504 20328 7504 0 _0280_
rlabel metal2 9576 8456 9576 8456 0 _0281_
rlabel metal2 7672 8176 7672 8176 0 _0282_
rlabel metal2 8008 8344 8008 8344 0 _0283_
rlabel metal2 8400 7448 8400 7448 0 _0284_
rlabel metal3 11424 8232 11424 8232 0 _0285_
rlabel metal2 16632 11312 16632 11312 0 _0286_
rlabel metal3 19824 15288 19824 15288 0 _0287_
rlabel metal2 21392 14728 21392 14728 0 _0288_
rlabel metal2 22344 16856 22344 16856 0 _0289_
rlabel metal3 25088 17640 25088 17640 0 _0290_
rlabel metal2 26040 21168 26040 21168 0 _0291_
rlabel metal2 25760 21672 25760 21672 0 _0292_
rlabel metal2 24136 23856 24136 23856 0 _0293_
rlabel metal2 23240 26096 23240 26096 0 _0294_
rlabel metal2 33992 25928 33992 25928 0 _0295_
rlabel metal2 42224 26488 42224 26488 0 _0296_
rlabel metal2 23800 25816 23800 25816 0 _0297_
rlabel metal2 25816 18704 25816 18704 0 _0298_
rlabel metal2 25424 19096 25424 19096 0 _0299_
rlabel metal2 28168 19600 28168 19600 0 _0300_
rlabel metal2 28056 20384 28056 20384 0 _0301_
rlabel metal3 25816 18424 25816 18424 0 _0302_
rlabel metal2 14952 15008 14952 15008 0 _0303_
rlabel metal3 18424 14728 18424 14728 0 _0304_
rlabel metal2 20664 16296 20664 16296 0 _0305_
rlabel metal2 23296 17752 23296 17752 0 _0306_
rlabel metal3 22568 17640 22568 17640 0 _0307_
rlabel metal2 26152 17360 26152 17360 0 _0308_
rlabel metal2 24136 16240 24136 16240 0 _0309_
rlabel metal3 24696 16072 24696 16072 0 _0310_
rlabel metal2 22456 15624 22456 15624 0 _0311_
rlabel metal2 23128 14728 23128 14728 0 _0312_
rlabel metal2 22568 15736 22568 15736 0 _0313_
rlabel metal2 21784 12320 21784 12320 0 _0314_
rlabel metal3 19320 12264 19320 12264 0 _0315_
rlabel metal2 14392 11424 14392 11424 0 _0316_
rlabel metal2 14560 16744 14560 16744 0 _0317_
rlabel metal2 10472 10024 10472 10024 0 _0318_
rlabel metal2 13048 10472 13048 10472 0 _0319_
rlabel metal2 15288 11480 15288 11480 0 _0320_
rlabel metal2 18536 11256 18536 11256 0 _0321_
rlabel metal2 17080 10864 17080 10864 0 _0322_
rlabel metal2 18200 12544 18200 12544 0 _0323_
rlabel metal2 19208 12432 19208 12432 0 _0324_
rlabel metal2 17976 8904 17976 8904 0 _0325_
rlabel metal2 14560 8344 14560 8344 0 _0326_
rlabel metal3 16408 9688 16408 9688 0 _0327_
rlabel metal2 15400 9016 15400 9016 0 _0328_
rlabel metal2 16912 8232 16912 8232 0 _0329_
rlabel metal2 14168 7840 14168 7840 0 _0330_
rlabel metal2 10472 7728 10472 7728 0 _0331_
rlabel metal2 25536 7672 25536 7672 0 _0332_
rlabel metal2 11312 7448 11312 7448 0 _0333_
rlabel metal2 11592 6888 11592 6888 0 _0334_
rlabel metal2 10920 6888 10920 6888 0 _0335_
rlabel metal2 11368 6664 11368 6664 0 _0336_
rlabel metal3 12656 6776 12656 6776 0 _0337_
rlabel metal2 8904 8344 8904 8344 0 _0338_
rlabel metal2 11256 8288 11256 8288 0 _0339_
rlabel metal2 15176 6552 15176 6552 0 _0340_
rlabel metal2 15512 7504 15512 7504 0 _0341_
rlabel metal2 19320 9128 19320 9128 0 _0342_
rlabel metal3 21784 13608 21784 13608 0 _0343_
rlabel metal3 25312 15176 25312 15176 0 _0344_
rlabel metal2 27552 19208 27552 19208 0 _0345_
rlabel metal2 28280 21224 28280 21224 0 _0346_
rlabel metal2 28056 18984 28056 18984 0 _0347_
rlabel metal2 28728 21840 28728 21840 0 _0348_
rlabel metal3 23968 22456 23968 22456 0 _0349_
rlabel metal2 24584 23184 24584 23184 0 _0350_
rlabel metal3 29008 22456 29008 22456 0 _0351_
rlabel metal2 27608 22624 27608 22624 0 _0352_
rlabel metal3 27776 28056 27776 28056 0 _0353_
rlabel metal2 27832 23912 27832 23912 0 _0354_
rlabel metal2 37184 23800 37184 23800 0 _0355_
rlabel metal2 35448 25200 35448 25200 0 _0356_
rlabel metal2 26488 18424 26488 18424 0 _0357_
rlabel metal2 28840 18816 28840 18816 0 _0358_
rlabel metal2 26040 15456 26040 15456 0 _0359_
rlabel metal2 23688 10192 23688 10192 0 _0360_
rlabel metal2 23912 14224 23912 14224 0 _0361_
rlabel metal3 23744 13720 23744 13720 0 _0362_
rlabel metal2 24584 14224 24584 14224 0 _0363_
rlabel metal2 26936 13440 26936 13440 0 _0364_
rlabel metal2 24360 11648 24360 11648 0 _0365_
rlabel metal2 22848 8344 22848 8344 0 _0366_
rlabel metal2 21000 11312 21000 11312 0 _0367_
rlabel metal2 20552 10080 20552 10080 0 _0368_
rlabel metal3 21168 11368 21168 11368 0 _0369_
rlabel metal2 22120 11648 22120 11648 0 _0370_
rlabel metal2 23800 12544 23800 12544 0 _0371_
rlabel metal2 21560 9464 21560 9464 0 _0372_
rlabel metal2 21224 9296 21224 9296 0 _0373_
rlabel metal2 17752 9296 17752 9296 0 _0374_
rlabel metal2 15960 8624 15960 8624 0 _0375_
rlabel metal2 18760 9520 18760 9520 0 _0376_
rlabel metal2 20104 8344 20104 8344 0 _0377_
rlabel metal2 20888 6608 20888 6608 0 _0378_
rlabel metal2 13888 5992 13888 5992 0 _0379_
rlabel metal3 15596 7448 15596 7448 0 _0380_
rlabel metal3 17416 7448 17416 7448 0 _0381_
rlabel metal2 16408 6720 16408 6720 0 _0382_
rlabel metal2 12208 6104 12208 6104 0 _0383_
rlabel metal2 16520 6720 16520 6720 0 _0384_
rlabel metal3 19096 6664 19096 6664 0 _0385_
rlabel metal2 20776 5600 20776 5600 0 _0386_
rlabel metal2 23016 10640 23016 10640 0 _0387_
rlabel metal2 25592 16072 25592 16072 0 _0388_
rlabel metal2 28280 16912 28280 16912 0 _0389_
rlabel metal2 29624 20048 29624 20048 0 _0390_
rlabel metal3 31472 23352 31472 23352 0 _0391_
rlabel metal2 28952 19096 28952 19096 0 _0392_
rlabel metal2 30072 23408 30072 23408 0 _0393_
rlabel metal3 13104 25256 13104 25256 0 _0394_
rlabel metal2 15008 25480 15008 25480 0 _0395_
rlabel metal2 23576 24752 23576 24752 0 _0396_
rlabel metal2 31640 24472 31640 24472 0 _0397_
rlabel metal2 30072 24136 30072 24136 0 _0398_
rlabel metal2 35336 31192 35336 31192 0 _0399_
rlabel metal2 37016 24192 37016 24192 0 _0400_
rlabel metal2 27720 18480 27720 18480 0 _0401_
rlabel metal2 26880 16072 26880 16072 0 _0402_
rlabel metal3 28896 16632 28896 16632 0 _0403_
rlabel metal2 26712 13328 26712 13328 0 _0404_
rlabel metal2 25928 12152 25928 12152 0 _0405_
rlabel metal3 24920 12152 24920 12152 0 _0406_
rlabel metal2 24696 12768 24696 12768 0 _0407_
rlabel metal2 27272 12488 27272 12488 0 _0408_
rlabel metal2 24584 8848 24584 8848 0 _0409_
rlabel metal2 21056 8232 21056 8232 0 _0410_
rlabel metal3 22904 9016 22904 9016 0 _0411_
rlabel metal2 24136 8960 24136 8960 0 _0412_
rlabel metal2 23576 7784 23576 7784 0 _0413_
rlabel metal2 22792 7728 22792 7728 0 _0414_
rlabel metal2 19208 6552 19208 6552 0 _0415_
rlabel metal2 19096 6160 19096 6160 0 _0416_
rlabel metal2 22456 6832 22456 6832 0 _0417_
rlabel metal2 21896 5376 21896 5376 0 _0418_
rlabel metal2 16520 6272 16520 6272 0 _0419_
rlabel metal3 20160 6776 20160 6776 0 _0420_
rlabel metal2 24360 6664 24360 6664 0 _0421_
rlabel metal2 24472 8288 24472 8288 0 _0422_
rlabel metal2 27608 10584 27608 10584 0 _0423_
rlabel metal2 29288 16576 29288 16576 0 _0424_
rlabel metal2 29904 16632 29904 16632 0 _0425_
rlabel metal2 29288 18312 29288 18312 0 _0426_
rlabel metal2 29624 24304 29624 24304 0 _0427_
rlabel metal3 13552 26488 13552 26488 0 _0428_
rlabel metal2 15288 25368 15288 25368 0 _0429_
rlabel metal2 30632 25480 30632 25480 0 _0430_
rlabel metal3 31136 26264 31136 26264 0 _0431_
rlabel metal2 30296 26264 30296 26264 0 _0432_
rlabel metal2 31304 25872 31304 25872 0 _0433_
rlabel metal3 30352 26376 30352 26376 0 _0434_
rlabel metal3 36736 23688 36736 23688 0 _0435_
rlabel metal2 28000 13720 28000 13720 0 _0436_
rlabel metal3 29960 14280 29960 14280 0 _0437_
rlabel metal2 30296 13328 30296 13328 0 _0438_
rlabel metal3 25312 9688 25312 9688 0 _0439_
rlabel metal2 26152 9296 26152 9296 0 _0440_
rlabel metal2 26992 10024 26992 10024 0 _0441_
rlabel metal2 29288 12432 29288 12432 0 _0442_
rlabel metal2 29512 9800 29512 9800 0 _0443_
rlabel metal2 25480 7056 25480 7056 0 _0444_
rlabel metal2 27608 8624 27608 8624 0 _0445_
rlabel metal2 28392 9800 28392 9800 0 _0446_
rlabel metal2 26040 7448 26040 7448 0 _0447_
rlabel metal3 28672 7448 28672 7448 0 _0448_
rlabel metal2 22456 5544 22456 5544 0 _0449_
rlabel metal2 26376 7112 26376 7112 0 _0450_
rlabel metal2 30184 7616 30184 7616 0 _0451_
rlabel metal2 31416 11368 31416 11368 0 _0452_
rlabel metal3 31416 14504 31416 14504 0 _0453_
rlabel metal2 30912 18200 30912 18200 0 _0454_
rlabel metal4 30184 19376 30184 19376 0 _0455_
rlabel metal2 31024 23352 31024 23352 0 _0456_
rlabel metal2 19544 25760 19544 25760 0 _0457_
rlabel metal2 23240 24528 23240 24528 0 _0458_
rlabel metal2 31752 24360 31752 24360 0 _0459_
rlabel metal2 35952 23912 35952 23912 0 _0460_
rlabel metal2 29456 9016 29456 9016 0 _0461_
rlabel metal2 30632 11312 30632 11312 0 _0462_
rlabel metal2 31024 12264 31024 12264 0 _0463_
rlabel metal2 31304 17584 31304 17584 0 _0464_
rlabel metal2 31080 17584 31080 17584 0 _0465_
rlabel metal3 29624 8344 29624 8344 0 _0466_
rlabel metal2 28504 10248 28504 10248 0 _0467_
rlabel metal3 31080 15176 31080 15176 0 _0468_
rlabel metal2 29288 15456 29288 15456 0 _0469_
rlabel metal2 26824 7896 26824 7896 0 _0470_
rlabel metal2 29792 15512 29792 15512 0 _0471_
rlabel metal3 31136 15288 31136 15288 0 _0472_
rlabel metal2 31192 18032 31192 18032 0 _0473_
rlabel metal2 31752 19712 31752 19712 0 _0474_
rlabel metal3 30296 19992 30296 19992 0 _0475_
rlabel metal3 31024 20104 31024 20104 0 _0476_
rlabel metal2 30240 20104 30240 20104 0 _0477_
rlabel metal3 24304 24920 24304 24920 0 _0478_
rlabel metal2 21336 24696 21336 24696 0 _0479_
rlabel metal2 21112 22568 21112 22568 0 _0480_
rlabel metal2 31192 21952 31192 21952 0 _0481_
rlabel metal3 35000 23800 35000 23800 0 _0482_
rlabel metal2 33824 26488 33824 26488 0 _0483_
rlabel metal2 30968 22680 30968 22680 0 _0484_
rlabel metal3 31640 22344 31640 22344 0 _0485_
rlabel metal2 30632 18200 30632 18200 0 _0486_
rlabel metal3 32032 19096 32032 19096 0 _0487_
rlabel metal2 31416 17584 31416 17584 0 _0488_
rlabel metal2 31864 15568 31864 15568 0 _0489_
rlabel metal2 31528 16800 31528 16800 0 _0490_
rlabel metal3 32200 19208 32200 19208 0 _0491_
rlabel metal2 32088 19824 32088 19824 0 _0492_
rlabel metal2 33096 19712 33096 19712 0 _0493_
rlabel metal2 23128 23408 23128 23408 0 _0494_
rlabel metal2 22792 21336 22792 21336 0 _0495_
rlabel metal2 33992 20888 33992 20888 0 _0496_
rlabel metal2 33768 21840 33768 21840 0 _0497_
rlabel metal2 36232 21280 36232 21280 0 _0498_
rlabel metal2 32424 19712 32424 19712 0 _0499_
rlabel metal2 27552 21000 27552 21000 0 _0500_
rlabel metal2 31304 21056 31304 21056 0 _0501_
rlabel metal2 35112 21224 35112 21224 0 _0502_
rlabel metal2 35000 21784 35000 21784 0 _0503_
rlabel metal2 35672 21616 35672 21616 0 _0504_
rlabel metal2 31192 51464 31192 51464 0 _0505_
rlabel metal3 34104 41048 34104 41048 0 _0506_
rlabel metal2 40264 34440 40264 34440 0 _0507_
rlabel metal2 45416 34384 45416 34384 0 _0508_
rlabel metal2 38360 37184 38360 37184 0 _0509_
rlabel metal2 19152 27272 19152 27272 0 _0510_
rlabel metal2 48888 39144 48888 39144 0 _0511_
rlabel metal2 37072 38920 37072 38920 0 _0512_
rlabel metal2 43792 43848 43792 43848 0 _0513_
rlabel metal2 33880 40712 33880 40712 0 _0514_
rlabel metal2 39592 47208 39592 47208 0 _0515_
rlabel metal2 31696 42056 31696 42056 0 _0516_
rlabel metal2 30296 52192 30296 52192 0 _0517_
rlabel metal2 30800 51912 30800 51912 0 _0518_
rlabel metal2 31416 52864 31416 52864 0 _0519_
rlabel metal3 30072 49784 30072 49784 0 _0520_
rlabel metal2 18760 28112 18760 28112 0 _0521_
rlabel metal3 31780 51464 31780 51464 0 _0522_
rlabel metal2 36120 51688 36120 51688 0 _0523_
rlabel metal2 31528 52640 31528 52640 0 _0524_
rlabel metal2 34888 50904 34888 50904 0 _0525_
rlabel metal2 35448 50624 35448 50624 0 _0526_
rlabel metal2 34216 50960 34216 50960 0 _0527_
rlabel metal3 32592 51240 32592 51240 0 _0528_
rlabel metal2 31304 48440 31304 48440 0 _0529_
rlabel metal2 30408 47488 30408 47488 0 _0530_
rlabel metal2 31080 46760 31080 46760 0 _0531_
rlabel metal2 19656 28280 19656 28280 0 _0532_
rlabel metal2 41496 49392 41496 49392 0 _0533_
rlabel metal2 32088 48104 32088 48104 0 _0534_
rlabel metal2 31416 43344 31416 43344 0 _0535_
rlabel metal2 29792 46760 29792 46760 0 _0536_
rlabel metal3 35000 48888 35000 48888 0 _0537_
rlabel metal2 32424 52416 32424 52416 0 _0538_
rlabel metal2 33880 51688 33880 51688 0 _0539_
rlabel metal2 35560 52248 35560 52248 0 _0540_
rlabel metal3 31472 46760 31472 46760 0 _0541_
rlabel metal3 33376 46536 33376 46536 0 _0542_
rlabel metal2 21336 27328 21336 27328 0 _0543_
rlabel metal2 30520 42280 30520 42280 0 _0544_
rlabel metal2 32200 42504 32200 42504 0 _0545_
rlabel metal2 37800 39368 37800 39368 0 _0546_
rlabel metal3 33992 44184 33992 44184 0 _0547_
rlabel metal2 32648 51352 32648 51352 0 _0548_
rlabel metal2 33544 52976 33544 52976 0 _0549_
rlabel metal2 35784 50960 35784 50960 0 _0550_
rlabel metal2 33152 45864 33152 45864 0 _0551_
rlabel metal2 33544 46368 33544 46368 0 _0552_
rlabel metal2 32312 46368 32312 46368 0 _0553_
rlabel metal2 22456 28616 22456 28616 0 _0554_
rlabel metal2 35000 46984 35000 46984 0 _0555_
rlabel metal2 32648 49168 32648 49168 0 _0556_
rlabel metal2 32760 49392 32760 49392 0 _0557_
rlabel metal2 35784 52920 35784 52920 0 _0558_
rlabel metal2 35672 54824 35672 54824 0 _0559_
rlabel metal2 35112 52472 35112 52472 0 _0560_
rlabel metal2 35504 47432 35504 47432 0 _0561_
rlabel metal2 32424 42336 32424 42336 0 _0562_
rlabel metal2 34104 40824 34104 40824 0 _0563_
rlabel metal2 35336 40880 35336 40880 0 _0564_
rlabel metal3 21952 27944 21952 27944 0 _0565_
rlabel metal3 36400 42616 36400 42616 0 _0566_
rlabel metal3 33936 42840 33936 42840 0 _0567_
rlabel metal2 35448 44044 35448 44044 0 _0568_
rlabel metal2 34048 41832 34048 41832 0 _0569_
rlabel metal3 36624 45640 36624 45640 0 _0570_
rlabel metal2 36232 44856 36232 44856 0 _0571_
rlabel metal2 36904 49840 36904 49840 0 _0572_
rlabel metal3 34048 51464 34048 51464 0 _0573_
rlabel metal2 36288 54488 36288 54488 0 _0574_
rlabel metal3 36568 53032 36568 53032 0 _0575_
rlabel metal2 25816 28672 25816 28672 0 _0576_
rlabel metal3 35672 49000 35672 49000 0 _0577_
rlabel metal2 36344 48104 36344 48104 0 _0578_
rlabel metal2 39480 49952 39480 49952 0 _0579_
rlabel metal2 37520 50456 37520 50456 0 _0580_
rlabel metal2 38360 50848 38360 50848 0 _0581_
rlabel metal2 38024 52696 38024 52696 0 _0582_
rlabel metal3 44856 50344 44856 50344 0 _0583_
rlabel metal2 38360 51800 38360 51800 0 _0584_
rlabel metal2 38920 52248 38920 52248 0 _0585_
rlabel metal2 37240 54096 37240 54096 0 _0586_
rlabel metal2 38920 29680 38920 29680 0 _0587_
rlabel metal2 36792 53984 36792 53984 0 _0588_
rlabel metal2 38808 54824 38808 54824 0 _0589_
rlabel metal2 39144 49896 39144 49896 0 _0590_
rlabel metal2 36456 42728 36456 42728 0 _0591_
rlabel metal2 35896 41720 35896 41720 0 _0592_
rlabel metal2 36848 38920 36848 38920 0 _0593_
rlabel metal3 37128 38808 37128 38808 0 _0594_
rlabel metal2 38360 40712 38360 40712 0 _0595_
rlabel metal2 37800 42672 37800 42672 0 _0596_
rlabel metal2 37912 43064 37912 43064 0 _0597_
rlabel metal2 36568 41832 36568 41832 0 _0598_
rlabel metal2 39256 41216 39256 41216 0 _0599_
rlabel metal2 40376 46592 40376 46592 0 _0600_
rlabel metal2 40824 43960 40824 43960 0 _0601_
rlabel metal2 47992 46928 47992 46928 0 _0602_
rlabel metal2 31416 46536 31416 46536 0 _0603_
rlabel metal2 33432 48216 33432 48216 0 _0604_
rlabel metal2 34216 48496 34216 48496 0 _0605_
rlabel metal2 34440 48104 34440 48104 0 _0606_
rlabel metal3 36008 48216 36008 48216 0 _0607_
rlabel metal2 11704 32144 11704 32144 0 _0608_
rlabel metal2 37352 48440 37352 48440 0 _0609_
rlabel metal2 36680 48888 36680 48888 0 _0610_
rlabel metal2 37912 48328 37912 48328 0 _0611_
rlabel metal3 39536 46760 39536 46760 0 _0612_
rlabel metal2 39592 46144 39592 46144 0 _0613_
rlabel metal2 38808 45808 38808 45808 0 _0614_
rlabel metal2 38696 44352 38696 44352 0 _0615_
rlabel metal2 38808 48608 38808 48608 0 _0616_
rlabel metal2 40096 52920 40096 52920 0 _0617_
rlabel metal2 41944 50960 41944 50960 0 _0618_
rlabel metal3 15736 36344 15736 36344 0 _0619_
rlabel metal2 37632 52696 37632 52696 0 _0620_
rlabel metal2 38248 50456 38248 50456 0 _0621_
rlabel metal2 39256 49728 39256 49728 0 _0622_
rlabel metal2 36568 51296 36568 51296 0 _0623_
rlabel metal2 49336 48776 49336 48776 0 _0624_
rlabel metal2 42784 52920 42784 52920 0 _0625_
rlabel metal2 43064 53368 43064 53368 0 _0626_
rlabel metal2 41384 51800 41384 51800 0 _0627_
rlabel metal3 41888 52136 41888 52136 0 _0628_
rlabel metal2 41944 47936 41944 47936 0 _0629_
rlabel metal2 22120 42672 22120 42672 0 _0630_
rlabel metal2 41384 47376 41384 47376 0 _0631_
rlabel metal2 39704 43876 39704 43876 0 _0632_
rlabel metal2 37296 40376 37296 40376 0 _0633_
rlabel metal2 39144 37296 39144 37296 0 _0634_
rlabel metal2 39480 36736 39480 36736 0 _0635_
rlabel metal2 39704 34664 39704 34664 0 _0636_
rlabel metal3 40600 38024 40600 38024 0 _0637_
rlabel metal3 36120 40600 36120 40600 0 _0638_
rlabel metal2 42392 42504 42392 42504 0 _0639_
rlabel metal2 39144 52752 39144 52752 0 _0640_
rlabel metal3 18648 38920 18648 38920 0 _0641_
rlabel metal2 38920 48160 38920 48160 0 _0642_
rlabel metal2 42168 46368 42168 46368 0 _0643_
rlabel metal2 42952 43932 42952 43932 0 _0644_
rlabel metal2 39816 40040 39816 40040 0 _0645_
rlabel metal2 38920 41048 38920 41048 0 _0646_
rlabel metal2 43736 39256 43736 39256 0 _0647_
rlabel metal3 42280 40376 42280 40376 0 _0648_
rlabel metal2 41048 41384 41048 41384 0 _0649_
rlabel metal2 43624 45696 43624 45696 0 _0650_
rlabel metal2 41944 46200 41944 46200 0 _0651_
rlabel metal2 18984 36848 18984 36848 0 _0652_
rlabel metal2 41496 45640 41496 45640 0 _0653_
rlabel metal2 41664 45080 41664 45080 0 _0654_
rlabel metal2 45248 45192 45248 45192 0 _0655_
rlabel metal2 39704 43008 39704 43008 0 _0656_
rlabel metal2 40264 42616 40264 42616 0 _0657_
rlabel metal2 44968 42448 44968 42448 0 _0658_
rlabel metal2 43848 45640 43848 45640 0 _0659_
rlabel metal2 43736 45192 43736 45192 0 _0660_
rlabel metal2 42728 46256 42728 46256 0 _0661_
rlabel metal2 45528 44688 45528 44688 0 _0662_
rlabel metal2 15512 43624 15512 43624 0 _0663_
rlabel metal2 42056 43400 42056 43400 0 _0664_
rlabel metal2 43960 47040 43960 47040 0 _0665_
rlabel metal2 44184 47880 44184 47880 0 _0666_
rlabel metal2 41888 50008 41888 50008 0 _0667_
rlabel metal2 44968 50064 44968 50064 0 _0668_
rlabel metal2 44520 53032 44520 53032 0 _0669_
rlabel metal2 43792 51464 43792 51464 0 _0670_
rlabel metal3 42448 51352 42448 51352 0 _0671_
rlabel metal2 43288 48720 43288 48720 0 _0672_
rlabel metal2 43736 48496 43736 48496 0 _0673_
rlabel metal2 10696 33824 10696 33824 0 _0674_
rlabel metal3 47880 50456 47880 50456 0 _0675_
rlabel metal2 45416 51296 45416 51296 0 _0676_
rlabel metal2 45192 53144 45192 53144 0 _0677_
rlabel metal2 51016 51856 51016 51856 0 _0678_
rlabel metal2 50904 52304 50904 52304 0 _0679_
rlabel metal2 48888 52528 48888 52528 0 _0680_
rlabel metal2 46984 52080 46984 52080 0 _0681_
rlabel metal2 46872 48440 46872 48440 0 _0682_
rlabel metal2 45080 44296 45080 44296 0 _0683_
rlabel metal2 44968 41552 44968 41552 0 _0684_
rlabel metal2 15176 32172 15176 32172 0 _0685_
rlabel metal2 43568 39592 43568 39592 0 _0686_
rlabel metal2 41720 37408 41720 37408 0 _0687_
rlabel metal2 40880 34888 40880 34888 0 _0688_
rlabel metal2 41216 33432 41216 33432 0 _0689_
rlabel metal2 41048 33824 41048 33824 0 _0690_
rlabel metal2 39872 35112 39872 35112 0 _0691_
rlabel metal2 41944 39256 41944 39256 0 _0692_
rlabel metal2 40488 37016 40488 37016 0 _0693_
rlabel metal2 42728 36008 42728 36008 0 _0694_
rlabel metal3 44016 38920 44016 38920 0 _0695_
rlabel metal2 3024 35448 3024 35448 0 _0696_
rlabel metal2 49112 41272 49112 41272 0 _0697_
rlabel metal2 45416 41552 45416 41552 0 _0698_
rlabel metal2 44856 40880 44856 40880 0 _0699_
rlabel metal2 43960 40656 43960 40656 0 _0700_
rlabel metal2 44072 40096 44072 40096 0 _0701_
rlabel metal2 44408 40096 44408 40096 0 _0702_
rlabel metal2 46872 39144 46872 39144 0 _0703_
rlabel metal2 45080 46144 45080 46144 0 _0704_
rlabel metal3 42840 45752 42840 45752 0 _0705_
rlabel metal2 42952 50792 42952 50792 0 _0706_
rlabel metal3 1904 44408 1904 44408 0 _0707_
rlabel metal2 44184 50456 44184 50456 0 _0708_
rlabel metal3 44184 48104 44184 48104 0 _0709_
rlabel metal2 45416 47152 45416 47152 0 _0710_
rlabel metal3 45472 45304 45472 45304 0 _0711_
rlabel metal3 45136 44968 45136 44968 0 _0712_
rlabel metal2 46144 44072 46144 44072 0 _0713_
rlabel metal2 44072 43400 44072 43400 0 _0714_
rlabel metal3 47880 41832 47880 41832 0 _0715_
rlabel metal2 52808 42280 52808 42280 0 _0716_
rlabel metal2 47656 45920 47656 45920 0 _0717_
rlabel metal2 2744 34048 2744 34048 0 _0718_
rlabel metal3 49504 43288 49504 43288 0 _0719_
rlabel metal3 51912 45752 51912 45752 0 _0720_
rlabel metal2 47432 46088 47432 46088 0 _0721_
rlabel metal2 46984 44912 46984 44912 0 _0722_
rlabel metal2 47320 44408 47320 44408 0 _0723_
rlabel metal2 47880 47544 47880 47544 0 _0724_
rlabel metal3 49336 46760 49336 46760 0 _0725_
rlabel metal3 47208 51352 47208 51352 0 _0726_
rlabel metal2 51912 50624 51912 50624 0 _0727_
rlabel metal3 48104 50568 48104 50568 0 _0728_
rlabel metal2 17416 32760 17416 32760 0 _0729_
rlabel metal2 46760 49112 46760 49112 0 _0730_
rlabel metal2 47544 47992 47544 47992 0 _0731_
rlabel metal2 51016 48440 51016 48440 0 _0732_
rlabel metal2 50568 48440 50568 48440 0 _0733_
rlabel metal2 51128 50904 51128 50904 0 _0734_
rlabel metal2 49000 50456 49000 50456 0 _0735_
rlabel metal2 50456 49504 50456 49504 0 _0736_
rlabel metal2 51016 49280 51016 49280 0 _0737_
rlabel metal2 50008 46200 50008 46200 0 _0738_
rlabel metal3 47992 40264 47992 40264 0 _0739_
rlabel metal2 3472 30968 3472 30968 0 _0740_
rlabel metal2 46424 39536 46424 39536 0 _0741_
rlabel metal2 43680 38808 43680 38808 0 _0742_
rlabel metal2 42616 35336 42616 35336 0 _0743_
rlabel metal3 42504 34216 42504 34216 0 _0744_
rlabel metal3 36288 33992 36288 33992 0 _0745_
rlabel metal3 35728 34216 35728 34216 0 _0746_
rlabel metal2 32088 34216 32088 34216 0 _0747_
rlabel metal2 32424 39480 32424 39480 0 _0748_
rlabel metal2 31640 40432 31640 40432 0 _0749_
rlabel metal2 2520 49448 2520 49448 0 _0750_
rlabel metal3 36456 34664 36456 34664 0 _0751_
rlabel metal2 49336 34496 49336 34496 0 _0752_
rlabel metal2 43176 34608 43176 34608 0 _0753_
rlabel metal2 42952 33824 42952 33824 0 _0754_
rlabel metal3 42336 33320 42336 33320 0 _0755_
rlabel metal2 44240 34888 44240 34888 0 _0756_
rlabel metal2 43624 42448 43624 42448 0 _0757_
rlabel metal2 46592 39592 46592 39592 0 _0758_
rlabel metal2 45416 39872 45416 39872 0 _0759_
rlabel metal2 48048 39592 48048 39592 0 _0760_
rlabel metal2 7112 33040 7112 33040 0 _0761_
rlabel metal2 44072 37688 44072 37688 0 _0762_
rlabel metal2 45752 35392 45752 35392 0 _0763_
rlabel metal2 49672 35560 49672 35560 0 _0764_
rlabel metal2 46200 34608 46200 34608 0 _0765_
rlabel metal2 46872 36680 46872 36680 0 _0766_
rlabel metal2 47880 39256 47880 39256 0 _0767_
rlabel metal2 47656 38360 47656 38360 0 _0768_
rlabel metal2 49280 38808 49280 38808 0 _0769_
rlabel metal2 49168 39032 49168 39032 0 _0770_
rlabel metal2 48328 45416 48328 45416 0 _0771_
rlabel metal3 7560 31752 7560 31752 0 _0772_
rlabel metal2 45080 44912 45080 44912 0 _0773_
rlabel metal2 47656 51296 47656 51296 0 _0774_
rlabel metal2 50568 48944 50568 48944 0 _0775_
rlabel metal2 49672 46368 49672 46368 0 _0776_
rlabel metal2 49000 43176 49000 43176 0 _0777_
rlabel metal2 49896 42224 49896 42224 0 _0778_
rlabel metal2 49448 41440 49448 41440 0 _0779_
rlabel metal2 49112 39984 49112 39984 0 _0780_
rlabel metal2 51464 43176 51464 43176 0 _0781_
rlabel metal2 51688 46592 51688 46592 0 _0782_
rlabel metal3 7784 31864 7784 31864 0 _0783_
rlabel metal2 51688 45248 51688 45248 0 _0784_
rlabel metal2 50680 44576 50680 44576 0 _0785_
rlabel metal2 51016 43876 51016 43876 0 _0786_
rlabel metal2 53816 46536 53816 46536 0 _0787_
rlabel metal2 52136 49896 52136 49896 0 _0788_
rlabel metal2 52696 49168 52696 49168 0 _0789_
rlabel metal2 53032 50064 53032 50064 0 _0790_
rlabel metal2 53816 49168 53816 49168 0 _0791_
rlabel metal2 53928 50176 53928 50176 0 _0792_
rlabel metal3 53536 49224 53536 49224 0 _0793_
rlabel metal2 9688 32032 9688 32032 0 _0794_
rlabel metal2 52752 46648 52752 46648 0 _0795_
rlabel metal2 51800 50064 51800 50064 0 _0796_
rlabel metal2 51576 49168 51576 49168 0 _0797_
rlabel metal3 52304 48440 52304 48440 0 _0798_
rlabel metal2 52472 45136 52472 45136 0 _0799_
rlabel metal2 51576 41888 51576 41888 0 _0800_
rlabel metal2 48328 40208 48328 40208 0 _0801_
rlabel metal3 48832 34888 48832 34888 0 _0802_
rlabel metal2 43960 33824 43960 33824 0 _0803_
rlabel metal2 42224 32760 42224 32760 0 _0804_
rlabel metal2 20664 31080 20664 31080 0 _0805_
rlabel metal2 43848 33824 43848 33824 0 _0806_
rlabel metal2 42504 32536 42504 32536 0 _0807_
rlabel metal2 42056 32144 42056 32144 0 _0808_
rlabel metal2 34664 35336 34664 35336 0 _0809_
rlabel metal2 35000 32088 35000 32088 0 _0810_
rlabel metal2 36008 32648 36008 32648 0 _0811_
rlabel metal2 39200 28056 39200 28056 0 _0812_
rlabel metal2 44632 34496 44632 34496 0 _0813_
rlabel metal2 43680 34216 43680 34216 0 _0814_
rlabel metal3 11872 32536 11872 32536 0 _0815_
rlabel metal2 47544 34440 47544 34440 0 _0816_
rlabel metal2 47264 37128 47264 37128 0 _0817_
rlabel metal2 50288 39592 50288 39592 0 _0818_
rlabel metal3 48440 39368 48440 39368 0 _0819_
rlabel metal2 48328 36456 48328 36456 0 _0820_
rlabel metal2 49000 35952 49000 35952 0 _0821_
rlabel metal2 49896 37968 49896 37968 0 _0822_
rlabel metal3 51408 38584 51408 38584 0 _0823_
rlabel metal2 49672 43064 49672 43064 0 _0824_
rlabel metal2 50456 41440 50456 41440 0 _0825_
rlabel metal3 8232 50568 8232 50568 0 _0826_
rlabel metal2 51352 39536 51352 39536 0 _0827_
rlabel metal2 50008 39144 50008 39144 0 _0828_
rlabel metal2 50904 39368 50904 39368 0 _0829_
rlabel metal3 52472 39480 52472 39480 0 _0830_
rlabel metal2 53256 40432 53256 40432 0 _0831_
rlabel metal2 52584 45192 52584 45192 0 _0832_
rlabel metal2 51240 43456 51240 43456 0 _0833_
rlabel metal2 51688 41832 51688 41832 0 _0834_
rlabel metal2 54712 40656 54712 40656 0 _0835_
rlabel metal2 54936 42000 54936 42000 0 _0836_
rlabel metal2 8120 31752 8120 31752 0 _0837_
rlabel metal2 53312 46536 53312 46536 0 _0838_
rlabel metal2 53536 45080 53536 45080 0 _0839_
rlabel metal3 54208 45080 54208 45080 0 _0840_
rlabel metal2 54376 46312 54376 46312 0 _0841_
rlabel metal2 53704 48496 53704 48496 0 _0842_
rlabel metal2 54152 46816 54152 46816 0 _0843_
rlabel metal2 54824 45640 54824 45640 0 _0844_
rlabel metal2 54264 40768 54264 40768 0 _0845_
rlabel metal3 52696 39144 52696 39144 0 _0846_
rlabel metal2 48440 33992 48440 33992 0 _0847_
rlabel metal2 2352 39256 2352 39256 0 _0848_
rlabel metal3 45080 34104 45080 34104 0 _0849_
rlabel metal3 39480 34328 39480 34328 0 _0850_
rlabel metal2 43960 32648 43960 32648 0 _0851_
rlabel metal2 37128 33488 37128 33488 0 _0852_
rlabel metal3 34384 38696 34384 38696 0 _0853_
rlabel metal2 35000 34440 35000 34440 0 _0854_
rlabel metal2 35560 33600 35560 33600 0 _0855_
rlabel metal2 36344 32032 36344 32032 0 _0856_
rlabel metal2 34832 37352 34832 37352 0 _0857_
rlabel metal2 33544 38724 33544 38724 0 _0858_
rlabel metal3 2184 35896 2184 35896 0 _0859_
rlabel metal2 29960 34832 29960 34832 0 _0860_
rlabel metal3 42672 33208 42672 33208 0 _0861_
rlabel metal2 47376 33320 47376 33320 0 _0862_
rlabel metal2 45864 33040 45864 33040 0 _0863_
rlabel metal2 49616 32760 49616 32760 0 _0864_
rlabel metal2 52248 37464 52248 37464 0 _0865_
rlabel metal2 52696 36960 52696 36960 0 _0866_
rlabel metal2 50232 36512 50232 36512 0 _0867_
rlabel metal2 50344 35560 50344 35560 0 _0868_
rlabel metal3 4368 30856 4368 30856 0 _0869_
rlabel metal2 52304 34888 52304 34888 0 _0870_
rlabel metal2 53368 40320 53368 40320 0 _0871_
rlabel metal2 54264 36904 54264 36904 0 _0872_
rlabel metal2 55216 35672 55216 35672 0 _0873_
rlabel metal2 53536 38808 53536 38808 0 _0874_
rlabel metal2 53816 38416 53816 38416 0 _0875_
rlabel metal2 57176 43064 57176 43064 0 _0876_
rlabel metal2 54712 43008 54712 43008 0 _0877_
rlabel metal2 54488 40936 54488 40936 0 _0878_
rlabel metal2 54152 40096 54152 40096 0 _0879_
rlabel metal2 4984 32984 4984 32984 0 _0880_
rlabel metal2 54264 45752 54264 45752 0 _0881_
rlabel metal2 54488 44520 54488 44520 0 _0882_
rlabel metal2 54824 39144 54824 39144 0 _0883_
rlabel metal2 55272 36568 55272 36568 0 _0884_
rlabel metal2 49896 33712 49896 33712 0 _0885_
rlabel metal2 46648 32816 46648 32816 0 _0886_
rlabel metal2 44968 31472 44968 31472 0 _0887_
rlabel metal2 49000 31472 49000 31472 0 _0888_
rlabel metal3 33544 31752 33544 31752 0 _0889_
rlabel metal3 31416 41160 31416 41160 0 _0890_
rlabel metal2 5992 29568 5992 29568 0 _0891_
rlabel metal2 31976 40376 31976 40376 0 _0892_
rlabel metal2 34664 32368 34664 32368 0 _0893_
rlabel metal3 32312 33432 32312 33432 0 _0894_
rlabel metal3 38808 30968 38808 30968 0 _0895_
rlabel metal2 49784 33320 49784 33320 0 _0896_
rlabel metal2 49672 31976 49672 31976 0 _0897_
rlabel metal2 49896 30996 49896 30996 0 _0898_
rlabel metal2 51576 33152 51576 33152 0 _0899_
rlabel metal3 53704 34888 53704 34888 0 _0900_
rlabel metal2 4648 30296 4648 30296 0 _0901_
rlabel metal2 53088 34104 53088 34104 0 _0902_
rlabel metal2 53032 31360 53032 31360 0 _0903_
rlabel metal2 53816 31080 53816 31080 0 _0904_
rlabel metal2 53816 33992 53816 33992 0 _0905_
rlabel metal3 55272 33096 55272 33096 0 _0906_
rlabel metal2 54152 31808 54152 31808 0 _0907_
rlabel metal2 53256 38920 53256 38920 0 _0908_
rlabel metal3 54152 33320 54152 33320 0 _0909_
rlabel metal2 55496 39088 55496 39088 0 _0910_
rlabel metal2 54936 34608 54936 34608 0 _0911_
rlabel metal2 7112 31024 7112 31024 0 _0912_
rlabel metal2 54152 32872 54152 32872 0 _0913_
rlabel metal2 50232 31248 50232 31248 0 _0914_
rlabel metal2 48776 31416 48776 31416 0 _0915_
rlabel metal3 40264 33096 40264 33096 0 _0916_
rlabel metal2 49000 30408 49000 30408 0 _0917_
rlabel metal2 37576 32256 37576 32256 0 _0918_
rlabel metal2 33824 39592 33824 39592 0 _0919_
rlabel metal2 34832 39368 34832 39368 0 _0920_
rlabel metal3 37184 33320 37184 33320 0 _0921_
rlabel metal2 38248 32032 38248 32032 0 _0922_
rlabel metal2 3752 32088 3752 32088 0 _0923_
rlabel metal2 38080 29624 38080 29624 0 _0924_
rlabel metal3 54208 30744 54208 30744 0 _0925_
rlabel metal3 51968 30296 51968 30296 0 _0926_
rlabel metal2 50176 30184 50176 30184 0 _0927_
rlabel metal3 47712 29960 47712 29960 0 _0928_
rlabel metal2 45752 30296 45752 30296 0 _0929_
rlabel metal3 55440 30968 55440 30968 0 _0930_
rlabel metal2 54376 30912 54376 30912 0 _0931_
rlabel metal2 47768 30464 47768 30464 0 _0932_
rlabel metal2 7448 30464 7448 30464 0 _0933_
rlabel metal2 47600 30968 47600 30968 0 _0934_
rlabel metal2 52136 31920 52136 31920 0 _0935_
rlabel metal2 48104 31080 48104 31080 0 _0936_
rlabel metal2 47208 30520 47208 30520 0 _0937_
rlabel metal2 46200 29680 46200 29680 0 _0938_
rlabel metal2 45192 30296 45192 30296 0 _0939_
rlabel metal2 46648 29736 46648 29736 0 _0940_
rlabel metal3 40992 30296 40992 30296 0 _0941_
rlabel metal2 37632 29512 37632 29512 0 _0942_
rlabel metal3 36792 38024 36792 38024 0 _0943_
rlabel metal2 10696 30576 10696 30576 0 _0944_
rlabel metal2 37128 30464 37128 30464 0 _0945_
rlabel metal2 37408 28056 37408 28056 0 _0946_
rlabel metal2 37128 28224 37128 28224 0 _0947_
rlabel metal2 38024 27832 38024 27832 0 _0948_
rlabel metal3 45472 29624 45472 29624 0 _0949_
rlabel metal2 43624 30688 43624 30688 0 _0950_
rlabel metal2 45808 31080 45808 31080 0 _0951_
rlabel metal2 46872 31304 46872 31304 0 _0952_
rlabel metal2 45584 30744 45584 30744 0 _0953_
rlabel metal2 15288 32144 15288 32144 0 _0954_
rlabel metal2 43400 30240 43400 30240 0 _0955_
rlabel metal2 41608 29288 41608 29288 0 _0956_
rlabel metal2 42728 29568 42728 29568 0 _0957_
rlabel metal2 38136 36960 38136 36960 0 _0958_
rlabel metal2 41272 28952 41272 28952 0 _0959_
rlabel metal3 42056 28392 42056 28392 0 _0960_
rlabel metal2 42168 28336 42168 28336 0 _0961_
rlabel metal2 42840 28616 42840 28616 0 _0962_
rlabel metal2 42840 30072 42840 30072 0 _0963_
rlabel metal3 16632 31696 16632 31696 0 _0964_
rlabel metal2 40376 34272 40376 34272 0 _0965_
rlabel metal2 41888 29400 41888 29400 0 _0966_
rlabel metal2 40040 28840 40040 28840 0 _0967_
rlabel metal2 39368 28112 39368 28112 0 _0968_
rlabel metal2 41608 26152 41608 26152 0 _0969_
rlabel metal2 18256 38920 18256 38920 0 _0970_
rlabel metal2 10472 34160 10472 34160 0 _0971_
rlabel metal3 7224 30968 7224 30968 0 _0972_
rlabel metal2 7896 29288 7896 29288 0 _0973_
rlabel metal2 7784 29680 7784 29680 0 _0974_
rlabel metal2 8232 30464 8232 30464 0 _0975_
rlabel metal3 9576 33432 9576 33432 0 _0976_
rlabel metal2 9576 37688 9576 37688 0 _0977_
rlabel metal2 7336 34608 7336 34608 0 _0978_
rlabel metal2 2408 36568 2408 36568 0 _0979_
rlabel metal2 3528 33600 3528 33600 0 _0980_
rlabel metal2 3640 36008 3640 36008 0 _0981_
rlabel metal2 4872 35280 4872 35280 0 _0982_
rlabel metal2 2744 36008 2744 36008 0 _0983_
rlabel metal2 4536 35672 4536 35672 0 _0984_
rlabel metal2 6888 35224 6888 35224 0 _0985_
rlabel metal2 11592 33656 11592 33656 0 _0986_
rlabel metal3 13664 33432 13664 33432 0 _0987_
rlabel metal2 15568 36456 15568 36456 0 _0988_
rlabel metal3 20776 34888 20776 34888 0 _0989_
rlabel metal2 13944 34496 13944 34496 0 _0990_
rlabel metal2 8344 40880 8344 40880 0 _0991_
rlabel metal2 12488 33656 12488 33656 0 _0992_
rlabel metal2 8904 31136 8904 31136 0 _0993_
rlabel metal2 9072 29624 9072 29624 0 _0994_
rlabel via2 9912 34104 9912 34104 0 _0995_
rlabel metal2 11984 33992 11984 33992 0 _0996_
rlabel metal2 13608 33264 13608 33264 0 _0997_
rlabel metal2 7448 36568 7448 36568 0 _0998_
rlabel metal2 8344 35056 8344 35056 0 _0999_
rlabel metal2 6888 37184 6888 37184 0 _1000_
rlabel metal2 6440 40320 6440 40320 0 _1001_
rlabel metal2 4816 37016 4816 37016 0 _1002_
rlabel metal2 2632 40264 2632 40264 0 _1003_
rlabel metal2 2128 36344 2128 36344 0 _1004_
rlabel metal2 3080 38808 3080 38808 0 _1005_
rlabel metal2 2856 39172 2856 39172 0 _1006_
rlabel metal2 2744 38136 2744 38136 0 _1007_
rlabel metal2 7896 37632 7896 37632 0 _1008_
rlabel metal2 14168 34496 14168 34496 0 _1009_
rlabel metal3 16632 34888 16632 34888 0 _1010_
rlabel metal3 18424 35112 18424 35112 0 _1011_
rlabel metal2 19320 36008 19320 36008 0 _1012_
rlabel metal2 18088 37016 18088 37016 0 _1013_
rlabel metal2 14504 35056 14504 35056 0 _1014_
rlabel metal2 14392 34944 14392 34944 0 _1015_
rlabel metal3 14616 35672 14616 35672 0 _1016_
rlabel metal2 15736 36456 15736 36456 0 _1017_
rlabel metal2 16296 39256 16296 39256 0 _1018_
rlabel metal2 15960 37744 15960 37744 0 _1019_
rlabel metal2 6440 46368 6440 46368 0 _1020_
rlabel metal2 8680 34496 8680 34496 0 _1021_
rlabel metal2 8120 34776 8120 34776 0 _1022_
rlabel metal2 8344 37520 8344 37520 0 _1023_
rlabel metal2 8624 39480 8624 39480 0 _1024_
rlabel metal3 10360 37800 10360 37800 0 _1025_
rlabel metal2 10696 39088 10696 39088 0 _1026_
rlabel metal2 11032 37240 11032 37240 0 _1027_
rlabel metal2 6888 40656 6888 40656 0 _1028_
rlabel metal2 6440 39648 6440 39648 0 _1029_
rlabel metal2 5208 38080 5208 38080 0 _1030_
rlabel metal2 5712 38696 5712 38696 0 _1031_
rlabel metal2 9576 43792 9576 43792 0 _1032_
rlabel metal2 6104 42112 6104 42112 0 _1033_
rlabel metal3 4648 44072 4648 44072 0 _1034_
rlabel metal2 3304 46256 3304 46256 0 _1035_
rlabel metal2 6888 44072 6888 44072 0 _1036_
rlabel metal2 5656 44744 5656 44744 0 _1037_
rlabel metal2 2744 43568 2744 43568 0 _1038_
rlabel metal2 3920 39592 3920 39592 0 _1039_
rlabel metal2 2968 41608 2968 41608 0 _1040_
rlabel metal2 3976 42672 3976 42672 0 _1041_
rlabel metal2 6216 41496 6216 41496 0 _1042_
rlabel metal2 10136 39256 10136 39256 0 _1043_
rlabel metal2 15624 37520 15624 37520 0 _1044_
rlabel metal3 19376 36568 19376 36568 0 _1045_
rlabel metal3 22736 37240 22736 37240 0 _1046_
rlabel metal2 22568 37016 22568 37016 0 _1047_
rlabel metal2 20328 38808 20328 38808 0 _1048_
rlabel metal2 21168 38696 21168 38696 0 _1049_
rlabel metal2 15064 35336 15064 35336 0 _1050_
rlabel metal3 14784 38808 14784 38808 0 _1051_
rlabel metal2 2296 37352 2296 37352 0 _1052_
rlabel metal2 7112 37352 7112 37352 0 _1053_
rlabel metal2 6776 41104 6776 41104 0 _1054_
rlabel metal2 11480 39536 11480 39536 0 _1055_
rlabel metal2 15288 38080 15288 38080 0 _1056_
rlabel metal2 15400 38080 15400 38080 0 _1057_
rlabel metal2 17976 37128 17976 37128 0 _1058_
rlabel metal2 19768 39480 19768 39480 0 _1059_
rlabel metal2 16072 39088 16072 39088 0 _1060_
rlabel metal3 10248 39592 10248 39592 0 _1061_
rlabel metal2 10640 39592 10640 39592 0 _1062_
rlabel metal2 11144 40824 11144 40824 0 _1063_
rlabel metal2 11816 40824 11816 40824 0 _1064_
rlabel metal2 17080 38360 17080 38360 0 _1065_
rlabel metal2 15176 37576 15176 37576 0 _1066_
rlabel metal2 15512 38416 15512 38416 0 _1067_
rlabel metal2 22680 42448 22680 42448 0 _1068_
rlabel metal2 14280 42336 14280 42336 0 _1069_
rlabel metal3 8960 44184 8960 44184 0 _1070_
rlabel metal2 9688 41384 9688 41384 0 _1071_
rlabel metal3 11760 41160 11760 41160 0 _1072_
rlabel metal2 12376 41608 12376 41608 0 _1073_
rlabel metal2 6664 41328 6664 41328 0 _1074_
rlabel metal2 5936 41160 5936 41160 0 _1075_
rlabel metal2 5880 42896 5880 42896 0 _1076_
rlabel metal3 5768 44296 5768 44296 0 _1077_
rlabel metal2 3752 45192 3752 45192 0 _1078_
rlabel metal2 3080 47152 3080 47152 0 _1079_
rlabel metal2 2408 47152 2408 47152 0 _1080_
rlabel metal2 2688 47432 2688 47432 0 _1081_
rlabel metal2 3080 46312 3080 46312 0 _1082_
rlabel metal2 4200 46312 4200 46312 0 _1083_
rlabel metal2 6776 43456 6776 43456 0 _1084_
rlabel metal2 10920 40768 10920 40768 0 _1085_
rlabel metal2 16184 39984 16184 39984 0 _1086_
rlabel metal2 19208 39144 19208 39144 0 _1087_
rlabel metal3 20776 38808 20776 38808 0 _1088_
rlabel metal2 24584 37800 24584 37800 0 _1089_
rlabel metal2 24360 38780 24360 38780 0 _1090_
rlabel metal2 24584 38724 24584 38724 0 _1091_
rlabel metal2 26488 40040 26488 40040 0 _1092_
rlabel metal2 25816 43624 25816 43624 0 _1093_
rlabel metal2 26096 46872 26096 46872 0 _1094_
rlabel metal2 24584 50960 24584 50960 0 _1095_
rlabel metal2 27104 40936 27104 40936 0 _1096_
rlabel metal2 21896 37912 21896 37912 0 _1097_
rlabel metal2 23352 37912 23352 37912 0 _1098_
rlabel metal2 22792 40824 22792 40824 0 _1099_
rlabel metal2 21560 39872 21560 39872 0 _1100_
rlabel metal2 22120 42056 22120 42056 0 _1101_
rlabel metal2 18480 49000 18480 49000 0 _1102_
rlabel metal2 15624 39256 15624 39256 0 _1103_
rlabel metal2 17640 41104 17640 41104 0 _1104_
rlabel metal3 19656 41048 19656 41048 0 _1105_
rlabel metal2 19544 39984 19544 39984 0 _1106_
rlabel metal2 19208 43008 19208 43008 0 _1107_
rlabel metal2 9912 42280 9912 42280 0 _1108_
rlabel metal3 10304 39368 10304 39368 0 _1109_
rlabel metal2 5208 40824 5208 40824 0 _1110_
rlabel metal2 4760 39816 4760 39816 0 _1111_
rlabel metal2 6888 42728 6888 42728 0 _1112_
rlabel metal3 11760 41944 11760 41944 0 _1113_
rlabel metal2 10808 44352 10808 44352 0 _1114_
rlabel metal2 14056 42336 14056 42336 0 _1115_
rlabel metal2 13832 42336 13832 42336 0 _1116_
rlabel metal2 14616 41832 14616 41832 0 _1117_
rlabel metal2 17528 41552 17528 41552 0 _1118_
rlabel metal2 16744 45472 16744 45472 0 _1119_
rlabel metal2 15848 44576 15848 44576 0 _1120_
rlabel metal2 9856 44296 9856 44296 0 _1121_
rlabel metal2 11088 45080 11088 45080 0 _1122_
rlabel metal2 12152 44184 12152 44184 0 _1123_
rlabel metal2 8568 45584 8568 45584 0 _1124_
rlabel metal2 6944 45752 6944 45752 0 _1125_
rlabel metal2 4536 45808 4536 45808 0 _1126_
rlabel metal2 5096 45304 5096 45304 0 _1127_
rlabel metal3 6552 45080 6552 45080 0 _1128_
rlabel metal2 7672 47824 7672 47824 0 _1129_
rlabel metal2 15400 49448 15400 49448 0 _1130_
rlabel metal2 5096 48496 5096 48496 0 _1131_
rlabel metal2 3416 46928 3416 46928 0 _1132_
rlabel metal2 3976 47432 3976 47432 0 _1133_
rlabel metal2 3976 48048 3976 48048 0 _1134_
rlabel metal2 4536 48160 4536 48160 0 _1135_
rlabel metal2 8008 46256 8008 46256 0 _1136_
rlabel metal2 11368 45360 11368 45360 0 _1137_
rlabel metal2 17640 42560 17640 42560 0 _1138_
rlabel metal2 19656 41496 19656 41496 0 _1139_
rlabel metal2 20552 42336 20552 42336 0 _1140_
rlabel metal3 21224 42504 21224 42504 0 _1141_
rlabel metal3 18816 40488 18816 40488 0 _1142_
rlabel metal3 19992 40376 19992 40376 0 _1143_
rlabel metal2 13384 42056 13384 42056 0 _1144_
rlabel metal2 15680 42840 15680 42840 0 _1145_
rlabel metal2 19096 40712 19096 40712 0 _1146_
rlabel metal2 21784 40880 21784 40880 0 _1147_
rlabel metal2 23800 40656 23800 40656 0 _1148_
rlabel metal2 25592 40264 25592 40264 0 _1149_
rlabel metal2 25256 33824 25256 33824 0 _1150_
rlabel via2 29176 29848 29176 29848 0 _1151_
rlabel metal2 30184 32144 30184 32144 0 _1152_
rlabel metal2 31080 32200 31080 32200 0 _1153_
rlabel metal2 20776 31136 20776 31136 0 _1154_
rlabel metal2 21672 31360 21672 31360 0 _1155_
rlabel metal2 28616 30856 28616 30856 0 _1156_
rlabel metal2 29512 31304 29512 31304 0 _1157_
rlabel metal2 28392 31360 28392 31360 0 _1158_
rlabel metal2 29624 30912 29624 30912 0 _1159_
rlabel metal2 23016 34888 23016 34888 0 _1160_
rlabel metal2 21448 33320 21448 33320 0 _1161_
rlabel metal2 16632 30408 16632 30408 0 _1162_
rlabel metal2 22568 28560 22568 28560 0 _1163_
rlabel metal3 21560 29512 21560 29512 0 _1164_
rlabel metal2 20328 29848 20328 29848 0 _1165_
rlabel metal3 15120 30184 15120 30184 0 _1166_
rlabel metal2 25816 41048 25816 41048 0 _1167_
rlabel metal2 25928 40712 25928 40712 0 _1168_
rlabel metal2 26376 42224 26376 42224 0 _1169_
rlabel metal2 24248 41216 24248 41216 0 _1170_
rlabel metal2 22568 41216 22568 41216 0 _1171_
rlabel metal2 23240 41440 23240 41440 0 _1172_
rlabel metal2 24024 41664 24024 41664 0 _1173_
rlabel metal2 21672 43176 21672 43176 0 _1174_
rlabel metal3 19040 43400 19040 43400 0 _1175_
rlabel metal2 20440 43456 20440 43456 0 _1176_
rlabel metal2 20888 43064 20888 43064 0 _1177_
rlabel metal3 17080 45304 17080 45304 0 _1178_
rlabel metal3 9240 47320 9240 47320 0 _1179_
rlabel metal2 10920 45584 10920 45584 0 _1180_
rlabel metal2 11704 42000 11704 42000 0 _1181_
rlabel metal2 12376 44744 12376 44744 0 _1182_
rlabel metal2 12040 47544 12040 47544 0 _1183_
rlabel metal2 13832 45080 13832 45080 0 _1184_
rlabel metal2 16856 44128 16856 44128 0 _1185_
rlabel metal2 17976 47376 17976 47376 0 _1186_
rlabel metal2 14952 52416 14952 52416 0 _1187_
rlabel metal2 16408 47152 16408 47152 0 _1188_
rlabel metal2 11704 49168 11704 49168 0 _1189_
rlabel metal2 9800 47824 9800 47824 0 _1190_
rlabel metal2 10248 46928 10248 46928 0 _1191_
rlabel metal2 11480 48440 11480 48440 0 _1192_
rlabel metal2 7560 49896 7560 49896 0 _1193_
rlabel metal2 7112 50540 7112 50540 0 _1194_
rlabel metal2 6216 49056 6216 49056 0 _1195_
rlabel metal2 6888 50960 6888 50960 0 _1196_
rlabel metal2 7784 50904 7784 50904 0 _1197_
rlabel metal2 6048 47656 6048 47656 0 _1198_
rlabel metal2 8008 51688 8008 51688 0 _1199_
rlabel metal3 10920 48216 10920 48216 0 _1200_
rlabel metal2 17752 47600 17752 47600 0 _1201_
rlabel metal3 19824 43624 19824 43624 0 _1202_
rlabel metal2 23912 43960 23912 43960 0 _1203_
rlabel metal2 25816 42224 25816 42224 0 _1204_
rlabel metal3 25816 31752 25816 31752 0 _1205_
rlabel metal2 12152 33544 12152 33544 0 _1206_
rlabel metal2 17752 31416 17752 31416 0 _1207_
rlabel metal2 18088 30016 18088 30016 0 _1208_
rlabel metal2 16296 28280 16296 28280 0 _1209_
rlabel metal2 26936 43008 26936 43008 0 _1210_
rlabel metal2 24696 42728 24696 42728 0 _1211_
rlabel metal2 26264 42952 26264 42952 0 _1212_
rlabel metal2 26824 43176 26824 43176 0 _1213_
rlabel metal3 29008 43624 29008 43624 0 _1214_
rlabel metal2 21560 45808 21560 45808 0 _1215_
rlabel metal2 19880 44184 19880 44184 0 _1216_
rlabel metal2 19656 43736 19656 43736 0 _1217_
rlabel metal2 14280 44632 14280 44632 0 _1218_
rlabel metal2 15624 45976 15624 45976 0 _1219_
rlabel metal2 19432 44408 19432 44408 0 _1220_
rlabel metal3 20664 44296 20664 44296 0 _1221_
rlabel metal2 22512 44296 22512 44296 0 _1222_
rlabel metal2 23576 45920 23576 45920 0 _1223_
rlabel metal2 21896 50568 21896 50568 0 _1224_
rlabel metal2 22344 45752 22344 45752 0 _1225_
rlabel metal2 22792 46816 22792 46816 0 _1226_
rlabel metal2 19320 49392 19320 49392 0 _1227_
rlabel metal3 19264 47320 19264 47320 0 _1228_
rlabel metal2 21672 47376 21672 47376 0 _1229_
rlabel metal2 15624 47096 15624 47096 0 _1230_
rlabel metal2 11032 47768 11032 47768 0 _1231_
rlabel metal2 10808 46256 10808 46256 0 _1232_
rlabel metal2 12376 48608 12376 48608 0 _1233_
rlabel metal2 11816 50960 11816 50960 0 _1234_
rlabel metal2 13384 46984 13384 46984 0 _1235_
rlabel metal2 13832 47096 13832 47096 0 _1236_
rlabel metal2 15960 47936 15960 47936 0 _1237_
rlabel metal3 14952 52248 14952 52248 0 _1238_
rlabel metal2 8456 51408 8456 51408 0 _1239_
rlabel metal2 12040 50624 12040 50624 0 _1240_
rlabel metal2 12824 52808 12824 52808 0 _1241_
rlabel metal2 5992 50736 5992 50736 0 _1242_
rlabel metal2 10472 52528 10472 52528 0 _1243_
rlabel metal3 10808 51408 10808 51408 0 _1244_
rlabel metal2 12376 51296 12376 51296 0 _1245_
rlabel metal2 15960 51128 15960 51128 0 _1246_
rlabel metal3 19264 47432 19264 47432 0 _1247_
rlabel metal2 21784 47880 21784 47880 0 _1248_
rlabel metal2 22568 45864 22568 45864 0 _1249_
rlabel metal2 19600 46760 19600 46760 0 _1250_
rlabel metal2 20160 46648 20160 46648 0 _1251_
rlabel metal2 15176 49336 15176 49336 0 _1252_
rlabel metal3 15764 49000 15764 49000 0 _1253_
rlabel metal3 18088 46760 18088 46760 0 _1254_
rlabel metal3 22792 46648 22792 46648 0 _1255_
rlabel metal2 23744 45304 23744 45304 0 _1256_
rlabel metal2 25144 44688 25144 44688 0 _1257_
rlabel metal2 25256 31136 25256 31136 0 _1258_
rlabel metal3 30184 28616 30184 28616 0 _1259_
rlabel metal2 25704 26572 25704 26572 0 _1260_
rlabel metal2 30072 27440 30072 27440 0 _1261_
rlabel metal2 20776 29512 20776 29512 0 _1262_
rlabel metal2 21112 31304 21112 31304 0 _1263_
rlabel metal2 21448 31192 21448 31192 0 _1264_
rlabel metal2 20104 30464 20104 30464 0 _1265_
rlabel metal2 18312 30128 18312 30128 0 _1266_
rlabel metal3 15232 31752 15232 31752 0 _1267_
rlabel metal2 27496 43568 27496 43568 0 _1268_
rlabel metal2 28952 43456 28952 43456 0 _1269_
rlabel metal2 28280 44912 28280 44912 0 _1270_
rlabel metal2 27608 44744 27608 44744 0 _1271_
rlabel metal2 22456 46704 22456 46704 0 _1272_
rlabel metal2 23464 46928 23464 46928 0 _1273_
rlabel metal2 24248 48160 24248 48160 0 _1274_
rlabel metal2 22120 50456 22120 50456 0 _1275_
rlabel metal2 21672 50120 21672 50120 0 _1276_
rlabel metal2 20552 51352 20552 51352 0 _1277_
rlabel metal3 18312 48888 18312 48888 0 _1278_
rlabel metal3 21056 48440 21056 48440 0 _1279_
rlabel metal2 21000 48608 21000 48608 0 _1280_
rlabel metal3 24192 50568 24192 50568 0 _1281_
rlabel metal2 17976 50960 17976 50960 0 _1282_
rlabel metal2 13496 53312 13496 53312 0 _1283_
rlabel metal2 14280 52136 14280 52136 0 _1284_
rlabel metal2 13720 50848 13720 50848 0 _1285_
rlabel metal2 13944 51856 13944 51856 0 _1286_
rlabel metal3 20188 52136 20188 52136 0 _1287_
rlabel metal2 15736 51744 15736 51744 0 _1288_
rlabel metal2 11144 51856 11144 51856 0 _1289_
rlabel metal3 13776 52136 13776 52136 0 _1290_
rlabel metal2 17976 52584 17976 52584 0 _1291_
rlabel metal2 19320 51212 19320 51212 0 _1292_
rlabel metal2 24136 49336 24136 49336 0 _1293_
rlabel metal2 24808 46200 24808 46200 0 _1294_
rlabel metal2 26712 33208 26712 33208 0 _1295_
rlabel metal2 16744 30688 16744 30688 0 _1296_
rlabel metal3 15008 29400 15008 29400 0 _1297_
rlabel metal2 26544 31752 26544 31752 0 _1298_
rlabel metal2 26264 34552 26264 34552 0 _1299_
rlabel metal3 31472 32760 31472 32760 0 _1300_
rlabel metal2 26152 26628 26152 26628 0 _1301_
rlabel metal2 26936 45472 26936 45472 0 _1302_
rlabel metal2 27776 45304 27776 45304 0 _1303_
rlabel metal2 27384 47096 27384 47096 0 _1304_
rlabel metal2 22624 48440 22624 48440 0 _1305_
rlabel metal2 27048 47712 27048 47712 0 _1306_
rlabel metal2 24584 52920 24584 52920 0 _1307_
rlabel metal2 19992 49504 19992 49504 0 _1308_
rlabel metal2 19600 46536 19600 46536 0 _1309_
rlabel metal2 19208 50456 19208 50456 0 _1310_
rlabel metal2 21896 51968 21896 51968 0 _1311_
rlabel metal2 21896 49056 21896 49056 0 _1312_
rlabel metal2 23464 49000 23464 49000 0 _1313_
rlabel metal2 24248 51352 24248 51352 0 _1314_
rlabel metal2 23352 51464 23352 51464 0 _1315_
rlabel metal2 19992 51464 19992 51464 0 _1316_
rlabel metal2 21672 51800 21672 51800 0 _1317_
rlabel metal2 22120 52192 22120 52192 0 _1318_
rlabel metal2 20664 52472 20664 52472 0 _1319_
rlabel metal2 16744 52248 16744 52248 0 _1320_
rlabel metal2 21336 53200 21336 53200 0 _1321_
rlabel metal2 22680 53424 22680 53424 0 _1322_
rlabel metal2 24416 52136 24416 52136 0 _1323_
rlabel metal2 26824 48440 26824 48440 0 _1324_
rlabel metal2 25312 39144 25312 39144 0 _1325_
rlabel metal3 20664 35560 20664 35560 0 _1326_
rlabel metal2 24248 35168 24248 35168 0 _1327_
rlabel metal3 25200 34328 25200 34328 0 _1328_
rlabel metal2 23240 30688 23240 30688 0 _1329_
rlabel metal2 27944 37632 27944 37632 0 _1330_
rlabel metal2 26712 34384 26712 34384 0 _1331_
rlabel metal2 19600 34888 19600 34888 0 _1332_
rlabel metal3 26544 46648 26544 46648 0 _1333_
rlabel metal2 26376 47376 26376 47376 0 _1334_
rlabel metal2 26656 46872 26656 46872 0 _1335_
rlabel metal2 25816 49840 25816 49840 0 _1336_
rlabel metal2 21336 52304 21336 52304 0 _1337_
rlabel metal3 22344 51912 22344 51912 0 _1338_
rlabel metal2 22568 52808 22568 52808 0 _1339_
rlabel metal2 26040 52248 26040 52248 0 _1340_
rlabel metal2 22008 52976 22008 52976 0 _1341_
rlabel metal2 24808 53424 24808 53424 0 _1342_
rlabel metal2 22008 51352 22008 51352 0 _1343_
rlabel metal2 23912 53088 23912 53088 0 _1344_
rlabel metal2 26264 53256 26264 53256 0 _1345_
rlabel metal2 26600 52024 26600 52024 0 _1346_
rlabel metal2 20440 34944 20440 34944 0 _1347_
rlabel metal2 20552 33936 20552 33936 0 _1348_
rlabel metal2 20664 33264 20664 33264 0 _1349_
rlabel metal2 19544 33600 19544 33600 0 _1350_
rlabel metal2 26824 49336 26824 49336 0 _1351_
rlabel metal2 28168 49000 28168 49000 0 _1352_
rlabel metal2 27608 50960 27608 50960 0 _1353_
rlabel metal3 25200 51464 25200 51464 0 _1354_
rlabel metal2 25704 53200 25704 53200 0 _1355_
rlabel via2 26376 52136 26376 52136 0 _1356_
rlabel metal2 26040 50960 26040 50960 0 _1357_
rlabel metal2 23128 36792 23128 36792 0 _1358_
rlabel metal2 27720 36008 27720 36008 0 _1359_
rlabel metal2 28168 36064 28168 36064 0 _1360_
rlabel metal2 29960 36456 29960 36456 0 _1361_
rlabel metal2 27048 50848 27048 50848 0 _1362_
rlabel metal2 26768 50568 26768 50568 0 _1363_
rlabel metal2 26376 29008 26376 29008 0 _1364_
rlabel metal2 25144 37352 25144 37352 0 _1365_
rlabel metal2 25928 37576 25928 37576 0 _1366_
rlabel metal2 26712 37128 26712 37128 0 _1367_
rlabel metal2 27496 37240 27496 37240 0 _1368_
rlabel metal2 23688 25760 23688 25760 0 _1369_
rlabel metal2 25480 31976 25480 31976 0 _1370_
rlabel metal2 37240 31640 37240 31640 0 _1371_
rlabel metal3 30968 21448 30968 21448 0 _1372_
rlabel metal2 33880 15848 33880 15848 0 _1373_
rlabel metal3 37464 18536 37464 18536 0 _1374_
rlabel metal2 39536 21784 39536 21784 0 _1375_
rlabel metal2 39928 24192 39928 24192 0 _1376_
rlabel metal2 46088 22400 46088 22400 0 _1377_
rlabel metal2 41944 17248 41944 17248 0 _1378_
rlabel metal2 39144 18704 39144 18704 0 _1379_
rlabel metal3 44184 15960 44184 15960 0 _1380_
rlabel metal2 42952 12096 42952 12096 0 _1381_
rlabel metal3 39144 3192 39144 3192 0 _1382_
rlabel metal2 31752 8288 31752 8288 0 _1383_
rlabel metal2 32256 9016 32256 9016 0 _1384_
rlabel metal2 31864 8736 31864 8736 0 _1385_
rlabel metal3 39760 3304 39760 3304 0 _1386_
rlabel metal2 32760 6608 32760 6608 0 _1387_
rlabel metal3 42504 4312 42504 4312 0 _1388_
rlabel metal2 39144 4144 39144 4144 0 _1389_
rlabel metal2 38920 4256 38920 4256 0 _1390_
rlabel metal2 35896 5488 35896 5488 0 _1391_
rlabel metal2 33096 10136 33096 10136 0 _1392_
rlabel metal3 31920 17640 31920 17640 0 _1393_
rlabel metal2 32200 9800 32200 9800 0 _1394_
rlabel metal3 44352 8344 44352 8344 0 _1395_
rlabel metal2 34888 10248 34888 10248 0 _1396_
rlabel metal2 32984 10640 32984 10640 0 _1397_
rlabel metal2 31192 8512 31192 8512 0 _1398_
rlabel metal2 36568 9800 36568 9800 0 _1399_
rlabel metal2 39256 4760 39256 4760 0 _1400_
rlabel metal3 35952 7224 35952 7224 0 _1401_
rlabel metal2 33992 4368 33992 4368 0 _1402_
rlabel metal2 37800 5208 37800 5208 0 _1403_
rlabel metal2 32872 8456 32872 8456 0 _1404_
rlabel metal2 33544 9464 33544 9464 0 _1405_
rlabel metal2 32424 12544 32424 12544 0 _1406_
rlabel metal3 33432 15288 33432 15288 0 _1407_
rlabel metal2 36344 12320 36344 12320 0 _1408_
rlabel metal2 34104 11032 34104 11032 0 _1409_
rlabel metal3 37296 7448 37296 7448 0 _1410_
rlabel metal2 33768 9296 33768 9296 0 _1411_
rlabel metal2 33992 9184 33992 9184 0 _1412_
rlabel metal2 34384 9240 34384 9240 0 _1413_
rlabel metal2 37464 10584 37464 10584 0 _1414_
rlabel metal2 40712 6888 40712 6888 0 _1415_
rlabel metal2 39256 9912 39256 9912 0 _1416_
rlabel metal2 35000 5096 35000 5096 0 _1417_
rlabel metal2 36120 6216 36120 6216 0 _1418_
rlabel metal3 36568 6776 36568 6776 0 _1419_
rlabel metal3 36792 8344 36792 8344 0 _1420_
rlabel metal2 39368 5656 39368 5656 0 _1421_
rlabel metal3 43400 12432 43400 12432 0 _1422_
rlabel metal2 39592 4760 39592 4760 0 _1423_
rlabel metal2 38696 6440 38696 6440 0 _1424_
rlabel metal2 38136 10472 38136 10472 0 _1425_
rlabel metal2 35672 13664 35672 13664 0 _1426_
rlabel metal2 34384 15176 34384 15176 0 _1427_
rlabel metal3 36792 16072 36792 16072 0 _1428_
rlabel metal2 35056 16184 35056 16184 0 _1429_
rlabel metal2 35112 14000 35112 14000 0 _1430_
rlabel metal2 37800 14000 37800 14000 0 _1431_
rlabel metal2 34048 15400 34048 15400 0 _1432_
rlabel metal3 33768 13944 33768 13944 0 _1433_
rlabel metal2 38360 14560 38360 14560 0 _1434_
rlabel metal3 36960 11256 36960 11256 0 _1435_
rlabel metal2 41384 6048 41384 6048 0 _1436_
rlabel metal3 39424 9128 39424 9128 0 _1437_
rlabel metal2 40040 9912 40040 9912 0 _1438_
rlabel metal2 38836 10584 38836 10584 0 _1439_
rlabel metal2 41496 9632 41496 9632 0 _1440_
rlabel metal2 42952 7336 42952 7336 0 _1441_
rlabel metal2 43176 8400 43176 8400 0 _1442_
rlabel metal2 44632 5936 44632 5936 0 _1443_
rlabel metal2 45192 5152 45192 5152 0 _1444_
rlabel metal2 47096 9912 47096 9912 0 _1445_
rlabel metal3 42728 4200 42728 4200 0 _1446_
rlabel metal2 39032 7056 39032 7056 0 _1447_
rlabel metal2 41048 6048 41048 6048 0 _1448_
rlabel metal2 40600 5824 40600 5824 0 _1449_
rlabel metal2 40936 8960 40936 8960 0 _1450_
rlabel metal2 39872 13496 39872 13496 0 _1451_
rlabel metal2 37296 16632 37296 16632 0 _1452_
rlabel metal2 37464 17360 37464 17360 0 _1453_
rlabel metal2 37352 18760 37352 18760 0 _1454_
rlabel metal2 38696 22456 38696 22456 0 _1455_
rlabel metal2 41384 17976 41384 17976 0 _1456_
rlabel metal2 34720 16632 34720 16632 0 _1457_
rlabel metal3 37576 15288 37576 15288 0 _1458_
rlabel metal2 39480 15568 39480 15568 0 _1459_
rlabel metal2 41160 15680 41160 15680 0 _1460_
rlabel metal2 41832 16072 41832 16072 0 _1461_
rlabel metal3 40992 16744 40992 16744 0 _1462_
rlabel metal2 39368 12320 39368 12320 0 _1463_
rlabel metal3 33712 9800 33712 9800 0 _1464_
rlabel metal2 36120 9464 36120 9464 0 _1465_
rlabel metal3 37240 9576 37240 9576 0 _1466_
rlabel metal2 38808 9408 38808 9408 0 _1467_
rlabel metal2 39480 10080 39480 10080 0 _1468_
rlabel metal2 41160 10192 41160 10192 0 _1469_
rlabel metal2 40264 11816 40264 11816 0 _1470_
rlabel metal2 41496 12208 41496 12208 0 _1471_
rlabel metal3 40824 13608 40824 13608 0 _1472_
rlabel metal2 42504 13832 42504 13832 0 _1473_
rlabel metal2 40600 10192 40600 10192 0 _1474_
rlabel metal2 41944 5992 41944 5992 0 _1475_
rlabel metal3 40600 8232 40600 8232 0 _1476_
rlabel metal3 41944 7448 41944 7448 0 _1477_
rlabel metal2 40376 7168 40376 7168 0 _1478_
rlabel metal2 43960 9184 43960 9184 0 _1479_
rlabel metal2 42448 8456 42448 8456 0 _1480_
rlabel metal2 45976 5768 45976 5768 0 _1481_
rlabel metal2 46088 5376 46088 5376 0 _1482_
rlabel metal2 47488 5096 47488 5096 0 _1483_
rlabel metal2 45416 5544 45416 5544 0 _1484_
rlabel metal2 42728 6720 42728 6720 0 _1485_
rlabel metal2 41608 8288 41608 8288 0 _1486_
rlabel metal2 41720 11872 41720 11872 0 _1487_
rlabel metal2 41496 16800 41496 16800 0 _1488_
rlabel metal3 39816 17640 39816 17640 0 _1489_
rlabel metal2 39032 21672 39032 21672 0 _1490_
rlabel via2 40040 22120 40040 22120 0 _1491_
rlabel metal2 39480 20720 39480 20720 0 _1492_
rlabel metal2 42280 18032 42280 18032 0 _1493_
rlabel metal3 42504 17584 42504 17584 0 _1494_
rlabel metal2 37856 18312 37856 18312 0 _1495_
rlabel metal3 38808 17696 38808 17696 0 _1496_
rlabel metal3 40712 19992 40712 19992 0 _1497_
rlabel metal2 41608 16520 41608 16520 0 _1498_
rlabel metal2 40152 12656 40152 12656 0 _1499_
rlabel metal3 39144 12824 39144 12824 0 _1500_
rlabel metal2 43064 14056 43064 14056 0 _1501_
rlabel metal2 41384 9072 41384 9072 0 _1502_
rlabel metal2 41048 9184 41048 9184 0 _1503_
rlabel metal2 41944 11872 41944 11872 0 _1504_
rlabel metal3 42896 13496 42896 13496 0 _1505_
rlabel metal2 43624 15232 43624 15232 0 _1506_
rlabel metal2 44128 16072 44128 16072 0 _1507_
rlabel metal2 43400 16296 43400 16296 0 _1508_
rlabel metal3 46312 12264 46312 12264 0 _1509_
rlabel metal2 44072 11032 44072 11032 0 _1510_
rlabel metal2 43400 14616 43400 14616 0 _1511_
rlabel metal2 43176 13944 43176 13944 0 _1512_
rlabel metal2 48496 19208 48496 19208 0 _1513_
rlabel metal2 46760 11312 46760 11312 0 _1514_
rlabel metal2 46424 6216 46424 6216 0 _1515_
rlabel metal3 42896 8120 42896 8120 0 _1516_
rlabel metal2 43848 8064 43848 8064 0 _1517_
rlabel metal2 44296 8736 44296 8736 0 _1518_
rlabel metal2 44856 8960 44856 8960 0 _1519_
rlabel metal3 46648 9128 46648 9128 0 _1520_
rlabel metal2 48328 8232 48328 8232 0 _1521_
rlabel metal2 46872 6272 46872 6272 0 _1522_
rlabel metal2 49168 8344 49168 8344 0 _1523_
rlabel metal2 50344 5320 50344 5320 0 _1524_
rlabel metal2 51464 6608 51464 6608 0 _1525_
rlabel metal2 50008 5768 50008 5768 0 _1526_
rlabel metal2 47208 7896 47208 7896 0 _1527_
rlabel metal2 47488 10584 47488 10584 0 _1528_
rlabel metal2 44744 13160 44744 13160 0 _1529_
rlabel metal2 43064 17640 43064 17640 0 _1530_
rlabel metal2 42392 19936 42392 19936 0 _1531_
rlabel metal2 41328 22232 41328 22232 0 _1532_
rlabel metal2 39984 23240 39984 23240 0 _1533_
rlabel metal2 40600 25480 40600 25480 0 _1534_
rlabel metal2 41440 23128 41440 23128 0 _1535_
rlabel metal2 41496 24024 41496 24024 0 _1536_
rlabel metal2 40376 21000 40376 21000 0 _1537_
rlabel metal2 40936 20832 40936 20832 0 _1538_
rlabel metal2 41832 22008 41832 22008 0 _1539_
rlabel metal2 43736 21672 43736 21672 0 _1540_
rlabel metal2 43064 23464 43064 23464 0 _1541_
rlabel metal2 43624 21840 43624 21840 0 _1542_
rlabel metal3 42896 19208 42896 19208 0 _1543_
rlabel metal2 42784 18312 42784 18312 0 _1544_
rlabel metal2 45192 19152 45192 19152 0 _1545_
rlabel metal3 44296 18984 44296 18984 0 _1546_
rlabel metal2 44296 17248 44296 17248 0 _1547_
rlabel metal2 46200 18368 46200 18368 0 _1548_
rlabel metal2 45080 12656 45080 12656 0 _1549_
rlabel metal2 41944 13160 41944 13160 0 _1550_
rlabel metal2 44968 8680 44968 8680 0 _1551_
rlabel metal2 42616 9016 42616 9016 0 _1552_
rlabel metal3 46424 10584 46424 10584 0 _1553_
rlabel metal2 46312 11816 46312 11816 0 _1554_
rlabel metal2 45752 13776 45752 13776 0 _1555_
rlabel metal3 44352 14504 44352 14504 0 _1556_
rlabel metal3 46872 15288 46872 15288 0 _1557_
rlabel metal2 47320 16464 47320 16464 0 _1558_
rlabel metal3 49168 15960 49168 15960 0 _1559_
rlabel metal2 47544 11760 47544 11760 0 _1560_
rlabel metal2 48776 12768 48776 12768 0 _1561_
rlabel metal2 49224 16352 49224 16352 0 _1562_
rlabel metal2 49560 20272 49560 20272 0 _1563_
rlabel metal2 49672 12432 49672 12432 0 _1564_
rlabel metal3 48216 8792 48216 8792 0 _1565_
rlabel metal2 48776 8232 48776 8232 0 _1566_
rlabel metal3 48552 9240 48552 9240 0 _1567_
rlabel metal2 49896 10976 49896 10976 0 _1568_
rlabel metal2 51240 9296 51240 9296 0 _1569_
rlabel metal3 48552 6552 48552 6552 0 _1570_
rlabel metal2 53704 9856 53704 9856 0 _1571_
rlabel metal2 50848 6776 50848 6776 0 _1572_
rlabel metal2 51016 8064 51016 8064 0 _1573_
rlabel metal2 52472 7504 52472 7504 0 _1574_
rlabel metal2 50120 10136 50120 10136 0 _1575_
rlabel metal2 48440 12264 48440 12264 0 _1576_
rlabel metal3 46368 18424 46368 18424 0 _1577_
rlabel metal2 44968 18816 44968 18816 0 _1578_
rlabel metal3 45640 20664 45640 20664 0 _1579_
rlabel metal2 45080 21224 45080 21224 0 _1580_
rlabel metal2 42952 20132 42952 20132 0 _1581_
rlabel metal3 43400 19992 43400 19992 0 _1582_
rlabel metal2 49224 11368 49224 11368 0 _1583_
rlabel metal3 48328 15288 48328 15288 0 _1584_
rlabel metal2 46480 16296 46480 16296 0 _1585_
rlabel metal2 44184 19432 44184 19432 0 _1586_
rlabel metal2 43400 20328 43400 20328 0 _1587_
rlabel metal3 43736 22344 43736 22344 0 _1588_
rlabel metal2 41944 23184 41944 23184 0 _1589_
rlabel metal2 41552 24696 41552 24696 0 _1590_
rlabel metal3 34160 25480 34160 25480 0 _1591_
rlabel metal2 33600 24808 33600 24808 0 _1592_
rlabel metal2 33096 24976 33096 24976 0 _1593_
rlabel metal2 32368 30184 32368 30184 0 _1594_
rlabel metal2 32536 25928 32536 25928 0 _1595_
rlabel metal2 32648 25424 32648 25424 0 _1596_
rlabel metal2 33096 25760 33096 25760 0 _1597_
rlabel metal2 33544 34160 33544 34160 0 _1598_
rlabel metal2 30856 33208 30856 33208 0 _1599_
rlabel metal2 31528 33320 31528 33320 0 _1600_
rlabel metal2 25480 33880 25480 33880 0 _1601_
rlabel metal2 40376 29736 40376 29736 0 _1602_
rlabel metal2 42952 30632 42952 30632 0 _1603_
rlabel metal2 41720 25032 41720 25032 0 _1604_
rlabel metal3 41832 24696 41832 24696 0 _1605_
rlabel metal3 42952 26264 42952 26264 0 _1606_
rlabel metal2 44296 24304 44296 24304 0 _1607_
rlabel metal2 43960 21616 43960 21616 0 _1608_
rlabel metal2 44072 21280 44072 21280 0 _1609_
rlabel metal2 46312 23352 46312 23352 0 _1610_
rlabel metal3 46928 22344 46928 22344 0 _1611_
rlabel metal2 46928 19320 46928 19320 0 _1612_
rlabel metal2 46144 20664 46144 20664 0 _1613_
rlabel metal2 46088 21224 46088 21224 0 _1614_
rlabel metal2 48888 18424 48888 18424 0 _1615_
rlabel metal2 50792 14840 50792 14840 0 _1616_
rlabel metal2 48328 14224 48328 14224 0 _1617_
rlabel metal2 49112 18032 49112 18032 0 _1618_
rlabel metal2 50232 15904 50232 15904 0 _1619_
rlabel metal2 50848 15288 50848 15288 0 _1620_
rlabel metal2 50008 15792 50008 15792 0 _1621_
rlabel metal2 49896 14392 49896 14392 0 _1622_
rlabel metal2 50232 14448 50232 14448 0 _1623_
rlabel metal2 53592 12544 53592 12544 0 _1624_
rlabel metal2 49840 9128 49840 9128 0 _1625_
rlabel metal2 53144 8344 53144 8344 0 _1626_
rlabel metal3 53648 10808 53648 10808 0 _1627_
rlabel metal2 54040 10304 54040 10304 0 _1628_
rlabel metal2 53256 11704 53256 11704 0 _1629_
rlabel metal2 51464 7784 51464 7784 0 _1630_
rlabel metal2 49672 8288 49672 8288 0 _1631_
rlabel metal3 52024 8344 52024 8344 0 _1632_
rlabel metal3 52864 8232 52864 8232 0 _1633_
rlabel metal3 52248 9016 52248 9016 0 _1634_
rlabel metal2 52920 10360 52920 10360 0 _1635_
rlabel metal2 51296 15848 51296 15848 0 _1636_
rlabel metal2 50344 17976 50344 17976 0 _1637_
rlabel metal2 47320 19656 47320 19656 0 _1638_
rlabel metal2 47432 22624 47432 22624 0 _1639_
rlabel metal2 44184 24304 44184 24304 0 _1640_
rlabel metal3 44072 26152 44072 26152 0 _1641_
rlabel metal2 42840 26600 42840 26600 0 _1642_
rlabel metal3 34608 17640 34608 17640 0 _1643_
rlabel metal2 32760 18368 32760 18368 0 _1644_
rlabel metal2 20552 26152 20552 26152 0 _1645_
rlabel metal2 26600 32032 26600 32032 0 _1646_
rlabel metal2 25816 32256 25816 32256 0 _1647_
rlabel metal2 24024 32424 24024 32424 0 _1648_
rlabel metal2 45192 25872 45192 25872 0 _1649_
rlabel metal3 45472 26936 45472 26936 0 _1650_
rlabel metal3 49280 25480 49280 25480 0 _1651_
rlabel metal2 45976 25760 45976 25760 0 _1652_
rlabel metal2 47040 20552 47040 20552 0 _1653_
rlabel metal2 48888 19600 48888 19600 0 _1654_
rlabel metal2 48440 20328 48440 20328 0 _1655_
rlabel metal2 49336 19096 49336 19096 0 _1656_
rlabel metal2 48776 20160 48776 20160 0 _1657_
rlabel metal2 48048 22120 48048 22120 0 _1658_
rlabel metal2 50008 23576 50008 23576 0 _1659_
rlabel metal2 49728 24584 49728 24584 0 _1660_
rlabel metal2 50232 23520 50232 23520 0 _1661_
rlabel metal3 49560 24696 49560 24696 0 _1662_
rlabel metal3 55440 20664 55440 20664 0 _1663_
rlabel metal2 51352 20664 51352 20664 0 _1664_
rlabel metal2 51688 21056 51688 21056 0 _1665_
rlabel metal3 54320 19096 54320 19096 0 _1666_
rlabel metal3 52528 13496 52528 13496 0 _1667_
rlabel metal3 52248 14616 52248 14616 0 _1668_
rlabel metal2 52808 15008 52808 15008 0 _1669_
rlabel metal2 51688 15960 51688 15960 0 _1670_
rlabel metal2 52136 23968 52136 23968 0 _1671_
rlabel metal2 54096 15960 54096 15960 0 _1672_
rlabel metal2 53704 11760 53704 11760 0 _1673_
rlabel metal2 53704 13440 53704 13440 0 _1674_
rlabel metal2 53816 15148 53816 15148 0 _1675_
rlabel metal2 55720 20412 55720 20412 0 _1676_
rlabel metal2 54824 13384 54824 13384 0 _1677_
rlabel metal2 54208 10808 54208 10808 0 _1678_
rlabel metal2 54600 12432 54600 12432 0 _1679_
rlabel metal2 55160 15288 55160 15288 0 _1680_
rlabel metal3 55496 18312 55496 18312 0 _1681_
rlabel metal2 53368 17416 53368 17416 0 _1682_
rlabel metal2 52024 21840 52024 21840 0 _1683_
rlabel metal2 50344 24248 50344 24248 0 _1684_
rlabel metal2 50568 21000 50568 21000 0 _1685_
rlabel metal3 49448 20552 49448 20552 0 _1686_
rlabel metal2 50120 20328 50120 20328 0 _1687_
rlabel metal2 50456 21616 50456 21616 0 _1688_
rlabel metal2 50008 22792 50008 22792 0 _1689_
rlabel metal3 47936 25368 47936 25368 0 _1690_
rlabel metal2 45472 27720 45472 27720 0 _1691_
rlabel metal2 44520 28672 44520 28672 0 _1692_
rlabel metal2 34888 24416 34888 24416 0 _1693_
rlabel metal2 25816 30520 25816 30520 0 _1694_
rlabel metal3 24976 31080 24976 31080 0 _1695_
rlabel metal2 23576 29904 23576 29904 0 _1696_
rlabel metal2 37576 25592 37576 25592 0 _1697_
rlabel metal2 32704 35896 32704 35896 0 _1698_
rlabel metal3 22848 29960 22848 29960 0 _1699_
rlabel metal2 33936 35560 33936 35560 0 _1700_
rlabel metal2 34664 15736 34664 15736 0 _1701_
rlabel metal2 33488 26152 33488 26152 0 _1702_
rlabel metal3 34776 28504 34776 28504 0 _1703_
rlabel metal2 46984 26236 46984 26236 0 _1704_
rlabel metal3 47320 27048 47320 27048 0 _1705_
rlabel metal2 49784 25312 49784 25312 0 _1706_
rlabel metal3 48944 26264 48944 26264 0 _1707_
rlabel metal2 50568 23184 50568 23184 0 _1708_
rlabel metal2 50904 23408 50904 23408 0 _1709_
rlabel metal2 51128 22568 51128 22568 0 _1710_
rlabel metal2 49784 21952 49784 21952 0 _1711_
rlabel metal2 52304 22344 52304 22344 0 _1712_
rlabel metal3 53760 18536 53760 18536 0 _1713_
rlabel metal2 53032 20552 53032 20552 0 _1714_
rlabel metal2 51688 22680 51688 22680 0 _1715_
rlabel metal2 56728 19712 56728 19712 0 _1716_
rlabel metal2 56840 15204 56840 15204 0 _1717_
rlabel metal3 56112 15176 56112 15176 0 _1718_
rlabel metal2 56616 15680 56616 15680 0 _1719_
rlabel metal2 55384 15652 55384 15652 0 _1720_
rlabel metal2 56168 15792 56168 15792 0 _1721_
rlabel metal3 56504 16968 56504 16968 0 _1722_
rlabel metal3 56168 16856 56168 16856 0 _1723_
rlabel metal2 55720 13944 55720 13944 0 _1724_
rlabel metal2 55720 16352 55720 16352 0 _1725_
rlabel metal2 57848 16520 57848 16520 0 _1726_
rlabel metal2 53592 20496 53592 20496 0 _1727_
rlabel metal3 53480 23352 53480 23352 0 _1728_
rlabel metal2 47992 25536 47992 25536 0 _1729_
rlabel metal2 45976 27440 45976 27440 0 _1730_
rlabel metal2 32872 27104 32872 27104 0 _1731_
rlabel metal2 32536 27104 32536 27104 0 _1732_
rlabel metal2 30632 34160 30632 34160 0 _1733_
rlabel metal2 32536 35336 32536 35336 0 _1734_
rlabel metal2 47656 26600 47656 26600 0 _1735_
rlabel metal2 47600 25480 47600 25480 0 _1736_
rlabel metal3 49000 26936 49000 26936 0 _1737_
rlabel metal2 50344 25592 50344 25592 0 _1738_
rlabel metal2 47768 23632 47768 23632 0 _1739_
rlabel metal2 54936 19432 54936 19432 0 _1740_
rlabel metal2 51184 19992 51184 19992 0 _1741_
rlabel metal2 55104 19992 55104 19992 0 _1742_
rlabel metal3 55720 21560 55720 21560 0 _1743_
rlabel metal2 53368 22288 53368 22288 0 _1744_
rlabel metal2 54488 22624 54488 22624 0 _1745_
rlabel metal2 57176 22232 57176 22232 0 _1746_
rlabel metal3 54600 23800 54600 23800 0 _1747_
rlabel metal2 56728 18536 56728 18536 0 _1748_
rlabel metal2 56728 21728 56728 21728 0 _1749_
rlabel metal2 56168 24808 56168 24808 0 _1750_
rlabel metal2 56896 20776 56896 20776 0 _1751_
rlabel metal2 56392 16856 56392 16856 0 _1752_
rlabel metal2 57064 20720 57064 20720 0 _1753_
rlabel metal2 56728 23632 56728 23632 0 _1754_
rlabel metal2 57400 23464 57400 23464 0 _1755_
rlabel metal2 49448 26040 49448 26040 0 _1756_
rlabel metal2 49112 26880 49112 26880 0 _1757_
rlabel metal2 48776 28056 48776 28056 0 _1758_
rlabel metal2 34552 17920 34552 17920 0 _1759_
rlabel metal2 35168 24696 35168 24696 0 _1760_
rlabel metal2 31360 23128 31360 23128 0 _1761_
rlabel metal3 39844 28616 39844 28616 0 _1762_
rlabel metal2 26488 26992 26488 26992 0 _1763_
rlabel metal2 32536 30128 32536 30128 0 _1764_
rlabel metal2 27608 29344 27608 29344 0 _1765_
rlabel metal2 27160 29456 27160 29456 0 _1766_
rlabel metal2 40600 30296 40600 30296 0 active
rlabel metal2 24752 29624 24752 29624 0 clk
rlabel metal2 26824 32088 26824 32088 0 clknet_0_clk
rlabel metal2 24304 25480 24304 25480 0 clknet_2_0__leaf_clk
rlabel metal2 26096 39032 26096 39032 0 clknet_2_1__leaf_clk
rlabel metal3 39704 25256 39704 25256 0 clknet_2_2__leaf_clk
rlabel metal3 39144 35056 39144 35056 0 clknet_2_3__leaf_clk
rlabel metal3 1680 11256 1680 11256 0 net1
rlabel metal2 2800 28056 2800 28056 0 net10
rlabel metal2 37688 35504 37688 35504 0 net100
rlabel metal2 39648 45640 39648 45640 0 net101
rlabel metal2 27496 53032 27496 53032 0 net102
rlabel metal2 39928 31640 39928 31640 0 net103
rlabel metal2 39928 28168 39928 28168 0 net104
rlabel metal2 17416 31136 17416 31136 0 net105
rlabel metal3 45136 28504 45136 28504 0 net106
rlabel metal3 42504 26488 42504 26488 0 net107
rlabel metal2 13496 29344 13496 29344 0 net108
rlabel metal2 27888 54376 27888 54376 0 net109
rlabel metal2 2016 12376 2016 12376 0 net11
rlabel metal2 17640 34552 17640 34552 0 net110
rlabel metal3 31584 54376 31584 54376 0 net111
rlabel metal3 30632 53816 30632 53816 0 net112
rlabel metal2 21784 34160 21784 34160 0 net113
rlabel metal2 21728 32424 21728 32424 0 net114
rlabel metal2 42784 30968 42784 30968 0 net115
rlabel metal3 43176 29792 43176 29792 0 net116
rlabel metal2 18984 39480 18984 39480 0 net117
rlabel metal2 19544 2030 19544 2030 0 net118
rlabel metal3 20944 39480 20944 39480 0 net119
rlabel metal2 2072 18368 2072 18368 0 net12
rlabel metal2 19656 29232 19656 29232 0 net13
rlabel metal2 2800 12824 2800 12824 0 net14
rlabel metal2 2072 16296 2072 16296 0 net15
rlabel metal2 2744 26544 2744 26544 0 net16
rlabel metal4 2072 21560 2072 21560 0 net17
rlabel metal3 1680 39368 1680 39368 0 net18
rlabel metal2 42952 5432 42952 5432 0 net19
rlabel metal2 24752 51688 24752 51688 0 net2
rlabel metal2 39032 4032 39032 4032 0 net20
rlabel metal2 45640 4648 45640 4648 0 net21
rlabel metal3 44800 4424 44800 4424 0 net22
rlabel metal2 48104 5040 48104 5040 0 net23
rlabel metal2 50232 4648 50232 4648 0 net24
rlabel metal2 2856 23576 2856 23576 0 net25
rlabel metal2 2296 22960 2296 22960 0 net26
rlabel metal4 2856 17136 2856 17136 0 net27
rlabel metal3 3304 21504 3304 21504 0 net28
rlabel metal3 7448 40936 7448 40936 0 net29
rlabel metal2 27160 52472 27160 52472 0 net3
rlabel metal2 2744 14532 2744 14532 0 net30
rlabel metal2 2968 15176 2968 15176 0 net31
rlabel metal2 2072 10864 2072 10864 0 net32
rlabel metal2 7112 8680 7112 8680 0 net33
rlabel metal2 30072 53200 30072 53200 0 net34
rlabel metal2 30128 52136 30128 52136 0 net35
rlabel metal2 30968 53592 30968 53592 0 net36
rlabel metal2 31752 53816 31752 53816 0 net37
rlabel metal2 37296 52136 37296 52136 0 net38
rlabel metal2 37464 52080 37464 52080 0 net39
rlabel metal2 29120 54824 29120 54824 0 net4
rlabel metal2 2408 32088 2408 32088 0 net40
rlabel metal2 50288 52136 50288 52136 0 net41
rlabel metal2 51352 51464 51352 51464 0 net42
rlabel metal2 2520 32872 2520 32872 0 net43
rlabel metal2 2072 42952 2072 42952 0 net44
rlabel metal3 3192 44408 3192 44408 0 net45
rlabel metal2 2072 45752 2072 45752 0 net46
rlabel metal2 4872 49672 4872 49672 0 net47
rlabel metal2 32200 4816 32200 4816 0 net48
rlabel metal3 29568 4872 29568 4872 0 net49
rlabel metal2 18200 26572 18200 26572 0 net5
rlabel metal2 1736 35504 1736 35504 0 net50
rlabel metal3 40488 7000 40488 7000 0 net51
rlabel metal2 44744 5096 44744 5096 0 net52
rlabel metal3 40152 16856 40152 16856 0 net53
rlabel metal3 43344 19320 43344 19320 0 net54
rlabel metal2 42504 21392 42504 21392 0 net55
rlabel metal2 45416 24808 45416 24808 0 net56
rlabel metal2 2128 23912 2128 23912 0 net57
rlabel metal2 2128 17080 2128 17080 0 net58
rlabel metal2 2744 18480 2744 18480 0 net59
rlabel metal2 20104 27496 20104 27496 0 net6
rlabel metal2 2072 14336 2072 14336 0 net60
rlabel metal2 2744 29008 2744 29008 0 net61
rlabel metal2 2072 21000 2072 21000 0 net62
rlabel metal2 18984 21504 18984 21504 0 net63
rlabel metal3 24136 22344 24136 22344 0 net64
rlabel metal2 24472 19768 24472 19768 0 net65
rlabel metal3 28448 53144 28448 53144 0 net66
rlabel metal2 30520 53704 30520 53704 0 net67
rlabel metal2 34944 53816 34944 53816 0 net68
rlabel metal2 40600 48244 40600 48244 0 net69
rlabel metal2 2072 27048 2072 27048 0 net7
rlabel metal3 39144 52920 39144 52920 0 net70
rlabel metal2 41104 46088 41104 46088 0 net71
rlabel metal2 2072 40824 2072 40824 0 net72
rlabel metal2 45640 36736 45640 36736 0 net73
rlabel metal3 44520 35000 44520 35000 0 net74
rlabel metal3 8792 34888 8792 34888 0 net75
rlabel metal2 13888 37240 13888 37240 0 net76
rlabel metal2 16632 44240 16632 44240 0 net77
rlabel metal2 20664 39424 20664 39424 0 net78
rlabel metal2 25088 53480 25088 53480 0 net79
rlabel metal2 2968 27664 2968 27664 0 net8
rlabel metal2 31976 5152 31976 5152 0 net80
rlabel metal3 29792 5096 29792 5096 0 net81
rlabel metal2 2744 19264 2744 19264 0 net82
rlabel metal2 15344 30072 15344 30072 0 net83
rlabel metal2 17416 41720 17416 41720 0 net84
rlabel metal2 38584 56000 38584 56000 0 net85
rlabel metal2 22904 27216 22904 27216 0 net86
rlabel metal2 31696 50680 31696 50680 0 net87
rlabel metal2 28784 21224 28784 21224 0 net88
rlabel metal2 27048 24696 27048 24696 0 net89
rlabel metal3 1792 48776 1792 48776 0 net9
rlabel metal2 20776 24920 20776 24920 0 net90
rlabel metal2 28448 24024 28448 24024 0 net91
rlabel metal2 39256 24696 39256 24696 0 net92
rlabel metal3 32088 25256 32088 25256 0 net93
rlabel metal2 15176 28336 15176 28336 0 net94
rlabel metal3 46088 23968 46088 23968 0 net95
rlabel metal2 32368 21448 32368 21448 0 net96
rlabel metal2 36288 20552 36288 20552 0 net97
rlabel metal2 39032 17276 39032 17276 0 net98
rlabel metal3 32872 54488 32872 54488 0 net99
rlabel metal2 1736 11032 1736 11032 0 pcpi_insn[0]
rlabel metal2 24920 57778 24920 57778 0 pcpi_insn[12]
rlabel metal2 26376 54712 26376 54712 0 pcpi_insn[13]
rlabel metal2 29008 55272 29008 55272 0 pcpi_insn[14]
rlabel metal2 1848 26320 1848 26320 0 pcpi_insn[1]
rlabel metal2 1960 28448 1960 28448 0 pcpi_insn[25]
rlabel metal2 1736 28672 1736 28672 0 pcpi_insn[26]
rlabel metal3 1638 26264 1638 26264 0 pcpi_insn[27]
rlabel metal2 1680 48776 1680 48776 0 pcpi_insn[28]
rlabel metal2 2408 27720 2408 27720 0 pcpi_insn[29]
rlabel metal2 1736 11816 1736 11816 0 pcpi_insn[2]
rlabel metal2 1904 23016 1904 23016 0 pcpi_insn[30]
rlabel metal3 1848 25872 1848 25872 0 pcpi_insn[31]
rlabel metal3 1638 12152 1638 12152 0 pcpi_insn[3]
rlabel metal2 3248 13944 3248 13944 0 pcpi_insn[4]
rlabel metal2 2408 25144 2408 25144 0 pcpi_insn[5]
rlabel metal2 1736 18928 1736 18928 0 pcpi_insn[6]
rlabel metal3 1358 40376 1358 40376 0 pcpi_rd[0]
rlabel metal3 1358 42392 1358 42392 0 pcpi_rd[10]
rlabel metal2 34328 57610 34328 57610 0 pcpi_rd[11]
rlabel metal3 1358 24920 1358 24920 0 pcpi_rd[12]
rlabel metal3 32928 55384 32928 55384 0 pcpi_rd[13]
rlabel metal2 28952 2058 28952 2058 0 pcpi_rd[14]
rlabel metal2 26880 3640 26880 3640 0 pcpi_rd[15]
rlabel metal3 1358 14840 1358 14840 0 pcpi_rd[16]
rlabel metal2 28280 1414 28280 1414 0 pcpi_rd[17]
rlabel metal2 57960 24528 57960 24528 0 pcpi_rd[18]
rlabel metal3 31360 3640 31360 3640 0 pcpi_rd[19]
rlabel metal3 1358 28952 1358 28952 0 pcpi_rd[1]
rlabel metal2 55384 24360 55384 24360 0 pcpi_rd[20]
rlabel metal3 32928 5208 32928 5208 0 pcpi_rd[21]
rlabel metal3 36344 3640 36344 3640 0 pcpi_rd[22]
rlabel metal2 37016 854 37016 854 0 pcpi_rd[23]
rlabel metal3 33600 54712 33600 54712 0 pcpi_rd[24]
rlabel metal2 57960 36176 57960 36176 0 pcpi_rd[25]
rlabel metal3 36680 55384 36680 55384 0 pcpi_rd[26]
rlabel metal2 24248 58338 24248 58338 0 pcpi_rd[27]
rlabel metal2 57960 32088 57960 32088 0 pcpi_rd[28]
rlabel metal2 57512 26264 57512 26264 0 pcpi_rd[29]
rlabel metal3 1358 30968 1358 30968 0 pcpi_rd[2]
rlabel metal2 57960 28504 57960 28504 0 pcpi_rd[30]
rlabel metal2 57960 27440 57960 27440 0 pcpi_rd[31]
rlabel metal3 1638 29624 1638 29624 0 pcpi_rd[3]
rlabel metal2 25592 57610 25592 57610 0 pcpi_rd[4]
rlabel metal3 1358 39704 1358 39704 0 pcpi_rd[5]
rlabel metal2 31640 57778 31640 57778 0 pcpi_rd[6]
rlabel metal2 27608 57610 27608 57610 0 pcpi_rd[7]
rlabel metal3 1358 37016 1358 37016 0 pcpi_rd[8]
rlabel metal3 1358 33656 1358 33656 0 pcpi_rd[9]
rlabel metal2 57848 32200 57848 32200 0 pcpi_ready
rlabel metal2 1848 37240 1848 37240 0 pcpi_rs1[0]
rlabel metal2 34328 1638 34328 1638 0 pcpi_rs1[10]
rlabel metal2 42224 3528 42224 3528 0 pcpi_rs1[11]
rlabel metal2 39704 1694 39704 1694 0 pcpi_rs1[12]
rlabel metal2 43064 1302 43064 1302 0 pcpi_rs1[13]
rlabel metal2 47096 2058 47096 2058 0 pcpi_rs1[14]
rlabel metal2 49896 3528 49896 3528 0 pcpi_rs1[15]
rlabel metal3 1974 16856 1974 16856 0 pcpi_rs1[16]
rlabel metal2 2632 17472 2632 17472 0 pcpi_rs1[17]
rlabel metal3 1246 12824 1246 12824 0 pcpi_rs1[18]
rlabel metal2 1848 14224 1848 14224 0 pcpi_rs1[19]
rlabel metal2 4760 41104 4760 41104 0 pcpi_rs1[1]
rlabel metal2 2408 13608 2408 13608 0 pcpi_rs1[20]
rlabel metal3 1694 15512 1694 15512 0 pcpi_rs1[21]
rlabel metal2 1736 10360 1736 10360 0 pcpi_rs1[22]
rlabel metal2 1736 8904 1736 8904 0 pcpi_rs1[23]
rlabel metal2 28504 54936 28504 54936 0 pcpi_rs1[24]
rlabel metal2 28952 54880 28952 54880 0 pcpi_rs1[25]
rlabel metal2 30520 55328 30520 55328 0 pcpi_rs1[26]
rlabel metal2 38360 58002 38360 58002 0 pcpi_rs1[27]
rlabel metal2 37016 57722 37016 57722 0 pcpi_rs1[28]
rlabel metal2 37688 56938 37688 56938 0 pcpi_rs1[29]
rlabel metal2 6216 32032 6216 32032 0 pcpi_rs1[2]
rlabel metal2 49784 57778 49784 57778 0 pcpi_rs1[30]
rlabel metal2 51016 55412 51016 55412 0 pcpi_rs1[31]
rlabel metal3 1246 35672 1246 35672 0 pcpi_rs1[3]
rlabel metal2 1904 51240 1904 51240 0 pcpi_rs1[4]
rlabel metal2 2408 49280 2408 49280 0 pcpi_rs1[5]
rlabel metal2 1848 46312 1848 46312 0 pcpi_rs1[6]
rlabel metal3 1246 50456 1246 50456 0 pcpi_rs1[7]
rlabel metal2 41160 4200 41160 4200 0 pcpi_rs1[8]
rlabel metal3 29680 3416 29680 3416 0 pcpi_rs1[9]
rlabel metal3 2058 35000 2058 35000 0 pcpi_rs2[0]
rlabel metal2 44520 3696 44520 3696 0 pcpi_rs2[10]
rlabel metal2 44968 4144 44968 4144 0 pcpi_rs2[11]
rlabel metal3 45528 3304 45528 3304 0 pcpi_rs2[12]
rlabel metal2 48832 3304 48832 3304 0 pcpi_rs2[13]
rlabel metal2 58184 21168 58184 21168 0 pcpi_rs2[14]
rlabel metal2 58184 24920 58184 24920 0 pcpi_rs2[15]
rlabel metal2 1792 21784 1792 21784 0 pcpi_rs2[16]
rlabel metal2 1848 17080 1848 17080 0 pcpi_rs2[17]
rlabel metal2 2520 18368 2520 18368 0 pcpi_rs2[18]
rlabel metal2 3136 13048 3136 13048 0 pcpi_rs2[19]
rlabel metal2 3640 29736 3640 29736 0 pcpi_rs2[1]
rlabel metal2 1736 21056 1736 21056 0 pcpi_rs2[20]
rlabel metal2 3024 17640 3024 17640 0 pcpi_rs2[21]
rlabel metal2 22344 3416 22344 3416 0 pcpi_rs2[22]
rlabel metal2 25144 4200 25144 4200 0 pcpi_rs2[23]
rlabel metal2 27440 55384 27440 55384 0 pcpi_rs2[24]
rlabel metal2 31304 55412 31304 55412 0 pcpi_rs2[25]
rlabel metal3 34664 55384 34664 55384 0 pcpi_rs2[26]
rlabel metal2 36344 57778 36344 57778 0 pcpi_rs2[27]
rlabel metal2 35000 57274 35000 57274 0 pcpi_rs2[28]
rlabel metal2 40992 55272 40992 55272 0 pcpi_rs2[29]
rlabel metal3 2296 41944 2296 41944 0 pcpi_rs2[2]
rlabel metal2 58184 37128 58184 37128 0 pcpi_rs2[30]
rlabel metal2 58184 35336 58184 35336 0 pcpi_rs2[31]
rlabel metal2 6552 35616 6552 35616 0 pcpi_rs2[3]
rlabel metal3 1736 43960 1736 43960 0 pcpi_rs2[4]
rlabel metal2 1736 47992 1736 47992 0 pcpi_rs2[5]
rlabel metal2 5544 39704 5544 39704 0 pcpi_rs2[6]
rlabel metal2 23520 56280 23520 56280 0 pcpi_rs2[7]
rlabel metal2 29288 5264 29288 5264 0 pcpi_rs2[8]
rlabel metal3 33488 3528 33488 3528 0 pcpi_rs2[9]
rlabel metal3 1246 22232 1246 22232 0 pcpi_valid
rlabel metal2 57960 31024 57960 31024 0 pcpi_wr
<< properties >>
string FIXED_BBOX 0 0 60000 60000
<< end >>

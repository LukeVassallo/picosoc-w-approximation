magic
tech gf180mcuD
magscale 1 10
timestamp 1702208760
<< metal1 >>
rect 27570 46958 27582 47010
rect 27634 47007 27646 47010
rect 28242 47007 28254 47010
rect 27634 46961 28254 47007
rect 27634 46958 27646 46961
rect 28242 46958 28254 46961
rect 28306 46958 28318 47010
rect 30258 46622 30270 46674
rect 30322 46671 30334 46674
rect 31042 46671 31054 46674
rect 30322 46625 31054 46671
rect 30322 46622 30334 46625
rect 31042 46622 31054 46625
rect 31106 46671 31118 46674
rect 31490 46671 31502 46674
rect 31106 46625 31502 46671
rect 31106 46622 31118 46625
rect 31490 46622 31502 46625
rect 31554 46622 31566 46674
rect 10098 46510 10110 46562
rect 10162 46559 10174 46562
rect 10770 46559 10782 46562
rect 10162 46513 10782 46559
rect 10162 46510 10174 46513
rect 10770 46510 10782 46513
rect 10834 46510 10846 46562
rect 8754 46398 8766 46450
rect 8818 46447 8830 46450
rect 9090 46447 9102 46450
rect 8818 46401 9102 46447
rect 8818 46398 8830 46401
rect 9090 46398 9102 46401
rect 9154 46447 9166 46450
rect 9426 46447 9438 46450
rect 9154 46401 9438 46447
rect 9154 46398 9166 46401
rect 9426 46398 9438 46401
rect 9490 46398 9502 46450
rect 42354 46398 42366 46450
rect 42418 46447 42430 46450
rect 44930 46447 44942 46450
rect 42418 46401 44942 46447
rect 42418 46398 42430 46401
rect 44930 46398 44942 46401
rect 44994 46398 45006 46450
rect 1344 46282 58576 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 58576 46282
rect 1344 46196 58576 46230
rect 29374 46114 29426 46126
rect 29374 46050 29426 46062
rect 9662 46002 9714 46014
rect 9662 45938 9714 45950
rect 14478 46002 14530 46014
rect 14478 45938 14530 45950
rect 16046 46002 16098 46014
rect 16046 45938 16098 45950
rect 19182 46002 19234 46014
rect 19182 45938 19234 45950
rect 26798 46002 26850 46014
rect 26798 45938 26850 45950
rect 35086 46002 35138 46014
rect 35086 45938 35138 45950
rect 44606 46002 44658 46014
rect 53790 46002 53842 46014
rect 49970 45950 49982 46002
rect 50034 45950 50046 46002
rect 44606 45938 44658 45950
rect 53790 45938 53842 45950
rect 8766 45890 8818 45902
rect 11902 45890 11954 45902
rect 13134 45890 13186 45902
rect 16494 45890 16546 45902
rect 9986 45838 9998 45890
rect 10050 45838 10062 45890
rect 10770 45838 10782 45890
rect 10834 45838 10846 45890
rect 12338 45838 12350 45890
rect 12402 45838 12414 45890
rect 13794 45838 13806 45890
rect 13858 45838 13870 45890
rect 8766 45826 8818 45838
rect 11902 45826 11954 45838
rect 13134 45826 13186 45838
rect 16494 45826 16546 45838
rect 17054 45890 17106 45902
rect 17054 45826 17106 45838
rect 17726 45890 17778 45902
rect 21086 45890 21138 45902
rect 18610 45838 18622 45890
rect 18674 45838 18686 45890
rect 17726 45826 17778 45838
rect 21086 45826 21138 45838
rect 27134 45890 27186 45902
rect 36542 45890 36594 45902
rect 27570 45838 27582 45890
rect 27634 45838 27646 45890
rect 28354 45838 28366 45890
rect 28418 45838 28430 45890
rect 31490 45838 31502 45890
rect 31554 45838 31566 45890
rect 27134 45826 27186 45838
rect 36542 45826 36594 45838
rect 37214 45890 37266 45902
rect 40462 45890 40514 45902
rect 41806 45890 41858 45902
rect 38098 45838 38110 45890
rect 38162 45838 38174 45890
rect 38658 45838 38670 45890
rect 38722 45838 38734 45890
rect 40002 45838 40014 45890
rect 40066 45838 40078 45890
rect 41346 45838 41358 45890
rect 41410 45838 41422 45890
rect 37214 45826 37266 45838
rect 40462 45826 40514 45838
rect 41806 45826 41858 45838
rect 42254 45890 42306 45902
rect 43598 45890 43650 45902
rect 45502 45890 45554 45902
rect 54238 45890 54290 45902
rect 42802 45838 42814 45890
rect 42866 45838 42878 45890
rect 45042 45838 45054 45890
rect 45106 45838 45118 45890
rect 50082 45838 50094 45890
rect 50146 45838 50158 45890
rect 51426 45838 51438 45890
rect 51490 45838 51502 45890
rect 52098 45838 52110 45890
rect 52162 45838 52174 45890
rect 52770 45838 52782 45890
rect 52834 45838 52846 45890
rect 42254 45826 42306 45838
rect 43598 45826 43650 45838
rect 45502 45826 45554 45838
rect 54238 45826 54290 45838
rect 8206 45778 8258 45790
rect 12574 45778 12626 45790
rect 13470 45778 13522 45790
rect 11554 45726 11566 45778
rect 11618 45726 11630 45778
rect 13234 45726 13246 45778
rect 13298 45726 13310 45778
rect 8206 45714 8258 45726
rect 12574 45714 12626 45726
rect 13470 45714 13522 45726
rect 15374 45778 15426 45790
rect 15374 45714 15426 45726
rect 20750 45778 20802 45790
rect 20750 45714 20802 45726
rect 21310 45778 21362 45790
rect 21310 45714 21362 45726
rect 35534 45778 35586 45790
rect 35534 45714 35586 45726
rect 42366 45778 42418 45790
rect 46062 45778 46114 45790
rect 42578 45726 42590 45778
rect 42642 45726 42654 45778
rect 42366 45714 42418 45726
rect 46062 45714 46114 45726
rect 46734 45778 46786 45790
rect 46734 45714 46786 45726
rect 47406 45778 47458 45790
rect 47406 45714 47458 45726
rect 47742 45778 47794 45790
rect 47742 45714 47794 45726
rect 49646 45778 49698 45790
rect 49646 45714 49698 45726
rect 53342 45778 53394 45790
rect 53342 45714 53394 45726
rect 8430 45666 8482 45678
rect 10558 45666 10610 45678
rect 10210 45614 10222 45666
rect 10274 45614 10286 45666
rect 8430 45602 8482 45614
rect 10558 45602 10610 45614
rect 14142 45666 14194 45678
rect 14142 45602 14194 45614
rect 15038 45666 15090 45678
rect 15038 45602 15090 45614
rect 17390 45666 17442 45678
rect 21086 45666 21138 45678
rect 18050 45614 18062 45666
rect 18114 45614 18126 45666
rect 18386 45614 18398 45666
rect 18450 45614 18462 45666
rect 17390 45602 17442 45614
rect 21086 45602 21138 45614
rect 27806 45666 27858 45678
rect 27806 45602 27858 45614
rect 31278 45666 31330 45678
rect 31278 45602 31330 45614
rect 36878 45666 36930 45678
rect 38894 45666 38946 45678
rect 37538 45614 37550 45666
rect 37602 45614 37614 45666
rect 37874 45614 37886 45666
rect 37938 45614 37950 45666
rect 36878 45602 36930 45614
rect 38894 45602 38946 45614
rect 39790 45666 39842 45678
rect 39790 45602 39842 45614
rect 40798 45666 40850 45678
rect 40798 45602 40850 45614
rect 43150 45666 43202 45678
rect 43150 45602 43202 45614
rect 44158 45666 44210 45678
rect 44158 45602 44210 45614
rect 46398 45666 46450 45678
rect 48414 45666 48466 45678
rect 48066 45614 48078 45666
rect 48130 45614 48142 45666
rect 46398 45602 46450 45614
rect 48414 45602 48466 45614
rect 48750 45666 48802 45678
rect 51886 45666 51938 45678
rect 49074 45614 49086 45666
rect 49138 45614 49150 45666
rect 51202 45614 51214 45666
rect 51266 45614 51278 45666
rect 52546 45614 52558 45666
rect 52610 45614 52622 45666
rect 48750 45602 48802 45614
rect 51886 45602 51938 45614
rect 1344 45498 58576 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 50558 45498
rect 50610 45446 50662 45498
rect 50714 45446 50766 45498
rect 50818 45446 58576 45498
rect 1344 45412 58576 45446
rect 9102 45330 9154 45342
rect 9102 45266 9154 45278
rect 10446 45330 10498 45342
rect 10446 45266 10498 45278
rect 14814 45330 14866 45342
rect 14814 45266 14866 45278
rect 21086 45330 21138 45342
rect 21086 45266 21138 45278
rect 21870 45330 21922 45342
rect 21870 45266 21922 45278
rect 30046 45330 30098 45342
rect 30046 45266 30098 45278
rect 31054 45330 31106 45342
rect 31054 45266 31106 45278
rect 52222 45330 52274 45342
rect 52222 45266 52274 45278
rect 14142 45218 14194 45230
rect 9874 45166 9886 45218
rect 9938 45166 9950 45218
rect 11554 45166 11566 45218
rect 11618 45166 11630 45218
rect 12226 45166 12238 45218
rect 12290 45166 12302 45218
rect 13906 45166 13918 45218
rect 13970 45166 13982 45218
rect 14142 45154 14194 45166
rect 16606 45218 16658 45230
rect 22542 45218 22594 45230
rect 40238 45218 40290 45230
rect 17714 45166 17726 45218
rect 17778 45166 17790 45218
rect 30370 45166 30382 45218
rect 30434 45166 30446 45218
rect 16606 45154 16658 45166
rect 22542 45154 22594 45166
rect 40238 45154 40290 45166
rect 42254 45218 42306 45230
rect 43822 45218 43874 45230
rect 53230 45218 53282 45230
rect 43026 45166 43038 45218
rect 43090 45166 43102 45218
rect 44706 45166 44718 45218
rect 44770 45166 44782 45218
rect 50978 45166 50990 45218
rect 51042 45166 51054 45218
rect 42254 45154 42306 45166
rect 43822 45154 43874 45166
rect 53230 45154 53282 45166
rect 15598 45106 15650 45118
rect 20190 45106 20242 45118
rect 9650 45054 9662 45106
rect 9714 45054 9726 45106
rect 10210 45054 10222 45106
rect 10274 45054 10286 45106
rect 11106 45054 11118 45106
rect 11170 45054 11182 45106
rect 12114 45054 12126 45106
rect 12178 45054 12190 45106
rect 12674 45054 12686 45106
rect 12738 45054 12750 45106
rect 13346 45054 13358 45106
rect 13410 45054 13422 45106
rect 14354 45054 14366 45106
rect 14418 45054 14430 45106
rect 15362 45054 15374 45106
rect 15426 45054 15438 45106
rect 16818 45054 16830 45106
rect 16882 45054 16894 45106
rect 18162 45054 18174 45106
rect 18226 45054 18238 45106
rect 18946 45054 18958 45106
rect 19010 45054 19022 45106
rect 15598 45042 15650 45054
rect 20190 45042 20242 45054
rect 21758 45106 21810 45118
rect 21758 45042 21810 45054
rect 21982 45106 22034 45118
rect 21982 45042 22034 45054
rect 22430 45106 22482 45118
rect 22430 45042 22482 45054
rect 22766 45106 22818 45118
rect 40350 45106 40402 45118
rect 44158 45106 44210 45118
rect 51998 45106 52050 45118
rect 29250 45054 29262 45106
rect 29314 45054 29326 45106
rect 36642 45054 36654 45106
rect 36706 45054 36718 45106
rect 38210 45054 38222 45106
rect 38274 45054 38286 45106
rect 39554 45054 39566 45106
rect 39618 45054 39630 45106
rect 41010 45054 41022 45106
rect 41074 45054 41086 45106
rect 42018 45054 42030 45106
rect 42082 45054 42094 45106
rect 42914 45054 42926 45106
rect 42978 45054 42990 45106
rect 45378 45054 45390 45106
rect 45442 45054 45454 45106
rect 46274 45054 46286 45106
rect 46338 45054 46350 45106
rect 47618 45054 47630 45106
rect 47682 45054 47694 45106
rect 49858 45054 49870 45106
rect 49922 45054 49934 45106
rect 22766 45042 22818 45054
rect 40350 45042 40402 45054
rect 44158 45042 44210 45054
rect 51998 45042 52050 45054
rect 13806 44994 13858 45006
rect 11554 44942 11566 44994
rect 11618 44942 11630 44994
rect 13806 44930 13858 44942
rect 15710 44994 15762 45006
rect 15710 44930 15762 44942
rect 19630 44994 19682 45006
rect 19630 44930 19682 44942
rect 19966 44994 20018 45006
rect 19966 44930 20018 44942
rect 20638 44994 20690 45006
rect 20638 44930 20690 44942
rect 21310 44994 21362 45006
rect 21310 44930 21362 44942
rect 21534 44994 21586 45006
rect 21534 44930 21586 44942
rect 27358 44994 27410 45006
rect 27358 44930 27410 44942
rect 34750 44994 34802 45006
rect 52110 44994 52162 45006
rect 37426 44942 37438 44994
rect 37490 44942 37502 44994
rect 39106 44942 39118 44994
rect 39170 44942 39182 44994
rect 41346 44942 41358 44994
rect 41410 44942 41422 44994
rect 43362 44942 43374 44994
rect 43426 44942 43438 44994
rect 45266 44942 45278 44994
rect 45330 44942 45342 44994
rect 49074 44942 49086 44994
rect 49138 44942 49150 44994
rect 51538 44942 51550 44994
rect 51602 44942 51614 44994
rect 34750 44930 34802 44942
rect 52110 44930 52162 44942
rect 52782 44994 52834 45006
rect 52782 44930 52834 44942
rect 11902 44882 11954 44894
rect 11902 44818 11954 44830
rect 16494 44882 16546 44894
rect 16494 44818 16546 44830
rect 20414 44882 20466 44894
rect 20414 44818 20466 44830
rect 40238 44882 40290 44894
rect 40238 44818 40290 44830
rect 1344 44714 58576 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 58576 44714
rect 1344 44628 58576 44662
rect 16270 44546 16322 44558
rect 16270 44482 16322 44494
rect 36318 44546 36370 44558
rect 36318 44482 36370 44494
rect 52894 44546 52946 44558
rect 52894 44482 52946 44494
rect 10558 44434 10610 44446
rect 10558 44370 10610 44382
rect 12126 44434 12178 44446
rect 28702 44434 28754 44446
rect 15586 44382 15598 44434
rect 15650 44382 15662 44434
rect 12126 44370 12178 44382
rect 28702 44370 28754 44382
rect 30046 44434 30098 44446
rect 30046 44370 30098 44382
rect 30382 44434 30434 44446
rect 37214 44434 37266 44446
rect 44942 44434 44994 44446
rect 52670 44434 52722 44446
rect 32498 44382 32510 44434
rect 32562 44382 32574 44434
rect 44370 44382 44382 44434
rect 44434 44382 44446 44434
rect 49970 44382 49982 44434
rect 50034 44382 50046 44434
rect 50866 44382 50878 44434
rect 50930 44382 50942 44434
rect 30382 44370 30434 44382
rect 37214 44370 37266 44382
rect 44942 44370 44994 44382
rect 52670 44370 52722 44382
rect 9662 44322 9714 44334
rect 9662 44258 9714 44270
rect 9886 44322 9938 44334
rect 13806 44322 13858 44334
rect 10098 44270 10110 44322
rect 10162 44270 10174 44322
rect 11442 44270 11454 44322
rect 11506 44270 11518 44322
rect 12450 44270 12462 44322
rect 12514 44270 12526 44322
rect 9886 44258 9938 44270
rect 13806 44258 13858 44270
rect 16382 44322 16434 44334
rect 16382 44258 16434 44270
rect 17054 44322 17106 44334
rect 17054 44258 17106 44270
rect 17502 44322 17554 44334
rect 17502 44258 17554 44270
rect 18958 44322 19010 44334
rect 21310 44322 21362 44334
rect 33518 44322 33570 44334
rect 19730 44270 19742 44322
rect 19794 44270 19806 44322
rect 20402 44270 20414 44322
rect 20466 44270 20478 44322
rect 22082 44270 22094 44322
rect 22146 44270 22158 44322
rect 23202 44270 23214 44322
rect 23266 44270 23278 44322
rect 29362 44270 29374 44322
rect 29426 44270 29438 44322
rect 18958 44258 19010 44270
rect 21310 44258 21362 44270
rect 33518 44258 33570 44270
rect 34078 44322 34130 44334
rect 34078 44258 34130 44270
rect 36206 44322 36258 44334
rect 39678 44322 39730 44334
rect 38882 44270 38894 44322
rect 38946 44270 38958 44322
rect 39106 44270 39118 44322
rect 39170 44270 39182 44322
rect 36206 44258 36258 44270
rect 39678 44258 39730 44270
rect 40350 44322 40402 44334
rect 41458 44270 41470 44322
rect 41522 44270 41534 44322
rect 44258 44270 44270 44322
rect 44322 44270 44334 44322
rect 46274 44270 46286 44322
rect 46338 44270 46350 44322
rect 47282 44270 47294 44322
rect 47346 44270 47358 44322
rect 48850 44270 48862 44322
rect 48914 44270 48926 44322
rect 49074 44270 49086 44322
rect 49138 44270 49150 44322
rect 50194 44270 50206 44322
rect 50258 44270 50270 44322
rect 50642 44270 50654 44322
rect 50706 44270 50718 44322
rect 40350 44258 40402 44270
rect 1710 44210 1762 44222
rect 9774 44210 9826 44222
rect 15262 44210 15314 44222
rect 7970 44158 7982 44210
rect 8034 44158 8046 44210
rect 11778 44158 11790 44210
rect 11842 44158 11854 44210
rect 12114 44158 12126 44210
rect 12178 44158 12190 44210
rect 1710 44146 1762 44158
rect 9774 44146 9826 44158
rect 15262 44146 15314 44158
rect 15486 44210 15538 44222
rect 15486 44146 15538 44158
rect 17614 44210 17666 44222
rect 17614 44146 17666 44158
rect 17838 44210 17890 44222
rect 17838 44146 17890 44158
rect 19294 44210 19346 44222
rect 32174 44210 32226 44222
rect 20738 44158 20750 44210
rect 20802 44158 20814 44210
rect 22754 44158 22766 44210
rect 22818 44158 22830 44210
rect 19294 44146 19346 44158
rect 32174 44146 32226 44158
rect 33630 44210 33682 44222
rect 33630 44146 33682 44158
rect 36318 44210 36370 44222
rect 36318 44146 36370 44158
rect 37550 44210 37602 44222
rect 37550 44146 37602 44158
rect 37662 44210 37714 44222
rect 37662 44146 37714 44158
rect 39342 44210 39394 44222
rect 40674 44158 40686 44210
rect 40738 44158 40750 44210
rect 41906 44158 41918 44210
rect 41970 44158 41982 44210
rect 42802 44158 42814 44210
rect 42866 44158 42878 44210
rect 45826 44158 45838 44210
rect 45890 44158 45902 44210
rect 48066 44158 48078 44210
rect 48130 44158 48142 44210
rect 39342 44146 39394 44158
rect 2046 44098 2098 44110
rect 2046 44034 2098 44046
rect 2494 44098 2546 44110
rect 2494 44034 2546 44046
rect 7646 44098 7698 44110
rect 7646 44034 7698 44046
rect 8766 44098 8818 44110
rect 16270 44098 16322 44110
rect 29150 44098 29202 44110
rect 9090 44046 9102 44098
rect 9154 44046 9166 44098
rect 13458 44046 13470 44098
rect 13522 44046 13534 44098
rect 16706 44046 16718 44098
rect 16770 44046 16782 44098
rect 19730 44046 19742 44098
rect 19794 44046 19806 44098
rect 21634 44046 21646 44098
rect 21698 44046 21710 44098
rect 22194 44046 22206 44098
rect 22258 44046 22270 44098
rect 8766 44034 8818 44046
rect 16270 44034 16322 44046
rect 29150 44034 29202 44046
rect 37326 44098 37378 44110
rect 37326 44034 37378 44046
rect 40014 44098 40066 44110
rect 40014 44034 40066 44046
rect 51886 44098 51938 44110
rect 53218 44046 53230 44098
rect 53282 44046 53294 44098
rect 51886 44034 51938 44046
rect 1344 43930 58576 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 50558 43930
rect 50610 43878 50662 43930
rect 50714 43878 50766 43930
rect 50818 43878 58576 43930
rect 1344 43844 58576 43878
rect 7086 43762 7138 43774
rect 7086 43698 7138 43710
rect 9886 43762 9938 43774
rect 9886 43698 9938 43710
rect 13246 43762 13298 43774
rect 13246 43698 13298 43710
rect 39342 43762 39394 43774
rect 46274 43710 46286 43762
rect 46338 43710 46350 43762
rect 39342 43698 39394 43710
rect 34414 43650 34466 43662
rect 38110 43650 38162 43662
rect 39566 43650 39618 43662
rect 10210 43598 10222 43650
rect 10274 43598 10286 43650
rect 10658 43598 10670 43650
rect 10722 43598 10734 43650
rect 14354 43598 14366 43650
rect 14418 43598 14430 43650
rect 37762 43598 37774 43650
rect 37826 43598 37838 43650
rect 38434 43598 38446 43650
rect 38498 43598 38510 43650
rect 34414 43586 34466 43598
rect 38110 43586 38162 43598
rect 39566 43586 39618 43598
rect 40126 43650 40178 43662
rect 42030 43650 42082 43662
rect 47294 43650 47346 43662
rect 41010 43598 41022 43650
rect 41074 43598 41086 43650
rect 42914 43598 42926 43650
rect 42978 43598 42990 43650
rect 44146 43598 44158 43650
rect 44210 43598 44222 43650
rect 46050 43598 46062 43650
rect 46114 43598 46126 43650
rect 40126 43586 40178 43598
rect 42030 43586 42082 43598
rect 47294 43586 47346 43598
rect 47630 43650 47682 43662
rect 47630 43586 47682 43598
rect 48862 43650 48914 43662
rect 48862 43586 48914 43598
rect 49086 43650 49138 43662
rect 49086 43586 49138 43598
rect 7198 43538 7250 43550
rect 12798 43538 12850 43550
rect 7858 43486 7870 43538
rect 7922 43486 7934 43538
rect 10546 43486 10558 43538
rect 10610 43486 10622 43538
rect 11330 43486 11342 43538
rect 11394 43486 11406 43538
rect 11778 43486 11790 43538
rect 11842 43486 11854 43538
rect 7198 43474 7250 43486
rect 12798 43474 12850 43486
rect 13470 43538 13522 43550
rect 20526 43538 20578 43550
rect 15586 43486 15598 43538
rect 15650 43486 15662 43538
rect 17826 43486 17838 43538
rect 17890 43486 17902 43538
rect 13470 43474 13522 43486
rect 20526 43474 20578 43486
rect 20750 43538 20802 43550
rect 38782 43538 38834 43550
rect 22194 43486 22206 43538
rect 22258 43486 22270 43538
rect 23426 43486 23438 43538
rect 23490 43486 23502 43538
rect 35858 43486 35870 43538
rect 35922 43486 35934 43538
rect 37202 43486 37214 43538
rect 37266 43486 37278 43538
rect 20750 43474 20802 43486
rect 38782 43474 38834 43486
rect 39678 43538 39730 43550
rect 39678 43474 39730 43486
rect 40014 43538 40066 43550
rect 40014 43474 40066 43486
rect 41358 43538 41410 43550
rect 48750 43538 48802 43550
rect 41794 43486 41806 43538
rect 41858 43486 41870 43538
rect 42578 43486 42590 43538
rect 42642 43486 42654 43538
rect 45602 43486 45614 43538
rect 45666 43486 45678 43538
rect 46498 43486 46510 43538
rect 46562 43486 46574 43538
rect 46946 43486 46958 43538
rect 47010 43486 47022 43538
rect 47954 43486 47966 43538
rect 48018 43486 48030 43538
rect 41358 43474 41410 43486
rect 48750 43474 48802 43486
rect 49310 43538 49362 43550
rect 49310 43474 49362 43486
rect 49534 43538 49586 43550
rect 49534 43474 49586 43486
rect 49758 43538 49810 43550
rect 53342 43538 53394 43550
rect 51202 43486 51214 43538
rect 51266 43486 51278 43538
rect 51538 43486 51550 43538
rect 51602 43486 51614 43538
rect 52994 43486 53006 43538
rect 53058 43486 53070 43538
rect 49758 43474 49810 43486
rect 53342 43474 53394 43486
rect 53566 43538 53618 43550
rect 53566 43474 53618 43486
rect 2158 43426 2210 43438
rect 8542 43426 8594 43438
rect 8194 43374 8206 43426
rect 8258 43374 8270 43426
rect 2158 43362 2210 43374
rect 8542 43362 8594 43374
rect 13358 43426 13410 43438
rect 16270 43426 16322 43438
rect 22654 43426 22706 43438
rect 47182 43426 47234 43438
rect 14130 43374 14142 43426
rect 14194 43374 14206 43426
rect 17490 43374 17502 43426
rect 17554 43374 17566 43426
rect 21858 43374 21870 43426
rect 21922 43374 21934 43426
rect 23650 43374 23662 43426
rect 23714 43374 23726 43426
rect 34290 43374 34302 43426
rect 34354 43374 34366 43426
rect 35074 43374 35086 43426
rect 35138 43374 35150 43426
rect 37090 43374 37102 43426
rect 37154 43374 37166 43426
rect 45378 43374 45390 43426
rect 45442 43374 45454 43426
rect 13358 43362 13410 43374
rect 16270 43362 16322 43374
rect 22654 43362 22706 43374
rect 47182 43362 47234 43374
rect 47742 43426 47794 43438
rect 51650 43374 51662 43426
rect 51714 43374 51726 43426
rect 47742 43362 47794 43374
rect 7086 43314 7138 43326
rect 7086 43250 7138 43262
rect 11342 43314 11394 43326
rect 11342 43250 11394 43262
rect 20974 43314 21026 43326
rect 20974 43250 21026 43262
rect 21422 43314 21474 43326
rect 34638 43314 34690 43326
rect 23986 43262 23998 43314
rect 24050 43262 24062 43314
rect 21422 43250 21474 43262
rect 34638 43250 34690 43262
rect 40126 43314 40178 43326
rect 40126 43250 40178 43262
rect 50206 43314 50258 43326
rect 53890 43262 53902 43314
rect 53954 43262 53966 43314
rect 50206 43250 50258 43262
rect 1344 43146 58576 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 58576 43146
rect 1344 43060 58576 43094
rect 8206 42978 8258 42990
rect 8206 42914 8258 42926
rect 15038 42978 15090 42990
rect 15038 42914 15090 42926
rect 15262 42978 15314 42990
rect 15262 42914 15314 42926
rect 34414 42978 34466 42990
rect 37102 42978 37154 42990
rect 34738 42926 34750 42978
rect 34802 42926 34814 42978
rect 34414 42914 34466 42926
rect 37102 42914 37154 42926
rect 41134 42978 41186 42990
rect 41134 42914 41186 42926
rect 45390 42978 45442 42990
rect 45390 42914 45442 42926
rect 51326 42978 51378 42990
rect 51326 42914 51378 42926
rect 7982 42866 8034 42878
rect 14814 42866 14866 42878
rect 40686 42866 40738 42878
rect 11442 42814 11454 42866
rect 11506 42814 11518 42866
rect 33506 42814 33518 42866
rect 33570 42814 33582 42866
rect 47058 42814 47070 42866
rect 47122 42814 47134 42866
rect 49186 42814 49198 42866
rect 49250 42814 49262 42866
rect 50082 42814 50094 42866
rect 50146 42814 50158 42866
rect 52882 42814 52894 42866
rect 52946 42814 52958 42866
rect 7982 42802 8034 42814
rect 14814 42802 14866 42814
rect 40686 42802 40738 42814
rect 7646 42754 7698 42766
rect 1810 42702 1822 42754
rect 1874 42702 1886 42754
rect 7646 42690 7698 42702
rect 8878 42754 8930 42766
rect 10558 42754 10610 42766
rect 10098 42702 10110 42754
rect 10162 42702 10174 42754
rect 8878 42690 8930 42702
rect 10558 42690 10610 42702
rect 11118 42754 11170 42766
rect 13918 42754 13970 42766
rect 12114 42702 12126 42754
rect 12178 42702 12190 42754
rect 11118 42690 11170 42702
rect 13918 42690 13970 42702
rect 15710 42754 15762 42766
rect 15710 42690 15762 42702
rect 16158 42754 16210 42766
rect 19518 42754 19570 42766
rect 19170 42702 19182 42754
rect 19234 42702 19246 42754
rect 16158 42690 16210 42702
rect 19518 42690 19570 42702
rect 23326 42754 23378 42766
rect 23326 42690 23378 42702
rect 23662 42754 23714 42766
rect 34190 42754 34242 42766
rect 31938 42702 31950 42754
rect 32002 42702 32014 42754
rect 33618 42702 33630 42754
rect 33682 42702 33694 42754
rect 23662 42690 23714 42702
rect 34190 42690 34242 42702
rect 34974 42754 35026 42766
rect 34974 42690 35026 42702
rect 37214 42754 37266 42766
rect 37214 42690 37266 42702
rect 37550 42754 37602 42766
rect 37550 42690 37602 42702
rect 39006 42754 39058 42766
rect 39006 42690 39058 42702
rect 41022 42754 41074 42766
rect 41022 42690 41074 42702
rect 41806 42754 41858 42766
rect 41806 42690 41858 42702
rect 42142 42754 42194 42766
rect 42142 42690 42194 42702
rect 43038 42754 43090 42766
rect 43038 42690 43090 42702
rect 44046 42754 44098 42766
rect 46174 42754 46226 42766
rect 45042 42702 45054 42754
rect 45106 42702 45118 42754
rect 47842 42702 47854 42754
rect 47906 42702 47918 42754
rect 48738 42702 48750 42754
rect 48802 42702 48814 42754
rect 49522 42702 49534 42754
rect 49586 42702 49598 42754
rect 54338 42702 54350 42754
rect 54402 42702 54414 42754
rect 44046 42690 44098 42702
rect 46174 42690 46226 42702
rect 2382 42642 2434 42654
rect 2382 42578 2434 42590
rect 7310 42642 7362 42654
rect 7310 42578 7362 42590
rect 10894 42642 10946 42654
rect 10894 42578 10946 42590
rect 13582 42642 13634 42654
rect 13582 42578 13634 42590
rect 19630 42642 19682 42654
rect 19630 42578 19682 42590
rect 22990 42642 23042 42654
rect 22990 42578 23042 42590
rect 23438 42642 23490 42654
rect 23438 42578 23490 42590
rect 30046 42642 30098 42654
rect 30046 42578 30098 42590
rect 30158 42642 30210 42654
rect 35310 42642 35362 42654
rect 31714 42590 31726 42642
rect 31778 42590 31790 42642
rect 30158 42578 30210 42590
rect 35310 42578 35362 42590
rect 39342 42642 39394 42654
rect 39342 42578 39394 42590
rect 41918 42642 41970 42654
rect 41918 42578 41970 42590
rect 42702 42642 42754 42654
rect 42702 42578 42754 42590
rect 51550 42642 51602 42654
rect 53442 42590 53454 42642
rect 53506 42590 53518 42642
rect 55682 42590 55694 42642
rect 55746 42590 55758 42642
rect 51550 42578 51602 42590
rect 2046 42530 2098 42542
rect 2046 42466 2098 42478
rect 2718 42530 2770 42542
rect 2718 42466 2770 42478
rect 3166 42530 3218 42542
rect 3166 42466 3218 42478
rect 7534 42530 7586 42542
rect 11342 42530 11394 42542
rect 8530 42478 8542 42530
rect 8594 42478 8606 42530
rect 9202 42478 9214 42530
rect 9266 42478 9278 42530
rect 7534 42466 7586 42478
rect 11342 42466 11394 42478
rect 11454 42530 11506 42542
rect 13694 42530 13746 42542
rect 11890 42478 11902 42530
rect 11954 42478 11966 42530
rect 11454 42466 11506 42478
rect 13694 42466 13746 42478
rect 16270 42530 16322 42542
rect 16270 42466 16322 42478
rect 16382 42530 16434 42542
rect 16382 42466 16434 42478
rect 16494 42530 16546 42542
rect 16494 42466 16546 42478
rect 16606 42530 16658 42542
rect 16606 42466 16658 42478
rect 22654 42530 22706 42542
rect 22654 42466 22706 42478
rect 22878 42530 22930 42542
rect 22878 42466 22930 42478
rect 30382 42530 30434 42542
rect 30382 42466 30434 42478
rect 30718 42530 30770 42542
rect 30718 42466 30770 42478
rect 35198 42530 35250 42542
rect 35198 42466 35250 42478
rect 37102 42530 37154 42542
rect 37102 42466 37154 42478
rect 37662 42530 37714 42542
rect 37662 42466 37714 42478
rect 37886 42530 37938 42542
rect 37886 42466 37938 42478
rect 39230 42530 39282 42542
rect 40238 42530 40290 42542
rect 39890 42478 39902 42530
rect 39954 42478 39966 42530
rect 39230 42466 39282 42478
rect 40238 42466 40290 42478
rect 41134 42530 41186 42542
rect 43374 42530 43426 42542
rect 42354 42478 42366 42530
rect 42418 42478 42430 42530
rect 41134 42466 41186 42478
rect 43374 42466 43426 42478
rect 43710 42530 43762 42542
rect 43710 42466 43762 42478
rect 45278 42530 45330 42542
rect 45278 42466 45330 42478
rect 45838 42530 45890 42542
rect 45838 42466 45890 42478
rect 51438 42530 51490 42542
rect 51438 42466 51490 42478
rect 1344 42362 58576 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 50558 42362
rect 50610 42310 50662 42362
rect 50714 42310 50766 42362
rect 50818 42310 58576 42362
rect 1344 42276 58576 42310
rect 4398 42194 4450 42206
rect 4398 42130 4450 42142
rect 9774 42194 9826 42206
rect 9774 42130 9826 42142
rect 10558 42194 10610 42206
rect 14590 42194 14642 42206
rect 14018 42142 14030 42194
rect 14082 42142 14094 42194
rect 10558 42130 10610 42142
rect 14590 42130 14642 42142
rect 30046 42194 30098 42206
rect 30046 42130 30098 42142
rect 30494 42194 30546 42206
rect 30494 42130 30546 42142
rect 44606 42194 44658 42206
rect 44606 42130 44658 42142
rect 44830 42194 44882 42206
rect 50754 42142 50766 42194
rect 50818 42142 50830 42194
rect 44830 42130 44882 42142
rect 2046 42082 2098 42094
rect 2046 42018 2098 42030
rect 2718 42082 2770 42094
rect 2718 42018 2770 42030
rect 7646 42082 7698 42094
rect 14478 42082 14530 42094
rect 41358 42082 41410 42094
rect 11442 42030 11454 42082
rect 11506 42030 11518 42082
rect 12674 42030 12686 42082
rect 12738 42030 12750 42082
rect 13458 42030 13470 42082
rect 13522 42030 13534 42082
rect 15362 42030 15374 42082
rect 15426 42030 15438 42082
rect 19058 42030 19070 42082
rect 19122 42030 19134 42082
rect 29698 42030 29710 42082
rect 29762 42030 29774 42082
rect 37538 42030 37550 42082
rect 37602 42030 37614 42082
rect 39442 42030 39454 42082
rect 39506 42030 39518 42082
rect 7646 42018 7698 42030
rect 14478 42018 14530 42030
rect 41358 42018 41410 42030
rect 41470 42082 41522 42094
rect 41470 42018 41522 42030
rect 42254 42082 42306 42094
rect 47966 42082 48018 42094
rect 43362 42030 43374 42082
rect 43426 42030 43438 42082
rect 44146 42030 44158 42082
rect 44210 42030 44222 42082
rect 47058 42030 47070 42082
rect 47122 42030 47134 42082
rect 42254 42018 42306 42030
rect 47966 42018 48018 42030
rect 48078 42082 48130 42094
rect 48078 42018 48130 42030
rect 49198 42082 49250 42094
rect 49746 42030 49758 42082
rect 49810 42030 49822 42082
rect 49198 42018 49250 42030
rect 1710 41970 1762 41982
rect 1710 41906 1762 41918
rect 2382 41970 2434 41982
rect 2382 41906 2434 41918
rect 3614 41970 3666 41982
rect 3614 41906 3666 41918
rect 4510 41970 4562 41982
rect 9998 41970 10050 41982
rect 14814 41970 14866 41982
rect 20638 41970 20690 41982
rect 23326 41970 23378 41982
rect 30270 41970 30322 41982
rect 7410 41918 7422 41970
rect 7474 41918 7486 41970
rect 9538 41918 9550 41970
rect 9602 41918 9614 41970
rect 10210 41918 10222 41970
rect 10274 41918 10286 41970
rect 11666 41918 11678 41970
rect 11730 41918 11742 41970
rect 12450 41918 12462 41970
rect 12514 41918 12526 41970
rect 13346 41918 13358 41970
rect 13410 41918 13422 41970
rect 14018 41918 14030 41970
rect 14082 41918 14094 41970
rect 15586 41918 15598 41970
rect 15650 41918 15662 41970
rect 16146 41918 16158 41970
rect 16210 41918 16222 41970
rect 16706 41918 16718 41970
rect 16770 41918 16782 41970
rect 19954 41918 19966 41970
rect 20018 41918 20030 41970
rect 22194 41918 22206 41970
rect 22258 41918 22270 41970
rect 22642 41918 22654 41970
rect 22706 41918 22718 41970
rect 23650 41918 23662 41970
rect 23714 41918 23726 41970
rect 4510 41906 4562 41918
rect 9998 41906 10050 41918
rect 14814 41906 14866 41918
rect 20638 41906 20690 41918
rect 23326 41906 23378 41918
rect 30270 41906 30322 41918
rect 30606 41970 30658 41982
rect 30606 41906 30658 41918
rect 33182 41970 33234 41982
rect 40350 41970 40402 41982
rect 33394 41918 33406 41970
rect 33458 41918 33470 41970
rect 37426 41918 37438 41970
rect 37490 41918 37502 41970
rect 37650 41918 37662 41970
rect 37714 41918 37726 41970
rect 38546 41918 38558 41970
rect 38610 41918 38622 41970
rect 39666 41918 39678 41970
rect 39730 41918 39742 41970
rect 33182 41906 33234 41918
rect 40350 41906 40402 41918
rect 41694 41970 41746 41982
rect 42702 41970 42754 41982
rect 42018 41918 42030 41970
rect 42082 41918 42094 41970
rect 41694 41906 41746 41918
rect 42702 41906 42754 41918
rect 43150 41970 43202 41982
rect 43150 41906 43202 41918
rect 43822 41970 43874 41982
rect 43822 41906 43874 41918
rect 44494 41970 44546 41982
rect 48302 41970 48354 41982
rect 45602 41918 45614 41970
rect 45666 41918 45678 41970
rect 45826 41918 45838 41970
rect 45890 41918 45902 41970
rect 46610 41918 46622 41970
rect 46674 41918 46686 41970
rect 44494 41906 44546 41918
rect 48302 41906 48354 41918
rect 48862 41970 48914 41982
rect 52446 41970 52498 41982
rect 53342 41970 53394 41982
rect 54686 41970 54738 41982
rect 49970 41918 49982 41970
rect 50034 41918 50046 41970
rect 50642 41918 50654 41970
rect 50706 41918 50718 41970
rect 52994 41918 53006 41970
rect 53058 41918 53070 41970
rect 53554 41918 53566 41970
rect 53618 41918 53630 41970
rect 53778 41918 53790 41970
rect 53842 41918 53854 41970
rect 55122 41918 55134 41970
rect 55186 41918 55198 41970
rect 48862 41906 48914 41918
rect 52446 41906 52498 41918
rect 53342 41906 53394 41918
rect 54686 41906 54738 41918
rect 3166 41858 3218 41870
rect 3166 41794 3218 41806
rect 9886 41858 9938 41870
rect 9886 41794 9938 41806
rect 11118 41858 11170 41870
rect 11118 41794 11170 41806
rect 18622 41858 18674 41870
rect 18622 41794 18674 41806
rect 21982 41858 22034 41870
rect 21982 41794 22034 41806
rect 23438 41858 23490 41870
rect 23438 41794 23490 41806
rect 31054 41858 31106 41870
rect 31054 41794 31106 41806
rect 34078 41858 34130 41870
rect 34078 41794 34130 41806
rect 43486 41858 43538 41870
rect 43486 41794 43538 41806
rect 45054 41858 45106 41870
rect 46498 41806 46510 41858
rect 46562 41806 46574 41858
rect 45054 41794 45106 41806
rect 4398 41746 4450 41758
rect 4398 41682 4450 41694
rect 16942 41746 16994 41758
rect 16942 41682 16994 41694
rect 42478 41746 42530 41758
rect 42478 41682 42530 41694
rect 45278 41746 45330 41758
rect 45278 41682 45330 41694
rect 52670 41746 52722 41758
rect 54002 41694 54014 41746
rect 54066 41694 54078 41746
rect 52670 41682 52722 41694
rect 1344 41578 58576 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 58576 41578
rect 1344 41492 58576 41526
rect 10334 41410 10386 41422
rect 38558 41410 38610 41422
rect 45726 41410 45778 41422
rect 32946 41358 32958 41410
rect 33010 41358 33022 41410
rect 44146 41358 44158 41410
rect 44210 41358 44222 41410
rect 10334 41346 10386 41358
rect 38558 41346 38610 41358
rect 45726 41346 45778 41358
rect 45950 41410 46002 41422
rect 45950 41346 46002 41358
rect 50318 41410 50370 41422
rect 50318 41346 50370 41358
rect 51550 41410 51602 41422
rect 51550 41346 51602 41358
rect 53006 41410 53058 41422
rect 53006 41346 53058 41358
rect 10670 41298 10722 41310
rect 37662 41298 37714 41310
rect 44942 41298 44994 41310
rect 13570 41246 13582 41298
rect 13634 41246 13646 41298
rect 18050 41246 18062 41298
rect 18114 41246 18126 41298
rect 23202 41246 23214 41298
rect 23266 41246 23278 41298
rect 42578 41246 42590 41298
rect 42642 41246 42654 41298
rect 43138 41246 43150 41298
rect 43202 41246 43214 41298
rect 10670 41234 10722 41246
rect 37662 41234 37714 41246
rect 44942 41234 44994 41246
rect 45502 41298 45554 41310
rect 48078 41298 48130 41310
rect 47506 41246 47518 41298
rect 47570 41246 47582 41298
rect 45502 41234 45554 41246
rect 48078 41234 48130 41246
rect 51326 41298 51378 41310
rect 54226 41246 54238 41298
rect 54290 41246 54302 41298
rect 51326 41234 51378 41246
rect 2606 41186 2658 41198
rect 5966 41186 6018 41198
rect 6974 41186 7026 41198
rect 2258 41134 2270 41186
rect 2322 41134 2334 41186
rect 3378 41134 3390 41186
rect 3442 41134 3454 41186
rect 4834 41134 4846 41186
rect 4898 41134 4910 41186
rect 6402 41134 6414 41186
rect 6466 41134 6478 41186
rect 2606 41122 2658 41134
rect 5966 41122 6018 41134
rect 6974 41122 7026 41134
rect 7310 41186 7362 41198
rect 7310 41122 7362 41134
rect 8318 41186 8370 41198
rect 8318 41122 8370 41134
rect 8878 41186 8930 41198
rect 8878 41122 8930 41134
rect 8990 41186 9042 41198
rect 12910 41186 12962 41198
rect 19518 41186 19570 41198
rect 9426 41134 9438 41186
rect 9490 41134 9502 41186
rect 15026 41134 15038 41186
rect 15090 41134 15102 41186
rect 17378 41134 17390 41186
rect 17442 41134 17454 41186
rect 18498 41134 18510 41186
rect 18562 41134 18574 41186
rect 8990 41122 9042 41134
rect 12910 41122 12962 41134
rect 19518 41122 19570 41134
rect 19630 41186 19682 41198
rect 19630 41122 19682 41134
rect 19966 41186 20018 41198
rect 19966 41122 20018 41134
rect 21422 41186 21474 41198
rect 32510 41186 32562 41198
rect 37774 41186 37826 41198
rect 21634 41134 21646 41186
rect 21698 41134 21710 41186
rect 23090 41134 23102 41186
rect 23154 41134 23166 41186
rect 30034 41134 30046 41186
rect 30098 41134 30110 41186
rect 32162 41134 32174 41186
rect 32226 41134 32238 41186
rect 36194 41134 36206 41186
rect 36258 41134 36270 41186
rect 37314 41134 37326 41186
rect 37378 41134 37390 41186
rect 21422 41122 21474 41134
rect 32510 41122 32562 41134
rect 37774 41122 37826 41134
rect 38334 41186 38386 41198
rect 40462 41186 40514 41198
rect 38994 41134 39006 41186
rect 39058 41134 39070 41186
rect 39778 41134 39790 41186
rect 39842 41134 39854 41186
rect 38334 41122 38386 41134
rect 40462 41122 40514 41134
rect 40798 41186 40850 41198
rect 40798 41122 40850 41134
rect 42142 41186 42194 41198
rect 42142 41122 42194 41134
rect 42254 41186 42306 41198
rect 42254 41122 42306 41134
rect 42478 41186 42530 41198
rect 48750 41186 48802 41198
rect 43586 41134 43598 41186
rect 43650 41134 43662 41186
rect 43922 41134 43934 41186
rect 43986 41134 43998 41186
rect 47058 41134 47070 41186
rect 47122 41134 47134 41186
rect 42478 41122 42530 41134
rect 48750 41122 48802 41134
rect 49310 41186 49362 41198
rect 49310 41122 49362 41134
rect 49646 41186 49698 41198
rect 49646 41122 49698 41134
rect 50094 41186 50146 41198
rect 50094 41122 50146 41134
rect 51774 41186 51826 41198
rect 52658 41134 52670 41186
rect 52722 41134 52734 41186
rect 55682 41134 55694 41186
rect 55746 41134 55758 41186
rect 51774 41122 51826 41134
rect 4062 41074 4114 41086
rect 4062 41010 4114 41022
rect 5070 41074 5122 41086
rect 5070 41010 5122 41022
rect 7198 41074 7250 41086
rect 9774 41074 9826 41086
rect 9202 41022 9214 41074
rect 9266 41022 9278 41074
rect 7198 41010 7250 41022
rect 9774 41010 9826 41022
rect 10110 41074 10162 41086
rect 10110 41010 10162 41022
rect 12574 41074 12626 41086
rect 19182 41074 19234 41086
rect 13794 41022 13806 41074
rect 13858 41022 13870 41074
rect 16370 41022 16382 41074
rect 16434 41022 16446 41074
rect 18386 41022 18398 41074
rect 18450 41022 18462 41074
rect 12574 41010 12626 41022
rect 19182 41010 19234 41022
rect 19294 41074 19346 41086
rect 19294 41010 19346 41022
rect 22318 41074 22370 41086
rect 22318 41010 22370 41022
rect 23998 41074 24050 41086
rect 32398 41074 32450 41086
rect 29810 41022 29822 41074
rect 29874 41022 29886 41074
rect 31154 41022 31166 41074
rect 31218 41022 31230 41074
rect 23998 41010 24050 41022
rect 32398 41010 32450 41022
rect 37550 41074 37602 41086
rect 41694 41074 41746 41086
rect 38546 41022 38558 41074
rect 38610 41022 38622 41074
rect 37550 41010 37602 41022
rect 41694 41010 41746 41022
rect 46622 41074 46674 41086
rect 50654 41074 50706 41086
rect 49410 41022 49422 41074
rect 49474 41022 49486 41074
rect 54450 41022 54462 41074
rect 54514 41022 54526 41074
rect 46622 41010 46674 41022
rect 50654 41010 50706 41022
rect 12798 40962 12850 40974
rect 17054 40962 17106 40974
rect 5618 40910 5630 40962
rect 5682 40910 5694 40962
rect 6626 40910 6638 40962
rect 6690 40910 6702 40962
rect 7970 40910 7982 40962
rect 8034 40910 8046 40962
rect 16706 40910 16718 40962
rect 16770 40910 16782 40962
rect 12798 40898 12850 40910
rect 17054 40898 17106 40910
rect 19854 40962 19906 40974
rect 33406 40962 33458 40974
rect 37886 40962 37938 40974
rect 41134 40962 41186 40974
rect 31266 40910 31278 40962
rect 31330 40910 31342 40962
rect 36418 40910 36430 40962
rect 36482 40910 36494 40962
rect 40114 40910 40126 40962
rect 40178 40910 40190 40962
rect 19854 40898 19906 40910
rect 33406 40898 33458 40910
rect 37886 40898 37938 40910
rect 41134 40898 41186 40910
rect 41358 40962 41410 40974
rect 41358 40898 41410 40910
rect 41582 40962 41634 40974
rect 41582 40898 41634 40910
rect 42590 40962 42642 40974
rect 42590 40898 42642 40910
rect 46398 40962 46450 40974
rect 46398 40898 46450 40910
rect 48862 40962 48914 40974
rect 48862 40898 48914 40910
rect 49086 40962 49138 40974
rect 49086 40898 49138 40910
rect 52222 40962 52274 40974
rect 52222 40898 52274 40910
rect 52894 40962 52946 40974
rect 56018 40910 56030 40962
rect 56082 40910 56094 40962
rect 52894 40898 52946 40910
rect 1344 40794 58576 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 50558 40794
rect 50610 40742 50662 40794
rect 50714 40742 50766 40794
rect 50818 40742 58576 40794
rect 1344 40708 58576 40742
rect 4510 40626 4562 40638
rect 4510 40562 4562 40574
rect 4958 40626 5010 40638
rect 4958 40562 5010 40574
rect 5294 40626 5346 40638
rect 5294 40562 5346 40574
rect 5854 40626 5906 40638
rect 5854 40562 5906 40574
rect 10670 40626 10722 40638
rect 10670 40562 10722 40574
rect 18846 40626 18898 40638
rect 28478 40626 28530 40638
rect 22754 40574 22766 40626
rect 22818 40574 22830 40626
rect 18846 40562 18898 40574
rect 28478 40562 28530 40574
rect 36318 40626 36370 40638
rect 36318 40562 36370 40574
rect 37326 40626 37378 40638
rect 37326 40562 37378 40574
rect 37998 40626 38050 40638
rect 37998 40562 38050 40574
rect 43710 40626 43762 40638
rect 43710 40562 43762 40574
rect 44158 40626 44210 40638
rect 44158 40562 44210 40574
rect 44718 40626 44770 40638
rect 44718 40562 44770 40574
rect 45390 40626 45442 40638
rect 45390 40562 45442 40574
rect 45950 40626 46002 40638
rect 45950 40562 46002 40574
rect 3502 40514 3554 40526
rect 3502 40450 3554 40462
rect 5518 40514 5570 40526
rect 7870 40514 7922 40526
rect 6178 40462 6190 40514
rect 6242 40462 6254 40514
rect 7074 40462 7086 40514
rect 7138 40462 7150 40514
rect 5518 40450 5570 40462
rect 7870 40450 7922 40462
rect 7982 40514 8034 40526
rect 13134 40514 13186 40526
rect 12226 40462 12238 40514
rect 12290 40462 12302 40514
rect 7982 40450 8034 40462
rect 13134 40450 13186 40462
rect 13246 40514 13298 40526
rect 13246 40450 13298 40462
rect 13358 40514 13410 40526
rect 19518 40514 19570 40526
rect 18386 40462 18398 40514
rect 18450 40462 18462 40514
rect 13358 40450 13410 40462
rect 19518 40450 19570 40462
rect 19630 40514 19682 40526
rect 19630 40450 19682 40462
rect 19854 40514 19906 40526
rect 23550 40514 23602 40526
rect 21522 40462 21534 40514
rect 21586 40462 21598 40514
rect 19854 40450 19906 40462
rect 23550 40450 23602 40462
rect 23662 40514 23714 40526
rect 23662 40450 23714 40462
rect 28702 40514 28754 40526
rect 28702 40450 28754 40462
rect 28814 40514 28866 40526
rect 28814 40450 28866 40462
rect 31838 40514 31890 40526
rect 31838 40450 31890 40462
rect 35086 40514 35138 40526
rect 35086 40450 35138 40462
rect 36542 40514 36594 40526
rect 36542 40450 36594 40462
rect 36654 40514 36706 40526
rect 43038 40514 43090 40526
rect 36978 40462 36990 40514
rect 37042 40462 37054 40514
rect 37650 40462 37662 40514
rect 37714 40462 37726 40514
rect 41234 40462 41246 40514
rect 41298 40462 41310 40514
rect 42802 40462 42814 40514
rect 42866 40462 42878 40514
rect 46274 40462 46286 40514
rect 46338 40462 46350 40514
rect 47170 40462 47182 40514
rect 47234 40462 47246 40514
rect 51650 40462 51662 40514
rect 51714 40462 51726 40514
rect 36654 40450 36706 40462
rect 43038 40450 43090 40462
rect 2942 40402 2994 40414
rect 2594 40350 2606 40402
rect 2658 40350 2670 40402
rect 2942 40338 2994 40350
rect 3278 40402 3330 40414
rect 3278 40338 3330 40350
rect 3614 40402 3666 40414
rect 3614 40338 3666 40350
rect 5070 40402 5122 40414
rect 7646 40402 7698 40414
rect 11566 40402 11618 40414
rect 7298 40350 7310 40402
rect 7362 40350 7374 40402
rect 11106 40350 11118 40402
rect 11170 40350 11182 40402
rect 5070 40338 5122 40350
rect 7646 40338 7698 40350
rect 11566 40338 11618 40350
rect 11902 40402 11954 40414
rect 11902 40338 11954 40350
rect 12686 40402 12738 40414
rect 14590 40402 14642 40414
rect 13794 40350 13806 40402
rect 13858 40350 13870 40402
rect 14130 40350 14142 40402
rect 14194 40350 14206 40402
rect 12686 40338 12738 40350
rect 14590 40338 14642 40350
rect 14702 40402 14754 40414
rect 20190 40402 20242 40414
rect 23326 40402 23378 40414
rect 17378 40350 17390 40402
rect 17442 40350 17454 40402
rect 17938 40350 17950 40402
rect 18002 40350 18014 40402
rect 19058 40350 19070 40402
rect 19122 40350 19134 40402
rect 22418 40350 22430 40402
rect 22482 40350 22494 40402
rect 14702 40338 14754 40350
rect 20190 40338 20242 40350
rect 23326 40338 23378 40350
rect 29038 40402 29090 40414
rect 30158 40402 30210 40414
rect 29810 40350 29822 40402
rect 29874 40350 29886 40402
rect 29038 40338 29090 40350
rect 30158 40338 30210 40350
rect 30382 40402 30434 40414
rect 30382 40338 30434 40350
rect 31390 40402 31442 40414
rect 31390 40338 31442 40350
rect 31502 40402 31554 40414
rect 31502 40338 31554 40350
rect 33070 40402 33122 40414
rect 44606 40402 44658 40414
rect 33954 40350 33966 40402
rect 34018 40350 34030 40402
rect 35746 40350 35758 40402
rect 35810 40350 35822 40402
rect 41010 40350 41022 40402
rect 41074 40350 41086 40402
rect 43250 40350 43262 40402
rect 43314 40350 43326 40402
rect 33070 40338 33122 40350
rect 44606 40338 44658 40350
rect 44942 40402 44994 40414
rect 44942 40338 44994 40350
rect 46622 40402 46674 40414
rect 46622 40338 46674 40350
rect 46846 40402 46898 40414
rect 50206 40402 50258 40414
rect 47394 40350 47406 40402
rect 47458 40350 47470 40402
rect 49522 40350 49534 40402
rect 49586 40350 49598 40402
rect 51986 40350 51998 40402
rect 52050 40350 52062 40402
rect 52882 40350 52894 40402
rect 52946 40350 52958 40402
rect 54898 40350 54910 40402
rect 54962 40350 54974 40402
rect 46846 40338 46898 40350
rect 50206 40338 50258 40350
rect 2046 40290 2098 40302
rect 5182 40290 5234 40302
rect 14366 40290 14418 40302
rect 31726 40290 31778 40302
rect 42702 40290 42754 40302
rect 4050 40238 4062 40290
rect 4114 40238 4126 40290
rect 10210 40238 10222 40290
rect 10274 40238 10286 40290
rect 18386 40238 18398 40290
rect 18450 40238 18462 40290
rect 20962 40238 20974 40290
rect 21026 40238 21038 40290
rect 33842 40238 33854 40290
rect 33906 40238 33918 40290
rect 35858 40238 35870 40290
rect 35922 40238 35934 40290
rect 2046 40226 2098 40238
rect 5182 40226 5234 40238
rect 14366 40226 14418 40238
rect 31726 40226 31778 40238
rect 42702 40226 42754 40238
rect 44046 40290 44098 40302
rect 55582 40290 55634 40302
rect 49298 40238 49310 40290
rect 49362 40238 49374 40290
rect 55122 40238 55134 40290
rect 55186 40238 55198 40290
rect 44046 40226 44098 40238
rect 55582 40226 55634 40238
rect 12574 40178 12626 40190
rect 12574 40114 12626 40126
rect 43934 40178 43986 40190
rect 43934 40114 43986 40126
rect 54238 40178 54290 40190
rect 54238 40114 54290 40126
rect 1344 40010 58576 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 58576 40010
rect 1344 39924 58576 39958
rect 13918 39842 13970 39854
rect 13918 39778 13970 39790
rect 14366 39842 14418 39854
rect 14366 39778 14418 39790
rect 32286 39842 32338 39854
rect 32286 39778 32338 39790
rect 32846 39842 32898 39854
rect 32846 39778 32898 39790
rect 33854 39842 33906 39854
rect 33854 39778 33906 39790
rect 35870 39842 35922 39854
rect 35870 39778 35922 39790
rect 49870 39842 49922 39854
rect 49870 39778 49922 39790
rect 34078 39730 34130 39742
rect 49646 39730 49698 39742
rect 5730 39678 5742 39730
rect 5794 39678 5806 39730
rect 6514 39678 6526 39730
rect 6578 39678 6590 39730
rect 12674 39678 12686 39730
rect 12738 39678 12750 39730
rect 14690 39678 14702 39730
rect 14754 39678 14766 39730
rect 22530 39678 22542 39730
rect 22594 39678 22606 39730
rect 23426 39678 23438 39730
rect 23490 39678 23502 39730
rect 29474 39678 29486 39730
rect 29538 39678 29550 39730
rect 32050 39678 32062 39730
rect 32114 39678 32126 39730
rect 40674 39678 40686 39730
rect 40738 39678 40750 39730
rect 43698 39678 43710 39730
rect 43762 39678 43774 39730
rect 51538 39678 51550 39730
rect 51602 39678 51614 39730
rect 54226 39678 54238 39730
rect 54290 39678 54302 39730
rect 34078 39666 34130 39678
rect 49646 39666 49698 39678
rect 2270 39618 2322 39630
rect 5070 39618 5122 39630
rect 3826 39566 3838 39618
rect 3890 39566 3902 39618
rect 4386 39566 4398 39618
rect 4450 39566 4462 39618
rect 2270 39554 2322 39566
rect 5070 39554 5122 39566
rect 5182 39618 5234 39630
rect 8654 39618 8706 39630
rect 18286 39618 18338 39630
rect 5506 39566 5518 39618
rect 5570 39566 5582 39618
rect 6290 39566 6302 39618
rect 6354 39566 6366 39618
rect 9650 39566 9662 39618
rect 9714 39566 9726 39618
rect 11554 39566 11566 39618
rect 11618 39566 11630 39618
rect 5182 39554 5234 39566
rect 8654 39554 8706 39566
rect 18286 39554 18338 39566
rect 19070 39618 19122 39630
rect 28702 39618 28754 39630
rect 32622 39618 32674 39630
rect 22754 39566 22766 39618
rect 22818 39566 22830 39618
rect 23090 39566 23102 39618
rect 23154 39566 23166 39618
rect 29362 39566 29374 39618
rect 29426 39566 29438 39618
rect 31042 39566 31054 39618
rect 31106 39566 31118 39618
rect 31938 39566 31950 39618
rect 32002 39566 32014 39618
rect 19070 39554 19122 39566
rect 28702 39554 28754 39566
rect 32622 39554 32674 39566
rect 35982 39618 36034 39630
rect 35982 39554 36034 39566
rect 36430 39618 36482 39630
rect 36430 39554 36482 39566
rect 37438 39618 37490 39630
rect 37438 39554 37490 39566
rect 39566 39618 39618 39630
rect 39566 39554 39618 39566
rect 39678 39618 39730 39630
rect 42478 39618 42530 39630
rect 40338 39566 40350 39618
rect 40402 39566 40414 39618
rect 39678 39554 39730 39566
rect 42478 39554 42530 39566
rect 43598 39618 43650 39630
rect 43598 39554 43650 39566
rect 46286 39618 46338 39630
rect 46286 39554 46338 39566
rect 46958 39618 47010 39630
rect 55358 39618 55410 39630
rect 51090 39566 51102 39618
rect 51154 39566 51166 39618
rect 51426 39566 51438 39618
rect 51490 39566 51502 39618
rect 54002 39566 54014 39618
rect 54066 39566 54078 39618
rect 46958 39554 47010 39566
rect 55358 39554 55410 39566
rect 2942 39506 2994 39518
rect 2942 39442 2994 39454
rect 3054 39506 3106 39518
rect 14030 39506 14082 39518
rect 4834 39454 4846 39506
rect 4898 39454 4910 39506
rect 11106 39454 11118 39506
rect 11170 39454 11182 39506
rect 12002 39454 12014 39506
rect 12066 39454 12078 39506
rect 3054 39442 3106 39454
rect 14030 39442 14082 39454
rect 14590 39506 14642 39518
rect 14590 39442 14642 39454
rect 18622 39506 18674 39518
rect 18622 39442 18674 39454
rect 18958 39506 19010 39518
rect 18958 39442 19010 39454
rect 21870 39506 21922 39518
rect 21870 39442 21922 39454
rect 21982 39506 22034 39518
rect 21982 39442 22034 39454
rect 28366 39506 28418 39518
rect 28366 39442 28418 39454
rect 28478 39506 28530 39518
rect 28478 39442 28530 39454
rect 31502 39506 31554 39518
rect 31502 39442 31554 39454
rect 35870 39506 35922 39518
rect 35870 39442 35922 39454
rect 37326 39506 37378 39518
rect 37326 39442 37378 39454
rect 39790 39506 39842 39518
rect 39790 39442 39842 39454
rect 41134 39506 41186 39518
rect 41134 39442 41186 39454
rect 43150 39506 43202 39518
rect 43150 39442 43202 39454
rect 46622 39506 46674 39518
rect 54574 39506 54626 39518
rect 51762 39454 51774 39506
rect 51826 39454 51838 39506
rect 46622 39442 46674 39454
rect 54574 39442 54626 39454
rect 1710 39394 1762 39406
rect 1710 39330 1762 39342
rect 2718 39394 2770 39406
rect 13918 39394 13970 39406
rect 8306 39342 8318 39394
rect 8370 39342 8382 39394
rect 2718 39330 2770 39342
rect 13918 39330 13970 39342
rect 17950 39394 18002 39406
rect 17950 39330 18002 39342
rect 18174 39394 18226 39406
rect 18174 39330 18226 39342
rect 18846 39394 18898 39406
rect 18846 39330 18898 39342
rect 22206 39394 22258 39406
rect 22206 39330 22258 39342
rect 28142 39394 28194 39406
rect 37102 39394 37154 39406
rect 41470 39394 41522 39406
rect 33170 39342 33182 39394
rect 33234 39342 33246 39394
rect 33506 39342 33518 39394
rect 33570 39342 33582 39394
rect 39106 39342 39118 39394
rect 39170 39342 39182 39394
rect 28142 39330 28194 39342
rect 37102 39330 37154 39342
rect 41470 39330 41522 39342
rect 42254 39394 42306 39406
rect 43374 39394 43426 39406
rect 42802 39342 42814 39394
rect 42866 39342 42878 39394
rect 42254 39330 42306 39342
rect 43374 39330 43426 39342
rect 43710 39394 43762 39406
rect 46734 39394 46786 39406
rect 45938 39342 45950 39394
rect 46002 39342 46014 39394
rect 43710 39330 43762 39342
rect 46734 39330 46786 39342
rect 47294 39394 47346 39406
rect 55470 39394 55522 39406
rect 50194 39342 50206 39394
rect 50258 39342 50270 39394
rect 47294 39330 47346 39342
rect 55470 39330 55522 39342
rect 55694 39394 55746 39406
rect 55694 39330 55746 39342
rect 1344 39226 58576 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 50558 39226
rect 50610 39174 50662 39226
rect 50714 39174 50766 39226
rect 50818 39174 58576 39226
rect 1344 39140 58576 39174
rect 2046 39058 2098 39070
rect 3054 39058 3106 39070
rect 2706 39006 2718 39058
rect 2770 39006 2782 39058
rect 2046 38994 2098 39006
rect 3054 38994 3106 39006
rect 3726 39058 3778 39070
rect 3726 38994 3778 39006
rect 4734 39058 4786 39070
rect 4734 38994 4786 39006
rect 5854 39058 5906 39070
rect 5854 38994 5906 39006
rect 6974 39058 7026 39070
rect 6974 38994 7026 39006
rect 8430 39058 8482 39070
rect 10782 39058 10834 39070
rect 8754 39006 8766 39058
rect 8818 39006 8830 39058
rect 8430 38994 8482 39006
rect 10782 38994 10834 39006
rect 11006 39058 11058 39070
rect 11006 38994 11058 39006
rect 13246 39058 13298 39070
rect 13246 38994 13298 39006
rect 13470 39058 13522 39070
rect 28702 39058 28754 39070
rect 16818 39006 16830 39058
rect 16882 39006 16894 39058
rect 13470 38994 13522 39006
rect 28702 38994 28754 39006
rect 30382 39058 30434 39070
rect 44830 39058 44882 39070
rect 42914 39006 42926 39058
rect 42978 39006 42990 39058
rect 30382 38994 30434 39006
rect 44830 38994 44882 39006
rect 45166 39058 45218 39070
rect 45166 38994 45218 39006
rect 51102 39058 51154 39070
rect 51102 38994 51154 39006
rect 4622 38946 4674 38958
rect 4622 38882 4674 38894
rect 6414 38946 6466 38958
rect 6414 38882 6466 38894
rect 6526 38946 6578 38958
rect 6526 38882 6578 38894
rect 6862 38946 6914 38958
rect 6862 38882 6914 38894
rect 10110 38946 10162 38958
rect 10110 38882 10162 38894
rect 10222 38946 10274 38958
rect 10222 38882 10274 38894
rect 10558 38946 10610 38958
rect 25454 38946 25506 38958
rect 14130 38894 14142 38946
rect 14194 38894 14206 38946
rect 17938 38894 17950 38946
rect 18002 38894 18014 38946
rect 18610 38894 18622 38946
rect 18674 38894 18686 38946
rect 21970 38894 21982 38946
rect 22034 38894 22046 38946
rect 23650 38894 23662 38946
rect 23714 38894 23726 38946
rect 10558 38882 10610 38894
rect 25454 38882 25506 38894
rect 29038 38946 29090 38958
rect 29038 38882 29090 38894
rect 29374 38946 29426 38958
rect 29374 38882 29426 38894
rect 29822 38946 29874 38958
rect 29822 38882 29874 38894
rect 29934 38946 29986 38958
rect 29934 38882 29986 38894
rect 31502 38946 31554 38958
rect 42254 38946 42306 38958
rect 46734 38946 46786 38958
rect 37090 38894 37102 38946
rect 37154 38894 37166 38946
rect 38434 38894 38446 38946
rect 38498 38894 38510 38946
rect 39666 38894 39678 38946
rect 39730 38894 39742 38946
rect 41010 38894 41022 38946
rect 41074 38894 41086 38946
rect 45490 38894 45502 38946
rect 45554 38894 45566 38946
rect 31502 38882 31554 38894
rect 42254 38882 42306 38894
rect 46734 38882 46786 38894
rect 47070 38946 47122 38958
rect 51538 38894 51550 38946
rect 51602 38894 51614 38946
rect 47070 38882 47122 38894
rect 4286 38834 4338 38846
rect 1810 38782 1822 38834
rect 1874 38782 1886 38834
rect 4286 38770 4338 38782
rect 5742 38834 5794 38846
rect 5742 38770 5794 38782
rect 6078 38834 6130 38846
rect 12014 38834 12066 38846
rect 12798 38834 12850 38846
rect 20526 38834 20578 38846
rect 22318 38834 22370 38846
rect 11218 38782 11230 38834
rect 11282 38782 11294 38834
rect 12226 38782 12238 38834
rect 12290 38782 12302 38834
rect 15362 38782 15374 38834
rect 15426 38782 15438 38834
rect 16594 38782 16606 38834
rect 16658 38782 16670 38834
rect 17714 38782 17726 38834
rect 17778 38782 17790 38834
rect 19842 38782 19854 38834
rect 19906 38782 19918 38834
rect 20850 38782 20862 38834
rect 20914 38782 20926 38834
rect 21858 38782 21870 38834
rect 21922 38782 21934 38834
rect 6078 38770 6130 38782
rect 12014 38770 12066 38782
rect 12798 38770 12850 38782
rect 20526 38770 20578 38782
rect 22318 38770 22370 38782
rect 22542 38834 22594 38846
rect 22542 38770 22594 38782
rect 22766 38834 22818 38846
rect 22766 38770 22818 38782
rect 23214 38834 23266 38846
rect 31838 38834 31890 38846
rect 35198 38834 35250 38846
rect 23426 38782 23438 38834
rect 23490 38782 23502 38834
rect 35074 38782 35086 38834
rect 35138 38782 35150 38834
rect 23214 38770 23266 38782
rect 31838 38770 31890 38782
rect 35198 38770 35250 38782
rect 38670 38834 38722 38846
rect 41918 38834 41970 38846
rect 45838 38834 45890 38846
rect 38994 38782 39006 38834
rect 39058 38782 39070 38834
rect 39890 38782 39902 38834
rect 39954 38782 39966 38834
rect 40898 38782 40910 38834
rect 40962 38782 40974 38834
rect 43138 38782 43150 38834
rect 43202 38782 43214 38834
rect 38670 38770 38722 38782
rect 41918 38770 41970 38782
rect 45838 38770 45890 38782
rect 46062 38834 46114 38846
rect 50094 38834 50146 38846
rect 49186 38782 49198 38834
rect 49250 38782 49262 38834
rect 46062 38770 46114 38782
rect 50094 38770 50146 38782
rect 50318 38834 50370 38846
rect 50318 38770 50370 38782
rect 51774 38834 51826 38846
rect 51774 38770 51826 38782
rect 52222 38834 52274 38846
rect 53778 38782 53790 38834
rect 53842 38782 53854 38834
rect 55122 38782 55134 38834
rect 55186 38782 55198 38834
rect 52222 38770 52274 38782
rect 10894 38722 10946 38734
rect 10894 38658 10946 38670
rect 11902 38722 11954 38734
rect 11902 38658 11954 38670
rect 13358 38722 13410 38734
rect 16046 38722 16098 38734
rect 25230 38722 25282 38734
rect 13906 38670 13918 38722
rect 13970 38670 13982 38722
rect 18386 38670 18398 38722
rect 18450 38670 18462 38722
rect 21522 38670 21534 38722
rect 21586 38670 21598 38722
rect 23538 38670 23550 38722
rect 23602 38670 23614 38722
rect 13358 38658 13410 38670
rect 16046 38658 16098 38670
rect 25230 38658 25282 38670
rect 31614 38722 31666 38734
rect 31614 38658 31666 38670
rect 31950 38722 32002 38734
rect 48750 38722 48802 38734
rect 51438 38722 51490 38734
rect 57822 38722 57874 38734
rect 34738 38670 34750 38722
rect 34802 38670 34814 38722
rect 36530 38670 36542 38722
rect 36594 38670 36606 38722
rect 39442 38670 39454 38722
rect 39506 38670 39518 38722
rect 41458 38670 41470 38722
rect 41522 38670 41534 38722
rect 46386 38670 46398 38722
rect 46450 38670 46462 38722
rect 49522 38670 49534 38722
rect 49586 38670 49598 38722
rect 54002 38670 54014 38722
rect 54066 38670 54078 38722
rect 31950 38658 32002 38670
rect 48750 38658 48802 38670
rect 51438 38658 51490 38670
rect 57822 38658 57874 38670
rect 58270 38722 58322 38734
rect 58270 38658 58322 38670
rect 4734 38610 4786 38622
rect 4734 38546 4786 38558
rect 6414 38610 6466 38622
rect 6414 38546 6466 38558
rect 6974 38610 7026 38622
rect 6974 38546 7026 38558
rect 10110 38610 10162 38622
rect 10110 38546 10162 38558
rect 25566 38610 25618 38622
rect 25566 38546 25618 38558
rect 29822 38610 29874 38622
rect 52446 38610 52498 38622
rect 34514 38558 34526 38610
rect 34578 38558 34590 38610
rect 50642 38558 50654 38610
rect 50706 38558 50718 38610
rect 55794 38558 55806 38610
rect 55858 38558 55870 38610
rect 29822 38546 29874 38558
rect 52446 38546 52498 38558
rect 1344 38442 58576 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 58576 38442
rect 1344 38356 58576 38390
rect 14366 38274 14418 38286
rect 14366 38210 14418 38222
rect 14590 38274 14642 38286
rect 14590 38210 14642 38222
rect 24334 38274 24386 38286
rect 24334 38210 24386 38222
rect 39678 38274 39730 38286
rect 39678 38210 39730 38222
rect 41806 38274 41858 38286
rect 41806 38210 41858 38222
rect 50542 38274 50594 38286
rect 50542 38210 50594 38222
rect 54910 38274 54962 38286
rect 54910 38210 54962 38222
rect 1822 38162 1874 38174
rect 1822 38098 1874 38110
rect 2270 38162 2322 38174
rect 14142 38162 14194 38174
rect 21870 38162 21922 38174
rect 30158 38162 30210 38174
rect 6066 38110 6078 38162
rect 6130 38110 6142 38162
rect 8866 38110 8878 38162
rect 8930 38110 8942 38162
rect 11106 38110 11118 38162
rect 11170 38110 11182 38162
rect 18498 38110 18510 38162
rect 18562 38110 18574 38162
rect 21970 38110 21982 38162
rect 22034 38110 22046 38162
rect 25554 38110 25566 38162
rect 25618 38110 25630 38162
rect 29586 38110 29598 38162
rect 29650 38110 29662 38162
rect 2270 38098 2322 38110
rect 14142 38098 14194 38110
rect 21870 38098 21922 38110
rect 30158 38098 30210 38110
rect 45950 38162 46002 38174
rect 45950 38098 46002 38110
rect 51214 38162 51266 38174
rect 51214 38098 51266 38110
rect 54686 38162 54738 38174
rect 54686 38098 54738 38110
rect 3838 38050 3890 38062
rect 2146 37998 2158 38050
rect 2210 37998 2222 38050
rect 3378 37998 3390 38050
rect 3442 37998 3454 38050
rect 3838 37986 3890 37998
rect 4734 38050 4786 38062
rect 8206 38050 8258 38062
rect 9662 38050 9714 38062
rect 7634 37998 7646 38050
rect 7698 37998 7710 38050
rect 8754 37998 8766 38050
rect 8818 37998 8830 38050
rect 4734 37986 4786 37998
rect 8206 37986 8258 37998
rect 9662 37986 9714 37998
rect 9998 38050 10050 38062
rect 9998 37986 10050 37998
rect 10334 38050 10386 38062
rect 24110 38050 24162 38062
rect 28254 38050 28306 38062
rect 32734 38050 32786 38062
rect 10882 37998 10894 38050
rect 10946 37998 10958 38050
rect 16706 37998 16718 38050
rect 16770 37998 16782 38050
rect 17154 37998 17166 38050
rect 17218 37998 17230 38050
rect 18722 37998 18734 38050
rect 18786 37998 18798 38050
rect 22194 37998 22206 38050
rect 22258 37998 22270 38050
rect 23874 37998 23886 38050
rect 23938 37998 23950 38050
rect 24994 37998 25006 38050
rect 25058 37998 25070 38050
rect 29810 37998 29822 38050
rect 29874 37998 29886 38050
rect 10334 37986 10386 37998
rect 24110 37986 24162 37998
rect 28254 37986 28306 37998
rect 32734 37986 32786 37998
rect 33630 38050 33682 38062
rect 33630 37986 33682 37998
rect 33966 38050 34018 38062
rect 33966 37986 34018 37998
rect 34862 38050 34914 38062
rect 34862 37986 34914 37998
rect 35086 38050 35138 38062
rect 35086 37986 35138 37998
rect 35534 38050 35586 38062
rect 41582 38050 41634 38062
rect 39106 37998 39118 38050
rect 39170 37998 39182 38050
rect 39330 37998 39342 38050
rect 39394 37998 39406 38050
rect 40226 37998 40238 38050
rect 40290 37998 40302 38050
rect 41122 37998 41134 38050
rect 41186 37998 41198 38050
rect 35534 37986 35586 37998
rect 41582 37986 41634 37998
rect 43598 38050 43650 38062
rect 43598 37986 43650 37998
rect 46622 38050 46674 38062
rect 51438 38050 51490 38062
rect 48514 37998 48526 38050
rect 48578 37998 48590 38050
rect 53218 37998 53230 38050
rect 53282 37998 53294 38050
rect 54226 37998 54238 38050
rect 54290 37998 54302 38050
rect 58034 37998 58046 38050
rect 58098 37998 58110 38050
rect 46622 37986 46674 37998
rect 51438 37986 51490 37998
rect 3950 37938 4002 37950
rect 11566 37938 11618 37950
rect 19406 37938 19458 37950
rect 5058 37886 5070 37938
rect 5122 37886 5134 37938
rect 6402 37886 6414 37938
rect 6466 37886 6478 37938
rect 16258 37886 16270 37938
rect 16322 37886 16334 37938
rect 3950 37874 4002 37886
rect 11566 37874 11618 37886
rect 19406 37874 19458 37886
rect 24446 37938 24498 37950
rect 24446 37874 24498 37886
rect 25902 37938 25954 37950
rect 25902 37874 25954 37886
rect 33294 37938 33346 37950
rect 33294 37874 33346 37886
rect 34302 37938 34354 37950
rect 34302 37874 34354 37886
rect 39566 37938 39618 37950
rect 42478 37938 42530 37950
rect 41234 37886 41246 37938
rect 41298 37886 41310 37938
rect 39566 37874 39618 37886
rect 42478 37874 42530 37886
rect 42702 37938 42754 37950
rect 42702 37874 42754 37886
rect 44158 37938 44210 37950
rect 44158 37874 44210 37886
rect 46286 37938 46338 37950
rect 46286 37874 46338 37886
rect 46398 37938 46450 37950
rect 46398 37874 46450 37886
rect 47070 37938 47122 37950
rect 47070 37874 47122 37886
rect 47406 37938 47458 37950
rect 55806 37938 55858 37950
rect 48290 37886 48302 37938
rect 48354 37886 48366 37938
rect 49634 37886 49646 37938
rect 49698 37886 49710 37938
rect 54002 37886 54014 37938
rect 54066 37886 54078 37938
rect 47406 37874 47458 37886
rect 55806 37874 55858 37886
rect 55918 37938 55970 37950
rect 55918 37874 55970 37886
rect 57486 37938 57538 37950
rect 57486 37874 57538 37886
rect 57822 37938 57874 37950
rect 57822 37874 57874 37886
rect 2382 37826 2434 37838
rect 2382 37762 2434 37774
rect 2606 37826 2658 37838
rect 2606 37762 2658 37774
rect 10110 37826 10162 37838
rect 10110 37762 10162 37774
rect 15038 37826 15090 37838
rect 17502 37826 17554 37838
rect 17378 37774 17390 37826
rect 17442 37774 17454 37826
rect 15038 37762 15090 37774
rect 17502 37762 17554 37774
rect 28590 37826 28642 37838
rect 28590 37762 28642 37774
rect 33182 37826 33234 37838
rect 33182 37762 33234 37774
rect 33406 37826 33458 37838
rect 33406 37762 33458 37774
rect 33854 37826 33906 37838
rect 33854 37762 33906 37774
rect 34974 37826 35026 37838
rect 42590 37826 42642 37838
rect 40338 37774 40350 37826
rect 40402 37774 40414 37826
rect 42130 37774 42142 37826
rect 42194 37774 42206 37826
rect 34974 37762 35026 37774
rect 42590 37762 42642 37774
rect 43262 37826 43314 37838
rect 43262 37762 43314 37774
rect 43822 37826 43874 37838
rect 43822 37762 43874 37774
rect 44046 37826 44098 37838
rect 44046 37762 44098 37774
rect 44942 37826 44994 37838
rect 44942 37762 44994 37774
rect 47182 37826 47234 37838
rect 50318 37826 50370 37838
rect 49522 37774 49534 37826
rect 49586 37774 49598 37826
rect 47182 37762 47234 37774
rect 50318 37762 50370 37774
rect 50430 37826 50482 37838
rect 56142 37826 56194 37838
rect 51762 37774 51774 37826
rect 51826 37774 51838 37826
rect 53442 37774 53454 37826
rect 53506 37774 53518 37826
rect 55234 37774 55246 37826
rect 55298 37774 55310 37826
rect 50430 37762 50482 37774
rect 56142 37762 56194 37774
rect 56926 37826 56978 37838
rect 56926 37762 56978 37774
rect 57150 37826 57202 37838
rect 57150 37762 57202 37774
rect 1344 37658 58576 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 50558 37658
rect 50610 37606 50662 37658
rect 50714 37606 50766 37658
rect 50818 37606 58576 37658
rect 1344 37572 58576 37606
rect 2270 37490 2322 37502
rect 2270 37426 2322 37438
rect 6078 37490 6130 37502
rect 6078 37426 6130 37438
rect 6750 37490 6802 37502
rect 8542 37490 8594 37502
rect 7074 37438 7086 37490
rect 7138 37438 7150 37490
rect 13470 37490 13522 37502
rect 6750 37426 6802 37438
rect 8542 37426 8594 37438
rect 9774 37434 9826 37446
rect 2830 37378 2882 37390
rect 2830 37314 2882 37326
rect 2942 37378 2994 37390
rect 2942 37314 2994 37326
rect 3054 37378 3106 37390
rect 8766 37378 8818 37390
rect 9662 37378 9714 37390
rect 6402 37326 6414 37378
rect 6466 37326 6478 37378
rect 8866 37326 8878 37378
rect 8930 37375 8942 37378
rect 9090 37375 9102 37378
rect 8930 37329 9102 37375
rect 8930 37326 8942 37329
rect 9090 37326 9102 37329
rect 9154 37326 9166 37378
rect 13470 37426 13522 37438
rect 14478 37490 14530 37502
rect 14478 37426 14530 37438
rect 16494 37490 16546 37502
rect 16494 37426 16546 37438
rect 20078 37490 20130 37502
rect 20078 37426 20130 37438
rect 29598 37490 29650 37502
rect 29598 37426 29650 37438
rect 29822 37490 29874 37502
rect 29822 37426 29874 37438
rect 30494 37490 30546 37502
rect 30494 37426 30546 37438
rect 30942 37490 30994 37502
rect 30942 37426 30994 37438
rect 32062 37490 32114 37502
rect 32062 37426 32114 37438
rect 34414 37490 34466 37502
rect 34414 37426 34466 37438
rect 39790 37490 39842 37502
rect 39790 37426 39842 37438
rect 40462 37490 40514 37502
rect 40462 37426 40514 37438
rect 43486 37490 43538 37502
rect 43486 37426 43538 37438
rect 43934 37490 43986 37502
rect 43934 37426 43986 37438
rect 57822 37490 57874 37502
rect 57822 37426 57874 37438
rect 9774 37370 9826 37382
rect 12462 37378 12514 37390
rect 3054 37314 3106 37326
rect 8766 37314 8818 37326
rect 9662 37314 9714 37326
rect 12462 37314 12514 37326
rect 14590 37378 14642 37390
rect 14590 37314 14642 37326
rect 19966 37378 20018 37390
rect 28478 37378 28530 37390
rect 25890 37326 25902 37378
rect 25954 37326 25966 37378
rect 19966 37314 20018 37326
rect 28478 37314 28530 37326
rect 28814 37378 28866 37390
rect 28814 37314 28866 37326
rect 29262 37378 29314 37390
rect 29262 37314 29314 37326
rect 29374 37378 29426 37390
rect 29374 37314 29426 37326
rect 29934 37378 29986 37390
rect 29934 37314 29986 37326
rect 32398 37378 32450 37390
rect 32398 37314 32450 37326
rect 32510 37378 32562 37390
rect 32510 37314 32562 37326
rect 33630 37378 33682 37390
rect 33630 37314 33682 37326
rect 35534 37378 35586 37390
rect 35534 37314 35586 37326
rect 40126 37378 40178 37390
rect 40126 37314 40178 37326
rect 40238 37378 40290 37390
rect 43374 37378 43426 37390
rect 56590 37378 56642 37390
rect 41458 37326 41470 37378
rect 41522 37326 41534 37378
rect 44258 37326 44270 37378
rect 44322 37326 44334 37378
rect 52210 37326 52222 37378
rect 52274 37326 52286 37378
rect 40238 37314 40290 37326
rect 43374 37314 43426 37326
rect 56590 37314 56642 37326
rect 4174 37266 4226 37278
rect 4174 37202 4226 37214
rect 4398 37266 4450 37278
rect 14030 37266 14082 37278
rect 10322 37214 10334 37266
rect 10386 37214 10398 37266
rect 11666 37214 11678 37266
rect 11730 37214 11742 37266
rect 4398 37202 4450 37214
rect 14030 37202 14082 37214
rect 14254 37266 14306 37278
rect 14254 37202 14306 37214
rect 16158 37266 16210 37278
rect 16158 37202 16210 37214
rect 16270 37266 16322 37278
rect 16270 37202 16322 37214
rect 16606 37266 16658 37278
rect 19070 37266 19122 37278
rect 17490 37214 17502 37266
rect 17554 37214 17566 37266
rect 18386 37214 18398 37266
rect 18450 37214 18462 37266
rect 16606 37202 16658 37214
rect 19070 37202 19122 37214
rect 19294 37266 19346 37278
rect 19294 37202 19346 37214
rect 19518 37266 19570 37278
rect 19518 37202 19570 37214
rect 20302 37266 20354 37278
rect 20302 37202 20354 37214
rect 23326 37266 23378 37278
rect 33406 37266 33458 37278
rect 23538 37214 23550 37266
rect 23602 37214 23614 37266
rect 25218 37214 25230 37266
rect 25282 37214 25294 37266
rect 25778 37214 25790 37266
rect 25842 37214 25854 37266
rect 23326 37202 23378 37214
rect 33406 37202 33458 37214
rect 34302 37266 34354 37278
rect 43710 37266 43762 37278
rect 49198 37266 49250 37278
rect 55134 37266 55186 37278
rect 56814 37266 56866 37278
rect 34514 37214 34526 37266
rect 34578 37214 34590 37266
rect 36306 37214 36318 37266
rect 36370 37214 36382 37266
rect 37314 37214 37326 37266
rect 37378 37214 37390 37266
rect 41794 37214 41806 37266
rect 41858 37214 41870 37266
rect 42354 37214 42366 37266
rect 42418 37214 42430 37266
rect 45042 37214 45054 37266
rect 45106 37214 45118 37266
rect 46722 37214 46734 37266
rect 46786 37214 46798 37266
rect 49522 37214 49534 37266
rect 49586 37214 49598 37266
rect 50642 37214 50654 37266
rect 50706 37214 50718 37266
rect 51090 37214 51102 37266
rect 51154 37214 51166 37266
rect 52434 37214 52446 37266
rect 52498 37214 52510 37266
rect 53218 37214 53230 37266
rect 53282 37214 53294 37266
rect 55346 37214 55358 37266
rect 55410 37214 55422 37266
rect 34302 37202 34354 37214
rect 43710 37202 43762 37214
rect 49198 37202 49250 37214
rect 55134 37202 55186 37214
rect 56814 37202 56866 37214
rect 57150 37266 57202 37278
rect 57150 37202 57202 37214
rect 58158 37266 58210 37278
rect 58158 37202 58210 37214
rect 1822 37154 1874 37166
rect 1822 37090 1874 37102
rect 8654 37154 8706 37166
rect 16382 37154 16434 37166
rect 19182 37154 19234 37166
rect 45614 37154 45666 37166
rect 56702 37154 56754 37166
rect 10210 37102 10222 37154
rect 10274 37102 10286 37154
rect 17938 37102 17950 37154
rect 18002 37102 18014 37154
rect 26002 37102 26014 37154
rect 26066 37102 26078 37154
rect 37762 37102 37774 37154
rect 37826 37102 37838 37154
rect 41682 37102 41694 37154
rect 41746 37102 41758 37154
rect 44706 37102 44718 37154
rect 44770 37102 44782 37154
rect 47058 37102 47070 37154
rect 47122 37102 47134 37154
rect 50418 37102 50430 37154
rect 50482 37102 50494 37154
rect 54226 37102 54238 37154
rect 54290 37102 54302 37154
rect 8654 37090 8706 37102
rect 16382 37090 16434 37102
rect 19182 37090 19234 37102
rect 45614 37090 45666 37102
rect 56702 37090 56754 37102
rect 9662 37042 9714 37054
rect 29262 37042 29314 37054
rect 3490 36990 3502 37042
rect 3554 36990 3566 37042
rect 3826 36990 3838 37042
rect 3890 36990 3902 37042
rect 18386 36990 18398 37042
rect 18450 36990 18462 37042
rect 23986 36990 23998 37042
rect 24050 36990 24062 37042
rect 9662 36978 9714 36990
rect 29262 36978 29314 36990
rect 32398 37042 32450 37054
rect 32398 36978 32450 36990
rect 33070 37042 33122 37054
rect 33070 36978 33122 36990
rect 34078 37042 34130 37054
rect 46386 36990 46398 37042
rect 46450 36990 46462 37042
rect 50306 36990 50318 37042
rect 50370 36990 50382 37042
rect 55010 36990 55022 37042
rect 55074 36990 55086 37042
rect 34078 36978 34130 36990
rect 1344 36874 58576 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 58576 36874
rect 1344 36788 58576 36822
rect 10334 36706 10386 36718
rect 10334 36642 10386 36654
rect 23438 36706 23490 36718
rect 23438 36642 23490 36654
rect 24558 36706 24610 36718
rect 53006 36706 53058 36718
rect 33730 36654 33742 36706
rect 33794 36654 33806 36706
rect 24558 36642 24610 36654
rect 53006 36642 53058 36654
rect 54462 36706 54514 36718
rect 54462 36642 54514 36654
rect 20750 36594 20802 36606
rect 3826 36542 3838 36594
rect 3890 36542 3902 36594
rect 4386 36542 4398 36594
rect 4450 36542 4462 36594
rect 8866 36542 8878 36594
rect 8930 36542 8942 36594
rect 18610 36542 18622 36594
rect 18674 36542 18686 36594
rect 20750 36530 20802 36542
rect 21310 36594 21362 36606
rect 21310 36530 21362 36542
rect 23214 36594 23266 36606
rect 41470 36594 41522 36606
rect 25330 36542 25342 36594
rect 25394 36542 25406 36594
rect 29474 36542 29486 36594
rect 29538 36542 29550 36594
rect 23214 36530 23266 36542
rect 41470 36530 41522 36542
rect 53230 36594 53282 36606
rect 57026 36542 57038 36594
rect 57090 36542 57102 36594
rect 53230 36530 53282 36542
rect 2830 36482 2882 36494
rect 7422 36482 7474 36494
rect 9438 36482 9490 36494
rect 3490 36430 3502 36482
rect 3554 36430 3566 36482
rect 4162 36430 4174 36482
rect 4226 36430 4238 36482
rect 8306 36430 8318 36482
rect 8370 36430 8382 36482
rect 8642 36430 8654 36482
rect 8706 36430 8718 36482
rect 2830 36418 2882 36430
rect 7422 36418 7474 36430
rect 9438 36418 9490 36430
rect 10222 36482 10274 36494
rect 10222 36418 10274 36430
rect 12238 36482 12290 36494
rect 12238 36418 12290 36430
rect 12350 36482 12402 36494
rect 12350 36418 12402 36430
rect 12462 36482 12514 36494
rect 17950 36482 18002 36494
rect 21534 36482 21586 36494
rect 14242 36430 14254 36482
rect 14306 36430 14318 36482
rect 15138 36430 15150 36482
rect 15202 36430 15214 36482
rect 20178 36430 20190 36482
rect 20242 36430 20254 36482
rect 12462 36418 12514 36430
rect 17950 36418 18002 36430
rect 21534 36418 21586 36430
rect 21758 36482 21810 36494
rect 21758 36418 21810 36430
rect 22206 36482 22258 36494
rect 22206 36418 22258 36430
rect 22654 36482 22706 36494
rect 24782 36482 24834 36494
rect 32734 36482 32786 36494
rect 36430 36482 36482 36494
rect 24322 36430 24334 36482
rect 24386 36430 24398 36482
rect 25778 36430 25790 36482
rect 25842 36430 25854 36482
rect 29362 36430 29374 36482
rect 29426 36430 29438 36482
rect 30818 36430 30830 36482
rect 30882 36430 30894 36482
rect 32386 36430 32398 36482
rect 32450 36430 32462 36482
rect 33506 36430 33518 36482
rect 33570 36430 33582 36482
rect 22654 36418 22706 36430
rect 24782 36418 24834 36430
rect 32734 36418 32786 36430
rect 36430 36418 36482 36430
rect 37102 36482 37154 36494
rect 38334 36482 38386 36494
rect 37650 36430 37662 36482
rect 37714 36430 37726 36482
rect 37102 36418 37154 36430
rect 38334 36418 38386 36430
rect 38446 36482 38498 36494
rect 38446 36418 38498 36430
rect 39006 36482 39058 36494
rect 39006 36418 39058 36430
rect 40686 36482 40738 36494
rect 40686 36418 40738 36430
rect 41582 36482 41634 36494
rect 41582 36418 41634 36430
rect 41918 36482 41970 36494
rect 41918 36418 41970 36430
rect 44046 36482 44098 36494
rect 44046 36418 44098 36430
rect 44382 36482 44434 36494
rect 46286 36482 46338 36494
rect 44818 36430 44830 36482
rect 44882 36430 44894 36482
rect 45714 36430 45726 36482
rect 45778 36430 45790 36482
rect 44382 36418 44434 36430
rect 46286 36418 46338 36430
rect 46622 36482 46674 36494
rect 46622 36418 46674 36430
rect 47070 36482 47122 36494
rect 47070 36418 47122 36430
rect 50318 36482 50370 36494
rect 54574 36482 54626 36494
rect 51426 36430 51438 36482
rect 51490 36430 51502 36482
rect 51874 36430 51886 36482
rect 51938 36430 51950 36482
rect 50318 36418 50370 36430
rect 54574 36418 54626 36430
rect 1710 36370 1762 36382
rect 1710 36306 1762 36318
rect 2718 36370 2770 36382
rect 9662 36370 9714 36382
rect 8754 36318 8766 36370
rect 8818 36318 8830 36370
rect 2718 36306 2770 36318
rect 9662 36306 9714 36318
rect 9774 36370 9826 36382
rect 9774 36306 9826 36318
rect 10334 36370 10386 36382
rect 18062 36370 18114 36382
rect 14018 36318 14030 36370
rect 14082 36318 14094 36370
rect 16482 36318 16494 36370
rect 16546 36318 16558 36370
rect 10334 36306 10386 36318
rect 18062 36306 18114 36318
rect 18286 36370 18338 36382
rect 26238 36370 26290 36382
rect 18946 36318 18958 36370
rect 19010 36318 19022 36370
rect 23762 36318 23774 36370
rect 23826 36318 23838 36370
rect 23986 36318 23998 36370
rect 24050 36367 24062 36370
rect 24322 36367 24334 36370
rect 24050 36321 24334 36367
rect 24050 36318 24062 36321
rect 24322 36318 24334 36321
rect 24386 36318 24398 36370
rect 18286 36306 18338 36318
rect 26238 36306 26290 36318
rect 30270 36370 30322 36382
rect 30270 36306 30322 36318
rect 36990 36370 37042 36382
rect 36990 36306 37042 36318
rect 40574 36370 40626 36382
rect 40574 36306 40626 36318
rect 41134 36370 41186 36382
rect 41134 36306 41186 36318
rect 42030 36370 42082 36382
rect 42030 36306 42082 36318
rect 43486 36370 43538 36382
rect 43486 36306 43538 36318
rect 43598 36370 43650 36382
rect 48302 36370 48354 36382
rect 54462 36370 54514 36382
rect 58158 36370 58210 36382
rect 45266 36318 45278 36370
rect 45330 36318 45342 36370
rect 51202 36318 51214 36370
rect 51266 36318 51278 36370
rect 56466 36318 56478 36370
rect 56530 36318 56542 36370
rect 43598 36306 43650 36318
rect 48302 36306 48354 36318
rect 54462 36306 54514 36318
rect 58158 36306 58210 36318
rect 2046 36258 2098 36270
rect 2046 36194 2098 36206
rect 2494 36258 2546 36270
rect 2494 36194 2546 36206
rect 7086 36258 7138 36270
rect 7086 36194 7138 36206
rect 7310 36258 7362 36270
rect 7310 36194 7362 36206
rect 10894 36258 10946 36270
rect 22318 36258 22370 36270
rect 12898 36206 12910 36258
rect 12962 36206 12974 36258
rect 10894 36194 10946 36206
rect 22318 36194 22370 36206
rect 22542 36258 22594 36270
rect 22542 36194 22594 36206
rect 24446 36258 24498 36270
rect 36094 36258 36146 36270
rect 31042 36206 31054 36258
rect 31106 36206 31118 36258
rect 24446 36194 24498 36206
rect 36094 36194 36146 36206
rect 38558 36258 38610 36270
rect 38558 36194 38610 36206
rect 40350 36258 40402 36270
rect 40350 36194 40402 36206
rect 41358 36258 41410 36270
rect 41358 36194 41410 36206
rect 42254 36258 42306 36270
rect 42254 36194 42306 36206
rect 43262 36258 43314 36270
rect 43262 36194 43314 36206
rect 44158 36258 44210 36270
rect 46398 36258 46450 36270
rect 48414 36258 48466 36270
rect 45826 36206 45838 36258
rect 45890 36206 45902 36258
rect 47394 36206 47406 36258
rect 47458 36206 47470 36258
rect 44158 36194 44210 36206
rect 46398 36194 46450 36206
rect 48414 36194 48466 36206
rect 48526 36258 48578 36270
rect 55694 36258 55746 36270
rect 49970 36206 49982 36258
rect 50034 36206 50046 36258
rect 51986 36206 51998 36258
rect 52050 36206 52062 36258
rect 52658 36206 52670 36258
rect 52722 36206 52734 36258
rect 48526 36194 48578 36206
rect 55694 36194 55746 36206
rect 57822 36258 57874 36270
rect 57822 36194 57874 36206
rect 1344 36090 58576 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 50558 36090
rect 50610 36038 50662 36090
rect 50714 36038 50766 36090
rect 50818 36038 58576 36090
rect 1344 36004 58576 36038
rect 4734 35922 4786 35934
rect 17502 35922 17554 35934
rect 13906 35870 13918 35922
rect 13970 35870 13982 35922
rect 4734 35858 4786 35870
rect 17502 35858 17554 35870
rect 20638 35922 20690 35934
rect 20638 35858 20690 35870
rect 23438 35922 23490 35934
rect 23438 35858 23490 35870
rect 24558 35922 24610 35934
rect 24558 35858 24610 35870
rect 28254 35922 28306 35934
rect 28254 35858 28306 35870
rect 28478 35922 28530 35934
rect 28478 35858 28530 35870
rect 33742 35922 33794 35934
rect 44606 35922 44658 35934
rect 37874 35870 37886 35922
rect 37938 35870 37950 35922
rect 33742 35858 33794 35870
rect 44606 35858 44658 35870
rect 49086 35922 49138 35934
rect 49086 35858 49138 35870
rect 50766 35922 50818 35934
rect 50766 35858 50818 35870
rect 50990 35922 51042 35934
rect 50990 35858 51042 35870
rect 51326 35922 51378 35934
rect 51326 35858 51378 35870
rect 4958 35810 5010 35822
rect 8206 35810 8258 35822
rect 28926 35810 28978 35822
rect 2482 35758 2494 35810
rect 2546 35758 2558 35810
rect 6066 35758 6078 35810
rect 6130 35758 6142 35810
rect 13010 35758 13022 35810
rect 13074 35758 13086 35810
rect 16594 35758 16606 35810
rect 16658 35758 16670 35810
rect 17602 35758 17614 35810
rect 17666 35758 17678 35810
rect 22530 35758 22542 35810
rect 22594 35758 22606 35810
rect 4958 35746 5010 35758
rect 8206 35746 8258 35758
rect 28926 35746 28978 35758
rect 29822 35810 29874 35822
rect 29822 35746 29874 35758
rect 31838 35810 31890 35822
rect 31838 35746 31890 35758
rect 34190 35810 34242 35822
rect 34190 35746 34242 35758
rect 35422 35810 35474 35822
rect 35422 35746 35474 35758
rect 36318 35810 36370 35822
rect 36318 35746 36370 35758
rect 36542 35810 36594 35822
rect 36542 35746 36594 35758
rect 37326 35810 37378 35822
rect 37326 35746 37378 35758
rect 41246 35810 41298 35822
rect 41246 35746 41298 35758
rect 42478 35810 42530 35822
rect 42478 35746 42530 35758
rect 42590 35810 42642 35822
rect 45278 35810 45330 35822
rect 44930 35758 44942 35810
rect 44994 35758 45006 35810
rect 42590 35746 42642 35758
rect 45278 35746 45330 35758
rect 45390 35810 45442 35822
rect 45390 35746 45442 35758
rect 49310 35810 49362 35822
rect 49310 35746 49362 35758
rect 49646 35810 49698 35822
rect 49646 35746 49698 35758
rect 57822 35810 57874 35822
rect 57822 35746 57874 35758
rect 4398 35698 4450 35710
rect 2594 35646 2606 35698
rect 2658 35646 2670 35698
rect 3602 35646 3614 35698
rect 3666 35646 3678 35698
rect 4398 35634 4450 35646
rect 6414 35698 6466 35710
rect 6414 35634 6466 35646
rect 6638 35698 6690 35710
rect 14702 35698 14754 35710
rect 7298 35646 7310 35698
rect 7362 35646 7374 35698
rect 13234 35646 13246 35698
rect 13298 35646 13310 35698
rect 14130 35646 14142 35698
rect 14194 35646 14206 35698
rect 14466 35646 14478 35698
rect 14530 35646 14542 35698
rect 6638 35634 6690 35646
rect 14702 35634 14754 35646
rect 16270 35698 16322 35710
rect 16270 35634 16322 35646
rect 17390 35698 17442 35710
rect 20190 35698 20242 35710
rect 17938 35646 17950 35698
rect 18002 35646 18014 35698
rect 18610 35646 18622 35698
rect 18674 35646 18686 35698
rect 19506 35646 19518 35698
rect 19570 35646 19582 35698
rect 17390 35634 17442 35646
rect 20190 35634 20242 35646
rect 20526 35698 20578 35710
rect 20526 35634 20578 35646
rect 20862 35698 20914 35710
rect 23550 35698 23602 35710
rect 21746 35646 21758 35698
rect 21810 35646 21822 35698
rect 22082 35646 22094 35698
rect 22146 35646 22158 35698
rect 20862 35634 20914 35646
rect 23550 35634 23602 35646
rect 24446 35698 24498 35710
rect 24446 35634 24498 35646
rect 24782 35698 24834 35710
rect 28590 35698 28642 35710
rect 25330 35646 25342 35698
rect 25394 35646 25406 35698
rect 26114 35646 26126 35698
rect 26178 35646 26190 35698
rect 24782 35634 24834 35646
rect 28590 35634 28642 35646
rect 29262 35698 29314 35710
rect 29262 35634 29314 35646
rect 29710 35698 29762 35710
rect 29710 35634 29762 35646
rect 30046 35698 30098 35710
rect 31166 35698 31218 35710
rect 30482 35646 30494 35698
rect 30546 35646 30558 35698
rect 30046 35634 30098 35646
rect 31166 35634 31218 35646
rect 31614 35698 31666 35710
rect 31614 35634 31666 35646
rect 31950 35698 32002 35710
rect 31950 35634 32002 35646
rect 33630 35698 33682 35710
rect 33630 35634 33682 35646
rect 33966 35698 34018 35710
rect 36878 35698 36930 35710
rect 37438 35698 37490 35710
rect 35074 35646 35086 35698
rect 35138 35646 35150 35698
rect 37090 35646 37102 35698
rect 37154 35646 37166 35698
rect 33966 35634 34018 35646
rect 36878 35634 36930 35646
rect 37438 35634 37490 35646
rect 38110 35698 38162 35710
rect 38110 35634 38162 35646
rect 38446 35698 38498 35710
rect 38446 35634 38498 35646
rect 38782 35698 38834 35710
rect 38782 35634 38834 35646
rect 39230 35698 39282 35710
rect 45614 35698 45666 35710
rect 40114 35646 40126 35698
rect 40178 35646 40190 35698
rect 40898 35646 40910 35698
rect 40962 35646 40974 35698
rect 43250 35646 43262 35698
rect 43314 35646 43326 35698
rect 43922 35646 43934 35698
rect 43986 35646 43998 35698
rect 39230 35634 39282 35646
rect 45614 35634 45666 35646
rect 47406 35698 47458 35710
rect 47406 35634 47458 35646
rect 47630 35698 47682 35710
rect 47630 35634 47682 35646
rect 47854 35698 47906 35710
rect 47854 35634 47906 35646
rect 48638 35698 48690 35710
rect 48638 35634 48690 35646
rect 49982 35698 50034 35710
rect 49982 35634 50034 35646
rect 50654 35698 50706 35710
rect 50654 35634 50706 35646
rect 51214 35698 51266 35710
rect 51214 35634 51266 35646
rect 51550 35698 51602 35710
rect 57150 35698 57202 35710
rect 51986 35646 51998 35698
rect 52050 35646 52062 35698
rect 52210 35646 52222 35698
rect 52274 35646 52286 35698
rect 53666 35646 53678 35698
rect 53730 35646 53742 35698
rect 51550 35634 51602 35646
rect 57150 35634 57202 35646
rect 58158 35698 58210 35710
rect 58158 35634 58210 35646
rect 4174 35586 4226 35598
rect 14926 35586 14978 35598
rect 23998 35586 24050 35598
rect 32398 35586 32450 35598
rect 4946 35534 4958 35586
rect 5010 35534 5022 35586
rect 7410 35534 7422 35586
rect 7474 35534 7486 35586
rect 19282 35534 19294 35586
rect 19346 35534 19358 35586
rect 21970 35534 21982 35586
rect 22034 35534 22046 35586
rect 26002 35534 26014 35586
rect 26066 35534 26078 35586
rect 4174 35522 4226 35534
rect 14926 35522 14978 35534
rect 23998 35522 24050 35534
rect 32398 35522 32450 35534
rect 34414 35586 34466 35598
rect 34414 35522 34466 35534
rect 38334 35586 38386 35598
rect 41134 35586 41186 35598
rect 40002 35534 40014 35586
rect 40066 35534 40078 35586
rect 38334 35522 38386 35534
rect 41134 35522 41186 35534
rect 43150 35586 43202 35598
rect 43150 35522 43202 35534
rect 45950 35586 46002 35598
rect 45950 35522 46002 35534
rect 49198 35586 49250 35598
rect 57598 35586 57650 35598
rect 52658 35534 52670 35586
rect 52722 35534 52734 35586
rect 53442 35534 53454 35586
rect 53506 35534 53518 35586
rect 49198 35522 49250 35534
rect 57598 35522 57650 35534
rect 15038 35474 15090 35486
rect 15038 35410 15090 35422
rect 23438 35474 23490 35486
rect 23438 35410 23490 35422
rect 25566 35474 25618 35486
rect 34750 35474 34802 35486
rect 31266 35422 31278 35474
rect 31330 35422 31342 35474
rect 25566 35410 25618 35422
rect 34750 35410 34802 35422
rect 35086 35474 35138 35486
rect 35086 35410 35138 35422
rect 36654 35474 36706 35486
rect 48302 35474 48354 35486
rect 43474 35422 43486 35474
rect 43538 35422 43550 35474
rect 52322 35422 52334 35474
rect 52386 35422 52398 35474
rect 36654 35410 36706 35422
rect 48302 35410 48354 35422
rect 1344 35306 58576 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 58576 35306
rect 1344 35220 58576 35254
rect 3166 35138 3218 35150
rect 3166 35074 3218 35086
rect 9774 35138 9826 35150
rect 9774 35074 9826 35086
rect 33406 35138 33458 35150
rect 33406 35074 33458 35086
rect 53006 35138 53058 35150
rect 53006 35074 53058 35086
rect 9214 35026 9266 35038
rect 4498 34974 4510 35026
rect 4562 34974 4574 35026
rect 8418 34974 8430 35026
rect 8482 34974 8494 35026
rect 9214 34962 9266 34974
rect 11566 35026 11618 35038
rect 30382 35026 30434 35038
rect 17826 34974 17838 35026
rect 17890 34974 17902 35026
rect 22754 34974 22766 35026
rect 22818 34974 22830 35026
rect 25218 34974 25230 35026
rect 25282 34974 25294 35026
rect 11566 34962 11618 34974
rect 30382 34962 30434 34974
rect 33630 35026 33682 35038
rect 37102 35026 37154 35038
rect 34962 34974 34974 35026
rect 35026 34974 35038 35026
rect 33630 34962 33682 34974
rect 37102 34962 37154 34974
rect 39566 35026 39618 35038
rect 50990 35026 51042 35038
rect 40002 34974 40014 35026
rect 40066 34974 40078 35026
rect 47506 34974 47518 35026
rect 47570 34974 47582 35026
rect 53554 34974 53566 35026
rect 53618 34974 53630 35026
rect 39566 34962 39618 34974
rect 50990 34962 51042 34974
rect 5070 34914 5122 34926
rect 10670 34914 10722 34926
rect 14030 34914 14082 34926
rect 3042 34862 3054 34914
rect 3106 34862 3118 34914
rect 4162 34862 4174 34914
rect 4226 34862 4238 34914
rect 7074 34862 7086 34914
rect 7138 34862 7150 34914
rect 8754 34862 8766 34914
rect 8818 34862 8830 34914
rect 11106 34862 11118 34914
rect 11170 34862 11182 34914
rect 5070 34850 5122 34862
rect 10670 34850 10722 34862
rect 14030 34850 14082 34862
rect 14366 34914 14418 34926
rect 18846 34914 18898 34926
rect 17378 34862 17390 34914
rect 17442 34862 17454 34914
rect 17938 34862 17950 34914
rect 18002 34862 18014 34914
rect 14366 34850 14418 34862
rect 18846 34850 18898 34862
rect 19742 34914 19794 34926
rect 19742 34850 19794 34862
rect 22430 34914 22482 34926
rect 26014 34914 26066 34926
rect 23426 34862 23438 34914
rect 23490 34862 23502 34914
rect 23762 34862 23774 34914
rect 23826 34862 23838 34914
rect 24322 34862 24334 34914
rect 24386 34862 24398 34914
rect 25330 34862 25342 34914
rect 25394 34862 25406 34914
rect 22430 34850 22482 34862
rect 26014 34850 26066 34862
rect 26350 34914 26402 34926
rect 26350 34850 26402 34862
rect 26686 34914 26738 34926
rect 26686 34850 26738 34862
rect 26910 34914 26962 34926
rect 29374 34914 29426 34926
rect 29138 34862 29150 34914
rect 29202 34862 29214 34914
rect 26910 34850 26962 34862
rect 29374 34850 29426 34862
rect 29710 34914 29762 34926
rect 29710 34850 29762 34862
rect 31278 34914 31330 34926
rect 31278 34850 31330 34862
rect 31502 34914 31554 34926
rect 31502 34850 31554 34862
rect 31838 34914 31890 34926
rect 31838 34850 31890 34862
rect 32398 34914 32450 34926
rect 36094 34914 36146 34926
rect 37998 34914 38050 34926
rect 41358 34914 41410 34926
rect 32722 34862 32734 34914
rect 32786 34862 32798 34914
rect 33170 34862 33182 34914
rect 33234 34862 33246 34914
rect 34402 34862 34414 34914
rect 34466 34862 34478 34914
rect 35298 34862 35310 34914
rect 35362 34862 35374 34914
rect 37650 34862 37662 34914
rect 37714 34862 37726 34914
rect 40114 34862 40126 34914
rect 40178 34862 40190 34914
rect 32398 34850 32450 34862
rect 36094 34850 36146 34862
rect 37998 34850 38050 34862
rect 41358 34850 41410 34862
rect 43262 34914 43314 34926
rect 43262 34850 43314 34862
rect 43598 34914 43650 34926
rect 45266 34862 45278 34914
rect 45330 34862 45342 34914
rect 48962 34862 48974 34914
rect 49026 34862 49038 34914
rect 55010 34862 55022 34914
rect 55074 34862 55086 34914
rect 43598 34850 43650 34862
rect 2830 34802 2882 34814
rect 2830 34738 2882 34750
rect 3278 34802 3330 34814
rect 3278 34738 3330 34750
rect 6190 34802 6242 34814
rect 9886 34802 9938 34814
rect 19518 34802 19570 34814
rect 6850 34750 6862 34802
rect 6914 34750 6926 34802
rect 18274 34750 18286 34802
rect 18338 34750 18350 34802
rect 6190 34738 6242 34750
rect 9886 34738 9938 34750
rect 19518 34738 19570 34750
rect 20078 34802 20130 34814
rect 20078 34738 20130 34750
rect 22654 34802 22706 34814
rect 32286 34802 32338 34814
rect 23874 34750 23886 34802
rect 23938 34750 23950 34802
rect 22654 34738 22706 34750
rect 32286 34738 32338 34750
rect 33742 34802 33794 34814
rect 35982 34802 36034 34814
rect 34514 34750 34526 34802
rect 34578 34750 34590 34802
rect 33742 34738 33794 34750
rect 35982 34738 36034 34750
rect 37438 34802 37490 34814
rect 53006 34802 53058 34814
rect 47730 34750 47742 34802
rect 47794 34750 47806 34802
rect 50306 34750 50318 34802
rect 50370 34750 50382 34802
rect 37438 34738 37490 34750
rect 53006 34738 53058 34750
rect 53118 34802 53170 34814
rect 58158 34802 58210 34814
rect 53778 34750 53790 34802
rect 53842 34750 53854 34802
rect 53118 34738 53170 34750
rect 58158 34738 58210 34750
rect 6526 34690 6578 34702
rect 6526 34626 6578 34638
rect 9774 34690 9826 34702
rect 9774 34626 9826 34638
rect 14254 34690 14306 34702
rect 14254 34626 14306 34638
rect 18958 34690 19010 34702
rect 18958 34626 19010 34638
rect 19182 34690 19234 34702
rect 19182 34626 19234 34638
rect 19630 34690 19682 34702
rect 19630 34626 19682 34638
rect 22094 34690 22146 34702
rect 22094 34626 22146 34638
rect 26574 34690 26626 34702
rect 26574 34626 26626 34638
rect 29486 34690 29538 34702
rect 29486 34626 29538 34638
rect 29598 34690 29650 34702
rect 29598 34626 29650 34638
rect 31502 34690 31554 34702
rect 31502 34626 31554 34638
rect 32174 34690 32226 34702
rect 32174 34626 32226 34638
rect 35758 34690 35810 34702
rect 35758 34626 35810 34638
rect 37326 34690 37378 34702
rect 37326 34626 37378 34638
rect 38334 34690 38386 34702
rect 38334 34626 38386 34638
rect 41134 34690 41186 34702
rect 41134 34626 41186 34638
rect 41246 34690 41298 34702
rect 41246 34626 41298 34638
rect 41582 34690 41634 34702
rect 41582 34626 41634 34638
rect 43374 34690 43426 34702
rect 57598 34690 57650 34702
rect 45042 34638 45054 34690
rect 45106 34638 45118 34690
rect 55346 34638 55358 34690
rect 55410 34638 55422 34690
rect 43374 34626 43426 34638
rect 57598 34626 57650 34638
rect 57822 34690 57874 34702
rect 57822 34626 57874 34638
rect 1344 34522 58576 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 50558 34522
rect 50610 34470 50662 34522
rect 50714 34470 50766 34522
rect 50818 34470 58576 34522
rect 1344 34436 58576 34470
rect 2046 34354 2098 34366
rect 2046 34290 2098 34302
rect 6862 34354 6914 34366
rect 9774 34354 9826 34366
rect 21646 34354 21698 34366
rect 7186 34302 7198 34354
rect 7250 34302 7262 34354
rect 8082 34302 8094 34354
rect 8146 34302 8158 34354
rect 11218 34302 11230 34354
rect 11282 34302 11294 34354
rect 6862 34290 6914 34302
rect 9774 34290 9826 34302
rect 21646 34290 21698 34302
rect 22990 34354 23042 34366
rect 22990 34290 23042 34302
rect 25454 34354 25506 34366
rect 25454 34290 25506 34302
rect 27918 34354 27970 34366
rect 27918 34290 27970 34302
rect 29598 34354 29650 34366
rect 29598 34290 29650 34302
rect 31502 34354 31554 34366
rect 34862 34354 34914 34366
rect 34290 34302 34302 34354
rect 34354 34302 34366 34354
rect 31502 34290 31554 34302
rect 34862 34290 34914 34302
rect 35982 34354 36034 34366
rect 35982 34290 36034 34302
rect 38782 34354 38834 34366
rect 38782 34290 38834 34302
rect 42254 34354 42306 34366
rect 42254 34290 42306 34302
rect 43262 34354 43314 34366
rect 43262 34290 43314 34302
rect 47742 34354 47794 34366
rect 50754 34302 50766 34354
rect 50818 34302 50830 34354
rect 47742 34290 47794 34302
rect 8542 34242 8594 34254
rect 4162 34190 4174 34242
rect 4226 34190 4238 34242
rect 8542 34178 8594 34190
rect 8654 34242 8706 34254
rect 8654 34178 8706 34190
rect 9886 34242 9938 34254
rect 11678 34242 11730 34254
rect 10658 34190 10670 34242
rect 10722 34190 10734 34242
rect 9886 34178 9938 34190
rect 11678 34178 11730 34190
rect 11790 34242 11842 34254
rect 11790 34178 11842 34190
rect 16606 34242 16658 34254
rect 16606 34178 16658 34190
rect 18398 34242 18450 34254
rect 21534 34242 21586 34254
rect 19170 34190 19182 34242
rect 19234 34190 19246 34242
rect 18398 34178 18450 34190
rect 21534 34178 21586 34190
rect 22318 34242 22370 34254
rect 22318 34178 22370 34190
rect 22430 34242 22482 34254
rect 22430 34178 22482 34190
rect 26126 34242 26178 34254
rect 26126 34178 26178 34190
rect 27694 34242 27746 34254
rect 27694 34178 27746 34190
rect 28814 34242 28866 34254
rect 28814 34178 28866 34190
rect 28926 34242 28978 34254
rect 28926 34178 28978 34190
rect 29486 34242 29538 34254
rect 29486 34178 29538 34190
rect 31054 34242 31106 34254
rect 31054 34178 31106 34190
rect 33742 34242 33794 34254
rect 33742 34178 33794 34190
rect 36206 34242 36258 34254
rect 36206 34178 36258 34190
rect 36318 34242 36370 34254
rect 36318 34178 36370 34190
rect 37326 34242 37378 34254
rect 37326 34178 37378 34190
rect 39006 34242 39058 34254
rect 39006 34178 39058 34190
rect 40014 34242 40066 34254
rect 40014 34178 40066 34190
rect 42590 34242 42642 34254
rect 42590 34178 42642 34190
rect 45166 34242 45218 34254
rect 45166 34178 45218 34190
rect 45502 34242 45554 34254
rect 45502 34178 45554 34190
rect 45726 34242 45778 34254
rect 45726 34178 45778 34190
rect 45838 34242 45890 34254
rect 45838 34178 45890 34190
rect 47518 34242 47570 34254
rect 47518 34178 47570 34190
rect 47966 34242 48018 34254
rect 47966 34178 48018 34190
rect 48078 34242 48130 34254
rect 48078 34178 48130 34190
rect 48974 34242 49026 34254
rect 53342 34242 53394 34254
rect 49186 34190 49198 34242
rect 49250 34190 49262 34242
rect 51762 34190 51774 34242
rect 51826 34190 51838 34242
rect 48974 34178 49026 34190
rect 53342 34178 53394 34190
rect 57822 34242 57874 34254
rect 57822 34178 57874 34190
rect 1710 34130 1762 34142
rect 8766 34130 8818 34142
rect 4386 34078 4398 34130
rect 4450 34078 4462 34130
rect 5058 34078 5070 34130
rect 5122 34078 5134 34130
rect 5842 34078 5854 34130
rect 5906 34078 5918 34130
rect 1710 34066 1762 34078
rect 8766 34066 8818 34078
rect 9550 34130 9602 34142
rect 12014 34130 12066 34142
rect 13582 34130 13634 34142
rect 10546 34078 10558 34130
rect 10610 34078 10622 34130
rect 11106 34078 11118 34130
rect 11170 34078 11182 34130
rect 12674 34078 12686 34130
rect 12738 34078 12750 34130
rect 13122 34078 13134 34130
rect 13186 34078 13198 34130
rect 9550 34066 9602 34078
rect 12014 34066 12066 34078
rect 13582 34066 13634 34078
rect 13918 34130 13970 34142
rect 14702 34130 14754 34142
rect 14354 34078 14366 34130
rect 14418 34078 14430 34130
rect 13918 34066 13970 34078
rect 14702 34066 14754 34078
rect 16718 34130 16770 34142
rect 21422 34130 21474 34142
rect 17938 34078 17950 34130
rect 18002 34078 18014 34130
rect 20290 34078 20302 34130
rect 20354 34078 20366 34130
rect 16718 34066 16770 34078
rect 21422 34066 21474 34078
rect 21982 34130 22034 34142
rect 21982 34066 22034 34078
rect 23438 34130 23490 34142
rect 24334 34130 24386 34142
rect 23650 34078 23662 34130
rect 23714 34078 23726 34130
rect 23438 34066 23490 34078
rect 24334 34066 24386 34078
rect 25230 34130 25282 34142
rect 25230 34066 25282 34078
rect 25902 34130 25954 34142
rect 25902 34066 25954 34078
rect 26350 34130 26402 34142
rect 29150 34130 29202 34142
rect 27458 34078 27470 34130
rect 27522 34078 27534 34130
rect 28578 34078 28590 34130
rect 28642 34078 28654 34130
rect 26350 34066 26402 34078
rect 29150 34066 29202 34078
rect 29822 34130 29874 34142
rect 29822 34066 29874 34078
rect 30382 34130 30434 34142
rect 30382 34066 30434 34078
rect 30830 34130 30882 34142
rect 30830 34066 30882 34078
rect 31390 34130 31442 34142
rect 31390 34066 31442 34078
rect 31614 34130 31666 34142
rect 31614 34066 31666 34078
rect 32062 34130 32114 34142
rect 32062 34066 32114 34078
rect 33966 34130 34018 34142
rect 33966 34066 34018 34078
rect 34638 34130 34690 34142
rect 34638 34066 34690 34078
rect 36542 34130 36594 34142
rect 36542 34066 36594 34078
rect 36878 34130 36930 34142
rect 36878 34066 36930 34078
rect 37102 34130 37154 34142
rect 37102 34066 37154 34078
rect 37886 34130 37938 34142
rect 37886 34066 37938 34078
rect 38446 34130 38498 34142
rect 40910 34130 40962 34142
rect 40338 34078 40350 34130
rect 40402 34078 40414 34130
rect 38446 34066 38498 34078
rect 40910 34066 40962 34078
rect 41134 34130 41186 34142
rect 41134 34066 41186 34078
rect 41358 34130 41410 34142
rect 41358 34066 41410 34078
rect 41806 34130 41858 34142
rect 41806 34066 41858 34078
rect 42030 34130 42082 34142
rect 42030 34066 42082 34078
rect 42254 34130 42306 34142
rect 42254 34066 42306 34078
rect 43038 34130 43090 34142
rect 43038 34066 43090 34078
rect 43150 34130 43202 34142
rect 45054 34130 45106 34142
rect 43586 34078 43598 34130
rect 43650 34078 43662 34130
rect 43150 34066 43202 34078
rect 45054 34066 45106 34078
rect 48750 34130 48802 34142
rect 49758 34130 49810 34142
rect 54238 34130 54290 34142
rect 49298 34078 49310 34130
rect 49362 34078 49374 34130
rect 50642 34078 50654 34130
rect 50706 34078 50718 34130
rect 51650 34078 51662 34130
rect 51714 34078 51726 34130
rect 53778 34078 53790 34130
rect 53842 34078 53854 34130
rect 48750 34066 48802 34078
rect 49758 34066 49810 34078
rect 54238 34066 54290 34078
rect 55694 34130 55746 34142
rect 55694 34066 55746 34078
rect 58158 34130 58210 34142
rect 58158 34066 58210 34078
rect 2494 34018 2546 34030
rect 6302 34018 6354 34030
rect 4498 33966 4510 34018
rect 4562 33966 4574 34018
rect 2494 33954 2546 33966
rect 6302 33954 6354 33966
rect 14926 34018 14978 34030
rect 20974 34018 21026 34030
rect 17490 33966 17502 34018
rect 17554 33966 17566 34018
rect 18834 33966 18846 34018
rect 18898 33966 18910 34018
rect 14926 33954 14978 33966
rect 20974 33954 21026 33966
rect 25342 34018 25394 34030
rect 25342 33954 25394 33966
rect 30606 34018 30658 34030
rect 30606 33954 30658 33966
rect 34750 34018 34802 34030
rect 34750 33954 34802 33966
rect 37214 34018 37266 34030
rect 37214 33954 37266 33966
rect 37662 34018 37714 34030
rect 37662 33954 37714 33966
rect 40126 34018 40178 34030
rect 40126 33954 40178 33966
rect 57598 34018 57650 34030
rect 57598 33954 57650 33966
rect 16606 33906 16658 33918
rect 16606 33842 16658 33854
rect 22318 33906 22370 33918
rect 22318 33842 22370 33854
rect 26686 33906 26738 33918
rect 26686 33842 26738 33854
rect 28030 33906 28082 33918
rect 28030 33842 28082 33854
rect 28142 33906 28194 33918
rect 38670 33906 38722 33918
rect 38210 33854 38222 33906
rect 38274 33854 38286 33906
rect 28142 33842 28194 33854
rect 38670 33842 38722 33854
rect 45166 33906 45218 33918
rect 45166 33842 45218 33854
rect 47406 33906 47458 33918
rect 47406 33842 47458 33854
rect 54798 33906 54850 33918
rect 54798 33842 54850 33854
rect 55246 33906 55298 33918
rect 55246 33842 55298 33854
rect 55470 33906 55522 33918
rect 55470 33842 55522 33854
rect 1344 33738 58576 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 58576 33738
rect 1344 33652 58576 33686
rect 27806 33570 27858 33582
rect 4050 33518 4062 33570
rect 4114 33518 4126 33570
rect 15698 33518 15710 33570
rect 15762 33518 15774 33570
rect 17378 33518 17390 33570
rect 17442 33518 17454 33570
rect 27806 33506 27858 33518
rect 28254 33570 28306 33582
rect 28254 33506 28306 33518
rect 28478 33570 28530 33582
rect 28478 33506 28530 33518
rect 39566 33570 39618 33582
rect 44158 33570 44210 33582
rect 41122 33518 41134 33570
rect 41186 33518 41198 33570
rect 39566 33506 39618 33518
rect 44158 33506 44210 33518
rect 31838 33458 31890 33470
rect 39678 33458 39730 33470
rect 45838 33458 45890 33470
rect 5954 33406 5966 33458
rect 6018 33406 6030 33458
rect 13570 33406 13582 33458
rect 13634 33406 13646 33458
rect 16482 33406 16494 33458
rect 16546 33406 16558 33458
rect 17826 33406 17838 33458
rect 17890 33406 17902 33458
rect 37090 33406 37102 33458
rect 37154 33406 37166 33458
rect 42802 33406 42814 33458
rect 42866 33406 42878 33458
rect 45378 33406 45390 33458
rect 45442 33406 45454 33458
rect 31838 33394 31890 33406
rect 39678 33394 39730 33406
rect 45838 33394 45890 33406
rect 48750 33458 48802 33470
rect 48750 33394 48802 33406
rect 50318 33458 50370 33470
rect 50318 33394 50370 33406
rect 53342 33458 53394 33470
rect 53342 33394 53394 33406
rect 2718 33346 2770 33358
rect 7982 33346 8034 33358
rect 2370 33294 2382 33346
rect 2434 33294 2446 33346
rect 3714 33294 3726 33346
rect 3778 33294 3790 33346
rect 6402 33294 6414 33346
rect 6466 33294 6478 33346
rect 6962 33294 6974 33346
rect 7026 33294 7038 33346
rect 2718 33282 2770 33294
rect 7982 33282 8034 33294
rect 8990 33346 9042 33358
rect 11006 33346 11058 33358
rect 18846 33346 18898 33358
rect 10546 33294 10558 33346
rect 10610 33294 10622 33346
rect 14018 33294 14030 33346
rect 14082 33294 14094 33346
rect 15026 33294 15038 33346
rect 15090 33294 15102 33346
rect 16818 33294 16830 33346
rect 16882 33294 16894 33346
rect 17266 33294 17278 33346
rect 17330 33294 17342 33346
rect 17938 33294 17950 33346
rect 18002 33294 18014 33346
rect 8990 33282 9042 33294
rect 11006 33282 11058 33294
rect 18846 33282 18898 33294
rect 19182 33346 19234 33358
rect 19182 33282 19234 33294
rect 19406 33346 19458 33358
rect 22542 33346 22594 33358
rect 22306 33294 22318 33346
rect 22370 33294 22382 33346
rect 19406 33282 19458 33294
rect 22542 33282 22594 33294
rect 24894 33346 24946 33358
rect 24894 33282 24946 33294
rect 25454 33346 25506 33358
rect 25454 33282 25506 33294
rect 32062 33346 32114 33358
rect 32062 33282 32114 33294
rect 34302 33346 34354 33358
rect 34302 33282 34354 33294
rect 34638 33346 34690 33358
rect 34638 33282 34690 33294
rect 34974 33346 35026 33358
rect 34974 33282 35026 33294
rect 35086 33346 35138 33358
rect 35086 33282 35138 33294
rect 35534 33346 35586 33358
rect 35534 33282 35586 33294
rect 35646 33346 35698 33358
rect 35646 33282 35698 33294
rect 35758 33346 35810 33358
rect 47182 33346 47234 33358
rect 38658 33294 38670 33346
rect 38722 33294 38734 33346
rect 41010 33294 41022 33346
rect 41074 33294 41086 33346
rect 42578 33294 42590 33346
rect 42642 33294 42654 33346
rect 45266 33294 45278 33346
rect 45330 33294 45342 33346
rect 35758 33282 35810 33294
rect 47182 33282 47234 33294
rect 47406 33346 47458 33358
rect 47406 33282 47458 33294
rect 47742 33346 47794 33358
rect 49982 33346 50034 33358
rect 51998 33346 52050 33358
rect 48178 33294 48190 33346
rect 48242 33294 48254 33346
rect 48962 33294 48974 33346
rect 49026 33294 49038 33346
rect 50642 33294 50654 33346
rect 50706 33294 50718 33346
rect 51762 33294 51774 33346
rect 51826 33294 51838 33346
rect 47742 33282 47794 33294
rect 49982 33282 50034 33294
rect 51998 33282 52050 33294
rect 55246 33346 55298 33358
rect 55246 33282 55298 33294
rect 55470 33346 55522 33358
rect 55470 33282 55522 33294
rect 22766 33234 22818 33246
rect 5954 33182 5966 33234
rect 6018 33182 6030 33234
rect 8642 33182 8654 33234
rect 8706 33182 8718 33234
rect 22766 33170 22818 33182
rect 25342 33234 25394 33246
rect 25342 33170 25394 33182
rect 27694 33234 27746 33246
rect 27694 33170 27746 33182
rect 27918 33234 27970 33246
rect 27918 33170 27970 33182
rect 32846 33234 32898 33246
rect 32846 33170 32898 33182
rect 32958 33234 33010 33246
rect 44158 33234 44210 33246
rect 37314 33182 37326 33234
rect 37378 33182 37390 33234
rect 32958 33170 33010 33182
rect 44158 33170 44210 33182
rect 44270 33234 44322 33246
rect 49870 33234 49922 33246
rect 51102 33234 51154 33246
rect 48402 33182 48414 33234
rect 48466 33182 48478 33234
rect 50082 33182 50094 33234
rect 50146 33182 50158 33234
rect 44270 33170 44322 33182
rect 49870 33170 49922 33182
rect 51102 33170 51154 33182
rect 52670 33234 52722 33246
rect 52670 33170 52722 33182
rect 52782 33234 52834 33246
rect 52782 33170 52834 33182
rect 55022 33234 55074 33246
rect 55022 33170 55074 33182
rect 58158 33234 58210 33246
rect 58158 33170 58210 33182
rect 7310 33122 7362 33134
rect 7310 33058 7362 33070
rect 7422 33122 7474 33134
rect 7422 33058 7474 33070
rect 7534 33122 7586 33134
rect 7534 33058 7586 33070
rect 9662 33122 9714 33134
rect 19070 33122 19122 33134
rect 9986 33070 9998 33122
rect 10050 33070 10062 33122
rect 9662 33058 9714 33070
rect 19070 33058 19122 33070
rect 25118 33122 25170 33134
rect 25118 33058 25170 33070
rect 29374 33122 29426 33134
rect 29374 33058 29426 33070
rect 30382 33122 30434 33134
rect 32622 33122 32674 33134
rect 32386 33070 32398 33122
rect 32450 33070 32462 33122
rect 30382 33058 30434 33070
rect 32622 33058 32674 33070
rect 34750 33122 34802 33134
rect 47518 33122 47570 33134
rect 53006 33122 53058 33134
rect 38994 33070 39006 33122
rect 39058 33070 39070 33122
rect 48514 33070 48526 33122
rect 48578 33070 48590 33122
rect 34750 33058 34802 33070
rect 47518 33058 47570 33070
rect 53006 33058 53058 33070
rect 55358 33122 55410 33134
rect 55358 33058 55410 33070
rect 57598 33122 57650 33134
rect 57598 33058 57650 33070
rect 57822 33122 57874 33134
rect 57822 33058 57874 33070
rect 1344 32954 58576 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 50558 32954
rect 50610 32902 50662 32954
rect 50714 32902 50766 32954
rect 50818 32902 58576 32954
rect 1344 32868 58576 32902
rect 7982 32786 8034 32798
rect 3602 32734 3614 32786
rect 3666 32734 3678 32786
rect 6178 32734 6190 32786
rect 6242 32734 6254 32786
rect 7982 32722 8034 32734
rect 9662 32786 9714 32798
rect 9662 32722 9714 32734
rect 18398 32786 18450 32798
rect 37550 32786 37602 32798
rect 31042 32734 31054 32786
rect 31106 32734 31118 32786
rect 18398 32722 18450 32734
rect 37550 32722 37602 32734
rect 39678 32786 39730 32798
rect 39678 32722 39730 32734
rect 46286 32786 46338 32798
rect 46286 32722 46338 32734
rect 46734 32786 46786 32798
rect 46734 32722 46786 32734
rect 49422 32786 49474 32798
rect 49422 32722 49474 32734
rect 7758 32674 7810 32686
rect 2370 32622 2382 32674
rect 2434 32622 2446 32674
rect 3714 32622 3726 32674
rect 3778 32622 3790 32674
rect 6066 32622 6078 32674
rect 6130 32622 6142 32674
rect 7758 32610 7810 32622
rect 10334 32674 10386 32686
rect 10334 32610 10386 32622
rect 10670 32674 10722 32686
rect 10670 32610 10722 32622
rect 11118 32674 11170 32686
rect 15262 32674 15314 32686
rect 17390 32674 17442 32686
rect 13682 32622 13694 32674
rect 13746 32622 13758 32674
rect 14914 32622 14926 32674
rect 14978 32622 14990 32674
rect 16370 32622 16382 32674
rect 16434 32622 16446 32674
rect 11118 32610 11170 32622
rect 15262 32610 15314 32622
rect 17390 32610 17442 32622
rect 18286 32674 18338 32686
rect 18286 32610 18338 32622
rect 20078 32674 20130 32686
rect 20078 32610 20130 32622
rect 23214 32674 23266 32686
rect 28366 32674 28418 32686
rect 26114 32622 26126 32674
rect 26178 32622 26190 32674
rect 26898 32622 26910 32674
rect 26962 32622 26974 32674
rect 23214 32610 23266 32622
rect 28366 32610 28418 32622
rect 32062 32674 32114 32686
rect 32062 32610 32114 32622
rect 42702 32674 42754 32686
rect 42702 32610 42754 32622
rect 43262 32674 43314 32686
rect 43262 32610 43314 32622
rect 48862 32674 48914 32686
rect 48862 32610 48914 32622
rect 49534 32674 49586 32686
rect 49534 32610 49586 32622
rect 57822 32674 57874 32686
rect 57822 32610 57874 32622
rect 6750 32562 6802 32574
rect 2594 32510 2606 32562
rect 2658 32510 2670 32562
rect 6290 32510 6302 32562
rect 6354 32510 6366 32562
rect 6750 32498 6802 32510
rect 7086 32562 7138 32574
rect 7086 32498 7138 32510
rect 7422 32562 7474 32574
rect 7422 32498 7474 32510
rect 9774 32562 9826 32574
rect 9774 32498 9826 32510
rect 11230 32562 11282 32574
rect 17726 32562 17778 32574
rect 15698 32510 15710 32562
rect 15762 32510 15774 32562
rect 16258 32510 16270 32562
rect 16322 32510 16334 32562
rect 11230 32498 11282 32510
rect 17726 32498 17778 32510
rect 17838 32562 17890 32574
rect 17838 32498 17890 32510
rect 19966 32562 20018 32574
rect 19966 32498 20018 32510
rect 20302 32562 20354 32574
rect 30046 32562 30098 32574
rect 22306 32510 22318 32562
rect 22370 32510 22382 32562
rect 22530 32510 22542 32562
rect 22594 32510 22606 32562
rect 24210 32510 24222 32562
rect 24274 32510 24286 32562
rect 26226 32510 26238 32562
rect 26290 32510 26302 32562
rect 26674 32510 26686 32562
rect 26738 32510 26750 32562
rect 27570 32510 27582 32562
rect 27634 32510 27646 32562
rect 28578 32510 28590 32562
rect 28642 32510 28654 32562
rect 29810 32510 29822 32562
rect 29874 32510 29886 32562
rect 20302 32498 20354 32510
rect 30046 32498 30098 32510
rect 30718 32562 30770 32574
rect 32622 32562 32674 32574
rect 37662 32562 37714 32574
rect 32274 32510 32286 32562
rect 32338 32510 32350 32562
rect 33618 32510 33630 32562
rect 33682 32510 33694 32562
rect 30718 32498 30770 32510
rect 32622 32498 32674 32510
rect 37662 32498 37714 32510
rect 37774 32562 37826 32574
rect 37774 32498 37826 32510
rect 38222 32562 38274 32574
rect 42366 32562 42418 32574
rect 38882 32510 38894 32562
rect 38946 32510 38958 32562
rect 41458 32510 41470 32562
rect 41522 32510 41534 32562
rect 38222 32498 38274 32510
rect 42366 32498 42418 32510
rect 42926 32562 42978 32574
rect 42926 32498 42978 32510
rect 43150 32562 43202 32574
rect 46398 32562 46450 32574
rect 45378 32510 45390 32562
rect 45442 32510 45454 32562
rect 45826 32510 45838 32562
rect 45890 32510 45902 32562
rect 43150 32498 43202 32510
rect 46398 32498 46450 32510
rect 46510 32562 46562 32574
rect 46510 32498 46562 32510
rect 48750 32562 48802 32574
rect 48750 32498 48802 32510
rect 50766 32562 50818 32574
rect 50766 32498 50818 32510
rect 50990 32562 51042 32574
rect 58158 32562 58210 32574
rect 51874 32510 51886 32562
rect 51938 32510 51950 32562
rect 52882 32510 52894 32562
rect 52946 32510 52958 32562
rect 50990 32498 51042 32510
rect 58158 32498 58210 32510
rect 6974 32450 7026 32462
rect 6974 32386 7026 32398
rect 7870 32450 7922 32462
rect 18062 32450 18114 32462
rect 13122 32398 13134 32450
rect 13186 32398 13198 32450
rect 16706 32398 16718 32450
rect 16770 32398 16782 32450
rect 7870 32386 7922 32398
rect 18062 32386 18114 32398
rect 22766 32450 22818 32462
rect 22766 32386 22818 32398
rect 23326 32450 23378 32462
rect 24670 32450 24722 32462
rect 31726 32450 31778 32462
rect 34078 32450 34130 32462
rect 43710 32450 43762 32462
rect 57150 32450 57202 32462
rect 23762 32398 23774 32450
rect 23826 32398 23838 32450
rect 26338 32398 26350 32450
rect 26402 32398 26414 32450
rect 28690 32398 28702 32450
rect 28754 32398 28766 32450
rect 32050 32398 32062 32450
rect 32114 32398 32126 32450
rect 33170 32398 33182 32450
rect 33234 32398 33246 32450
rect 38994 32398 39006 32450
rect 39058 32398 39070 32450
rect 41570 32398 41582 32450
rect 41634 32398 41646 32450
rect 44370 32398 44382 32450
rect 44434 32398 44446 32450
rect 51762 32398 51774 32450
rect 51826 32398 51838 32450
rect 23326 32386 23378 32398
rect 24670 32386 24722 32398
rect 31726 32386 31778 32398
rect 34078 32386 34130 32398
rect 43710 32386 43762 32398
rect 57150 32386 57202 32398
rect 57598 32450 57650 32462
rect 57598 32386 57650 32398
rect 9662 32338 9714 32350
rect 9662 32274 9714 32286
rect 11118 32338 11170 32350
rect 48862 32338 48914 32350
rect 38546 32286 38558 32338
rect 38610 32286 38622 32338
rect 11118 32274 11170 32286
rect 48862 32274 48914 32286
rect 49422 32338 49474 32350
rect 50418 32286 50430 32338
rect 50482 32286 50494 32338
rect 53554 32286 53566 32338
rect 53618 32286 53630 32338
rect 49422 32274 49474 32286
rect 1344 32170 58576 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 58576 32170
rect 1344 32084 58576 32118
rect 39790 32002 39842 32014
rect 25106 31950 25118 32002
rect 25170 31950 25182 32002
rect 48738 31950 48750 32002
rect 48802 31950 48814 32002
rect 39790 31938 39842 31950
rect 4174 31890 4226 31902
rect 7198 31890 7250 31902
rect 26126 31890 26178 31902
rect 34526 31890 34578 31902
rect 40350 31890 40402 31902
rect 46846 31890 46898 31902
rect 6626 31838 6638 31890
rect 6690 31838 6702 31890
rect 11330 31838 11342 31890
rect 11394 31838 11406 31890
rect 17378 31838 17390 31890
rect 17442 31838 17454 31890
rect 19618 31838 19630 31890
rect 19682 31838 19694 31890
rect 33170 31838 33182 31890
rect 33234 31838 33246 31890
rect 34850 31838 34862 31890
rect 34914 31838 34926 31890
rect 36082 31838 36094 31890
rect 36146 31838 36158 31890
rect 36978 31838 36990 31890
rect 37042 31838 37054 31890
rect 39218 31838 39230 31890
rect 39282 31838 39294 31890
rect 42354 31838 42366 31890
rect 42418 31838 42430 31890
rect 49298 31838 49310 31890
rect 49362 31838 49374 31890
rect 4174 31826 4226 31838
rect 7198 31826 7250 31838
rect 26126 31826 26178 31838
rect 34526 31826 34578 31838
rect 40350 31826 40402 31838
rect 46846 31826 46898 31838
rect 3614 31778 3666 31790
rect 3266 31726 3278 31778
rect 3330 31726 3342 31778
rect 3614 31714 3666 31726
rect 3726 31778 3778 31790
rect 3726 31714 3778 31726
rect 3950 31778 4002 31790
rect 3950 31714 4002 31726
rect 5070 31778 5122 31790
rect 5070 31714 5122 31726
rect 6078 31778 6130 31790
rect 6078 31714 6130 31726
rect 6974 31778 7026 31790
rect 11790 31778 11842 31790
rect 11106 31726 11118 31778
rect 11170 31726 11182 31778
rect 6974 31714 7026 31726
rect 11790 31714 11842 31726
rect 12126 31778 12178 31790
rect 12126 31714 12178 31726
rect 12574 31778 12626 31790
rect 18174 31778 18226 31790
rect 16706 31726 16718 31778
rect 16770 31726 16782 31778
rect 17714 31726 17726 31778
rect 17778 31726 17790 31778
rect 12574 31714 12626 31726
rect 18174 31714 18226 31726
rect 18510 31778 18562 31790
rect 18510 31714 18562 31726
rect 18846 31778 18898 31790
rect 18846 31714 18898 31726
rect 19966 31778 20018 31790
rect 19966 31714 20018 31726
rect 20190 31778 20242 31790
rect 20190 31714 20242 31726
rect 24110 31778 24162 31790
rect 25342 31778 25394 31790
rect 24882 31726 24894 31778
rect 24946 31726 24958 31778
rect 24110 31714 24162 31726
rect 25342 31714 25394 31726
rect 25678 31778 25730 31790
rect 25678 31714 25730 31726
rect 26574 31778 26626 31790
rect 26574 31714 26626 31726
rect 27806 31778 27858 31790
rect 30942 31778 30994 31790
rect 31838 31778 31890 31790
rect 45502 31778 45554 31790
rect 28242 31726 28254 31778
rect 28306 31726 28318 31778
rect 29362 31726 29374 31778
rect 29426 31726 29438 31778
rect 31378 31726 31390 31778
rect 31442 31726 31454 31778
rect 33506 31726 33518 31778
rect 33570 31726 33582 31778
rect 35186 31726 35198 31778
rect 35250 31726 35262 31778
rect 38098 31726 38110 31778
rect 38162 31726 38174 31778
rect 38546 31726 38558 31778
rect 38610 31726 38622 31778
rect 39442 31726 39454 31778
rect 39506 31726 39518 31778
rect 42466 31726 42478 31778
rect 42530 31726 42542 31778
rect 43698 31726 43710 31778
rect 43762 31726 43774 31778
rect 27806 31714 27858 31726
rect 30942 31714 30994 31726
rect 31838 31714 31890 31726
rect 45502 31714 45554 31726
rect 45838 31778 45890 31790
rect 48638 31778 48690 31790
rect 54574 31778 54626 31790
rect 47954 31726 47966 31778
rect 48018 31726 48030 31778
rect 49410 31726 49422 31778
rect 49474 31726 49486 31778
rect 50754 31726 50766 31778
rect 50818 31726 50830 31778
rect 45838 31714 45890 31726
rect 48638 31714 48690 31726
rect 54574 31714 54626 31726
rect 55134 31778 55186 31790
rect 55134 31714 55186 31726
rect 4510 31666 4562 31678
rect 4510 31602 4562 31614
rect 7870 31666 7922 31678
rect 7870 31602 7922 31614
rect 7982 31666 8034 31678
rect 7982 31602 8034 31614
rect 8654 31666 8706 31678
rect 8654 31602 8706 31614
rect 11566 31666 11618 31678
rect 11566 31602 11618 31614
rect 14142 31666 14194 31678
rect 14142 31602 14194 31614
rect 14926 31666 14978 31678
rect 14926 31602 14978 31614
rect 15038 31666 15090 31678
rect 15038 31602 15090 31614
rect 15486 31666 15538 31678
rect 15486 31602 15538 31614
rect 18622 31666 18674 31678
rect 18622 31602 18674 31614
rect 19294 31666 19346 31678
rect 19294 31602 19346 31614
rect 19518 31666 19570 31678
rect 19518 31602 19570 31614
rect 20414 31666 20466 31678
rect 20414 31602 20466 31614
rect 24446 31666 24498 31678
rect 24446 31602 24498 31614
rect 26014 31666 26066 31678
rect 26014 31602 26066 31614
rect 26350 31666 26402 31678
rect 36206 31666 36258 31678
rect 29138 31614 29150 31666
rect 29202 31614 29214 31666
rect 26350 31602 26402 31614
rect 36206 31602 36258 31614
rect 36430 31666 36482 31678
rect 36430 31602 36482 31614
rect 37102 31666 37154 31678
rect 37102 31602 37154 31614
rect 37326 31666 37378 31678
rect 37326 31602 37378 31614
rect 39678 31666 39730 31678
rect 39678 31602 39730 31614
rect 39790 31666 39842 31678
rect 44942 31666 44994 31678
rect 43362 31614 43374 31666
rect 43426 31614 43438 31666
rect 39790 31602 39842 31614
rect 44942 31602 44994 31614
rect 45166 31666 45218 31678
rect 45166 31602 45218 31614
rect 45950 31666 46002 31678
rect 45950 31602 46002 31614
rect 46286 31666 46338 31678
rect 46286 31602 46338 31614
rect 51550 31666 51602 31678
rect 51550 31602 51602 31614
rect 53342 31666 53394 31678
rect 53342 31602 53394 31614
rect 53678 31666 53730 31678
rect 53678 31602 53730 31614
rect 53902 31666 53954 31678
rect 56926 31666 56978 31678
rect 54226 31614 54238 31666
rect 54290 31614 54302 31666
rect 53902 31602 53954 31614
rect 56926 31602 56978 31614
rect 57486 31666 57538 31678
rect 57486 31602 57538 31614
rect 4286 31554 4338 31566
rect 4286 31490 4338 31502
rect 4734 31554 4786 31566
rect 4734 31490 4786 31502
rect 4958 31554 5010 31566
rect 4958 31490 5010 31502
rect 6190 31554 6242 31566
rect 6190 31490 6242 31502
rect 6414 31554 6466 31566
rect 6414 31490 6466 31502
rect 7646 31554 7698 31566
rect 7646 31490 7698 31502
rect 8318 31554 8370 31566
rect 8318 31490 8370 31502
rect 8542 31554 8594 31566
rect 8542 31490 8594 31502
rect 9550 31554 9602 31566
rect 12014 31554 12066 31566
rect 9874 31502 9886 31554
rect 9938 31502 9950 31554
rect 9550 31490 9602 31502
rect 12014 31490 12066 31502
rect 13918 31554 13970 31566
rect 13918 31490 13970 31502
rect 14030 31554 14082 31566
rect 14030 31490 14082 31502
rect 14366 31554 14418 31566
rect 14366 31490 14418 31502
rect 14702 31554 14754 31566
rect 14702 31490 14754 31502
rect 16494 31554 16546 31566
rect 16494 31490 16546 31502
rect 20078 31554 20130 31566
rect 20078 31490 20130 31502
rect 24222 31554 24274 31566
rect 30382 31554 30434 31566
rect 25442 31502 25454 31554
rect 25506 31502 25518 31554
rect 24222 31490 24274 31502
rect 30382 31490 30434 31502
rect 42590 31554 42642 31566
rect 44158 31554 44210 31566
rect 43138 31502 43150 31554
rect 43202 31502 43214 31554
rect 42590 31490 42642 31502
rect 44158 31490 44210 31502
rect 44830 31554 44882 31566
rect 44830 31490 44882 31502
rect 46062 31554 46114 31566
rect 46062 31490 46114 31502
rect 53454 31554 53506 31566
rect 53454 31490 53506 31502
rect 54798 31554 54850 31566
rect 54798 31490 54850 31502
rect 55022 31554 55074 31566
rect 55022 31490 55074 31502
rect 57150 31554 57202 31566
rect 58158 31554 58210 31566
rect 57810 31502 57822 31554
rect 57874 31502 57886 31554
rect 57150 31490 57202 31502
rect 58158 31490 58210 31502
rect 1344 31386 58576 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 50558 31386
rect 50610 31334 50662 31386
rect 50714 31334 50766 31386
rect 50818 31334 58576 31386
rect 1344 31300 58576 31334
rect 2718 31218 2770 31230
rect 2718 31154 2770 31166
rect 10894 31218 10946 31230
rect 15934 31218 15986 31230
rect 11218 31166 11230 31218
rect 11282 31166 11294 31218
rect 10894 31154 10946 31166
rect 15934 31154 15986 31166
rect 17614 31218 17666 31230
rect 17614 31154 17666 31166
rect 23214 31218 23266 31230
rect 27918 31218 27970 31230
rect 26226 31166 26238 31218
rect 26290 31166 26302 31218
rect 23214 31154 23266 31166
rect 27918 31154 27970 31166
rect 28926 31218 28978 31230
rect 28926 31154 28978 31166
rect 30046 31218 30098 31230
rect 30046 31154 30098 31166
rect 37214 31218 37266 31230
rect 39790 31218 39842 31230
rect 38098 31166 38110 31218
rect 38162 31166 38174 31218
rect 37214 31154 37266 31166
rect 39790 31154 39842 31166
rect 2830 31106 2882 31118
rect 7198 31106 7250 31118
rect 4610 31054 4622 31106
rect 4674 31054 4686 31106
rect 2830 31042 2882 31054
rect 7198 31042 7250 31054
rect 11678 31106 11730 31118
rect 11678 31042 11730 31054
rect 11790 31106 11842 31118
rect 11790 31042 11842 31054
rect 12350 31106 12402 31118
rect 12350 31042 12402 31054
rect 12462 31106 12514 31118
rect 12462 31042 12514 31054
rect 13918 31106 13970 31118
rect 13918 31042 13970 31054
rect 15598 31106 15650 31118
rect 15598 31042 15650 31054
rect 17390 31106 17442 31118
rect 21982 31106 22034 31118
rect 20066 31054 20078 31106
rect 20130 31054 20142 31106
rect 17390 31042 17442 31054
rect 21982 31042 22034 31054
rect 22094 31106 22146 31118
rect 22094 31042 22146 31054
rect 23550 31106 23602 31118
rect 23550 31042 23602 31054
rect 24558 31106 24610 31118
rect 24558 31042 24610 31054
rect 28478 31106 28530 31118
rect 36990 31106 37042 31118
rect 46174 31106 46226 31118
rect 49198 31106 49250 31118
rect 32498 31054 32510 31106
rect 32562 31054 32574 31106
rect 43810 31054 43822 31106
rect 43874 31054 43886 31106
rect 44594 31054 44606 31106
rect 44658 31054 44670 31106
rect 47954 31054 47966 31106
rect 48018 31054 48030 31106
rect 28478 31042 28530 31054
rect 36990 31042 37042 31054
rect 46174 31042 46226 31054
rect 49198 31042 49250 31054
rect 49422 31106 49474 31118
rect 49422 31042 49474 31054
rect 50094 31106 50146 31118
rect 52434 31054 52446 31106
rect 52498 31054 52510 31106
rect 57810 31054 57822 31106
rect 57874 31054 57886 31106
rect 50094 31042 50146 31054
rect 2494 30994 2546 31006
rect 2494 30930 2546 30942
rect 3502 30994 3554 31006
rect 3502 30930 3554 30942
rect 3726 30994 3778 31006
rect 3726 30930 3778 30942
rect 4062 30994 4114 31006
rect 4062 30930 4114 30942
rect 4286 30994 4338 31006
rect 4286 30930 4338 30942
rect 5406 30994 5458 31006
rect 9550 30994 9602 31006
rect 6290 30942 6302 30994
rect 6354 30942 6366 30994
rect 6850 30942 6862 30994
rect 6914 30942 6926 30994
rect 7970 30942 7982 30994
rect 8034 30942 8046 30994
rect 8642 30942 8654 30994
rect 8706 30942 8718 30994
rect 5406 30930 5458 30942
rect 9550 30930 9602 30942
rect 9662 30994 9714 31006
rect 9662 30930 9714 30942
rect 11454 30994 11506 31006
rect 16270 30994 16322 31006
rect 13010 30942 13022 30994
rect 13074 30942 13086 30994
rect 14690 30942 14702 30994
rect 14754 30942 14766 30994
rect 11454 30930 11506 30942
rect 16270 30930 16322 30942
rect 17838 30994 17890 31006
rect 17838 30930 17890 30942
rect 17950 30994 18002 31006
rect 22878 30994 22930 31006
rect 20962 30942 20974 30994
rect 21026 30942 21038 30994
rect 17950 30930 18002 30942
rect 22878 30930 22930 30942
rect 23326 30994 23378 31006
rect 23326 30930 23378 30942
rect 25902 30994 25954 31006
rect 28926 30994 28978 31006
rect 38446 30994 38498 31006
rect 26898 30942 26910 30994
rect 26962 30942 26974 30994
rect 28242 30942 28254 30994
rect 28306 30942 28318 30994
rect 29810 30942 29822 30994
rect 29874 30942 29886 30994
rect 32274 30942 32286 30994
rect 32338 30942 32350 30994
rect 36082 30942 36094 30994
rect 36146 30942 36158 30994
rect 25902 30930 25954 30942
rect 28926 30930 28978 30942
rect 38446 30930 38498 30942
rect 38670 30994 38722 31006
rect 42814 30994 42866 31006
rect 46062 30994 46114 31006
rect 49310 30994 49362 31006
rect 41346 30942 41358 30994
rect 41410 30942 41422 30994
rect 43138 30942 43150 30994
rect 43202 30942 43214 30994
rect 45266 30942 45278 30994
rect 45330 30942 45342 30994
rect 45826 30942 45838 30994
rect 45890 30942 45902 30994
rect 47282 30942 47294 30994
rect 47346 30942 47358 30994
rect 48178 30942 48190 30994
rect 48242 30942 48254 30994
rect 38670 30930 38722 30942
rect 42814 30930 42866 30942
rect 46062 30930 46114 30942
rect 49310 30930 49362 30942
rect 50206 30994 50258 31006
rect 50206 30930 50258 30942
rect 50430 30994 50482 31006
rect 50430 30930 50482 30942
rect 50878 30994 50930 31006
rect 58158 30994 58210 31006
rect 51538 30942 51550 30994
rect 51602 30942 51614 30994
rect 52322 30942 52334 30994
rect 52386 30942 52398 30994
rect 52882 30942 52894 30994
rect 52946 30942 52958 30994
rect 54338 30942 54350 30994
rect 54402 30942 54414 30994
rect 50878 30930 50930 30942
rect 58158 30930 58210 30942
rect 3838 30882 3890 30894
rect 15262 30882 15314 30894
rect 6178 30830 6190 30882
rect 6242 30830 6254 30882
rect 8530 30830 8542 30882
rect 8594 30830 8606 30882
rect 13122 30830 13134 30882
rect 13186 30830 13198 30882
rect 14354 30830 14366 30882
rect 14418 30830 14430 30882
rect 3838 30818 3890 30830
rect 15262 30818 15314 30830
rect 17726 30882 17778 30894
rect 21646 30882 21698 30894
rect 19506 30830 19518 30882
rect 19570 30830 19582 30882
rect 17726 30818 17778 30830
rect 21646 30818 21698 30830
rect 24334 30882 24386 30894
rect 25678 30882 25730 30894
rect 24658 30830 24670 30882
rect 24722 30830 24734 30882
rect 24334 30818 24386 30830
rect 25678 30818 25730 30830
rect 26574 30882 26626 30894
rect 26574 30818 26626 30830
rect 26686 30882 26738 30894
rect 26686 30818 26738 30830
rect 30494 30882 30546 30894
rect 30494 30818 30546 30830
rect 31838 30882 31890 30894
rect 31838 30818 31890 30830
rect 35422 30882 35474 30894
rect 35422 30818 35474 30830
rect 39342 30882 39394 30894
rect 51102 30882 51154 30894
rect 47618 30830 47630 30882
rect 47682 30830 47694 30882
rect 39342 30818 39394 30830
rect 51102 30818 51154 30830
rect 51326 30882 51378 30894
rect 57598 30882 57650 30894
rect 53890 30830 53902 30882
rect 53954 30830 53966 30882
rect 51326 30818 51378 30830
rect 57598 30818 57650 30830
rect 6862 30770 6914 30782
rect 12350 30770 12402 30782
rect 8642 30718 8654 30770
rect 8706 30718 8718 30770
rect 6862 30706 6914 30718
rect 12350 30706 12402 30718
rect 16494 30770 16546 30782
rect 22094 30770 22146 30782
rect 16818 30718 16830 30770
rect 16882 30718 16894 30770
rect 16494 30706 16546 30718
rect 22094 30706 22146 30718
rect 29038 30770 29090 30782
rect 29038 30706 29090 30718
rect 29262 30770 29314 30782
rect 29262 30706 29314 30718
rect 34862 30770 34914 30782
rect 34862 30706 34914 30718
rect 35198 30770 35250 30782
rect 35198 30706 35250 30718
rect 35758 30770 35810 30782
rect 35758 30706 35810 30718
rect 36094 30770 36146 30782
rect 36094 30706 36146 30718
rect 37326 30770 37378 30782
rect 50094 30770 50146 30782
rect 46610 30718 46622 30770
rect 46674 30718 46686 30770
rect 48738 30718 48750 30770
rect 48802 30718 48814 30770
rect 53554 30718 53566 30770
rect 53618 30718 53630 30770
rect 37326 30706 37378 30718
rect 50094 30706 50146 30718
rect 1344 30602 58576 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 58576 30602
rect 1344 30516 58576 30550
rect 4510 30434 4562 30446
rect 4510 30370 4562 30382
rect 4734 30434 4786 30446
rect 4734 30370 4786 30382
rect 7086 30434 7138 30446
rect 21422 30434 21474 30446
rect 28590 30434 28642 30446
rect 8978 30382 8990 30434
rect 9042 30382 9054 30434
rect 24658 30382 24670 30434
rect 24722 30382 24734 30434
rect 7086 30370 7138 30382
rect 21422 30370 21474 30382
rect 28590 30370 28642 30382
rect 30494 30434 30546 30446
rect 30494 30370 30546 30382
rect 32398 30434 32450 30446
rect 32398 30370 32450 30382
rect 38894 30434 38946 30446
rect 38894 30370 38946 30382
rect 39902 30434 39954 30446
rect 39902 30370 39954 30382
rect 44046 30434 44098 30446
rect 44046 30370 44098 30382
rect 44830 30434 44882 30446
rect 44830 30370 44882 30382
rect 45390 30434 45442 30446
rect 45390 30370 45442 30382
rect 45614 30434 45666 30446
rect 45614 30370 45666 30382
rect 46398 30434 46450 30446
rect 46398 30370 46450 30382
rect 17614 30322 17666 30334
rect 29710 30322 29762 30334
rect 6066 30270 6078 30322
rect 6130 30270 6142 30322
rect 9874 30270 9886 30322
rect 9938 30270 9950 30322
rect 20178 30270 20190 30322
rect 20242 30270 20254 30322
rect 21746 30270 21758 30322
rect 21810 30270 21822 30322
rect 23538 30270 23550 30322
rect 23602 30270 23614 30322
rect 17614 30258 17666 30270
rect 29710 30258 29762 30270
rect 29934 30322 29986 30334
rect 29934 30258 29986 30270
rect 31614 30322 31666 30334
rect 31614 30258 31666 30270
rect 39230 30322 39282 30334
rect 39230 30258 39282 30270
rect 40126 30322 40178 30334
rect 40126 30258 40178 30270
rect 42590 30322 42642 30334
rect 43822 30322 43874 30334
rect 43362 30270 43374 30322
rect 43426 30270 43438 30322
rect 47842 30270 47854 30322
rect 47906 30270 47918 30322
rect 42590 30258 42642 30270
rect 43822 30258 43874 30270
rect 6302 30210 6354 30222
rect 2482 30158 2494 30210
rect 2546 30158 2558 30210
rect 3490 30158 3502 30210
rect 3554 30158 3566 30210
rect 4274 30158 4286 30210
rect 4338 30158 4350 30210
rect 6302 30146 6354 30158
rect 6638 30210 6690 30222
rect 6638 30146 6690 30158
rect 7198 30210 7250 30222
rect 12686 30210 12738 30222
rect 7970 30158 7982 30210
rect 8034 30158 8046 30210
rect 8642 30158 8654 30210
rect 8706 30158 8718 30210
rect 9202 30158 9214 30210
rect 9266 30158 9278 30210
rect 10322 30158 10334 30210
rect 10386 30158 10398 30210
rect 7198 30146 7250 30158
rect 12686 30146 12738 30158
rect 13022 30210 13074 30222
rect 13022 30146 13074 30158
rect 13470 30210 13522 30222
rect 13470 30146 13522 30158
rect 13806 30210 13858 30222
rect 13806 30146 13858 30158
rect 13918 30210 13970 30222
rect 13918 30146 13970 30158
rect 14366 30210 14418 30222
rect 14366 30146 14418 30158
rect 16606 30210 16658 30222
rect 16606 30146 16658 30158
rect 16942 30210 16994 30222
rect 16942 30146 16994 30158
rect 17166 30210 17218 30222
rect 17166 30146 17218 30158
rect 17390 30210 17442 30222
rect 22094 30210 22146 30222
rect 23102 30210 23154 30222
rect 24110 30210 24162 30222
rect 25230 30210 25282 30222
rect 29486 30210 29538 30222
rect 36990 30210 37042 30222
rect 19730 30158 19742 30210
rect 19794 30158 19806 30210
rect 22306 30158 22318 30210
rect 22370 30158 22382 30210
rect 23314 30158 23326 30210
rect 23378 30158 23390 30210
rect 24322 30158 24334 30210
rect 24386 30158 24398 30210
rect 24882 30158 24894 30210
rect 24946 30158 24958 30210
rect 26114 30158 26126 30210
rect 26178 30158 26190 30210
rect 27010 30158 27022 30210
rect 27074 30158 27086 30210
rect 27794 30158 27806 30210
rect 27858 30158 27870 30210
rect 31266 30158 31278 30210
rect 31330 30158 31342 30210
rect 32498 30158 32510 30210
rect 32562 30158 32574 30210
rect 34066 30158 34078 30210
rect 34130 30158 34142 30210
rect 35074 30158 35086 30210
rect 35138 30158 35150 30210
rect 36194 30158 36206 30210
rect 36258 30158 36270 30210
rect 17390 30146 17442 30158
rect 22094 30146 22146 30158
rect 23102 30146 23154 30158
rect 24110 30146 24162 30158
rect 25230 30146 25282 30158
rect 29486 30146 29538 30158
rect 36990 30146 37042 30158
rect 37662 30210 37714 30222
rect 39790 30210 39842 30222
rect 38658 30158 38670 30210
rect 38722 30158 38734 30210
rect 37662 30146 37714 30158
rect 39790 30146 39842 30158
rect 41470 30210 41522 30222
rect 41470 30146 41522 30158
rect 41918 30210 41970 30222
rect 41918 30146 41970 30158
rect 42142 30210 42194 30222
rect 42142 30146 42194 30158
rect 43710 30210 43762 30222
rect 44942 30210 44994 30222
rect 44258 30158 44270 30210
rect 44322 30158 44334 30210
rect 43710 30146 43762 30158
rect 44942 30146 44994 30158
rect 46622 30210 46674 30222
rect 46622 30146 46674 30158
rect 47630 30210 47682 30222
rect 55570 30158 55582 30210
rect 55634 30158 55646 30210
rect 47630 30146 47682 30158
rect 4846 30098 4898 30110
rect 2370 30046 2382 30098
rect 2434 30046 2446 30098
rect 4846 30034 4898 30046
rect 7086 30098 7138 30110
rect 7086 30034 7138 30046
rect 10782 30098 10834 30110
rect 10782 30034 10834 30046
rect 14590 30098 14642 30110
rect 14590 30034 14642 30046
rect 17950 30098 18002 30110
rect 17950 30034 18002 30046
rect 19294 30098 19346 30110
rect 19294 30034 19346 30046
rect 25342 30098 25394 30110
rect 28478 30098 28530 30110
rect 26338 30046 26350 30098
rect 26402 30046 26414 30098
rect 26898 30046 26910 30098
rect 26962 30046 26974 30098
rect 25342 30034 25394 30046
rect 28478 30034 28530 30046
rect 30270 30098 30322 30110
rect 30270 30034 30322 30046
rect 31502 30098 31554 30110
rect 31502 30034 31554 30046
rect 31950 30098 32002 30110
rect 37326 30098 37378 30110
rect 39342 30098 39394 30110
rect 32162 30046 32174 30098
rect 32226 30046 32238 30098
rect 35298 30046 35310 30098
rect 35362 30046 35374 30098
rect 36082 30046 36094 30098
rect 36146 30046 36158 30098
rect 39106 30046 39118 30098
rect 39170 30046 39182 30098
rect 31950 30034 32002 30046
rect 37326 30034 37378 30046
rect 39342 30034 39394 30046
rect 40238 30098 40290 30110
rect 40238 30034 40290 30046
rect 41134 30098 41186 30110
rect 41134 30034 41186 30046
rect 41246 30098 41298 30110
rect 41246 30034 41298 30046
rect 42478 30098 42530 30110
rect 42478 30034 42530 30046
rect 43038 30098 43090 30110
rect 43038 30034 43090 30046
rect 43262 30098 43314 30110
rect 43262 30034 43314 30046
rect 45166 30098 45218 30110
rect 45166 30034 45218 30046
rect 47294 30098 47346 30110
rect 57250 30046 57262 30098
rect 57314 30046 57326 30098
rect 47294 30034 47346 30046
rect 12798 29986 12850 29998
rect 3602 29934 3614 29986
rect 3666 29934 3678 29986
rect 12798 29922 12850 29934
rect 13582 29986 13634 29998
rect 13582 29922 13634 29934
rect 14254 29986 14306 29998
rect 14254 29922 14306 29934
rect 17054 29986 17106 29998
rect 17054 29922 17106 29934
rect 17726 29986 17778 29998
rect 17726 29922 17778 29934
rect 21646 29986 21698 29998
rect 21646 29922 21698 29934
rect 24222 29986 24274 29998
rect 24222 29922 24274 29934
rect 25566 29986 25618 29998
rect 25566 29922 25618 29934
rect 28254 29986 28306 29998
rect 28254 29922 28306 29934
rect 29038 29986 29090 29998
rect 32734 29986 32786 29998
rect 30818 29934 30830 29986
rect 30882 29934 30894 29986
rect 29038 29922 29090 29934
rect 32734 29922 32786 29934
rect 33742 29986 33794 29998
rect 37214 29986 37266 29998
rect 35186 29934 35198 29986
rect 35250 29934 35262 29986
rect 33742 29922 33794 29934
rect 37214 29922 37266 29934
rect 37774 29986 37826 29998
rect 37774 29922 37826 29934
rect 37886 29986 37938 29998
rect 37886 29922 37938 29934
rect 38110 29986 38162 29998
rect 38110 29922 38162 29934
rect 40910 29986 40962 29998
rect 40910 29922 40962 29934
rect 41694 29986 41746 29998
rect 46050 29934 46062 29986
rect 46114 29934 46126 29986
rect 41694 29922 41746 29934
rect 1344 29818 58576 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 50558 29818
rect 50610 29766 50662 29818
rect 50714 29766 50766 29818
rect 50818 29766 58576 29818
rect 1344 29732 58576 29766
rect 15038 29650 15090 29662
rect 3826 29598 3838 29650
rect 3890 29598 3902 29650
rect 11442 29598 11454 29650
rect 11506 29598 11518 29650
rect 14590 29594 14642 29606
rect 3166 29538 3218 29550
rect 3166 29474 3218 29486
rect 3278 29538 3330 29550
rect 3278 29474 3330 29486
rect 3390 29538 3442 29550
rect 14478 29538 14530 29550
rect 4386 29486 4398 29538
rect 4450 29486 4462 29538
rect 10658 29486 10670 29538
rect 10722 29486 10734 29538
rect 15038 29586 15090 29598
rect 15598 29650 15650 29662
rect 15598 29586 15650 29598
rect 15934 29650 15986 29662
rect 15934 29586 15986 29598
rect 16606 29650 16658 29662
rect 16606 29586 16658 29598
rect 16830 29650 16882 29662
rect 16830 29586 16882 29598
rect 17614 29650 17666 29662
rect 17614 29586 17666 29598
rect 22206 29650 22258 29662
rect 22206 29586 22258 29598
rect 22542 29650 22594 29662
rect 22542 29586 22594 29598
rect 27134 29650 27186 29662
rect 27134 29586 27186 29598
rect 28142 29650 28194 29662
rect 30382 29650 30434 29662
rect 30034 29598 30046 29650
rect 30098 29598 30110 29650
rect 28142 29586 28194 29598
rect 30382 29586 30434 29598
rect 32062 29650 32114 29662
rect 35758 29650 35810 29662
rect 33506 29598 33518 29650
rect 33570 29598 33582 29650
rect 32062 29586 32114 29598
rect 35758 29586 35810 29598
rect 43822 29650 43874 29662
rect 43822 29586 43874 29598
rect 43934 29650 43986 29662
rect 43934 29586 43986 29598
rect 44718 29650 44770 29662
rect 44718 29586 44770 29598
rect 45390 29650 45442 29662
rect 45390 29586 45442 29598
rect 45950 29650 46002 29662
rect 45950 29586 46002 29598
rect 57598 29650 57650 29662
rect 57598 29586 57650 29598
rect 14590 29530 14642 29542
rect 16046 29538 16098 29550
rect 3390 29474 3442 29486
rect 14478 29474 14530 29486
rect 16046 29474 16098 29486
rect 21758 29538 21810 29550
rect 28478 29538 28530 29550
rect 26786 29486 26798 29538
rect 26850 29486 26862 29538
rect 21758 29474 21810 29486
rect 28478 29474 28530 29486
rect 28702 29538 28754 29550
rect 28702 29474 28754 29486
rect 31726 29538 31778 29550
rect 31726 29474 31778 29486
rect 35310 29538 35362 29550
rect 35310 29474 35362 29486
rect 35982 29538 36034 29550
rect 35982 29474 36034 29486
rect 36766 29538 36818 29550
rect 36766 29474 36818 29486
rect 37102 29538 37154 29550
rect 37102 29474 37154 29486
rect 37326 29538 37378 29550
rect 37326 29474 37378 29486
rect 45502 29538 45554 29550
rect 45502 29474 45554 29486
rect 57822 29538 57874 29550
rect 57822 29474 57874 29486
rect 58158 29538 58210 29550
rect 58158 29474 58210 29486
rect 15710 29426 15762 29438
rect 17390 29426 17442 29438
rect 4162 29374 4174 29426
rect 4226 29374 4238 29426
rect 5058 29374 5070 29426
rect 5122 29374 5134 29426
rect 7298 29374 7310 29426
rect 7362 29374 7374 29426
rect 7746 29374 7758 29426
rect 7810 29374 7822 29426
rect 8418 29374 8430 29426
rect 8482 29374 8494 29426
rect 10434 29374 10446 29426
rect 10498 29374 10510 29426
rect 11330 29374 11342 29426
rect 11394 29374 11406 29426
rect 16370 29374 16382 29426
rect 16434 29374 16446 29426
rect 15710 29362 15762 29374
rect 17390 29362 17442 29374
rect 18062 29426 18114 29438
rect 18062 29362 18114 29374
rect 18398 29426 18450 29438
rect 18398 29362 18450 29374
rect 18622 29426 18674 29438
rect 18622 29362 18674 29374
rect 18958 29426 19010 29438
rect 18958 29362 19010 29374
rect 19294 29426 19346 29438
rect 19294 29362 19346 29374
rect 19518 29426 19570 29438
rect 19518 29362 19570 29374
rect 19966 29426 20018 29438
rect 22430 29426 22482 29438
rect 21410 29374 21422 29426
rect 21474 29374 21486 29426
rect 19966 29362 20018 29374
rect 22430 29362 22482 29374
rect 22654 29426 22706 29438
rect 22654 29362 22706 29374
rect 29150 29426 29202 29438
rect 31390 29426 31442 29438
rect 29586 29374 29598 29426
rect 29650 29374 29662 29426
rect 29150 29362 29202 29374
rect 31390 29362 31442 29374
rect 32398 29426 32450 29438
rect 33854 29426 33906 29438
rect 34862 29426 34914 29438
rect 33058 29374 33070 29426
rect 33122 29374 33134 29426
rect 33618 29374 33630 29426
rect 33682 29374 33694 29426
rect 34738 29374 34750 29426
rect 34802 29374 34814 29426
rect 32398 29362 32450 29374
rect 33854 29362 33906 29374
rect 34862 29362 34914 29374
rect 34974 29426 35026 29438
rect 34974 29362 35026 29374
rect 35646 29426 35698 29438
rect 35646 29362 35698 29374
rect 36206 29426 36258 29438
rect 36206 29362 36258 29374
rect 38670 29426 38722 29438
rect 38670 29362 38722 29374
rect 39118 29426 39170 29438
rect 39118 29362 39170 29374
rect 40910 29426 40962 29438
rect 43710 29426 43762 29438
rect 44942 29426 44994 29438
rect 41682 29374 41694 29426
rect 41746 29374 41758 29426
rect 43026 29374 43038 29426
rect 43090 29374 43102 29426
rect 44258 29374 44270 29426
rect 44322 29374 44334 29426
rect 40910 29362 40962 29374
rect 43710 29362 43762 29374
rect 44942 29362 44994 29374
rect 13134 29314 13186 29326
rect 17502 29314 17554 29326
rect 4722 29262 4734 29314
rect 4786 29262 4798 29314
rect 7410 29262 7422 29314
rect 7474 29262 7486 29314
rect 8530 29262 8542 29314
rect 8594 29262 8606 29314
rect 16706 29262 16718 29314
rect 16770 29262 16782 29314
rect 13134 29250 13186 29262
rect 17502 29250 17554 29262
rect 18510 29314 18562 29326
rect 18510 29250 18562 29262
rect 19406 29314 19458 29326
rect 19406 29250 19458 29262
rect 20638 29314 20690 29326
rect 20638 29250 20690 29262
rect 21086 29314 21138 29326
rect 21086 29250 21138 29262
rect 21646 29314 21698 29326
rect 35198 29314 35250 29326
rect 28802 29262 28814 29314
rect 28866 29262 28878 29314
rect 21646 29250 21698 29262
rect 35198 29250 35250 29262
rect 36878 29314 36930 29326
rect 42914 29262 42926 29314
rect 42978 29262 42990 29314
rect 36878 29250 36930 29262
rect 14478 29202 14530 29214
rect 44606 29202 44658 29214
rect 8306 29150 8318 29202
rect 8370 29150 8382 29202
rect 33282 29150 33294 29202
rect 33346 29150 33358 29202
rect 38434 29150 38446 29202
rect 38498 29150 38510 29202
rect 14478 29138 14530 29150
rect 44606 29138 44658 29150
rect 45390 29202 45442 29214
rect 45390 29138 45442 29150
rect 1344 29034 58576 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 58576 29034
rect 1344 28948 58576 28982
rect 8766 28866 8818 28878
rect 8766 28802 8818 28814
rect 9102 28866 9154 28878
rect 9102 28802 9154 28814
rect 15262 28866 15314 28878
rect 15262 28802 15314 28814
rect 18174 28866 18226 28878
rect 18174 28802 18226 28814
rect 21758 28866 21810 28878
rect 21758 28802 21810 28814
rect 29486 28866 29538 28878
rect 29486 28802 29538 28814
rect 30046 28866 30098 28878
rect 30046 28802 30098 28814
rect 4958 28754 5010 28766
rect 4162 28702 4174 28754
rect 4226 28702 4238 28754
rect 4958 28690 5010 28702
rect 8430 28754 8482 28766
rect 15710 28754 15762 28766
rect 10770 28702 10782 28754
rect 10834 28702 10846 28754
rect 14130 28702 14142 28754
rect 14194 28702 14206 28754
rect 8430 28690 8482 28702
rect 15710 28690 15762 28702
rect 16382 28754 16434 28766
rect 16382 28690 16434 28702
rect 18734 28754 18786 28766
rect 18734 28690 18786 28702
rect 20190 28754 20242 28766
rect 20190 28690 20242 28702
rect 21982 28754 22034 28766
rect 29710 28754 29762 28766
rect 39678 28754 39730 28766
rect 26786 28702 26798 28754
rect 26850 28702 26862 28754
rect 32274 28702 32286 28754
rect 32338 28702 32350 28754
rect 39218 28702 39230 28754
rect 39282 28702 39294 28754
rect 21982 28690 22034 28702
rect 29710 28690 29762 28702
rect 39678 28690 39730 28702
rect 43598 28754 43650 28766
rect 43598 28690 43650 28702
rect 44158 28754 44210 28766
rect 44158 28690 44210 28702
rect 44942 28754 44994 28766
rect 44942 28690 44994 28702
rect 57934 28754 57986 28766
rect 57934 28690 57986 28702
rect 11230 28642 11282 28654
rect 12798 28642 12850 28654
rect 17726 28642 17778 28654
rect 4274 28590 4286 28642
rect 4338 28590 4350 28642
rect 6962 28590 6974 28642
rect 7026 28590 7038 28642
rect 7858 28590 7870 28642
rect 7922 28590 7934 28642
rect 8754 28590 8766 28642
rect 8818 28590 8830 28642
rect 10546 28590 10558 28642
rect 10610 28590 10622 28642
rect 12562 28590 12574 28642
rect 12626 28590 12638 28642
rect 13906 28590 13918 28642
rect 13970 28590 13982 28642
rect 14354 28590 14366 28642
rect 14418 28590 14430 28642
rect 14914 28590 14926 28642
rect 14978 28590 14990 28642
rect 11230 28578 11282 28590
rect 12798 28578 12850 28590
rect 17726 28578 17778 28590
rect 20414 28642 20466 28654
rect 20414 28578 20466 28590
rect 20750 28642 20802 28654
rect 27022 28642 27074 28654
rect 30830 28642 30882 28654
rect 32734 28642 32786 28654
rect 37102 28642 37154 28654
rect 22866 28590 22878 28642
rect 22930 28590 22942 28642
rect 23986 28590 23998 28642
rect 24050 28590 24062 28642
rect 30370 28590 30382 28642
rect 30434 28590 30446 28642
rect 31042 28590 31054 28642
rect 31106 28590 31118 28642
rect 35298 28590 35310 28642
rect 35362 28590 35374 28642
rect 20750 28578 20802 28590
rect 27022 28578 27074 28590
rect 30830 28578 30882 28590
rect 32734 28578 32786 28590
rect 37102 28578 37154 28590
rect 37662 28642 37714 28654
rect 37662 28578 37714 28590
rect 38110 28642 38162 28654
rect 55246 28642 55298 28654
rect 38882 28590 38894 28642
rect 38946 28590 38958 28642
rect 55570 28590 55582 28642
rect 55634 28590 55646 28642
rect 38110 28578 38162 28590
rect 55246 28578 55298 28590
rect 12014 28530 12066 28542
rect 6514 28478 6526 28530
rect 6578 28478 6590 28530
rect 12014 28466 12066 28478
rect 12126 28530 12178 28542
rect 12126 28466 12178 28478
rect 12350 28530 12402 28542
rect 12350 28466 12402 28478
rect 12910 28530 12962 28542
rect 17502 28530 17554 28542
rect 13570 28478 13582 28530
rect 13634 28478 13646 28530
rect 12910 28466 12962 28478
rect 17502 28466 17554 28478
rect 18062 28530 18114 28542
rect 18062 28466 18114 28478
rect 20638 28530 20690 28542
rect 20638 28466 20690 28478
rect 22542 28530 22594 28542
rect 27246 28530 27298 28542
rect 24658 28478 24670 28530
rect 24722 28478 24734 28530
rect 22542 28466 22594 28478
rect 27246 28466 27298 28478
rect 27358 28530 27410 28542
rect 27358 28466 27410 28478
rect 27806 28530 27858 28542
rect 27806 28466 27858 28478
rect 30718 28530 30770 28542
rect 30718 28466 30770 28478
rect 34526 28530 34578 28542
rect 34526 28466 34578 28478
rect 35534 28530 35586 28542
rect 35534 28466 35586 28478
rect 36094 28530 36146 28542
rect 36094 28466 36146 28478
rect 36206 28530 36258 28542
rect 38994 28478 39006 28530
rect 39058 28478 39070 28530
rect 36206 28466 36258 28478
rect 11790 28418 11842 28430
rect 11790 28354 11842 28366
rect 15150 28418 15202 28430
rect 15150 28354 15202 28366
rect 16942 28418 16994 28430
rect 16942 28354 16994 28366
rect 17278 28418 17330 28430
rect 17278 28354 17330 28366
rect 17614 28418 17666 28430
rect 17614 28354 17666 28366
rect 18174 28418 18226 28430
rect 22318 28418 22370 28430
rect 21410 28366 21422 28418
rect 21474 28366 21486 28418
rect 18174 28354 18226 28366
rect 22318 28354 22370 28366
rect 22430 28418 22482 28430
rect 30158 28418 30210 28430
rect 29138 28366 29150 28418
rect 29202 28366 29214 28418
rect 22430 28354 22482 28366
rect 30158 28354 30210 28366
rect 34302 28418 34354 28430
rect 34302 28354 34354 28366
rect 34414 28418 34466 28430
rect 34414 28354 34466 28366
rect 34750 28418 34802 28430
rect 34750 28354 34802 28366
rect 36430 28418 36482 28430
rect 36430 28354 36482 28366
rect 38446 28418 38498 28430
rect 38446 28354 38498 28366
rect 38670 28418 38722 28430
rect 38670 28354 38722 28366
rect 1344 28250 58576 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 50558 28250
rect 50610 28198 50662 28250
rect 50714 28198 50766 28250
rect 50818 28198 58576 28250
rect 1344 28164 58576 28198
rect 16270 28082 16322 28094
rect 7410 28030 7422 28082
rect 7474 28030 7486 28082
rect 10882 28030 10894 28082
rect 10946 28030 10958 28082
rect 16270 28018 16322 28030
rect 17502 28082 17554 28094
rect 17502 28018 17554 28030
rect 20750 28082 20802 28094
rect 20750 28018 20802 28030
rect 21422 28082 21474 28094
rect 21422 28018 21474 28030
rect 25342 28082 25394 28094
rect 25342 28018 25394 28030
rect 25454 28082 25506 28094
rect 25454 28018 25506 28030
rect 25678 28082 25730 28094
rect 25678 28018 25730 28030
rect 27246 28082 27298 28094
rect 33182 28082 33234 28094
rect 30930 28030 30942 28082
rect 30994 28030 31006 28082
rect 27246 28018 27298 28030
rect 33182 28018 33234 28030
rect 33294 28082 33346 28094
rect 33294 28018 33346 28030
rect 34078 28082 34130 28094
rect 34078 28018 34130 28030
rect 38110 28082 38162 28094
rect 38110 28018 38162 28030
rect 38334 28082 38386 28094
rect 38334 28018 38386 28030
rect 38446 28082 38498 28094
rect 38446 28018 38498 28030
rect 41022 28082 41074 28094
rect 41022 28018 41074 28030
rect 43038 28082 43090 28094
rect 43038 28018 43090 28030
rect 43262 28082 43314 28094
rect 43262 28018 43314 28030
rect 45502 28082 45554 28094
rect 45502 28018 45554 28030
rect 46062 28082 46114 28094
rect 46062 28018 46114 28030
rect 15822 27970 15874 27982
rect 12562 27918 12574 27970
rect 12626 27918 12638 27970
rect 13906 27918 13918 27970
rect 13970 27918 13982 27970
rect 15822 27906 15874 27918
rect 18062 27970 18114 27982
rect 18062 27906 18114 27918
rect 18958 27970 19010 27982
rect 18958 27906 19010 27918
rect 21646 27970 21698 27982
rect 21646 27906 21698 27918
rect 29934 27970 29986 27982
rect 29934 27906 29986 27918
rect 33070 27970 33122 27982
rect 33070 27906 33122 27918
rect 33854 27970 33906 27982
rect 33854 27906 33906 27918
rect 34190 27970 34242 27982
rect 38670 27970 38722 27982
rect 35522 27918 35534 27970
rect 35586 27918 35598 27970
rect 34190 27906 34242 27918
rect 38670 27906 38722 27918
rect 38782 27970 38834 27982
rect 38782 27906 38834 27918
rect 39230 27970 39282 27982
rect 39230 27906 39282 27918
rect 39678 27970 39730 27982
rect 39678 27906 39730 27918
rect 40798 27970 40850 27982
rect 44718 27970 44770 27982
rect 44258 27918 44270 27970
rect 44322 27918 44334 27970
rect 40798 27906 40850 27918
rect 44718 27906 44770 27918
rect 44830 27970 44882 27982
rect 44830 27906 44882 27918
rect 57822 27970 57874 27982
rect 57822 27906 57874 27918
rect 6862 27858 6914 27870
rect 6862 27794 6914 27806
rect 7086 27858 7138 27870
rect 8990 27858 9042 27870
rect 8082 27806 8094 27858
rect 8146 27806 8158 27858
rect 7086 27794 7138 27806
rect 8990 27794 9042 27806
rect 10334 27858 10386 27870
rect 10334 27794 10386 27806
rect 10558 27858 10610 27870
rect 15598 27858 15650 27870
rect 12786 27806 12798 27858
rect 12850 27806 12862 27858
rect 14914 27806 14926 27858
rect 14978 27806 14990 27858
rect 10558 27794 10610 27806
rect 15598 27794 15650 27806
rect 17950 27858 18002 27870
rect 17950 27794 18002 27806
rect 18510 27858 18562 27870
rect 18510 27794 18562 27806
rect 18734 27858 18786 27870
rect 18734 27794 18786 27806
rect 18846 27858 18898 27870
rect 18846 27794 18898 27806
rect 19406 27858 19458 27870
rect 25230 27858 25282 27870
rect 22530 27806 22542 27858
rect 22594 27806 22606 27858
rect 19406 27794 19458 27806
rect 25230 27794 25282 27806
rect 28366 27858 28418 27870
rect 28366 27794 28418 27806
rect 28926 27858 28978 27870
rect 30606 27858 30658 27870
rect 30146 27806 30158 27858
rect 30210 27806 30222 27858
rect 28926 27794 28978 27806
rect 30606 27794 30658 27806
rect 33742 27858 33794 27870
rect 37998 27858 38050 27870
rect 34738 27806 34750 27858
rect 34802 27806 34814 27858
rect 33742 27794 33794 27806
rect 37998 27794 38050 27806
rect 39566 27858 39618 27870
rect 39566 27794 39618 27806
rect 39902 27858 39954 27870
rect 39902 27794 39954 27806
rect 41134 27858 41186 27870
rect 41134 27794 41186 27806
rect 42702 27858 42754 27870
rect 42702 27794 42754 27806
rect 42926 27858 42978 27870
rect 44046 27858 44098 27870
rect 58158 27858 58210 27870
rect 43810 27806 43822 27858
rect 43874 27806 43886 27858
rect 45042 27806 45054 27858
rect 45106 27806 45118 27858
rect 42926 27794 42978 27806
rect 44046 27794 44098 27806
rect 58158 27794 58210 27806
rect 14142 27746 14194 27758
rect 8418 27694 8430 27746
rect 8482 27694 8494 27746
rect 14142 27682 14194 27694
rect 18286 27746 18338 27758
rect 21534 27746 21586 27758
rect 31502 27746 31554 27758
rect 41582 27746 41634 27758
rect 20626 27694 20638 27746
rect 20690 27694 20702 27746
rect 22306 27694 22318 27746
rect 22370 27694 22382 27746
rect 37650 27694 37662 27746
rect 37714 27694 37726 27746
rect 18286 27682 18338 27694
rect 21534 27682 21586 27694
rect 31502 27682 31554 27694
rect 41582 27682 41634 27694
rect 44382 27746 44434 27758
rect 44382 27682 44434 27694
rect 57598 27746 57650 27758
rect 57598 27682 57650 27694
rect 20974 27634 21026 27646
rect 43374 27634 43426 27646
rect 22978 27582 22990 27634
rect 23042 27582 23054 27634
rect 20974 27570 21026 27582
rect 43374 27570 43426 27582
rect 1344 27466 58576 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 58576 27466
rect 1344 27380 58576 27414
rect 16270 27298 16322 27310
rect 16270 27234 16322 27246
rect 43598 27298 43650 27310
rect 43598 27234 43650 27246
rect 43822 27298 43874 27310
rect 43822 27234 43874 27246
rect 43934 27298 43986 27310
rect 43934 27234 43986 27246
rect 1934 27186 1986 27198
rect 1934 27122 1986 27134
rect 13918 27186 13970 27198
rect 21534 27186 21586 27198
rect 28030 27186 28082 27198
rect 30158 27186 30210 27198
rect 46510 27186 46562 27198
rect 14242 27134 14254 27186
rect 14306 27134 14318 27186
rect 16594 27134 16606 27186
rect 16658 27134 16670 27186
rect 17938 27134 17950 27186
rect 18002 27134 18014 27186
rect 27122 27134 27134 27186
rect 27186 27134 27198 27186
rect 29250 27134 29262 27186
rect 29314 27134 29326 27186
rect 32386 27134 32398 27186
rect 32450 27134 32462 27186
rect 34514 27134 34526 27186
rect 34578 27134 34590 27186
rect 40002 27134 40014 27186
rect 40066 27134 40078 27186
rect 42130 27134 42142 27186
rect 42194 27134 42206 27186
rect 45938 27134 45950 27186
rect 46002 27134 46014 27186
rect 13918 27122 13970 27134
rect 21534 27122 21586 27134
rect 28030 27122 28082 27134
rect 30158 27122 30210 27134
rect 46510 27122 46562 27134
rect 47070 27186 47122 27198
rect 47070 27122 47122 27134
rect 47518 27186 47570 27198
rect 47518 27122 47570 27134
rect 57934 27186 57986 27198
rect 57934 27122 57986 27134
rect 17054 27074 17106 27086
rect 20190 27074 20242 27086
rect 4274 27022 4286 27074
rect 4338 27022 4350 27074
rect 14690 27022 14702 27074
rect 14754 27022 14766 27074
rect 15138 27022 15150 27074
rect 15202 27022 15214 27074
rect 18162 27022 18174 27074
rect 18226 27022 18238 27074
rect 18610 27022 18622 27074
rect 18674 27022 18686 27074
rect 19282 27022 19294 27074
rect 19346 27022 19358 27074
rect 19842 27022 19854 27074
rect 19906 27022 19918 27074
rect 17054 27010 17106 27022
rect 20190 27010 20242 27022
rect 20750 27074 20802 27086
rect 28590 27074 28642 27086
rect 30494 27074 30546 27086
rect 21858 27022 21870 27074
rect 21922 27022 21934 27074
rect 24210 27022 24222 27074
rect 24274 27022 24286 27074
rect 29586 27022 29598 27074
rect 29650 27022 29662 27074
rect 20750 27010 20802 27022
rect 28590 27010 28642 27022
rect 30494 27010 30546 27022
rect 31054 27074 31106 27086
rect 31602 27022 31614 27074
rect 31666 27022 31678 27074
rect 39218 27022 39230 27074
rect 39282 27022 39294 27074
rect 45490 27022 45502 27074
rect 45554 27022 45566 27074
rect 45714 27022 45726 27074
rect 45778 27022 45790 27074
rect 55570 27022 55582 27074
rect 55634 27022 55646 27074
rect 31054 27010 31106 27022
rect 12014 26962 12066 26974
rect 12014 26898 12066 26910
rect 12350 26962 12402 26974
rect 16494 26962 16546 26974
rect 14466 26910 14478 26962
rect 14530 26910 14542 26962
rect 17390 26962 17442 26974
rect 21646 26962 21698 26974
rect 12350 26898 12402 26910
rect 16494 26898 16546 26910
rect 17166 26906 17218 26918
rect 12238 26850 12290 26862
rect 17602 26910 17614 26962
rect 17666 26910 17678 26962
rect 17390 26898 17442 26910
rect 21646 26898 21698 26910
rect 22878 26962 22930 26974
rect 22878 26898 22930 26910
rect 23102 26962 23154 26974
rect 23102 26898 23154 26910
rect 23214 26962 23266 26974
rect 23214 26898 23266 26910
rect 23774 26962 23826 26974
rect 27358 26962 27410 26974
rect 24994 26910 25006 26962
rect 25058 26910 25070 26962
rect 23774 26898 23826 26910
rect 27358 26898 27410 26910
rect 27582 26962 27634 26974
rect 42590 26962 42642 26974
rect 27582 26898 27634 26910
rect 27694 26906 27746 26918
rect 37426 26910 37438 26962
rect 37490 26910 37502 26962
rect 17166 26842 17218 26854
rect 23438 26850 23490 26862
rect 12238 26786 12290 26798
rect 42590 26898 42642 26910
rect 27694 26842 27746 26854
rect 35086 26850 35138 26862
rect 23438 26786 23490 26798
rect 35086 26786 35138 26798
rect 37774 26850 37826 26862
rect 37774 26786 37826 26798
rect 38222 26850 38274 26862
rect 38222 26786 38274 26798
rect 43038 26850 43090 26862
rect 43038 26786 43090 26798
rect 43934 26850 43986 26862
rect 43934 26786 43986 26798
rect 44718 26850 44770 26862
rect 44718 26786 44770 26798
rect 46398 26850 46450 26862
rect 46398 26786 46450 26798
rect 1344 26682 58576 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 50558 26682
rect 50610 26630 50662 26682
rect 50714 26630 50766 26682
rect 50818 26630 58576 26682
rect 1344 26596 58576 26630
rect 23774 26514 23826 26526
rect 23774 26450 23826 26462
rect 28926 26514 28978 26526
rect 28926 26450 28978 26462
rect 29150 26514 29202 26526
rect 29150 26450 29202 26462
rect 34862 26514 34914 26526
rect 34862 26450 34914 26462
rect 37102 26514 37154 26526
rect 37102 26450 37154 26462
rect 38446 26514 38498 26526
rect 57598 26514 57650 26526
rect 44930 26462 44942 26514
rect 44994 26462 45006 26514
rect 49074 26462 49086 26514
rect 49138 26462 49150 26514
rect 38446 26450 38498 26462
rect 57598 26450 57650 26462
rect 16270 26402 16322 26414
rect 11666 26350 11678 26402
rect 11730 26350 11742 26402
rect 16270 26338 16322 26350
rect 16830 26402 16882 26414
rect 28366 26402 28418 26414
rect 17714 26350 17726 26402
rect 17778 26350 17790 26402
rect 27906 26350 27918 26402
rect 27970 26350 27982 26402
rect 16830 26338 16882 26350
rect 28366 26338 28418 26350
rect 28590 26402 28642 26414
rect 28590 26338 28642 26350
rect 29262 26402 29314 26414
rect 40126 26402 40178 26414
rect 29474 26350 29486 26402
rect 29538 26350 29550 26402
rect 30370 26350 30382 26402
rect 30434 26350 30446 26402
rect 31042 26350 31054 26402
rect 31106 26350 31118 26402
rect 29262 26338 29314 26350
rect 40126 26338 40178 26350
rect 44382 26402 44434 26414
rect 44382 26338 44434 26350
rect 57822 26402 57874 26414
rect 57822 26338 57874 26350
rect 58158 26402 58210 26414
rect 58158 26338 58210 26350
rect 16046 26290 16098 26302
rect 4274 26238 4286 26290
rect 4338 26238 4350 26290
rect 12450 26238 12462 26290
rect 12514 26238 12526 26290
rect 15698 26238 15710 26290
rect 15762 26238 15774 26290
rect 16046 26226 16098 26238
rect 16382 26290 16434 26302
rect 23550 26290 23602 26302
rect 26350 26290 26402 26302
rect 28254 26290 28306 26302
rect 34638 26290 34690 26302
rect 39006 26290 39058 26302
rect 18274 26238 18286 26290
rect 18338 26238 18350 26290
rect 18610 26238 18622 26290
rect 18674 26238 18686 26290
rect 19730 26238 19742 26290
rect 19794 26238 19806 26290
rect 19954 26238 19966 26290
rect 20018 26238 20030 26290
rect 23090 26238 23102 26290
rect 23154 26238 23166 26290
rect 24098 26238 24110 26290
rect 24162 26238 24174 26290
rect 26114 26238 26126 26290
rect 26178 26238 26190 26290
rect 26674 26238 26686 26290
rect 26738 26238 26750 26290
rect 27682 26238 27694 26290
rect 27746 26238 27758 26290
rect 30706 26238 30718 26290
rect 30770 26238 30782 26290
rect 31154 26238 31166 26290
rect 31218 26238 31230 26290
rect 32050 26238 32062 26290
rect 32114 26238 32126 26290
rect 35186 26238 35198 26290
rect 35250 26238 35262 26290
rect 16382 26226 16434 26238
rect 23550 26226 23602 26238
rect 26350 26226 26402 26238
rect 28254 26226 28306 26238
rect 34638 26226 34690 26238
rect 39006 26226 39058 26238
rect 39566 26290 39618 26302
rect 44494 26290 44546 26302
rect 39890 26238 39902 26290
rect 39954 26238 39966 26290
rect 41010 26238 41022 26290
rect 41074 26238 41086 26290
rect 44146 26238 44158 26290
rect 44210 26238 44222 26290
rect 45378 26238 45390 26290
rect 45442 26238 45454 26290
rect 48850 26238 48862 26290
rect 48914 26238 48926 26290
rect 39566 26226 39618 26238
rect 44494 26226 44546 26238
rect 1934 26178 1986 26190
rect 23662 26178 23714 26190
rect 33406 26178 33458 26190
rect 9538 26126 9550 26178
rect 9602 26126 9614 26178
rect 12898 26126 12910 26178
rect 12962 26126 12974 26178
rect 15026 26126 15038 26178
rect 15090 26126 15102 26178
rect 18722 26126 18734 26178
rect 18786 26126 18798 26178
rect 20290 26126 20302 26178
rect 20354 26126 20366 26178
rect 22418 26126 22430 26178
rect 22482 26126 22494 26178
rect 29698 26126 29710 26178
rect 29762 26126 29774 26178
rect 30258 26126 30270 26178
rect 30322 26126 30334 26178
rect 1934 26114 1986 26126
rect 23662 26114 23714 26126
rect 33406 26114 33458 26126
rect 34750 26178 34802 26190
rect 34750 26114 34802 26126
rect 36766 26178 36818 26190
rect 36766 26114 36818 26126
rect 39790 26178 39842 26190
rect 41682 26126 41694 26178
rect 41746 26126 41758 26178
rect 43810 26126 43822 26178
rect 43874 26126 43886 26178
rect 46050 26126 46062 26178
rect 46114 26126 46126 26178
rect 48178 26126 48190 26178
rect 48242 26126 48254 26178
rect 39790 26114 39842 26126
rect 25666 26014 25678 26066
rect 25730 26014 25742 26066
rect 32946 26014 32958 26066
rect 33010 26063 33022 26066
rect 33394 26063 33406 26066
rect 33010 26017 33406 26063
rect 33010 26014 33022 26017
rect 33394 26014 33406 26017
rect 33458 26014 33470 26066
rect 1344 25898 58576 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 58576 25898
rect 1344 25812 58576 25846
rect 12126 25730 12178 25742
rect 12126 25666 12178 25678
rect 13582 25730 13634 25742
rect 13582 25666 13634 25678
rect 37102 25730 37154 25742
rect 37102 25666 37154 25678
rect 42030 25730 42082 25742
rect 42030 25666 42082 25678
rect 1934 25618 1986 25630
rect 14142 25618 14194 25630
rect 27918 25618 27970 25630
rect 8642 25566 8654 25618
rect 8706 25566 8718 25618
rect 17378 25566 17390 25618
rect 17442 25566 17454 25618
rect 19618 25566 19630 25618
rect 19682 25566 19694 25618
rect 21858 25566 21870 25618
rect 21922 25566 21934 25618
rect 1934 25554 1986 25566
rect 14142 25554 14194 25566
rect 27918 25554 27970 25566
rect 30046 25618 30098 25630
rect 31390 25618 31442 25630
rect 30482 25566 30494 25618
rect 30546 25566 30558 25618
rect 30046 25554 30098 25566
rect 31390 25554 31442 25566
rect 31950 25618 32002 25630
rect 40798 25618 40850 25630
rect 34290 25566 34302 25618
rect 34354 25566 34366 25618
rect 36418 25566 36430 25618
rect 36482 25566 36494 25618
rect 31950 25554 32002 25566
rect 40798 25554 40850 25566
rect 41470 25618 41522 25630
rect 41470 25554 41522 25566
rect 45054 25618 45106 25630
rect 45054 25554 45106 25566
rect 45502 25618 45554 25630
rect 45502 25554 45554 25566
rect 57934 25618 57986 25630
rect 57934 25554 57986 25566
rect 12798 25506 12850 25518
rect 4274 25454 4286 25506
rect 4338 25454 4350 25506
rect 11554 25454 11566 25506
rect 11618 25454 11630 25506
rect 12798 25442 12850 25454
rect 13694 25506 13746 25518
rect 13694 25442 13746 25454
rect 14926 25506 14978 25518
rect 14926 25442 14978 25454
rect 15262 25506 15314 25518
rect 18622 25506 18674 25518
rect 32510 25506 32562 25518
rect 38110 25506 38162 25518
rect 40014 25506 40066 25518
rect 17266 25454 17278 25506
rect 17330 25454 17342 25506
rect 18274 25454 18286 25506
rect 18338 25454 18350 25506
rect 18722 25454 18734 25506
rect 18786 25454 18798 25506
rect 19730 25454 19742 25506
rect 19794 25454 19806 25506
rect 26562 25454 26574 25506
rect 26626 25454 26638 25506
rect 29362 25454 29374 25506
rect 29426 25454 29438 25506
rect 32946 25454 32958 25506
rect 33010 25454 33022 25506
rect 33618 25454 33630 25506
rect 33682 25454 33694 25506
rect 38994 25454 39006 25506
rect 39058 25454 39070 25506
rect 15262 25442 15314 25454
rect 18622 25442 18674 25454
rect 32510 25442 32562 25454
rect 38110 25442 38162 25454
rect 40014 25442 40066 25454
rect 40350 25506 40402 25518
rect 41918 25506 41970 25518
rect 41346 25454 41358 25506
rect 41410 25454 41422 25506
rect 40350 25442 40402 25454
rect 41918 25442 41970 25454
rect 42366 25506 42418 25518
rect 42366 25442 42418 25454
rect 42702 25506 42754 25518
rect 46286 25506 46338 25518
rect 44258 25454 44270 25506
rect 44322 25454 44334 25506
rect 55570 25454 55582 25506
rect 55634 25454 55646 25506
rect 42702 25442 42754 25454
rect 46286 25442 46338 25454
rect 12238 25394 12290 25406
rect 10770 25342 10782 25394
rect 10834 25342 10846 25394
rect 12238 25330 12290 25342
rect 12462 25394 12514 25406
rect 12462 25330 12514 25342
rect 12686 25394 12738 25406
rect 12686 25330 12738 25342
rect 13582 25394 13634 25406
rect 20078 25394 20130 25406
rect 17154 25342 17166 25394
rect 17218 25342 17230 25394
rect 13582 25330 13634 25342
rect 20078 25330 20130 25342
rect 20190 25394 20242 25406
rect 37102 25394 37154 25406
rect 39454 25394 39506 25406
rect 28242 25342 28254 25394
rect 28306 25342 28318 25394
rect 32722 25342 32734 25394
rect 32786 25342 32798 25394
rect 20190 25330 20242 25342
rect 37102 25330 37154 25342
rect 37214 25338 37266 25350
rect 38770 25342 38782 25394
rect 38834 25342 38846 25394
rect 12126 25282 12178 25294
rect 12126 25218 12178 25230
rect 15150 25282 15202 25294
rect 15150 25218 15202 25230
rect 16606 25282 16658 25294
rect 16606 25218 16658 25230
rect 20414 25282 20466 25294
rect 27022 25282 27074 25294
rect 26562 25230 26574 25282
rect 26626 25279 26638 25282
rect 26786 25279 26798 25282
rect 26626 25233 26798 25279
rect 26626 25230 26638 25233
rect 26786 25230 26798 25233
rect 26850 25230 26862 25282
rect 20414 25218 20466 25230
rect 27022 25218 27074 25230
rect 28590 25282 28642 25294
rect 28590 25218 28642 25230
rect 29150 25282 29202 25294
rect 29150 25218 29202 25230
rect 30942 25282 30994 25294
rect 30942 25218 30994 25230
rect 31838 25282 31890 25294
rect 31838 25218 31890 25230
rect 32062 25282 32114 25294
rect 39454 25330 39506 25342
rect 39790 25394 39842 25406
rect 39790 25330 39842 25342
rect 41582 25394 41634 25406
rect 41582 25330 41634 25342
rect 42030 25394 42082 25406
rect 42030 25330 42082 25342
rect 42590 25394 42642 25406
rect 42590 25330 42642 25342
rect 43038 25394 43090 25406
rect 45838 25394 45890 25406
rect 43362 25342 43374 25394
rect 43426 25342 43438 25394
rect 44146 25342 44158 25394
rect 44210 25342 44222 25394
rect 43038 25330 43090 25342
rect 45838 25330 45890 25342
rect 37214 25274 37266 25286
rect 40238 25282 40290 25294
rect 37762 25230 37774 25282
rect 37826 25230 37838 25282
rect 32062 25218 32114 25230
rect 40238 25218 40290 25230
rect 41134 25282 41186 25294
rect 41134 25218 41186 25230
rect 1344 25114 58576 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 50558 25114
rect 50610 25062 50662 25114
rect 50714 25062 50766 25114
rect 50818 25062 58576 25114
rect 1344 25028 58576 25062
rect 4734 24946 4786 24958
rect 4734 24882 4786 24894
rect 13134 24946 13186 24958
rect 13134 24882 13186 24894
rect 23214 24946 23266 24958
rect 23214 24882 23266 24894
rect 23326 24946 23378 24958
rect 23326 24882 23378 24894
rect 24222 24946 24274 24958
rect 24222 24882 24274 24894
rect 24446 24946 24498 24958
rect 24446 24882 24498 24894
rect 24558 24946 24610 24958
rect 24558 24882 24610 24894
rect 25902 24946 25954 24958
rect 25902 24882 25954 24894
rect 26014 24946 26066 24958
rect 26014 24882 26066 24894
rect 30046 24946 30098 24958
rect 30046 24882 30098 24894
rect 33182 24946 33234 24958
rect 33182 24882 33234 24894
rect 33518 24946 33570 24958
rect 33518 24882 33570 24894
rect 38894 24946 38946 24958
rect 38894 24882 38946 24894
rect 41358 24946 41410 24958
rect 41358 24882 41410 24894
rect 41582 24946 41634 24958
rect 41582 24882 41634 24894
rect 44270 24946 44322 24958
rect 44270 24882 44322 24894
rect 47854 24946 47906 24958
rect 47854 24882 47906 24894
rect 18846 24834 18898 24846
rect 18846 24770 18898 24782
rect 18958 24834 19010 24846
rect 18958 24770 19010 24782
rect 20302 24834 20354 24846
rect 20302 24770 20354 24782
rect 20526 24834 20578 24846
rect 20526 24770 20578 24782
rect 20638 24834 20690 24846
rect 20638 24770 20690 24782
rect 21086 24834 21138 24846
rect 21086 24770 21138 24782
rect 22654 24834 22706 24846
rect 22654 24770 22706 24782
rect 22766 24834 22818 24846
rect 22766 24770 22818 24782
rect 26910 24834 26962 24846
rect 37550 24834 37602 24846
rect 41806 24834 41858 24846
rect 28018 24782 28030 24834
rect 28082 24782 28094 24834
rect 28802 24782 28814 24834
rect 28866 24782 28878 24834
rect 31714 24782 31726 24834
rect 31778 24782 31790 24834
rect 32050 24782 32062 24834
rect 32114 24782 32126 24834
rect 39218 24782 39230 24834
rect 39282 24782 39294 24834
rect 26910 24770 26962 24782
rect 37550 24770 37602 24782
rect 41806 24770 41858 24782
rect 43934 24834 43986 24846
rect 47518 24834 47570 24846
rect 46386 24782 46398 24834
rect 46450 24782 46462 24834
rect 43934 24770 43986 24782
rect 47518 24770 47570 24782
rect 15262 24722 15314 24734
rect 4274 24670 4286 24722
rect 4338 24670 4350 24722
rect 11890 24670 11902 24722
rect 11954 24670 11966 24722
rect 14578 24670 14590 24722
rect 14642 24670 14654 24722
rect 15262 24658 15314 24670
rect 15710 24722 15762 24734
rect 15710 24658 15762 24670
rect 18622 24722 18674 24734
rect 18622 24658 18674 24670
rect 19294 24722 19346 24734
rect 19294 24658 19346 24670
rect 19854 24722 19906 24734
rect 19854 24658 19906 24670
rect 21534 24722 21586 24734
rect 21534 24658 21586 24670
rect 22990 24722 23042 24734
rect 22990 24658 23042 24670
rect 23438 24722 23490 24734
rect 24670 24722 24722 24734
rect 23762 24670 23774 24722
rect 23826 24670 23838 24722
rect 23438 24658 23490 24670
rect 24670 24658 24722 24670
rect 25790 24722 25842 24734
rect 25790 24658 25842 24670
rect 26462 24722 26514 24734
rect 31838 24722 31890 24734
rect 33070 24722 33122 24734
rect 27122 24670 27134 24722
rect 27186 24670 27198 24722
rect 27346 24670 27358 24722
rect 27410 24670 27422 24722
rect 27906 24670 27918 24722
rect 27970 24670 27982 24722
rect 28578 24670 28590 24722
rect 28642 24670 28654 24722
rect 29474 24670 29486 24722
rect 29538 24670 29550 24722
rect 30706 24670 30718 24722
rect 30770 24670 30782 24722
rect 31266 24670 31278 24722
rect 31330 24670 31342 24722
rect 32386 24670 32398 24722
rect 32450 24670 32462 24722
rect 26462 24658 26514 24670
rect 31838 24658 31890 24670
rect 33070 24658 33122 24670
rect 33294 24722 33346 24734
rect 37662 24722 37714 24734
rect 41918 24722 41970 24734
rect 46958 24722 47010 24734
rect 34178 24670 34190 24722
rect 34242 24670 34254 24722
rect 40898 24670 40910 24722
rect 40962 24670 40974 24722
rect 41122 24670 41134 24722
rect 41186 24670 41198 24722
rect 44482 24670 44494 24722
rect 44546 24670 44558 24722
rect 46498 24670 46510 24722
rect 46562 24670 46574 24722
rect 53442 24670 53454 24722
rect 53506 24670 53518 24722
rect 33294 24658 33346 24670
rect 37662 24658 37714 24670
rect 41918 24658 41970 24670
rect 46958 24658 47010 24670
rect 1934 24610 1986 24622
rect 1934 24546 1986 24558
rect 5294 24610 5346 24622
rect 5294 24546 5346 24558
rect 10334 24610 10386 24622
rect 12574 24610 12626 24622
rect 25342 24610 25394 24622
rect 38110 24610 38162 24622
rect 12114 24558 12126 24610
rect 12178 24558 12190 24610
rect 14354 24558 14366 24610
rect 14418 24558 14430 24610
rect 34962 24558 34974 24610
rect 35026 24558 35038 24610
rect 37090 24558 37102 24610
rect 37154 24558 37166 24610
rect 10334 24546 10386 24558
rect 12574 24546 12626 24558
rect 25342 24546 25394 24558
rect 38110 24546 38162 24558
rect 40462 24610 40514 24622
rect 40462 24546 40514 24558
rect 42366 24610 42418 24622
rect 42366 24546 42418 24558
rect 10558 24498 10610 24510
rect 15598 24498 15650 24510
rect 10882 24446 10894 24498
rect 10946 24446 10958 24498
rect 10558 24434 10610 24446
rect 15598 24434 15650 24446
rect 27246 24498 27298 24510
rect 27246 24434 27298 24446
rect 37550 24498 37602 24510
rect 37550 24434 37602 24446
rect 41470 24498 41522 24510
rect 41470 24434 41522 24446
rect 42254 24498 42306 24510
rect 55346 24446 55358 24498
rect 55410 24446 55422 24498
rect 42254 24434 42306 24446
rect 1344 24330 58576 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 58576 24330
rect 1344 24244 58576 24278
rect 1934 24162 1986 24174
rect 1934 24098 1986 24110
rect 29710 24162 29762 24174
rect 29710 24098 29762 24110
rect 45726 24162 45778 24174
rect 45726 24098 45778 24110
rect 57934 24162 57986 24174
rect 57934 24098 57986 24110
rect 33854 24050 33906 24062
rect 4946 23998 4958 24050
rect 5010 23998 5022 24050
rect 10098 23998 10110 24050
rect 10162 23998 10174 24050
rect 15250 23998 15262 24050
rect 15314 23998 15326 24050
rect 16706 23998 16718 24050
rect 16770 23998 16782 24050
rect 18498 23998 18510 24050
rect 18562 23998 18574 24050
rect 20626 23998 20638 24050
rect 20690 23998 20702 24050
rect 21298 23998 21310 24050
rect 21362 23998 21374 24050
rect 23426 23998 23438 24050
rect 23490 23998 23502 24050
rect 33394 23998 33406 24050
rect 33458 23998 33470 24050
rect 33854 23986 33906 23998
rect 35646 24050 35698 24062
rect 35646 23986 35698 23998
rect 46846 24050 46898 24062
rect 46846 23986 46898 23998
rect 47294 24050 47346 24062
rect 47294 23986 47346 23998
rect 55358 24050 55410 24062
rect 55358 23986 55410 23998
rect 14030 23938 14082 23950
rect 24446 23938 24498 23950
rect 4274 23886 4286 23938
rect 4338 23886 4350 23938
rect 6402 23886 6414 23938
rect 6466 23886 6478 23938
rect 7858 23886 7870 23938
rect 7922 23886 7934 23938
rect 8306 23886 8318 23938
rect 8370 23886 8382 23938
rect 9986 23886 9998 23938
rect 10050 23886 10062 23938
rect 15138 23886 15150 23938
rect 15202 23886 15214 23938
rect 16818 23886 16830 23938
rect 16882 23886 16894 23938
rect 17826 23886 17838 23938
rect 17890 23886 17902 23938
rect 24098 23886 24110 23938
rect 24162 23886 24174 23938
rect 14030 23874 14082 23886
rect 24446 23874 24498 23886
rect 24782 23938 24834 23950
rect 24782 23874 24834 23886
rect 25118 23938 25170 23950
rect 25118 23874 25170 23886
rect 25454 23938 25506 23950
rect 33742 23938 33794 23950
rect 26338 23886 26350 23938
rect 26402 23886 26414 23938
rect 27234 23886 27246 23938
rect 27298 23886 27310 23938
rect 27794 23886 27806 23938
rect 27858 23886 27870 23938
rect 29138 23886 29150 23938
rect 29202 23886 29214 23938
rect 30034 23886 30046 23938
rect 30098 23886 30110 23938
rect 31602 23886 31614 23938
rect 31666 23886 31678 23938
rect 32162 23886 32174 23938
rect 32226 23886 32238 23938
rect 33058 23886 33070 23938
rect 33122 23886 33134 23938
rect 25454 23874 25506 23886
rect 33742 23874 33794 23886
rect 33966 23938 34018 23950
rect 33966 23874 34018 23886
rect 34526 23938 34578 23950
rect 34526 23874 34578 23886
rect 35086 23938 35138 23950
rect 35086 23874 35138 23886
rect 35534 23938 35586 23950
rect 35534 23874 35586 23886
rect 35758 23938 35810 23950
rect 35758 23874 35810 23886
rect 36206 23938 36258 23950
rect 36206 23874 36258 23886
rect 38558 23938 38610 23950
rect 45614 23938 45666 23950
rect 40226 23886 40238 23938
rect 40290 23886 40302 23938
rect 45154 23886 45166 23938
rect 45218 23886 45230 23938
rect 55570 23886 55582 23938
rect 55634 23886 55646 23938
rect 38558 23874 38610 23886
rect 45614 23874 45666 23886
rect 4622 23826 4674 23838
rect 4622 23762 4674 23774
rect 5630 23826 5682 23838
rect 5630 23762 5682 23774
rect 6638 23826 6690 23838
rect 6638 23762 6690 23774
rect 6750 23826 6802 23838
rect 6750 23762 6802 23774
rect 8542 23826 8594 23838
rect 8542 23762 8594 23774
rect 10670 23826 10722 23838
rect 10670 23762 10722 23774
rect 11006 23826 11058 23838
rect 11006 23762 11058 23774
rect 14254 23826 14306 23838
rect 14254 23762 14306 23774
rect 14366 23826 14418 23838
rect 14366 23762 14418 23774
rect 24670 23826 24722 23838
rect 24670 23762 24722 23774
rect 25678 23826 25730 23838
rect 34190 23826 34242 23838
rect 26114 23774 26126 23826
rect 26178 23774 26190 23826
rect 27010 23774 27022 23826
rect 27074 23774 27086 23826
rect 32610 23774 32622 23826
rect 32674 23774 32686 23826
rect 32946 23774 32958 23826
rect 33010 23774 33022 23826
rect 25678 23762 25730 23774
rect 34190 23762 34242 23774
rect 34974 23826 35026 23838
rect 44942 23826 44994 23838
rect 41234 23774 41246 23826
rect 41298 23774 41310 23826
rect 34974 23762 35026 23774
rect 44942 23762 44994 23774
rect 46398 23826 46450 23838
rect 46398 23762 46450 23774
rect 46622 23826 46674 23838
rect 46622 23762 46674 23774
rect 46958 23826 47010 23838
rect 46958 23762 47010 23774
rect 4846 23714 4898 23726
rect 4846 23650 4898 23662
rect 5070 23714 5122 23726
rect 5070 23650 5122 23662
rect 5742 23714 5794 23726
rect 5742 23650 5794 23662
rect 5966 23714 6018 23726
rect 11118 23714 11170 23726
rect 7186 23662 7198 23714
rect 7250 23662 7262 23714
rect 5966 23650 6018 23662
rect 11118 23650 11170 23662
rect 25342 23714 25394 23726
rect 25342 23650 25394 23662
rect 28366 23714 28418 23726
rect 28366 23650 28418 23662
rect 29374 23714 29426 23726
rect 29374 23650 29426 23662
rect 29598 23714 29650 23726
rect 30830 23714 30882 23726
rect 30258 23662 30270 23714
rect 30322 23662 30334 23714
rect 29598 23650 29650 23662
rect 30830 23650 30882 23662
rect 35198 23714 35250 23726
rect 35198 23650 35250 23662
rect 45726 23714 45778 23726
rect 45726 23650 45778 23662
rect 47406 23714 47458 23726
rect 47406 23650 47458 23662
rect 1344 23546 58576 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 50558 23546
rect 50610 23494 50662 23546
rect 50714 23494 50766 23546
rect 50818 23494 58576 23546
rect 1344 23460 58576 23494
rect 13806 23378 13858 23390
rect 13806 23314 13858 23326
rect 24222 23378 24274 23390
rect 24222 23314 24274 23326
rect 24782 23378 24834 23390
rect 24782 23314 24834 23326
rect 25230 23378 25282 23390
rect 31614 23378 31666 23390
rect 25554 23326 25566 23378
rect 25618 23326 25630 23378
rect 25230 23314 25282 23326
rect 31614 23314 31666 23326
rect 37662 23378 37714 23390
rect 37662 23314 37714 23326
rect 38558 23378 38610 23390
rect 38558 23314 38610 23326
rect 6974 23266 7026 23278
rect 16158 23266 16210 23278
rect 7858 23214 7870 23266
rect 7922 23214 7934 23266
rect 12002 23214 12014 23266
rect 12066 23214 12078 23266
rect 6974 23202 7026 23214
rect 16158 23202 16210 23214
rect 18062 23266 18114 23278
rect 24446 23266 24498 23278
rect 21634 23214 21646 23266
rect 21698 23214 21710 23266
rect 18062 23202 18114 23214
rect 24446 23202 24498 23214
rect 24558 23266 24610 23278
rect 32398 23266 32450 23278
rect 29810 23214 29822 23266
rect 29874 23214 29886 23266
rect 31938 23214 31950 23266
rect 32002 23214 32014 23266
rect 42018 23214 42030 23266
rect 42082 23214 42094 23266
rect 45378 23214 45390 23266
rect 45442 23214 45454 23266
rect 24558 23202 24610 23214
rect 32398 23202 32450 23214
rect 15262 23154 15314 23166
rect 17950 23154 18002 23166
rect 4274 23102 4286 23154
rect 4338 23102 4350 23154
rect 5170 23102 5182 23154
rect 5234 23102 5246 23154
rect 6178 23102 6190 23154
rect 6242 23102 6254 23154
rect 8306 23102 8318 23154
rect 8370 23102 8382 23154
rect 8978 23102 8990 23154
rect 9042 23102 9054 23154
rect 10770 23102 10782 23154
rect 10834 23102 10846 23154
rect 11778 23102 11790 23154
rect 11842 23102 11854 23154
rect 13458 23102 13470 23154
rect 13522 23102 13534 23154
rect 14242 23102 14254 23154
rect 14306 23102 14318 23154
rect 15474 23102 15486 23154
rect 15538 23102 15550 23154
rect 15262 23090 15314 23102
rect 17950 23090 18002 23102
rect 18286 23154 18338 23166
rect 18286 23090 18338 23102
rect 19182 23154 19234 23166
rect 22430 23154 22482 23166
rect 21522 23102 21534 23154
rect 21586 23102 21598 23154
rect 19182 23090 19234 23102
rect 22430 23090 22482 23102
rect 22766 23154 22818 23166
rect 22766 23090 22818 23102
rect 22990 23154 23042 23166
rect 38334 23154 38386 23166
rect 26786 23102 26798 23154
rect 26850 23102 26862 23154
rect 37874 23102 37886 23154
rect 37938 23102 37950 23154
rect 22990 23090 23042 23102
rect 38334 23090 38386 23102
rect 38670 23154 38722 23166
rect 39454 23154 39506 23166
rect 38994 23102 39006 23154
rect 39058 23102 39070 23154
rect 38670 23090 38722 23102
rect 39454 23090 39506 23102
rect 39790 23154 39842 23166
rect 47966 23154 48018 23166
rect 41234 23102 41246 23154
rect 41298 23102 41310 23154
rect 44594 23102 44606 23154
rect 44658 23102 44670 23154
rect 53442 23102 53454 23154
rect 53506 23102 53518 23154
rect 39790 23090 39842 23102
rect 47966 23090 48018 23102
rect 1934 23042 1986 23054
rect 18510 23042 18562 23054
rect 22654 23042 22706 23054
rect 4722 22990 4734 23042
rect 4786 22990 4798 23042
rect 8530 22990 8542 23042
rect 8594 22990 8606 23042
rect 10994 22990 11006 23042
rect 11058 22990 11070 23042
rect 22194 22990 22206 23042
rect 22258 22990 22270 23042
rect 1934 22978 1986 22990
rect 18510 22978 18562 22990
rect 22654 22978 22706 22990
rect 23662 23042 23714 23054
rect 23662 22978 23714 22990
rect 39678 23042 39730 23054
rect 44146 22990 44158 23042
rect 44210 22990 44222 23042
rect 47506 22990 47518 23042
rect 47570 22990 47582 23042
rect 39678 22978 39730 22990
rect 14254 22930 14306 22942
rect 11106 22878 11118 22930
rect 11170 22878 11182 22930
rect 14254 22866 14306 22878
rect 14590 22930 14642 22942
rect 14590 22866 14642 22878
rect 18622 22930 18674 22942
rect 18622 22866 18674 22878
rect 19294 22930 19346 22942
rect 38098 22878 38110 22930
rect 38162 22878 38174 22930
rect 39218 22878 39230 22930
rect 39282 22878 39294 22930
rect 55346 22878 55358 22930
rect 55410 22878 55422 22930
rect 19294 22866 19346 22878
rect 1344 22762 58576 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 58576 22762
rect 1344 22676 58576 22710
rect 3054 22594 3106 22606
rect 8990 22594 9042 22606
rect 3378 22542 3390 22594
rect 3442 22542 3454 22594
rect 3054 22530 3106 22542
rect 8990 22530 9042 22542
rect 12014 22594 12066 22606
rect 37102 22594 37154 22606
rect 22082 22542 22094 22594
rect 22146 22542 22158 22594
rect 12014 22530 12066 22542
rect 37102 22530 37154 22542
rect 37550 22594 37602 22606
rect 37550 22530 37602 22542
rect 38334 22594 38386 22606
rect 38334 22530 38386 22542
rect 39790 22594 39842 22606
rect 39790 22530 39842 22542
rect 57934 22594 57986 22606
rect 57934 22530 57986 22542
rect 8094 22482 8146 22494
rect 16606 22482 16658 22494
rect 4498 22430 4510 22482
rect 4562 22430 4574 22482
rect 4834 22430 4846 22482
rect 4898 22430 4910 22482
rect 5954 22430 5966 22482
rect 6018 22430 6030 22482
rect 9874 22430 9886 22482
rect 9938 22430 9950 22482
rect 12114 22430 12126 22482
rect 12178 22430 12190 22482
rect 13570 22430 13582 22482
rect 13634 22430 13646 22482
rect 15250 22430 15262 22482
rect 15314 22430 15326 22482
rect 15698 22430 15710 22482
rect 15762 22430 15774 22482
rect 8094 22418 8146 22430
rect 16606 22418 16658 22430
rect 19070 22482 19122 22494
rect 25678 22482 25730 22494
rect 24882 22430 24894 22482
rect 24946 22430 24958 22482
rect 19070 22418 19122 22430
rect 25678 22418 25730 22430
rect 29374 22482 29426 22494
rect 36990 22482 37042 22494
rect 33506 22430 33518 22482
rect 33570 22430 33582 22482
rect 29374 22418 29426 22430
rect 36990 22418 37042 22430
rect 42590 22482 42642 22494
rect 42590 22418 42642 22430
rect 43038 22482 43090 22494
rect 55022 22482 55074 22494
rect 47618 22430 47630 22482
rect 47682 22430 47694 22482
rect 49746 22430 49758 22482
rect 49810 22430 49822 22482
rect 43038 22418 43090 22430
rect 55022 22418 55074 22430
rect 2830 22370 2882 22382
rect 8654 22370 8706 22382
rect 2258 22318 2270 22370
rect 2322 22318 2334 22370
rect 4050 22318 4062 22370
rect 4114 22318 4126 22370
rect 4946 22318 4958 22370
rect 5010 22318 5022 22370
rect 7410 22318 7422 22370
rect 7474 22318 7486 22370
rect 8418 22318 8430 22370
rect 8482 22318 8494 22370
rect 2830 22306 2882 22318
rect 8654 22306 8706 22318
rect 8878 22370 8930 22382
rect 8878 22306 8930 22318
rect 11342 22370 11394 22382
rect 14478 22370 14530 22382
rect 18174 22370 18226 22382
rect 21422 22370 21474 22382
rect 23438 22370 23490 22382
rect 37214 22370 37266 22382
rect 11554 22318 11566 22370
rect 11618 22318 11630 22370
rect 12562 22318 12574 22370
rect 12626 22318 12638 22370
rect 14018 22318 14030 22370
rect 14082 22318 14094 22370
rect 15922 22318 15934 22370
rect 15986 22318 15998 22370
rect 18386 22318 18398 22370
rect 18450 22318 18462 22370
rect 21634 22318 21646 22370
rect 21698 22318 21710 22370
rect 23090 22318 23102 22370
rect 23154 22318 23166 22370
rect 24098 22318 24110 22370
rect 24162 22318 24174 22370
rect 26786 22318 26798 22370
rect 26850 22318 26862 22370
rect 27234 22318 27246 22370
rect 27298 22318 27310 22370
rect 28242 22318 28254 22370
rect 28306 22318 28318 22370
rect 29586 22318 29598 22370
rect 29650 22318 29662 22370
rect 35410 22318 35422 22370
rect 35474 22318 35486 22370
rect 11342 22306 11394 22318
rect 14478 22306 14530 22318
rect 18174 22306 18226 22318
rect 21422 22306 21474 22318
rect 23438 22306 23490 22318
rect 37214 22306 37266 22318
rect 37774 22370 37826 22382
rect 37774 22306 37826 22318
rect 39230 22370 39282 22382
rect 39230 22306 39282 22318
rect 39566 22370 39618 22382
rect 39566 22306 39618 22318
rect 40238 22370 40290 22382
rect 40238 22306 40290 22318
rect 40910 22370 40962 22382
rect 40910 22306 40962 22318
rect 42142 22370 42194 22382
rect 42142 22306 42194 22318
rect 42478 22370 42530 22382
rect 42478 22306 42530 22318
rect 42702 22370 42754 22382
rect 46062 22370 46114 22382
rect 44034 22318 44046 22370
rect 44098 22318 44110 22370
rect 42702 22306 42754 22318
rect 46062 22306 46114 22318
rect 46398 22370 46450 22382
rect 46834 22318 46846 22370
rect 46898 22318 46910 22370
rect 52658 22318 52670 22370
rect 52722 22318 52734 22370
rect 55570 22318 55582 22370
rect 55634 22318 55646 22370
rect 46398 22306 46450 22318
rect 9550 22258 9602 22270
rect 2482 22206 2494 22258
rect 2546 22206 2558 22258
rect 6514 22206 6526 22258
rect 6578 22206 6590 22258
rect 9550 22194 9602 22206
rect 11006 22258 11058 22270
rect 11006 22194 11058 22206
rect 14926 22258 14978 22270
rect 14926 22194 14978 22206
rect 17726 22258 17778 22270
rect 17726 22194 17778 22206
rect 25342 22258 25394 22270
rect 25342 22194 25394 22206
rect 25790 22258 25842 22270
rect 35982 22258 36034 22270
rect 26450 22206 26462 22258
rect 26514 22206 26526 22258
rect 27458 22206 27470 22258
rect 27522 22206 27534 22258
rect 25790 22194 25842 22206
rect 35982 22194 36034 22206
rect 36094 22258 36146 22270
rect 36094 22194 36146 22206
rect 38222 22258 38274 22270
rect 38222 22194 38274 22206
rect 38894 22258 38946 22270
rect 38894 22194 38946 22206
rect 40350 22258 40402 22270
rect 40350 22194 40402 22206
rect 40574 22258 40626 22270
rect 40574 22194 40626 22206
rect 41246 22258 41298 22270
rect 41246 22194 41298 22206
rect 41470 22258 41522 22270
rect 41470 22194 41522 22206
rect 41806 22258 41858 22270
rect 45502 22258 45554 22270
rect 45154 22206 45166 22258
rect 45218 22206 45230 22258
rect 41806 22194 41858 22206
rect 45502 22194 45554 22206
rect 46286 22258 46338 22270
rect 46286 22194 46338 22206
rect 9774 22146 9826 22158
rect 9774 22082 9826 22094
rect 11118 22146 11170 22158
rect 11118 22082 11170 22094
rect 15150 22146 15202 22158
rect 15150 22082 15202 22094
rect 17390 22146 17442 22158
rect 17390 22082 17442 22094
rect 17614 22146 17666 22158
rect 17614 22082 17666 22094
rect 25566 22146 25618 22158
rect 25566 22082 25618 22094
rect 28702 22146 28754 22158
rect 35758 22146 35810 22158
rect 35186 22094 35198 22146
rect 35250 22094 35262 22146
rect 28702 22082 28754 22094
rect 35758 22082 35810 22094
rect 38334 22146 38386 22158
rect 38334 22082 38386 22094
rect 39006 22146 39058 22158
rect 39006 22082 39058 22094
rect 39454 22146 39506 22158
rect 39454 22082 39506 22094
rect 40798 22146 40850 22158
rect 40798 22082 40850 22094
rect 41694 22146 41746 22158
rect 41694 22082 41746 22094
rect 43598 22146 43650 22158
rect 43598 22082 43650 22094
rect 44270 22146 44322 22158
rect 44270 22082 44322 22094
rect 44830 22146 44882 22158
rect 44830 22082 44882 22094
rect 45838 22146 45890 22158
rect 45838 22082 45890 22094
rect 1344 21978 58576 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 50558 21978
rect 50610 21926 50662 21978
rect 50714 21926 50766 21978
rect 50818 21926 58576 21978
rect 1344 21892 58576 21926
rect 3950 21810 4002 21822
rect 3950 21746 4002 21758
rect 4734 21810 4786 21822
rect 4734 21746 4786 21758
rect 5070 21810 5122 21822
rect 10222 21810 10274 21822
rect 23886 21810 23938 21822
rect 8082 21758 8094 21810
rect 8146 21758 8158 21810
rect 22530 21758 22542 21810
rect 22594 21758 22606 21810
rect 5070 21746 5122 21758
rect 10222 21746 10274 21758
rect 23886 21746 23938 21758
rect 24334 21810 24386 21822
rect 40002 21758 40014 21810
rect 40066 21758 40078 21810
rect 24334 21746 24386 21758
rect 2270 21698 2322 21710
rect 2270 21634 2322 21646
rect 4062 21698 4114 21710
rect 11230 21698 11282 21710
rect 7186 21646 7198 21698
rect 7250 21646 7262 21698
rect 4062 21634 4114 21646
rect 11230 21634 11282 21646
rect 13582 21698 13634 21710
rect 13582 21634 13634 21646
rect 14590 21698 14642 21710
rect 14590 21634 14642 21646
rect 16494 21698 16546 21710
rect 23102 21698 23154 21710
rect 19506 21646 19518 21698
rect 19570 21646 19582 21698
rect 20738 21646 20750 21698
rect 20802 21646 20814 21698
rect 22418 21646 22430 21698
rect 22482 21646 22494 21698
rect 16494 21634 16546 21646
rect 23102 21634 23154 21646
rect 32062 21698 32114 21710
rect 32062 21634 32114 21646
rect 32510 21698 32562 21710
rect 39678 21698 39730 21710
rect 37090 21646 37102 21698
rect 37154 21646 37166 21698
rect 32510 21634 32562 21646
rect 39678 21634 39730 21646
rect 2718 21586 2770 21598
rect 2718 21522 2770 21534
rect 3166 21586 3218 21598
rect 3166 21522 3218 21534
rect 3614 21586 3666 21598
rect 3614 21522 3666 21534
rect 4286 21586 4338 21598
rect 4286 21522 4338 21534
rect 4622 21586 4674 21598
rect 4622 21522 4674 21534
rect 4846 21586 4898 21598
rect 9886 21586 9938 21598
rect 14702 21586 14754 21598
rect 15598 21586 15650 21598
rect 7074 21534 7086 21586
rect 7138 21534 7150 21586
rect 7970 21534 7982 21586
rect 8034 21534 8046 21586
rect 10322 21534 10334 21586
rect 10386 21534 10398 21586
rect 12338 21534 12350 21586
rect 12402 21534 12414 21586
rect 15138 21534 15150 21586
rect 15202 21534 15214 21586
rect 15810 21534 15822 21586
rect 15874 21534 15886 21586
rect 17602 21534 17614 21586
rect 17666 21534 17678 21586
rect 19170 21534 19182 21586
rect 19234 21534 19246 21586
rect 21298 21534 21310 21586
rect 21362 21534 21374 21586
rect 25330 21534 25342 21586
rect 25394 21534 25406 21586
rect 28802 21534 28814 21586
rect 28866 21534 28878 21586
rect 33058 21534 33070 21586
rect 33122 21534 33134 21586
rect 36306 21534 36318 21586
rect 36370 21534 36382 21586
rect 40226 21534 40238 21586
rect 40290 21534 40302 21586
rect 40898 21534 40910 21586
rect 40962 21534 40974 21586
rect 53442 21534 53454 21586
rect 53506 21534 53518 21586
rect 4846 21522 4898 21534
rect 9886 21522 9938 21534
rect 14702 21522 14754 21534
rect 15598 21522 15650 21534
rect 2942 21474 2994 21486
rect 23214 21474 23266 21486
rect 12450 21422 12462 21474
rect 12514 21422 12526 21474
rect 17714 21422 17726 21474
rect 17778 21422 17790 21474
rect 2942 21410 2994 21422
rect 23214 21410 23266 21422
rect 24670 21474 24722 21486
rect 46622 21474 46674 21486
rect 26002 21422 26014 21474
rect 26066 21422 26078 21474
rect 28130 21422 28142 21474
rect 28194 21422 28206 21474
rect 29474 21422 29486 21474
rect 29538 21422 29550 21474
rect 31602 21422 31614 21474
rect 31666 21422 31678 21474
rect 33842 21422 33854 21474
rect 33906 21422 33918 21474
rect 35970 21422 35982 21474
rect 36034 21422 36046 21474
rect 39218 21422 39230 21474
rect 39282 21422 39294 21474
rect 43698 21422 43710 21474
rect 43762 21422 43774 21474
rect 24670 21410 24722 21422
rect 46622 21410 46674 21422
rect 10110 21362 10162 21374
rect 10110 21298 10162 21310
rect 11006 21362 11058 21374
rect 11006 21298 11058 21310
rect 11342 21362 11394 21374
rect 11342 21298 11394 21310
rect 14926 21362 14978 21374
rect 14926 21298 14978 21310
rect 23326 21362 23378 21374
rect 55346 21310 55358 21362
rect 55410 21310 55422 21362
rect 23326 21298 23378 21310
rect 1344 21194 58576 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 58576 21194
rect 1344 21108 58576 21142
rect 3390 21026 3442 21038
rect 16158 21026 16210 21038
rect 4946 20974 4958 21026
rect 5010 20974 5022 21026
rect 12338 20974 12350 21026
rect 12402 20974 12414 21026
rect 3390 20962 3442 20974
rect 16158 20962 16210 20974
rect 17502 21026 17554 21038
rect 17502 20962 17554 20974
rect 19182 21026 19234 21038
rect 19182 20962 19234 20974
rect 27022 21026 27074 21038
rect 27022 20962 27074 20974
rect 28142 21026 28194 21038
rect 28142 20962 28194 20974
rect 28478 21026 28530 21038
rect 28478 20962 28530 20974
rect 30046 21026 30098 21038
rect 30046 20962 30098 20974
rect 33518 21026 33570 21038
rect 33518 20962 33570 20974
rect 34078 21026 34130 21038
rect 43822 21026 43874 21038
rect 37538 20974 37550 21026
rect 37602 20974 37614 21026
rect 34078 20962 34130 20974
rect 43822 20962 43874 20974
rect 44158 21026 44210 21038
rect 44158 20962 44210 20974
rect 57934 21026 57986 21038
rect 57934 20962 57986 20974
rect 3166 20914 3218 20926
rect 3166 20850 3218 20862
rect 6750 20914 6802 20926
rect 13806 20914 13858 20926
rect 15262 20914 15314 20926
rect 8754 20862 8766 20914
rect 8818 20862 8830 20914
rect 12226 20862 12238 20914
rect 12290 20862 12302 20914
rect 14354 20862 14366 20914
rect 14418 20862 14430 20914
rect 6750 20850 6802 20862
rect 13806 20850 13858 20862
rect 15262 20850 15314 20862
rect 32062 20914 32114 20926
rect 35982 20914 36034 20926
rect 33842 20862 33854 20914
rect 33906 20862 33918 20914
rect 32062 20850 32114 20862
rect 35982 20850 36034 20862
rect 36990 20914 37042 20926
rect 36990 20850 37042 20862
rect 38334 20914 38386 20926
rect 45838 20914 45890 20926
rect 39554 20862 39566 20914
rect 39618 20862 39630 20914
rect 41682 20862 41694 20914
rect 41746 20862 41758 20914
rect 45266 20862 45278 20914
rect 45330 20862 45342 20914
rect 49746 20862 49758 20914
rect 49810 20862 49822 20914
rect 38334 20850 38386 20862
rect 45838 20850 45890 20862
rect 3614 20802 3666 20814
rect 3614 20738 3666 20750
rect 4062 20802 4114 20814
rect 4062 20738 4114 20750
rect 4398 20802 4450 20814
rect 4398 20738 4450 20750
rect 4622 20802 4674 20814
rect 6638 20802 6690 20814
rect 6290 20750 6302 20802
rect 6354 20750 6366 20802
rect 4622 20738 4674 20750
rect 6638 20738 6690 20750
rect 7982 20802 8034 20814
rect 9886 20802 9938 20814
rect 10670 20802 10722 20814
rect 15822 20802 15874 20814
rect 8866 20750 8878 20802
rect 8930 20750 8942 20802
rect 10098 20750 10110 20802
rect 10162 20750 10174 20802
rect 11106 20750 11118 20802
rect 11170 20750 11182 20802
rect 11554 20750 11566 20802
rect 11618 20750 11630 20802
rect 12450 20750 12462 20802
rect 12514 20750 12526 20802
rect 13570 20750 13582 20802
rect 13634 20750 13646 20802
rect 14578 20750 14590 20802
rect 14642 20750 14654 20802
rect 15586 20750 15598 20802
rect 15650 20750 15662 20802
rect 7982 20738 8034 20750
rect 9886 20738 9938 20750
rect 10670 20738 10722 20750
rect 15822 20738 15874 20750
rect 16046 20802 16098 20814
rect 16046 20738 16098 20750
rect 17166 20802 17218 20814
rect 17166 20738 17218 20750
rect 17390 20802 17442 20814
rect 27246 20802 27298 20814
rect 18498 20750 18510 20802
rect 18562 20750 18574 20802
rect 22418 20750 22430 20802
rect 22482 20750 22494 20802
rect 23986 20750 23998 20802
rect 24050 20750 24062 20802
rect 26002 20750 26014 20802
rect 26066 20750 26078 20802
rect 17390 20738 17442 20750
rect 27246 20738 27298 20750
rect 29822 20802 29874 20814
rect 29822 20738 29874 20750
rect 30382 20802 30434 20814
rect 30382 20738 30434 20750
rect 33294 20802 33346 20814
rect 33294 20738 33346 20750
rect 33966 20802 34018 20814
rect 34862 20802 34914 20814
rect 35758 20802 35810 20814
rect 34402 20750 34414 20802
rect 34466 20750 34478 20802
rect 35410 20750 35422 20802
rect 35474 20750 35486 20802
rect 33966 20738 34018 20750
rect 34862 20738 34914 20750
rect 35758 20738 35810 20750
rect 37214 20802 37266 20814
rect 37214 20738 37266 20750
rect 37886 20802 37938 20814
rect 42590 20802 42642 20814
rect 44830 20802 44882 20814
rect 38770 20750 38782 20802
rect 38834 20750 38846 20802
rect 43138 20750 43150 20802
rect 43202 20750 43214 20802
rect 46834 20750 46846 20802
rect 46898 20750 46910 20802
rect 55570 20750 55582 20802
rect 55634 20750 55646 20802
rect 37886 20738 37938 20750
rect 42590 20738 42642 20750
rect 44830 20738 44882 20750
rect 10222 20690 10274 20702
rect 10222 20626 10274 20638
rect 13918 20690 13970 20702
rect 13918 20626 13970 20638
rect 16830 20690 16882 20702
rect 16830 20626 16882 20638
rect 19070 20690 19122 20702
rect 19070 20626 19122 20638
rect 21198 20690 21250 20702
rect 21198 20626 21250 20638
rect 21422 20690 21474 20702
rect 21422 20626 21474 20638
rect 21534 20690 21586 20702
rect 27582 20690 27634 20702
rect 22194 20638 22206 20690
rect 22258 20638 22270 20690
rect 24098 20638 24110 20690
rect 24162 20638 24174 20690
rect 25442 20638 25454 20690
rect 25506 20638 25518 20690
rect 21534 20626 21586 20638
rect 27582 20626 27634 20638
rect 27806 20690 27858 20702
rect 27806 20626 27858 20638
rect 29038 20690 29090 20702
rect 29038 20626 29090 20638
rect 29374 20690 29426 20702
rect 29374 20626 29426 20638
rect 30606 20690 30658 20702
rect 30606 20626 30658 20638
rect 30830 20690 30882 20702
rect 30830 20626 30882 20638
rect 31166 20690 31218 20702
rect 31166 20626 31218 20638
rect 38110 20690 38162 20702
rect 38110 20626 38162 20638
rect 38446 20690 38498 20702
rect 38446 20626 38498 20638
rect 42030 20690 42082 20702
rect 55358 20690 55410 20702
rect 43026 20638 43038 20690
rect 43090 20638 43102 20690
rect 47618 20638 47630 20690
rect 47682 20638 47694 20690
rect 42030 20626 42082 20638
rect 55358 20626 55410 20638
rect 16942 20578 16994 20590
rect 16942 20514 16994 20526
rect 17502 20578 17554 20590
rect 19182 20578 19234 20590
rect 18722 20526 18734 20578
rect 18786 20526 18798 20578
rect 17502 20514 17554 20526
rect 19182 20514 19234 20526
rect 26910 20578 26962 20590
rect 26910 20514 26962 20526
rect 28254 20578 28306 20590
rect 28254 20514 28306 20526
rect 29262 20578 29314 20590
rect 29262 20514 29314 20526
rect 29710 20578 29762 20590
rect 29710 20514 29762 20526
rect 31054 20578 31106 20590
rect 31054 20514 31106 20526
rect 31614 20578 31666 20590
rect 31614 20514 31666 20526
rect 34638 20578 34690 20590
rect 34638 20514 34690 20526
rect 34750 20578 34802 20590
rect 34750 20514 34802 20526
rect 34974 20578 35026 20590
rect 34974 20514 35026 20526
rect 36542 20578 36594 20590
rect 36542 20514 36594 20526
rect 46510 20578 46562 20590
rect 46510 20514 46562 20526
rect 1344 20410 58576 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 50558 20410
rect 50610 20358 50662 20410
rect 50714 20358 50766 20410
rect 50818 20358 58576 20410
rect 1344 20324 58576 20358
rect 14590 20242 14642 20254
rect 12450 20190 12462 20242
rect 12514 20190 12526 20242
rect 14590 20178 14642 20190
rect 25902 20242 25954 20254
rect 25902 20178 25954 20190
rect 40462 20242 40514 20254
rect 40462 20178 40514 20190
rect 47630 20242 47682 20254
rect 47630 20178 47682 20190
rect 5182 20130 5234 20142
rect 5182 20066 5234 20078
rect 5406 20130 5458 20142
rect 5406 20066 5458 20078
rect 6526 20130 6578 20142
rect 6526 20066 6578 20078
rect 8206 20130 8258 20142
rect 14254 20130 14306 20142
rect 11106 20078 11118 20130
rect 11170 20078 11182 20130
rect 8206 20066 8258 20078
rect 14254 20066 14306 20078
rect 14478 20130 14530 20142
rect 14478 20066 14530 20078
rect 15262 20130 15314 20142
rect 15262 20066 15314 20078
rect 15374 20130 15426 20142
rect 15374 20066 15426 20078
rect 17502 20130 17554 20142
rect 17502 20066 17554 20078
rect 20414 20130 20466 20142
rect 25678 20130 25730 20142
rect 22530 20078 22542 20130
rect 22594 20078 22606 20130
rect 24546 20078 24558 20130
rect 24610 20078 24622 20130
rect 20414 20066 20466 20078
rect 25678 20066 25730 20078
rect 26238 20130 26290 20142
rect 26238 20066 26290 20078
rect 27694 20130 27746 20142
rect 27694 20066 27746 20078
rect 28478 20130 28530 20142
rect 28478 20066 28530 20078
rect 29710 20130 29762 20142
rect 29710 20066 29762 20078
rect 31726 20130 31778 20142
rect 39454 20130 39506 20142
rect 34290 20078 34302 20130
rect 34354 20078 34366 20130
rect 31726 20066 31778 20078
rect 39454 20066 39506 20078
rect 40910 20130 40962 20142
rect 40910 20066 40962 20078
rect 42030 20130 42082 20142
rect 47070 20130 47122 20142
rect 45826 20078 45838 20130
rect 45890 20078 45902 20130
rect 48962 20078 48974 20130
rect 49026 20078 49038 20130
rect 42030 20066 42082 20078
rect 47070 20066 47122 20078
rect 4734 20018 4786 20030
rect 2706 19966 2718 20018
rect 2770 19966 2782 20018
rect 3938 19966 3950 20018
rect 4002 19966 4014 20018
rect 4734 19954 4786 19966
rect 5518 20018 5570 20030
rect 14702 20018 14754 20030
rect 17614 20018 17666 20030
rect 7746 19966 7758 20018
rect 7810 19966 7822 20018
rect 11330 19966 11342 20018
rect 11394 19966 11406 20018
rect 12002 19966 12014 20018
rect 12066 19966 12078 20018
rect 14914 19966 14926 20018
rect 14978 19966 14990 20018
rect 5518 19954 5570 19966
rect 14702 19954 14754 19966
rect 17614 19954 17666 19966
rect 20190 20018 20242 20030
rect 20190 19954 20242 19966
rect 20526 20018 20578 20030
rect 22766 20018 22818 20030
rect 26014 20018 26066 20030
rect 29934 20018 29986 20030
rect 21298 19966 21310 20018
rect 21362 19966 21374 20018
rect 23650 19966 23662 20018
rect 23714 19966 23726 20018
rect 27234 19966 27246 20018
rect 27298 19966 27310 20018
rect 29026 19966 29038 20018
rect 29090 19966 29102 20018
rect 20526 19954 20578 19966
rect 22766 19954 22818 19966
rect 26014 19954 26066 19966
rect 29934 19954 29986 19966
rect 30382 20018 30434 20030
rect 30382 19954 30434 19966
rect 30606 20018 30658 20030
rect 30606 19954 30658 19966
rect 32062 20018 32114 20030
rect 32062 19954 32114 19966
rect 33182 20018 33234 20030
rect 39902 20018 39954 20030
rect 34178 19966 34190 20018
rect 34242 19966 34254 20018
rect 35634 19966 35646 20018
rect 35698 19966 35710 20018
rect 33182 19954 33234 19966
rect 39902 19954 39954 19966
rect 41246 20018 41298 20030
rect 47966 20018 48018 20030
rect 49982 20018 50034 20030
rect 46498 19966 46510 20018
rect 46562 19966 46574 20018
rect 48850 19966 48862 20018
rect 48914 19966 48926 20018
rect 53666 19966 53678 20018
rect 53730 19966 53742 20018
rect 41246 19954 41298 19966
rect 47966 19954 48018 19966
rect 49982 19954 50034 19966
rect 13246 19906 13298 19918
rect 2818 19854 2830 19906
rect 2882 19854 2894 19906
rect 6402 19854 6414 19906
rect 6466 19854 6478 19906
rect 7410 19854 7422 19906
rect 7474 19854 7486 19906
rect 13246 19842 13298 19854
rect 15934 19906 15986 19918
rect 23214 19906 23266 19918
rect 30494 19906 30546 19918
rect 21522 19854 21534 19906
rect 21586 19854 21598 19906
rect 27010 19854 27022 19906
rect 27074 19854 27086 19906
rect 28802 19854 28814 19906
rect 28866 19854 28878 19906
rect 15934 19842 15986 19854
rect 23214 19842 23266 19854
rect 30494 19842 30546 19854
rect 35198 19906 35250 19918
rect 38894 19906 38946 19918
rect 36306 19854 36318 19906
rect 36370 19854 36382 19906
rect 38434 19854 38446 19906
rect 38498 19854 38510 19906
rect 35198 19842 35250 19854
rect 38894 19842 38946 19854
rect 42926 19906 42978 19918
rect 43698 19854 43710 19906
rect 43762 19854 43774 19906
rect 42926 19842 42978 19854
rect 6750 19794 6802 19806
rect 6750 19730 6802 19742
rect 15374 19794 15426 19806
rect 15374 19730 15426 19742
rect 17502 19794 17554 19806
rect 33518 19794 33570 19806
rect 24098 19742 24110 19794
rect 24162 19742 24174 19794
rect 17502 19730 17554 19742
rect 33518 19730 33570 19742
rect 49646 19794 49698 19806
rect 55346 19742 55358 19794
rect 55410 19742 55422 19794
rect 49646 19730 49698 19742
rect 1344 19626 58576 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 58576 19626
rect 1344 19540 58576 19574
rect 8318 19458 8370 19470
rect 12126 19458 12178 19470
rect 2482 19406 2494 19458
rect 2546 19406 2558 19458
rect 6626 19406 6638 19458
rect 6690 19406 6702 19458
rect 8642 19406 8654 19458
rect 8706 19455 8718 19458
rect 8978 19455 8990 19458
rect 8706 19409 8990 19455
rect 8706 19406 8718 19409
rect 8978 19406 8990 19409
rect 9042 19406 9054 19458
rect 8318 19394 8370 19406
rect 12126 19394 12178 19406
rect 22766 19458 22818 19470
rect 22766 19394 22818 19406
rect 25790 19458 25842 19470
rect 25790 19394 25842 19406
rect 57934 19458 57986 19470
rect 57934 19394 57986 19406
rect 8990 19346 9042 19358
rect 3602 19294 3614 19346
rect 3666 19294 3678 19346
rect 8990 19282 9042 19294
rect 19294 19346 19346 19358
rect 19294 19282 19346 19294
rect 21310 19346 21362 19358
rect 21310 19282 21362 19294
rect 23438 19346 23490 19358
rect 23438 19282 23490 19294
rect 25454 19346 25506 19358
rect 38782 19346 38834 19358
rect 42814 19346 42866 19358
rect 29138 19294 29150 19346
rect 29202 19294 29214 19346
rect 31266 19294 31278 19346
rect 31330 19294 31342 19346
rect 33394 19294 33406 19346
rect 33458 19294 33470 19346
rect 40226 19294 40238 19346
rect 40290 19294 40302 19346
rect 42354 19294 42366 19346
rect 42418 19294 42430 19346
rect 25454 19282 25506 19294
rect 38782 19282 38834 19294
rect 42814 19282 42866 19294
rect 44270 19346 44322 19358
rect 53230 19346 53282 19358
rect 47730 19294 47742 19346
rect 47794 19294 47806 19346
rect 44270 19282 44322 19294
rect 53230 19282 53282 19294
rect 2830 19234 2882 19246
rect 2830 19170 2882 19182
rect 3054 19234 3106 19246
rect 4174 19234 4226 19246
rect 3714 19182 3726 19234
rect 3778 19182 3790 19234
rect 3054 19170 3106 19182
rect 4174 19170 4226 19182
rect 4510 19234 4562 19246
rect 4510 19170 4562 19182
rect 6974 19234 7026 19246
rect 6974 19170 7026 19182
rect 7198 19234 7250 19246
rect 7198 19170 7250 19182
rect 9662 19234 9714 19246
rect 12574 19234 12626 19246
rect 17502 19234 17554 19246
rect 19406 19234 19458 19246
rect 21422 19234 21474 19246
rect 28142 19234 28194 19246
rect 10658 19182 10670 19234
rect 10722 19182 10734 19234
rect 11330 19182 11342 19234
rect 11394 19182 11406 19234
rect 11554 19182 11566 19234
rect 11618 19182 11630 19234
rect 16930 19182 16942 19234
rect 16994 19182 17006 19234
rect 18162 19182 18174 19234
rect 18226 19182 18238 19234
rect 19730 19182 19742 19234
rect 19794 19182 19806 19234
rect 21746 19182 21758 19234
rect 21810 19182 21822 19234
rect 26114 19182 26126 19234
rect 26178 19182 26190 19234
rect 27010 19182 27022 19234
rect 27074 19182 27086 19234
rect 9662 19170 9714 19182
rect 12574 19170 12626 19182
rect 17502 19170 17554 19182
rect 19406 19170 19458 19182
rect 21422 19170 21474 19182
rect 28142 19170 28194 19182
rect 28254 19234 28306 19246
rect 37438 19234 37490 19246
rect 30482 19182 30494 19234
rect 30546 19182 30558 19234
rect 38210 19182 38222 19234
rect 38274 19182 38286 19234
rect 39442 19182 39454 19234
rect 39506 19182 39518 19234
rect 44818 19182 44830 19234
rect 44882 19182 44894 19234
rect 55570 19182 55582 19234
rect 55634 19182 55646 19234
rect 28254 19170 28306 19182
rect 37438 19170 37490 19182
rect 1710 19122 1762 19134
rect 1710 19058 1762 19070
rect 3390 19122 3442 19134
rect 3390 19058 3442 19070
rect 4398 19122 4450 19134
rect 4398 19058 4450 19070
rect 5630 19122 5682 19134
rect 5630 19058 5682 19070
rect 8430 19122 8482 19134
rect 8430 19058 8482 19070
rect 9998 19122 10050 19134
rect 12238 19122 12290 19134
rect 11666 19070 11678 19122
rect 11730 19070 11742 19122
rect 9998 19058 10050 19070
rect 12238 19058 12290 19070
rect 12686 19122 12738 19134
rect 22878 19122 22930 19134
rect 25902 19122 25954 19134
rect 28478 19122 28530 19134
rect 16258 19070 16270 19122
rect 16322 19070 16334 19122
rect 18722 19070 18734 19122
rect 18786 19070 18798 19122
rect 23538 19070 23550 19122
rect 23602 19070 23614 19122
rect 25218 19070 25230 19122
rect 25282 19070 25294 19122
rect 27234 19070 27246 19122
rect 27298 19070 27310 19122
rect 27682 19070 27694 19122
rect 27746 19070 27758 19122
rect 12686 19058 12738 19070
rect 22878 19058 22930 19070
rect 25902 19058 25954 19070
rect 28478 19058 28530 19070
rect 28590 19122 28642 19134
rect 29598 19122 29650 19134
rect 29474 19070 29486 19122
rect 29538 19070 29550 19122
rect 28590 19058 28642 19070
rect 29598 19058 29650 19070
rect 29710 19122 29762 19134
rect 29710 19058 29762 19070
rect 36094 19122 36146 19134
rect 36094 19058 36146 19070
rect 36430 19122 36482 19134
rect 36430 19058 36482 19070
rect 37102 19122 37154 19134
rect 52782 19122 52834 19134
rect 37986 19070 37998 19122
rect 38050 19070 38062 19122
rect 45602 19070 45614 19122
rect 45666 19070 45678 19122
rect 37102 19058 37154 19070
rect 52782 19058 52834 19070
rect 2046 19010 2098 19022
rect 2046 18946 2098 18958
rect 5070 19010 5122 19022
rect 5070 18946 5122 18958
rect 5966 19010 6018 19022
rect 5966 18946 6018 18958
rect 7534 19010 7586 19022
rect 8318 19010 8370 19022
rect 7858 18958 7870 19010
rect 7922 18958 7934 19010
rect 7534 18946 7586 18958
rect 8318 18946 8370 18958
rect 9886 19010 9938 19022
rect 9886 18946 9938 18958
rect 12126 19010 12178 19022
rect 12126 18946 12178 18958
rect 15934 19010 15986 19022
rect 15934 18946 15986 18958
rect 22766 19010 22818 19022
rect 22766 18946 22818 18958
rect 29934 19010 29986 19022
rect 29934 18946 29986 18958
rect 52670 19010 52722 19022
rect 52670 18946 52722 18958
rect 1344 18842 58576 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 50558 18842
rect 50610 18790 50662 18842
rect 50714 18790 50766 18842
rect 50818 18790 58576 18842
rect 1344 18756 58576 18790
rect 1822 18674 1874 18686
rect 7310 18674 7362 18686
rect 4834 18622 4846 18674
rect 4898 18622 4910 18674
rect 1822 18610 1874 18622
rect 7310 18610 7362 18622
rect 13470 18674 13522 18686
rect 16942 18674 16994 18686
rect 14242 18622 14254 18674
rect 14306 18622 14318 18674
rect 13470 18610 13522 18622
rect 16942 18610 16994 18622
rect 18174 18674 18226 18686
rect 18174 18610 18226 18622
rect 18622 18674 18674 18686
rect 18622 18610 18674 18622
rect 18846 18674 18898 18686
rect 18846 18610 18898 18622
rect 19182 18674 19234 18686
rect 19182 18610 19234 18622
rect 19406 18674 19458 18686
rect 19406 18610 19458 18622
rect 19966 18674 20018 18686
rect 19966 18610 20018 18622
rect 23662 18674 23714 18686
rect 23662 18610 23714 18622
rect 24446 18674 24498 18686
rect 24446 18610 24498 18622
rect 30606 18674 30658 18686
rect 30606 18610 30658 18622
rect 37886 18674 37938 18686
rect 37886 18610 37938 18622
rect 45166 18674 45218 18686
rect 45166 18610 45218 18622
rect 2942 18562 2994 18574
rect 5630 18562 5682 18574
rect 4162 18510 4174 18562
rect 4226 18510 4238 18562
rect 4946 18510 4958 18562
rect 5010 18510 5022 18562
rect 2942 18498 2994 18510
rect 5630 18498 5682 18510
rect 5742 18562 5794 18574
rect 5742 18498 5794 18510
rect 6190 18562 6242 18574
rect 6190 18498 6242 18510
rect 6750 18562 6802 18574
rect 6750 18498 6802 18510
rect 7534 18562 7586 18574
rect 7534 18498 7586 18510
rect 9998 18562 10050 18574
rect 9998 18498 10050 18510
rect 10110 18562 10162 18574
rect 13358 18562 13410 18574
rect 11778 18510 11790 18562
rect 11842 18510 11854 18562
rect 10110 18498 10162 18510
rect 13358 18498 13410 18510
rect 16718 18562 16770 18574
rect 16718 18498 16770 18510
rect 17838 18562 17890 18574
rect 17838 18498 17890 18510
rect 17950 18562 18002 18574
rect 17950 18498 18002 18510
rect 18510 18562 18562 18574
rect 18510 18498 18562 18510
rect 19518 18562 19570 18574
rect 19518 18498 19570 18510
rect 19854 18562 19906 18574
rect 19854 18498 19906 18510
rect 23774 18562 23826 18574
rect 23774 18498 23826 18510
rect 27918 18562 27970 18574
rect 27918 18498 27970 18510
rect 28030 18562 28082 18574
rect 48750 18562 48802 18574
rect 41122 18510 41134 18562
rect 41186 18510 41198 18562
rect 45714 18510 45726 18562
rect 45778 18510 45790 18562
rect 28030 18498 28082 18510
rect 48750 18498 48802 18510
rect 2718 18450 2770 18462
rect 2718 18386 2770 18398
rect 3054 18450 3106 18462
rect 6526 18450 6578 18462
rect 4050 18398 4062 18450
rect 4114 18398 4126 18450
rect 3054 18386 3106 18398
rect 6526 18386 6578 18398
rect 6862 18450 6914 18462
rect 6862 18386 6914 18398
rect 7646 18450 7698 18462
rect 7646 18386 7698 18398
rect 10558 18450 10610 18462
rect 11454 18450 11506 18462
rect 11106 18398 11118 18450
rect 11170 18398 11182 18450
rect 10558 18386 10610 18398
rect 11454 18386 11506 18398
rect 13918 18450 13970 18462
rect 15598 18450 15650 18462
rect 15138 18398 15150 18450
rect 15202 18398 15214 18450
rect 13918 18386 13970 18398
rect 15598 18386 15650 18398
rect 16606 18450 16658 18462
rect 16606 18386 16658 18398
rect 20190 18450 20242 18462
rect 24334 18450 24386 18462
rect 20738 18398 20750 18450
rect 20802 18398 20814 18450
rect 21298 18398 21310 18450
rect 21362 18398 21374 18450
rect 22082 18398 22094 18450
rect 22146 18398 22158 18450
rect 20190 18386 20242 18398
rect 24334 18386 24386 18398
rect 24670 18450 24722 18462
rect 28254 18450 28306 18462
rect 27122 18398 27134 18450
rect 27186 18398 27198 18450
rect 24670 18386 24722 18398
rect 28254 18386 28306 18398
rect 28590 18450 28642 18462
rect 28590 18386 28642 18398
rect 30270 18450 30322 18462
rect 30270 18386 30322 18398
rect 37326 18450 37378 18462
rect 37326 18386 37378 18398
rect 37774 18450 37826 18462
rect 37774 18386 37826 18398
rect 37998 18450 38050 18462
rect 42142 18450 42194 18462
rect 46734 18450 46786 18462
rect 41346 18398 41358 18450
rect 41410 18398 41422 18450
rect 44930 18398 44942 18450
rect 44994 18398 45006 18450
rect 45938 18398 45950 18450
rect 46002 18398 46014 18450
rect 37998 18386 38050 18398
rect 42142 18386 42194 18398
rect 46734 18386 46786 18398
rect 49086 18450 49138 18462
rect 51650 18398 51662 18450
rect 51714 18398 51726 18450
rect 52098 18398 52110 18450
rect 52162 18398 52174 18450
rect 53442 18398 53454 18450
rect 53506 18398 53518 18450
rect 49086 18386 49138 18398
rect 2270 18338 2322 18350
rect 2270 18274 2322 18286
rect 8094 18338 8146 18350
rect 8094 18274 8146 18286
rect 12350 18338 12402 18350
rect 27470 18338 27522 18350
rect 15250 18286 15262 18338
rect 15314 18286 15326 18338
rect 22530 18286 22542 18338
rect 22594 18286 22606 18338
rect 27346 18286 27358 18338
rect 27410 18286 27422 18338
rect 12350 18274 12402 18286
rect 27470 18274 27522 18286
rect 38558 18338 38610 18350
rect 38558 18274 38610 18286
rect 39006 18338 39058 18350
rect 39006 18274 39058 18286
rect 46398 18338 46450 18350
rect 51986 18286 51998 18338
rect 52050 18286 52062 18338
rect 46398 18274 46450 18286
rect 5630 18226 5682 18238
rect 1698 18174 1710 18226
rect 1762 18223 1774 18226
rect 2258 18223 2270 18226
rect 1762 18177 2270 18223
rect 1762 18174 1774 18177
rect 2258 18174 2270 18177
rect 2322 18174 2334 18226
rect 5630 18162 5682 18174
rect 10110 18226 10162 18238
rect 10110 18162 10162 18174
rect 10782 18226 10834 18238
rect 10782 18162 10834 18174
rect 13470 18226 13522 18238
rect 13470 18162 13522 18174
rect 23550 18226 23602 18238
rect 23550 18162 23602 18174
rect 41806 18226 41858 18238
rect 41806 18162 41858 18174
rect 51550 18226 51602 18238
rect 55346 18174 55358 18226
rect 55410 18174 55422 18226
rect 51550 18162 51602 18174
rect 1344 18058 58576 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 58576 18058
rect 1344 17972 58576 18006
rect 16270 17890 16322 17902
rect 3714 17838 3726 17890
rect 3778 17838 3790 17890
rect 15250 17838 15262 17890
rect 15314 17838 15326 17890
rect 16270 17826 16322 17838
rect 26574 17890 26626 17902
rect 26574 17826 26626 17838
rect 50766 17890 50818 17902
rect 50766 17826 50818 17838
rect 51102 17890 51154 17902
rect 51102 17826 51154 17838
rect 51214 17890 51266 17902
rect 51214 17826 51266 17838
rect 57934 17890 57986 17902
rect 57934 17826 57986 17838
rect 5854 17778 5906 17790
rect 5854 17714 5906 17726
rect 7870 17778 7922 17790
rect 27918 17778 27970 17790
rect 35310 17778 35362 17790
rect 10770 17726 10782 17778
rect 10834 17726 10846 17778
rect 13570 17726 13582 17778
rect 13634 17726 13646 17778
rect 31938 17726 31950 17778
rect 32002 17726 32014 17778
rect 7870 17714 7922 17726
rect 27918 17714 27970 17726
rect 35310 17714 35362 17726
rect 35758 17778 35810 17790
rect 35758 17714 35810 17726
rect 39230 17778 39282 17790
rect 39230 17714 39282 17726
rect 46958 17778 47010 17790
rect 51662 17778 51714 17790
rect 48066 17726 48078 17778
rect 48130 17726 48142 17778
rect 50194 17726 50206 17778
rect 50258 17726 50270 17778
rect 46958 17714 47010 17726
rect 51662 17714 51714 17726
rect 55022 17778 55074 17790
rect 55022 17714 55074 17726
rect 2606 17666 2658 17678
rect 4398 17666 4450 17678
rect 8318 17666 8370 17678
rect 2258 17614 2270 17666
rect 2322 17614 2334 17666
rect 3378 17614 3390 17666
rect 3442 17614 3454 17666
rect 7298 17614 7310 17666
rect 7362 17614 7374 17666
rect 2606 17602 2658 17614
rect 4398 17602 4450 17614
rect 8318 17602 8370 17614
rect 10334 17666 10386 17678
rect 10334 17602 10386 17614
rect 11118 17666 11170 17678
rect 11118 17602 11170 17614
rect 13022 17666 13074 17678
rect 18622 17666 18674 17678
rect 13682 17614 13694 17666
rect 13746 17614 13758 17666
rect 15026 17614 15038 17666
rect 15090 17614 15102 17666
rect 13022 17602 13074 17614
rect 18622 17602 18674 17614
rect 18846 17666 18898 17678
rect 27022 17666 27074 17678
rect 30718 17666 30770 17678
rect 37662 17666 37714 17678
rect 19506 17614 19518 17666
rect 19570 17614 19582 17666
rect 21858 17614 21870 17666
rect 21922 17614 21934 17666
rect 23202 17614 23214 17666
rect 23266 17614 23278 17666
rect 25106 17614 25118 17666
rect 25170 17614 25182 17666
rect 27234 17614 27246 17666
rect 27298 17614 27310 17666
rect 31378 17614 31390 17666
rect 31442 17614 31454 17666
rect 34850 17614 34862 17666
rect 34914 17614 34926 17666
rect 36306 17614 36318 17666
rect 36370 17614 36382 17666
rect 37202 17614 37214 17666
rect 37266 17614 37278 17666
rect 18846 17602 18898 17614
rect 27022 17602 27074 17614
rect 30718 17602 30770 17614
rect 37662 17602 37714 17614
rect 38334 17666 38386 17678
rect 39790 17666 39842 17678
rect 39442 17614 39454 17666
rect 39506 17614 39518 17666
rect 38334 17602 38386 17614
rect 39790 17602 39842 17614
rect 40126 17666 40178 17678
rect 40126 17602 40178 17614
rect 40350 17666 40402 17678
rect 40350 17602 40402 17614
rect 45278 17666 45330 17678
rect 50878 17666 50930 17678
rect 45938 17614 45950 17666
rect 46002 17614 46014 17666
rect 47282 17614 47294 17666
rect 47346 17614 47358 17666
rect 45278 17602 45330 17614
rect 50878 17602 50930 17614
rect 52222 17666 52274 17678
rect 52658 17614 52670 17666
rect 52722 17614 52734 17666
rect 55570 17614 55582 17666
rect 55634 17614 55646 17666
rect 52222 17602 52274 17614
rect 9886 17554 9938 17566
rect 4722 17502 4734 17554
rect 4786 17502 4798 17554
rect 6178 17502 6190 17554
rect 6242 17502 6254 17554
rect 9886 17490 9938 17502
rect 9998 17554 10050 17566
rect 9998 17490 10050 17502
rect 11454 17554 11506 17566
rect 11454 17490 11506 17502
rect 11678 17554 11730 17566
rect 11678 17490 11730 17502
rect 11902 17554 11954 17566
rect 11902 17490 11954 17502
rect 12014 17554 12066 17566
rect 12014 17490 12066 17502
rect 12686 17554 12738 17566
rect 12686 17490 12738 17502
rect 16382 17554 16434 17566
rect 26462 17554 26514 17566
rect 20626 17502 20638 17554
rect 20690 17502 20702 17554
rect 22082 17502 22094 17554
rect 22146 17502 22158 17554
rect 24770 17502 24782 17554
rect 24834 17502 24846 17554
rect 16382 17490 16434 17502
rect 26462 17490 26514 17502
rect 29934 17554 29986 17566
rect 29934 17490 29986 17502
rect 30382 17554 30434 17566
rect 40574 17554 40626 17566
rect 31490 17502 31502 17554
rect 31554 17502 31566 17554
rect 34066 17502 34078 17554
rect 34130 17502 34142 17554
rect 37986 17502 37998 17554
rect 38050 17502 38062 17554
rect 30382 17490 30434 17502
rect 40574 17490 40626 17502
rect 43822 17554 43874 17566
rect 43822 17490 43874 17502
rect 44942 17554 44994 17566
rect 51550 17554 51602 17566
rect 45826 17502 45838 17554
rect 45890 17502 45902 17554
rect 44942 17490 44994 17502
rect 51550 17490 51602 17502
rect 10222 17442 10274 17454
rect 8642 17390 8654 17442
rect 8706 17390 8718 17442
rect 10222 17378 10274 17390
rect 10670 17442 10722 17454
rect 10670 17378 10722 17390
rect 10894 17442 10946 17454
rect 10894 17378 10946 17390
rect 11342 17442 11394 17454
rect 11342 17378 11394 17390
rect 12798 17442 12850 17454
rect 12798 17378 12850 17390
rect 16270 17442 16322 17454
rect 25566 17442 25618 17454
rect 18274 17390 18286 17442
rect 18338 17390 18350 17442
rect 16270 17378 16322 17390
rect 25566 17378 25618 17390
rect 29598 17442 29650 17454
rect 39118 17442 39170 17454
rect 36082 17390 36094 17442
rect 36146 17390 36158 17442
rect 36978 17390 36990 17442
rect 37042 17390 37054 17442
rect 38658 17390 38670 17442
rect 38722 17390 38734 17442
rect 29598 17378 29650 17390
rect 39118 17378 39170 17390
rect 39342 17442 39394 17454
rect 39342 17378 39394 17390
rect 40686 17442 40738 17454
rect 40686 17378 40738 17390
rect 40798 17442 40850 17454
rect 40798 17378 40850 17390
rect 42142 17442 42194 17454
rect 42142 17378 42194 17390
rect 43486 17442 43538 17454
rect 43486 17378 43538 17390
rect 51774 17442 51826 17454
rect 51774 17378 51826 17390
rect 1344 17274 58576 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 50558 17274
rect 50610 17222 50662 17274
rect 50714 17222 50766 17274
rect 50818 17222 58576 17274
rect 1344 17188 58576 17222
rect 1710 17106 1762 17118
rect 3950 17106 4002 17118
rect 2034 17054 2046 17106
rect 2098 17054 2110 17106
rect 1710 17042 1762 17054
rect 3950 17042 4002 17054
rect 5182 17106 5234 17118
rect 5182 17042 5234 17054
rect 5854 17106 5906 17118
rect 26574 17106 26626 17118
rect 6962 17054 6974 17106
rect 7026 17054 7038 17106
rect 14690 17054 14702 17106
rect 14754 17054 14766 17106
rect 5854 17042 5906 17054
rect 26574 17042 26626 17054
rect 26798 17106 26850 17118
rect 26798 17042 26850 17054
rect 33518 17106 33570 17118
rect 33518 17042 33570 17054
rect 36430 17106 36482 17118
rect 36430 17042 36482 17054
rect 36990 17106 37042 17118
rect 36990 17042 37042 17054
rect 38110 17106 38162 17118
rect 38110 17042 38162 17054
rect 39678 17106 39730 17118
rect 39678 17042 39730 17054
rect 41806 17106 41858 17118
rect 41806 17042 41858 17054
rect 45614 17106 45666 17118
rect 45614 17042 45666 17054
rect 49982 17106 50034 17118
rect 49982 17042 50034 17054
rect 3614 16994 3666 17006
rect 3614 16930 3666 16942
rect 6078 16994 6130 17006
rect 9774 16994 9826 17006
rect 8306 16942 8318 16994
rect 8370 16942 8382 16994
rect 6078 16930 6130 16942
rect 9774 16930 9826 16942
rect 10110 16994 10162 17006
rect 15038 16994 15090 17006
rect 17726 16994 17778 17006
rect 12002 16942 12014 16994
rect 12066 16942 12078 16994
rect 15362 16942 15374 16994
rect 15426 16942 15438 16994
rect 10110 16930 10162 16942
rect 15038 16930 15090 16942
rect 17726 16930 17778 16942
rect 17838 16994 17890 17006
rect 24670 16994 24722 17006
rect 18498 16942 18510 16994
rect 18562 16942 18574 16994
rect 19058 16942 19070 16994
rect 19122 16942 19134 16994
rect 20962 16942 20974 16994
rect 21026 16942 21038 16994
rect 23202 16942 23214 16994
rect 23266 16942 23278 16994
rect 17838 16930 17890 16942
rect 24670 16930 24722 16942
rect 26014 16994 26066 17006
rect 32062 16994 32114 17006
rect 35758 16994 35810 17006
rect 50654 16994 50706 17006
rect 29138 16942 29150 16994
rect 29202 16942 29214 16994
rect 35074 16942 35086 16994
rect 35138 16942 35150 16994
rect 43026 16942 43038 16994
rect 43090 16942 43102 16994
rect 49074 16942 49086 16994
rect 49138 16942 49150 16994
rect 52210 16942 52222 16994
rect 52274 16942 52286 16994
rect 26014 16930 26066 16942
rect 32062 16930 32114 16942
rect 35758 16930 35810 16942
rect 50654 16930 50706 16942
rect 4510 16882 4562 16894
rect 2930 16830 2942 16882
rect 2994 16830 3006 16882
rect 3378 16830 3390 16882
rect 3442 16830 3454 16882
rect 4510 16818 4562 16830
rect 4958 16882 5010 16894
rect 4958 16818 5010 16830
rect 5070 16882 5122 16894
rect 6190 16882 6242 16894
rect 5506 16830 5518 16882
rect 5570 16830 5582 16882
rect 5070 16818 5122 16830
rect 6190 16818 6242 16830
rect 7310 16882 7362 16894
rect 9550 16882 9602 16894
rect 14030 16882 14082 16894
rect 7970 16830 7982 16882
rect 8034 16830 8046 16882
rect 9090 16830 9102 16882
rect 9154 16830 9166 16882
rect 12226 16830 12238 16882
rect 12290 16830 12302 16882
rect 7310 16818 7362 16830
rect 9550 16818 9602 16830
rect 14030 16818 14082 16830
rect 14366 16882 14418 16894
rect 14366 16818 14418 16830
rect 18286 16882 18338 16894
rect 26462 16882 26514 16894
rect 34078 16882 34130 16894
rect 36206 16882 36258 16894
rect 21970 16830 21982 16882
rect 22034 16830 22046 16882
rect 23090 16830 23102 16882
rect 23154 16830 23166 16882
rect 23986 16830 23998 16882
rect 24050 16830 24062 16882
rect 28466 16830 28478 16882
rect 28530 16830 28542 16882
rect 33282 16830 33294 16882
rect 33346 16830 33358 16882
rect 35186 16830 35198 16882
rect 35250 16830 35262 16882
rect 18286 16818 18338 16830
rect 26462 16818 26514 16830
rect 34078 16818 34130 16830
rect 36206 16818 36258 16830
rect 36542 16882 36594 16894
rect 36542 16818 36594 16830
rect 37438 16882 37490 16894
rect 39902 16882 39954 16894
rect 39442 16830 39454 16882
rect 39506 16830 39518 16882
rect 37438 16818 37490 16830
rect 39902 16818 39954 16830
rect 40014 16882 40066 16894
rect 40014 16818 40066 16830
rect 41358 16882 41410 16894
rect 41358 16818 41410 16830
rect 41582 16882 41634 16894
rect 42242 16830 42254 16882
rect 42306 16830 42318 16882
rect 48850 16830 48862 16882
rect 48914 16830 48926 16882
rect 51314 16830 51326 16882
rect 51378 16830 51390 16882
rect 51986 16830 51998 16882
rect 52050 16830 52062 16882
rect 53554 16830 53566 16882
rect 53618 16830 53630 16882
rect 41582 16818 41634 16830
rect 7870 16770 7922 16782
rect 7870 16706 7922 16718
rect 9998 16770 10050 16782
rect 9998 16706 10050 16718
rect 16046 16770 16098 16782
rect 16046 16706 16098 16718
rect 18174 16770 18226 16782
rect 34414 16770 34466 16782
rect 23762 16718 23774 16770
rect 23826 16718 23838 16770
rect 31266 16718 31278 16770
rect 31330 16718 31342 16770
rect 18174 16706 18226 16718
rect 34414 16706 34466 16718
rect 39790 16770 39842 16782
rect 41682 16718 41694 16770
rect 41746 16718 41758 16770
rect 45154 16718 45166 16770
rect 45218 16718 45230 16770
rect 39790 16706 39842 16718
rect 16270 16658 16322 16670
rect 16270 16594 16322 16606
rect 16494 16658 16546 16670
rect 16494 16594 16546 16606
rect 16942 16658 16994 16670
rect 16942 16594 16994 16606
rect 17726 16658 17778 16670
rect 17726 16594 17778 16606
rect 25790 16658 25842 16670
rect 25790 16594 25842 16606
rect 26126 16658 26178 16670
rect 26126 16594 26178 16606
rect 31838 16658 31890 16670
rect 31838 16594 31890 16606
rect 32174 16658 32226 16670
rect 32174 16594 32226 16606
rect 40910 16658 40962 16670
rect 40910 16594 40962 16606
rect 41134 16658 41186 16670
rect 41134 16594 41186 16606
rect 49646 16658 49698 16670
rect 55346 16606 55358 16658
rect 55410 16606 55422 16658
rect 49646 16594 49698 16606
rect 1344 16490 58576 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 58576 16490
rect 1344 16404 58576 16438
rect 7982 16322 8034 16334
rect 7982 16258 8034 16270
rect 9550 16322 9602 16334
rect 17614 16322 17666 16334
rect 31614 16322 31666 16334
rect 9874 16270 9886 16322
rect 9938 16270 9950 16322
rect 15698 16270 15710 16322
rect 15762 16319 15774 16322
rect 16258 16319 16270 16322
rect 15762 16273 16270 16319
rect 15762 16270 15774 16273
rect 16258 16270 16270 16273
rect 16322 16270 16334 16322
rect 20626 16270 20638 16322
rect 20690 16270 20702 16322
rect 26898 16270 26910 16322
rect 26962 16270 26974 16322
rect 9550 16258 9602 16270
rect 17614 16258 17666 16270
rect 31614 16258 31666 16270
rect 32510 16322 32562 16334
rect 32510 16258 32562 16270
rect 40798 16322 40850 16334
rect 40798 16258 40850 16270
rect 51998 16322 52050 16334
rect 57934 16322 57986 16334
rect 52770 16270 52782 16322
rect 52834 16270 52846 16322
rect 51998 16258 52050 16270
rect 57934 16258 57986 16270
rect 2830 16210 2882 16222
rect 10446 16210 10498 16222
rect 30158 16210 30210 16222
rect 6738 16158 6750 16210
rect 6802 16158 6814 16210
rect 14802 16158 14814 16210
rect 14866 16158 14878 16210
rect 16818 16158 16830 16210
rect 16882 16158 16894 16210
rect 26226 16158 26238 16210
rect 26290 16158 26302 16210
rect 2830 16146 2882 16158
rect 10446 16146 10498 16158
rect 30158 16146 30210 16158
rect 31166 16210 31218 16222
rect 34526 16210 34578 16222
rect 42590 16210 42642 16222
rect 32946 16158 32958 16210
rect 33010 16158 33022 16210
rect 34178 16158 34190 16210
rect 34242 16158 34254 16210
rect 35186 16158 35198 16210
rect 35250 16158 35262 16210
rect 41346 16158 41358 16210
rect 41410 16158 41422 16210
rect 31166 16146 31218 16158
rect 34526 16146 34578 16158
rect 42590 16146 42642 16158
rect 46510 16210 46562 16222
rect 48626 16158 48638 16210
rect 48690 16158 48702 16210
rect 46510 16146 46562 16158
rect 1710 16098 1762 16110
rect 4622 16098 4674 16110
rect 9214 16098 9266 16110
rect 10222 16098 10274 16110
rect 12686 16098 12738 16110
rect 22430 16098 22482 16110
rect 29822 16098 29874 16110
rect 3378 16046 3390 16098
rect 3442 16046 3454 16098
rect 6178 16046 6190 16098
rect 6242 16046 6254 16098
rect 7298 16046 7310 16098
rect 7362 16046 7374 16098
rect 7858 16046 7870 16098
rect 7922 16046 7934 16098
rect 9538 16046 9550 16098
rect 9602 16046 9614 16098
rect 11778 16046 11790 16098
rect 11842 16046 11854 16098
rect 13794 16046 13806 16098
rect 13858 16046 13870 16098
rect 14578 16046 14590 16098
rect 14642 16046 14654 16098
rect 16706 16046 16718 16098
rect 16770 16046 16782 16098
rect 17714 16046 17726 16098
rect 17778 16046 17790 16098
rect 18162 16046 18174 16098
rect 18226 16046 18238 16098
rect 19170 16046 19182 16098
rect 19234 16046 19246 16098
rect 20514 16046 20526 16098
rect 20578 16046 20590 16098
rect 24098 16046 24110 16098
rect 24162 16046 24174 16098
rect 24994 16046 25006 16098
rect 25058 16046 25070 16098
rect 26338 16046 26350 16098
rect 26402 16046 26414 16098
rect 1710 16034 1762 16046
rect 4622 16034 4674 16046
rect 9214 16034 9266 16046
rect 10222 16034 10274 16046
rect 12686 16034 12738 16046
rect 22430 16034 22482 16046
rect 29822 16034 29874 16046
rect 31390 16098 31442 16110
rect 32286 16098 32338 16110
rect 33182 16098 33234 16110
rect 31938 16046 31950 16098
rect 32002 16046 32014 16098
rect 32834 16046 32846 16098
rect 32898 16046 32910 16098
rect 31390 16034 31442 16046
rect 32286 16034 32338 16046
rect 33182 16034 33234 16046
rect 34750 16098 34802 16110
rect 34750 16034 34802 16046
rect 34974 16098 35026 16110
rect 34974 16034 35026 16046
rect 35422 16098 35474 16110
rect 35422 16034 35474 16046
rect 39118 16098 39170 16110
rect 39118 16034 39170 16046
rect 39454 16098 39506 16110
rect 39454 16034 39506 16046
rect 39566 16098 39618 16110
rect 40350 16098 40402 16110
rect 39890 16046 39902 16098
rect 39954 16046 39966 16098
rect 39566 16034 39618 16046
rect 40350 16034 40402 16046
rect 40574 16098 40626 16110
rect 42478 16098 42530 16110
rect 41122 16046 41134 16098
rect 41186 16046 41198 16098
rect 42130 16046 42142 16098
rect 42194 16046 42206 16098
rect 40574 16034 40626 16046
rect 42478 16034 42530 16046
rect 42702 16098 42754 16110
rect 52894 16098 52946 16110
rect 47058 16046 47070 16098
rect 47122 16046 47134 16098
rect 53106 16046 53118 16098
rect 53170 16046 53182 16098
rect 55570 16046 55582 16098
rect 55634 16046 55646 16098
rect 42702 16034 42754 16046
rect 52894 16034 52946 16046
rect 2046 15986 2098 15998
rect 2046 15922 2098 15934
rect 2942 15986 2994 15998
rect 2942 15922 2994 15934
rect 4062 15986 4114 15998
rect 4062 15922 4114 15934
rect 4174 15986 4226 15998
rect 15262 15986 15314 15998
rect 6290 15934 6302 15986
rect 6354 15934 6366 15986
rect 8082 15934 8094 15986
rect 8146 15934 8158 15986
rect 12002 15934 12014 15986
rect 12066 15934 12078 15986
rect 14466 15934 14478 15986
rect 14530 15934 14542 15986
rect 4174 15922 4226 15934
rect 15262 15922 15314 15934
rect 22766 15986 22818 15998
rect 25678 15986 25730 15998
rect 23986 15934 23998 15986
rect 24050 15934 24062 15986
rect 22766 15922 22818 15934
rect 25678 15922 25730 15934
rect 30046 15986 30098 15998
rect 30046 15922 30098 15934
rect 30382 15986 30434 15998
rect 30382 15922 30434 15934
rect 30606 15986 30658 15998
rect 30606 15922 30658 15934
rect 33854 15986 33906 15998
rect 33854 15922 33906 15934
rect 35198 15986 35250 15998
rect 35198 15922 35250 15934
rect 38782 15986 38834 15998
rect 41470 15986 41522 15998
rect 39778 15934 39790 15986
rect 39842 15934 39854 15986
rect 38782 15922 38834 15934
rect 41470 15922 41522 15934
rect 45278 15986 45330 15998
rect 51662 15986 51714 15998
rect 48066 15934 48078 15986
rect 48130 15934 48142 15986
rect 45278 15922 45330 15934
rect 51662 15922 51714 15934
rect 55358 15986 55410 15998
rect 55358 15922 55410 15934
rect 2718 15874 2770 15886
rect 2718 15810 2770 15822
rect 3614 15874 3666 15886
rect 3614 15810 3666 15822
rect 3838 15874 3890 15886
rect 3838 15810 3890 15822
rect 12798 15874 12850 15886
rect 12798 15810 12850 15822
rect 13022 15874 13074 15886
rect 13022 15810 13074 15822
rect 15374 15874 15426 15886
rect 15374 15810 15426 15822
rect 15598 15874 15650 15886
rect 15598 15810 15650 15822
rect 15934 15874 15986 15886
rect 15934 15810 15986 15822
rect 22542 15874 22594 15886
rect 22542 15810 22594 15822
rect 23102 15874 23154 15886
rect 23102 15810 23154 15822
rect 29150 15874 29202 15886
rect 29150 15810 29202 15822
rect 29262 15874 29314 15886
rect 29262 15810 29314 15822
rect 29374 15874 29426 15886
rect 29374 15810 29426 15822
rect 32958 15874 33010 15886
rect 32958 15810 33010 15822
rect 34078 15874 34130 15886
rect 34078 15810 34130 15822
rect 38894 15874 38946 15886
rect 38894 15810 38946 15822
rect 41246 15874 41298 15886
rect 41246 15810 41298 15822
rect 45054 15874 45106 15886
rect 45054 15810 45106 15822
rect 45166 15874 45218 15886
rect 45166 15810 45218 15822
rect 51886 15874 51938 15886
rect 51886 15810 51938 15822
rect 54238 15874 54290 15886
rect 54238 15810 54290 15822
rect 1344 15706 58576 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 50558 15706
rect 50610 15654 50662 15706
rect 50714 15654 50766 15706
rect 50818 15654 58576 15706
rect 1344 15620 58576 15654
rect 4846 15538 4898 15550
rect 4846 15474 4898 15486
rect 4958 15538 5010 15550
rect 5742 15538 5794 15550
rect 5506 15486 5518 15538
rect 5570 15486 5582 15538
rect 4958 15474 5010 15486
rect 5742 15474 5794 15486
rect 5966 15538 6018 15550
rect 5966 15474 6018 15486
rect 6526 15538 6578 15550
rect 8094 15538 8146 15550
rect 9886 15538 9938 15550
rect 16158 15538 16210 15550
rect 23886 15538 23938 15550
rect 7298 15486 7310 15538
rect 7362 15486 7374 15538
rect 8866 15486 8878 15538
rect 8930 15486 8942 15538
rect 12450 15486 12462 15538
rect 12514 15486 12526 15538
rect 18386 15486 18398 15538
rect 18450 15486 18462 15538
rect 6526 15474 6578 15486
rect 8094 15474 8146 15486
rect 9886 15474 9938 15486
rect 16158 15474 16210 15486
rect 23886 15474 23938 15486
rect 25902 15538 25954 15550
rect 25902 15474 25954 15486
rect 26126 15538 26178 15550
rect 40126 15538 40178 15550
rect 34514 15486 34526 15538
rect 34578 15486 34590 15538
rect 37538 15486 37550 15538
rect 37602 15486 37614 15538
rect 38546 15486 38558 15538
rect 38610 15486 38622 15538
rect 26126 15474 26178 15486
rect 40126 15474 40178 15486
rect 42142 15538 42194 15550
rect 42142 15474 42194 15486
rect 47182 15538 47234 15550
rect 47182 15474 47234 15486
rect 51998 15538 52050 15550
rect 51998 15474 52050 15486
rect 6190 15426 6242 15438
rect 6190 15362 6242 15374
rect 15598 15426 15650 15438
rect 23662 15426 23714 15438
rect 17602 15374 17614 15426
rect 17666 15374 17678 15426
rect 15598 15362 15650 15374
rect 23662 15362 23714 15374
rect 23998 15426 24050 15438
rect 23998 15362 24050 15374
rect 29038 15426 29090 15438
rect 40238 15426 40290 15438
rect 30146 15374 30158 15426
rect 30210 15374 30222 15426
rect 30930 15374 30942 15426
rect 30994 15374 31006 15426
rect 33282 15374 33294 15426
rect 33346 15374 33358 15426
rect 35970 15374 35982 15426
rect 36034 15374 36046 15426
rect 29038 15362 29090 15374
rect 40238 15362 40290 15374
rect 41134 15426 41186 15438
rect 41134 15362 41186 15374
rect 42478 15426 42530 15438
rect 46398 15426 46450 15438
rect 43698 15374 43710 15426
rect 43762 15374 43774 15426
rect 42478 15362 42530 15374
rect 46398 15362 46450 15374
rect 48750 15426 48802 15438
rect 48750 15362 48802 15374
rect 2606 15314 2658 15326
rect 4734 15314 4786 15326
rect 5518 15314 5570 15326
rect 7870 15314 7922 15326
rect 2146 15262 2158 15314
rect 2210 15262 2222 15314
rect 3378 15262 3390 15314
rect 3442 15262 3454 15314
rect 4498 15262 4510 15314
rect 4562 15262 4574 15314
rect 5170 15262 5182 15314
rect 5234 15262 5246 15314
rect 6738 15262 6750 15314
rect 6802 15262 6814 15314
rect 7522 15262 7534 15314
rect 7586 15262 7598 15314
rect 2606 15250 2658 15262
rect 4734 15250 4786 15262
rect 5518 15250 5570 15262
rect 7870 15250 7922 15262
rect 8206 15314 8258 15326
rect 8206 15250 8258 15262
rect 8542 15314 8594 15326
rect 12126 15314 12178 15326
rect 15150 15314 15202 15326
rect 9650 15262 9662 15314
rect 9714 15262 9726 15314
rect 13122 15262 13134 15314
rect 13186 15262 13198 15314
rect 13682 15262 13694 15314
rect 13746 15262 13758 15314
rect 8542 15250 8594 15262
rect 12126 15250 12178 15262
rect 15150 15250 15202 15262
rect 15486 15314 15538 15326
rect 15486 15250 15538 15262
rect 15822 15314 15874 15326
rect 15822 15250 15874 15262
rect 16494 15314 16546 15326
rect 21310 15314 21362 15326
rect 16706 15262 16718 15314
rect 16770 15262 16782 15314
rect 17826 15262 17838 15314
rect 17890 15262 17902 15314
rect 18498 15262 18510 15314
rect 18562 15262 18574 15314
rect 19170 15262 19182 15314
rect 19234 15262 19246 15314
rect 20626 15262 20638 15314
rect 20690 15262 20702 15314
rect 16494 15250 16546 15262
rect 21310 15250 21362 15262
rect 22206 15314 22258 15326
rect 23102 15314 23154 15326
rect 22418 15262 22430 15314
rect 22482 15262 22494 15314
rect 22206 15250 22258 15262
rect 23102 15250 23154 15262
rect 23438 15314 23490 15326
rect 23438 15250 23490 15262
rect 25678 15314 25730 15326
rect 35086 15314 35138 15326
rect 39006 15314 39058 15326
rect 28578 15262 28590 15314
rect 28642 15262 28654 15314
rect 29474 15262 29486 15314
rect 29538 15262 29550 15314
rect 30482 15262 30494 15314
rect 30546 15262 30558 15314
rect 31490 15262 31502 15314
rect 31554 15262 31566 15314
rect 32050 15262 32062 15314
rect 32114 15262 32126 15314
rect 33506 15262 33518 15314
rect 33570 15262 33582 15314
rect 34178 15262 34190 15314
rect 34242 15262 34254 15314
rect 36306 15262 36318 15314
rect 36370 15262 36382 15314
rect 36978 15262 36990 15314
rect 37042 15262 37054 15314
rect 25678 15250 25730 15262
rect 35086 15250 35138 15262
rect 39006 15250 39058 15262
rect 39118 15314 39170 15326
rect 39678 15314 39730 15326
rect 39330 15262 39342 15314
rect 39394 15262 39406 15314
rect 39118 15250 39170 15262
rect 39678 15250 39730 15262
rect 39902 15314 39954 15326
rect 39902 15250 39954 15262
rect 41358 15314 41410 15326
rect 41358 15250 41410 15262
rect 41582 15314 41634 15326
rect 41582 15250 41634 15262
rect 41806 15314 41858 15326
rect 41806 15250 41858 15262
rect 42030 15314 42082 15326
rect 42030 15250 42082 15262
rect 42254 15314 42306 15326
rect 46174 15314 46226 15326
rect 44370 15262 44382 15314
rect 44434 15262 44446 15314
rect 45378 15262 45390 15314
rect 45442 15262 45454 15314
rect 42254 15250 42306 15262
rect 46174 15250 46226 15262
rect 46510 15314 46562 15326
rect 46510 15250 46562 15262
rect 47070 15314 47122 15326
rect 47070 15250 47122 15262
rect 47406 15314 47458 15326
rect 53118 15314 53170 15326
rect 47954 15262 47966 15314
rect 48018 15262 48030 15314
rect 49186 15262 49198 15314
rect 49250 15262 49262 15314
rect 50866 15262 50878 15314
rect 50930 15262 50942 15314
rect 53442 15262 53454 15314
rect 53506 15262 53518 15314
rect 47406 15250 47458 15262
rect 53118 15250 53170 15262
rect 25790 15202 25842 15214
rect 47630 15202 47682 15214
rect 52670 15202 52722 15214
rect 14690 15150 14702 15202
rect 14754 15150 14766 15202
rect 19282 15150 19294 15202
rect 19346 15150 19358 15202
rect 28130 15150 28142 15202
rect 28194 15150 28206 15202
rect 30034 15150 30046 15202
rect 30098 15150 30110 15202
rect 31602 15150 31614 15202
rect 31666 15150 31678 15202
rect 33170 15150 33182 15202
rect 33234 15150 33246 15202
rect 45266 15150 45278 15202
rect 45330 15150 45342 15202
rect 50978 15150 50990 15202
rect 51042 15150 51054 15202
rect 25790 15138 25842 15150
rect 47630 15138 47682 15150
rect 52670 15138 52722 15150
rect 52894 15202 52946 15214
rect 52894 15138 52946 15150
rect 34862 15090 34914 15102
rect 3490 15038 3502 15090
rect 3554 15038 3566 15090
rect 34862 15026 34914 15038
rect 47966 15090 48018 15102
rect 47966 15026 48018 15038
rect 52446 15090 52498 15102
rect 55346 15038 55358 15090
rect 55410 15038 55422 15090
rect 52446 15026 52498 15038
rect 1344 14922 58576 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 58576 14922
rect 1344 14836 58576 14870
rect 7198 14754 7250 14766
rect 2930 14702 2942 14754
rect 2994 14702 3006 14754
rect 7198 14690 7250 14702
rect 12798 14754 12850 14766
rect 29486 14754 29538 14766
rect 32174 14754 32226 14766
rect 57934 14754 57986 14766
rect 26226 14702 26238 14754
rect 26290 14702 26302 14754
rect 31602 14702 31614 14754
rect 31666 14702 31678 14754
rect 42018 14702 42030 14754
rect 42082 14702 42094 14754
rect 52994 14702 53006 14754
rect 53058 14702 53070 14754
rect 12798 14690 12850 14702
rect 29486 14690 29538 14702
rect 32174 14690 32226 14702
rect 57934 14690 57986 14702
rect 1822 14642 1874 14654
rect 22206 14642 22258 14654
rect 34414 14642 34466 14654
rect 54910 14642 54962 14654
rect 3042 14590 3054 14642
rect 3106 14590 3118 14642
rect 15698 14590 15710 14642
rect 15762 14590 15774 14642
rect 18386 14590 18398 14642
rect 18450 14590 18462 14642
rect 19058 14590 19070 14642
rect 19122 14590 19134 14642
rect 25666 14590 25678 14642
rect 25730 14590 25742 14642
rect 27906 14590 27918 14642
rect 27970 14590 27982 14642
rect 33506 14590 33518 14642
rect 33570 14590 33582 14642
rect 37762 14590 37774 14642
rect 37826 14590 37838 14642
rect 41458 14590 41470 14642
rect 41522 14590 41534 14642
rect 46050 14590 46062 14642
rect 46114 14590 46126 14642
rect 48402 14590 48414 14642
rect 48466 14590 48478 14642
rect 54114 14590 54126 14642
rect 54178 14590 54190 14642
rect 1822 14578 1874 14590
rect 22206 14578 22258 14590
rect 34414 14578 34466 14590
rect 54910 14578 54962 14590
rect 3502 14530 3554 14542
rect 2594 14478 2606 14530
rect 2658 14478 2670 14530
rect 3502 14466 3554 14478
rect 3838 14530 3890 14542
rect 3838 14466 3890 14478
rect 6302 14530 6354 14542
rect 10558 14530 10610 14542
rect 10098 14478 10110 14530
rect 10162 14478 10174 14530
rect 6302 14466 6354 14478
rect 10558 14466 10610 14478
rect 12126 14530 12178 14542
rect 12126 14466 12178 14478
rect 14702 14530 14754 14542
rect 24222 14530 24274 14542
rect 17378 14478 17390 14530
rect 17442 14478 17454 14530
rect 19282 14478 19294 14530
rect 19346 14478 19358 14530
rect 23538 14478 23550 14530
rect 23602 14478 23614 14530
rect 14702 14466 14754 14478
rect 24222 14466 24274 14478
rect 25006 14530 25058 14542
rect 30158 14530 30210 14542
rect 31502 14530 31554 14542
rect 36206 14530 36258 14542
rect 40910 14530 40962 14542
rect 25442 14478 25454 14530
rect 25506 14478 25518 14530
rect 27010 14478 27022 14530
rect 27074 14478 27086 14530
rect 27570 14478 27582 14530
rect 27634 14478 27646 14530
rect 29474 14478 29486 14530
rect 29538 14478 29550 14530
rect 30818 14478 30830 14530
rect 30882 14478 30894 14530
rect 33170 14478 33182 14530
rect 33234 14478 33246 14530
rect 35970 14478 35982 14530
rect 36034 14478 36046 14530
rect 36866 14478 36878 14530
rect 36930 14478 36942 14530
rect 37650 14478 37662 14530
rect 37714 14478 37726 14530
rect 39218 14478 39230 14530
rect 39282 14478 39294 14530
rect 41346 14478 41358 14530
rect 41410 14478 41422 14530
rect 45154 14478 45166 14530
rect 45218 14478 45230 14530
rect 45602 14478 45614 14530
rect 45666 14478 45678 14530
rect 47730 14478 47742 14530
rect 47794 14478 47806 14530
rect 48514 14478 48526 14530
rect 48578 14478 48590 14530
rect 50530 14478 50542 14530
rect 50594 14478 50606 14530
rect 51314 14478 51326 14530
rect 51378 14478 51390 14530
rect 51986 14478 51998 14530
rect 52050 14478 52062 14530
rect 52882 14478 52894 14530
rect 52946 14478 52958 14530
rect 53330 14478 53342 14530
rect 53394 14478 53406 14530
rect 53778 14478 53790 14530
rect 53842 14478 53854 14530
rect 55570 14478 55582 14530
rect 55634 14478 55646 14530
rect 25006 14466 25058 14478
rect 30158 14466 30210 14478
rect 31502 14466 31554 14478
rect 36206 14466 36258 14478
rect 40910 14466 40962 14478
rect 4622 14418 4674 14430
rect 4622 14354 4674 14366
rect 4958 14418 5010 14430
rect 7198 14418 7250 14430
rect 6626 14366 6638 14418
rect 6690 14366 6702 14418
rect 4958 14354 5010 14366
rect 7198 14354 7250 14366
rect 7310 14418 7362 14430
rect 12238 14418 12290 14430
rect 11218 14366 11230 14418
rect 11282 14366 11294 14418
rect 12798 14418 12850 14430
rect 7310 14354 7362 14366
rect 12238 14354 12290 14366
rect 12686 14362 12738 14374
rect 3726 14306 3778 14318
rect 3726 14242 3778 14254
rect 10894 14306 10946 14318
rect 10894 14242 10946 14254
rect 12462 14306 12514 14318
rect 12798 14354 12850 14366
rect 14478 14418 14530 14430
rect 14478 14354 14530 14366
rect 14590 14418 14642 14430
rect 19966 14418 20018 14430
rect 16146 14366 16158 14418
rect 16210 14366 16222 14418
rect 14590 14354 14642 14366
rect 19966 14354 20018 14366
rect 20302 14418 20354 14430
rect 20302 14354 20354 14366
rect 21422 14418 21474 14430
rect 21422 14354 21474 14366
rect 21758 14418 21810 14430
rect 24670 14418 24722 14430
rect 29150 14418 29202 14430
rect 22418 14366 22430 14418
rect 22482 14366 22494 14418
rect 28018 14366 28030 14418
rect 28082 14366 28094 14418
rect 21758 14354 21810 14366
rect 24670 14354 24722 14366
rect 29150 14354 29202 14366
rect 29822 14418 29874 14430
rect 29822 14354 29874 14366
rect 32174 14418 32226 14430
rect 32174 14354 32226 14366
rect 32286 14418 32338 14430
rect 32286 14354 32338 14366
rect 33854 14418 33906 14430
rect 33854 14354 33906 14366
rect 35534 14418 35586 14430
rect 35534 14354 35586 14366
rect 35646 14418 35698 14430
rect 35646 14354 35698 14366
rect 36318 14418 36370 14430
rect 39006 14418 39058 14430
rect 38322 14366 38334 14418
rect 38386 14366 38398 14418
rect 36318 14354 36370 14366
rect 39006 14354 39058 14366
rect 40574 14418 40626 14430
rect 54798 14418 54850 14430
rect 46162 14366 46174 14418
rect 46226 14366 46238 14418
rect 49186 14366 49198 14418
rect 49250 14366 49262 14418
rect 50418 14366 50430 14418
rect 50482 14366 50494 14418
rect 51762 14366 51774 14418
rect 51826 14366 51838 14418
rect 40574 14354 40626 14366
rect 54798 14354 54850 14366
rect 12686 14298 12738 14310
rect 20414 14306 20466 14318
rect 15138 14254 15150 14306
rect 15202 14254 15214 14306
rect 12462 14242 12514 14254
rect 20414 14242 20466 14254
rect 20638 14306 20690 14318
rect 20638 14242 20690 14254
rect 21534 14306 21586 14318
rect 21534 14242 21586 14254
rect 24782 14306 24834 14318
rect 24782 14242 24834 14254
rect 28590 14306 28642 14318
rect 28590 14242 28642 14254
rect 29934 14306 29986 14318
rect 29934 14242 29986 14254
rect 35310 14306 35362 14318
rect 35310 14242 35362 14254
rect 40686 14306 40738 14318
rect 55022 14306 55074 14318
rect 51202 14254 51214 14306
rect 51266 14254 51278 14306
rect 40686 14242 40738 14254
rect 55022 14242 55074 14254
rect 1344 14138 58576 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 50558 14138
rect 50610 14086 50662 14138
rect 50714 14086 50766 14138
rect 50818 14086 58576 14138
rect 1344 14052 58576 14086
rect 2718 13970 2770 13982
rect 2034 13918 2046 13970
rect 2098 13918 2110 13970
rect 2718 13906 2770 13918
rect 3166 13970 3218 13982
rect 6974 13970 7026 13982
rect 21646 13970 21698 13982
rect 3714 13918 3726 13970
rect 3778 13918 3790 13970
rect 4722 13918 4734 13970
rect 4786 13918 4798 13970
rect 15138 13918 15150 13970
rect 15202 13918 15214 13970
rect 3166 13906 3218 13918
rect 6974 13906 7026 13918
rect 21646 13906 21698 13918
rect 22542 13970 22594 13982
rect 22542 13906 22594 13918
rect 25454 13970 25506 13982
rect 25454 13906 25506 13918
rect 41246 13970 41298 13982
rect 41246 13906 41298 13918
rect 48862 13970 48914 13982
rect 55358 13970 55410 13982
rect 50306 13918 50318 13970
rect 50370 13918 50382 13970
rect 51202 13918 51214 13970
rect 51266 13918 51278 13970
rect 53890 13918 53902 13970
rect 53954 13918 53966 13970
rect 48862 13906 48914 13918
rect 55358 13906 55410 13918
rect 2382 13858 2434 13870
rect 2382 13794 2434 13806
rect 6526 13858 6578 13870
rect 6526 13794 6578 13806
rect 23102 13858 23154 13870
rect 23102 13794 23154 13806
rect 28142 13858 28194 13870
rect 28142 13794 28194 13806
rect 35646 13858 35698 13870
rect 40238 13858 40290 13870
rect 38546 13806 38558 13858
rect 38610 13806 38622 13858
rect 35646 13794 35698 13806
rect 40238 13794 40290 13806
rect 41022 13858 41074 13870
rect 41022 13794 41074 13806
rect 45054 13858 45106 13870
rect 45054 13794 45106 13806
rect 47406 13858 47458 13870
rect 47406 13794 47458 13806
rect 47854 13858 47906 13870
rect 47854 13794 47906 13806
rect 49086 13858 49138 13870
rect 49086 13794 49138 13806
rect 49758 13858 49810 13870
rect 49758 13794 49810 13806
rect 53566 13858 53618 13870
rect 53566 13794 53618 13806
rect 56590 13858 56642 13870
rect 56590 13794 56642 13806
rect 4398 13746 4450 13758
rect 6862 13746 6914 13758
rect 12686 13746 12738 13758
rect 14142 13746 14194 13758
rect 1810 13694 1822 13746
rect 1874 13694 1886 13746
rect 3938 13694 3950 13746
rect 4002 13694 4014 13746
rect 6290 13694 6302 13746
rect 6354 13694 6366 13746
rect 11330 13694 11342 13746
rect 11394 13694 11406 13746
rect 12898 13694 12910 13746
rect 12962 13694 12974 13746
rect 4398 13682 4450 13694
rect 6862 13682 6914 13694
rect 12686 13682 12738 13694
rect 14142 13682 14194 13694
rect 14814 13746 14866 13758
rect 16606 13746 16658 13758
rect 15698 13694 15710 13746
rect 15762 13694 15774 13746
rect 16146 13694 16158 13746
rect 16210 13694 16222 13746
rect 14814 13682 14866 13694
rect 16606 13682 16658 13694
rect 16942 13746 16994 13758
rect 16942 13682 16994 13694
rect 18062 13746 18114 13758
rect 22206 13746 22258 13758
rect 18722 13694 18734 13746
rect 18786 13694 18798 13746
rect 19730 13694 19742 13746
rect 19794 13694 19806 13746
rect 20066 13694 20078 13746
rect 20130 13694 20142 13746
rect 18062 13682 18114 13694
rect 22206 13682 22258 13694
rect 22318 13746 22370 13758
rect 22318 13682 22370 13694
rect 22654 13746 22706 13758
rect 22654 13682 22706 13694
rect 25118 13746 25170 13758
rect 25118 13682 25170 13694
rect 25454 13746 25506 13758
rect 25454 13682 25506 13694
rect 25678 13746 25730 13758
rect 40910 13746 40962 13758
rect 47742 13746 47794 13758
rect 27346 13694 27358 13746
rect 27410 13694 27422 13746
rect 30930 13694 30942 13746
rect 30994 13694 31006 13746
rect 35074 13694 35086 13746
rect 35138 13694 35150 13746
rect 38882 13694 38894 13746
rect 38946 13694 38958 13746
rect 39778 13694 39790 13746
rect 39842 13694 39854 13746
rect 44594 13694 44606 13746
rect 44658 13694 44670 13746
rect 46946 13694 46958 13746
rect 47010 13694 47022 13746
rect 25678 13682 25730 13694
rect 40910 13682 40962 13694
rect 47742 13682 47794 13694
rect 48078 13746 48130 13758
rect 48078 13682 48130 13694
rect 48750 13746 48802 13758
rect 48750 13682 48802 13694
rect 49982 13746 50034 13758
rect 49982 13682 50034 13694
rect 50654 13746 50706 13758
rect 53454 13746 53506 13758
rect 52882 13694 52894 13746
rect 52946 13694 52958 13746
rect 50654 13682 50706 13694
rect 53454 13682 53506 13694
rect 54238 13746 54290 13758
rect 57026 13694 57038 13746
rect 57090 13694 57102 13746
rect 54238 13682 54290 13694
rect 13582 13634 13634 13646
rect 10658 13582 10670 13634
rect 10722 13582 10734 13634
rect 13582 13570 13634 13582
rect 13918 13634 13970 13646
rect 13918 13570 13970 13582
rect 18286 13634 18338 13646
rect 29710 13634 29762 13646
rect 20850 13582 20862 13634
rect 20914 13582 20926 13634
rect 27906 13582 27918 13634
rect 27970 13582 27982 13634
rect 18286 13570 18338 13582
rect 29710 13570 29762 13582
rect 30158 13634 30210 13646
rect 41582 13634 41634 13646
rect 30594 13582 30606 13634
rect 30658 13582 30670 13634
rect 34738 13582 34750 13634
rect 34802 13582 34814 13634
rect 30158 13570 30210 13582
rect 41582 13570 41634 13582
rect 43038 13634 43090 13646
rect 54462 13634 54514 13646
rect 44258 13582 44270 13634
rect 44322 13582 44334 13634
rect 46498 13582 46510 13634
rect 46562 13582 46574 13634
rect 57362 13582 57374 13634
rect 57426 13582 57438 13634
rect 43038 13570 43090 13582
rect 54462 13570 54514 13582
rect 6974 13522 7026 13534
rect 14478 13522 14530 13534
rect 23326 13522 23378 13534
rect 10882 13470 10894 13522
rect 10946 13470 10958 13522
rect 17714 13470 17726 13522
rect 17778 13470 17790 13522
rect 6974 13458 7026 13470
rect 14478 13458 14530 13470
rect 23326 13458 23378 13470
rect 23662 13522 23714 13534
rect 23662 13458 23714 13470
rect 43262 13522 43314 13534
rect 50878 13522 50930 13534
rect 43586 13470 43598 13522
rect 43650 13470 43662 13522
rect 43262 13458 43314 13470
rect 50878 13458 50930 13470
rect 1344 13354 58576 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 58576 13354
rect 1344 13268 58576 13302
rect 3502 13186 3554 13198
rect 3502 13122 3554 13134
rect 25902 13186 25954 13198
rect 39790 13186 39842 13198
rect 31266 13134 31278 13186
rect 31330 13134 31342 13186
rect 25902 13122 25954 13134
rect 39790 13122 39842 13134
rect 46734 13186 46786 13198
rect 46734 13122 46786 13134
rect 4062 13074 4114 13086
rect 4062 13010 4114 13022
rect 15262 13074 15314 13086
rect 18734 13074 18786 13086
rect 16818 13022 16830 13074
rect 16882 13022 16894 13074
rect 15262 13010 15314 13022
rect 18734 13010 18786 13022
rect 22318 13074 22370 13086
rect 22318 13010 22370 13022
rect 23102 13074 23154 13086
rect 23102 13010 23154 13022
rect 26574 13074 26626 13086
rect 26574 13010 26626 13022
rect 33070 13074 33122 13086
rect 56814 13074 56866 13086
rect 52994 13022 53006 13074
rect 53058 13022 53070 13074
rect 33070 13010 33122 13022
rect 56814 13010 56866 13022
rect 1710 12962 1762 12974
rect 1710 12898 1762 12910
rect 6638 12962 6690 12974
rect 6638 12898 6690 12910
rect 7422 12962 7474 12974
rect 7422 12898 7474 12910
rect 8654 12962 8706 12974
rect 8654 12898 8706 12910
rect 8878 12962 8930 12974
rect 8878 12898 8930 12910
rect 9102 12962 9154 12974
rect 11790 12962 11842 12974
rect 20750 12962 20802 12974
rect 10434 12910 10446 12962
rect 10498 12910 10510 12962
rect 11330 12910 11342 12962
rect 11394 12910 11406 12962
rect 15698 12910 15710 12962
rect 15762 12910 15774 12962
rect 17378 12910 17390 12962
rect 17442 12910 17454 12962
rect 9102 12898 9154 12910
rect 11790 12898 11842 12910
rect 20750 12898 20802 12910
rect 21758 12962 21810 12974
rect 21758 12898 21810 12910
rect 23214 12962 23266 12974
rect 25790 12962 25842 12974
rect 31166 12962 31218 12974
rect 38558 12962 38610 12974
rect 23650 12910 23662 12962
rect 23714 12910 23726 12962
rect 30482 12910 30494 12962
rect 30546 12910 30558 12962
rect 34626 12910 34638 12962
rect 34690 12910 34702 12962
rect 23214 12898 23266 12910
rect 25790 12898 25842 12910
rect 31166 12898 31218 12910
rect 38558 12898 38610 12910
rect 38782 12962 38834 12974
rect 46286 12962 46338 12974
rect 42690 12910 42702 12962
rect 42754 12910 42766 12962
rect 43698 12910 43710 12962
rect 43762 12910 43774 12962
rect 45154 12910 45166 12962
rect 45218 12910 45230 12962
rect 38782 12898 38834 12910
rect 46286 12898 46338 12910
rect 47070 12962 47122 12974
rect 47070 12898 47122 12910
rect 48638 12962 48690 12974
rect 50430 12962 50482 12974
rect 49746 12910 49758 12962
rect 49810 12910 49822 12962
rect 48638 12898 48690 12910
rect 50430 12898 50482 12910
rect 50654 12962 50706 12974
rect 50654 12898 50706 12910
rect 51886 12962 51938 12974
rect 51886 12898 51938 12910
rect 52222 12962 52274 12974
rect 55582 12962 55634 12974
rect 52658 12910 52670 12962
rect 52722 12910 52734 12962
rect 53554 12910 53566 12962
rect 53618 12910 53630 12962
rect 52222 12898 52274 12910
rect 55582 12898 55634 12910
rect 56142 12962 56194 12974
rect 56142 12898 56194 12910
rect 56366 12962 56418 12974
rect 56366 12898 56418 12910
rect 56926 12962 56978 12974
rect 56926 12898 56978 12910
rect 57262 12962 57314 12974
rect 57262 12898 57314 12910
rect 2046 12850 2098 12862
rect 2046 12786 2098 12798
rect 2382 12850 2434 12862
rect 2382 12786 2434 12798
rect 3502 12850 3554 12862
rect 3502 12786 3554 12798
rect 3614 12850 3666 12862
rect 3614 12786 3666 12798
rect 4510 12850 4562 12862
rect 4510 12786 4562 12798
rect 5966 12850 6018 12862
rect 5966 12786 6018 12798
rect 6862 12850 6914 12862
rect 9550 12850 9602 12862
rect 12126 12850 12178 12862
rect 39006 12850 39058 12862
rect 7074 12798 7086 12850
rect 7138 12798 7150 12850
rect 10098 12798 10110 12850
rect 10162 12798 10174 12850
rect 10546 12798 10558 12850
rect 10610 12798 10622 12850
rect 15586 12798 15598 12850
rect 15650 12798 15662 12850
rect 19058 12798 19070 12850
rect 19122 12798 19134 12850
rect 20402 12798 20414 12850
rect 20466 12798 20478 12850
rect 26898 12798 26910 12850
rect 26962 12798 26974 12850
rect 28354 12798 28366 12850
rect 28418 12798 28430 12850
rect 33506 12798 33518 12850
rect 33570 12798 33582 12850
rect 6862 12786 6914 12798
rect 9550 12786 9602 12798
rect 12126 12786 12178 12798
rect 39006 12786 39058 12798
rect 39118 12850 39170 12862
rect 39118 12786 39170 12798
rect 39790 12850 39842 12862
rect 39790 12786 39842 12798
rect 39902 12850 39954 12862
rect 39902 12786 39954 12798
rect 41694 12850 41746 12862
rect 44270 12850 44322 12862
rect 42466 12798 42478 12850
rect 42530 12798 42542 12850
rect 41694 12786 41746 12798
rect 44270 12786 44322 12798
rect 44830 12850 44882 12862
rect 44830 12786 44882 12798
rect 46174 12850 46226 12862
rect 48302 12850 48354 12862
rect 47282 12798 47294 12850
rect 47346 12798 47358 12850
rect 47842 12798 47854 12850
rect 47906 12798 47918 12850
rect 46174 12786 46226 12798
rect 48302 12786 48354 12798
rect 51998 12850 52050 12862
rect 55246 12850 55298 12862
rect 53106 12798 53118 12850
rect 53170 12798 53182 12850
rect 51998 12786 52050 12798
rect 55246 12786 55298 12798
rect 55806 12850 55858 12862
rect 55806 12786 55858 12798
rect 56702 12850 56754 12862
rect 56702 12786 56754 12798
rect 4958 12738 5010 12750
rect 2706 12686 2718 12738
rect 2770 12686 2782 12738
rect 4958 12674 5010 12686
rect 6302 12738 6354 12750
rect 6302 12674 6354 12686
rect 7646 12738 7698 12750
rect 7646 12674 7698 12686
rect 9774 12738 9826 12750
rect 12014 12738 12066 12750
rect 11442 12686 11454 12738
rect 11506 12686 11518 12738
rect 9774 12674 9826 12686
rect 12014 12674 12066 12686
rect 14702 12738 14754 12750
rect 14702 12674 14754 12686
rect 25902 12738 25954 12750
rect 38110 12738 38162 12750
rect 28466 12686 28478 12738
rect 28530 12686 28542 12738
rect 34738 12686 34750 12738
rect 34802 12686 34814 12738
rect 25902 12674 25954 12686
rect 38110 12674 38162 12686
rect 38222 12738 38274 12750
rect 38222 12674 38274 12686
rect 38446 12738 38498 12750
rect 38446 12674 38498 12686
rect 41358 12738 41410 12750
rect 41358 12674 41410 12686
rect 41582 12738 41634 12750
rect 41582 12674 41634 12686
rect 44942 12738 44994 12750
rect 44942 12674 44994 12686
rect 48414 12738 48466 12750
rect 48414 12674 48466 12686
rect 55358 12738 55410 12750
rect 55358 12674 55410 12686
rect 56030 12738 56082 12750
rect 56030 12674 56082 12686
rect 1344 12570 58576 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 50558 12570
rect 50610 12518 50662 12570
rect 50714 12518 50766 12570
rect 50818 12518 58576 12570
rect 1344 12484 58576 12518
rect 1710 12402 1762 12414
rect 1710 12338 1762 12350
rect 4622 12402 4674 12414
rect 4622 12338 4674 12350
rect 8542 12402 8594 12414
rect 8542 12338 8594 12350
rect 8654 12402 8706 12414
rect 8654 12338 8706 12350
rect 9662 12402 9714 12414
rect 9662 12338 9714 12350
rect 10446 12402 10498 12414
rect 10446 12338 10498 12350
rect 10670 12402 10722 12414
rect 10670 12338 10722 12350
rect 13806 12402 13858 12414
rect 13806 12338 13858 12350
rect 15374 12402 15426 12414
rect 19742 12402 19794 12414
rect 18498 12350 18510 12402
rect 18562 12350 18574 12402
rect 15374 12338 15426 12350
rect 19742 12338 19794 12350
rect 20862 12402 20914 12414
rect 20862 12338 20914 12350
rect 23438 12402 23490 12414
rect 23438 12338 23490 12350
rect 26910 12402 26962 12414
rect 31166 12402 31218 12414
rect 30146 12350 30158 12402
rect 30210 12350 30222 12402
rect 26910 12338 26962 12350
rect 31166 12338 31218 12350
rect 31950 12402 32002 12414
rect 31950 12338 32002 12350
rect 33070 12402 33122 12414
rect 38222 12402 38274 12414
rect 35970 12350 35982 12402
rect 36034 12350 36046 12402
rect 33070 12338 33122 12350
rect 38222 12338 38274 12350
rect 38894 12402 38946 12414
rect 38894 12338 38946 12350
rect 47294 12402 47346 12414
rect 47294 12338 47346 12350
rect 47518 12402 47570 12414
rect 47518 12338 47570 12350
rect 47966 12402 48018 12414
rect 47966 12338 48018 12350
rect 50094 12402 50146 12414
rect 52098 12350 52110 12402
rect 52162 12350 52174 12402
rect 50094 12338 50146 12350
rect 2718 12290 2770 12302
rect 2034 12238 2046 12290
rect 2098 12238 2110 12290
rect 2718 12226 2770 12238
rect 5518 12290 5570 12302
rect 5518 12226 5570 12238
rect 5854 12290 5906 12302
rect 5854 12226 5906 12238
rect 6526 12290 6578 12302
rect 6526 12226 6578 12238
rect 8318 12290 8370 12302
rect 8318 12226 8370 12238
rect 9886 12290 9938 12302
rect 9886 12226 9938 12238
rect 10334 12290 10386 12302
rect 10334 12226 10386 12238
rect 16382 12290 16434 12302
rect 19518 12290 19570 12302
rect 17938 12238 17950 12290
rect 18002 12238 18014 12290
rect 18274 12238 18286 12290
rect 18338 12238 18350 12290
rect 16382 12226 16434 12238
rect 19518 12226 19570 12238
rect 19966 12290 20018 12302
rect 19966 12226 20018 12238
rect 20078 12290 20130 12302
rect 20078 12226 20130 12238
rect 20750 12290 20802 12302
rect 20750 12226 20802 12238
rect 22318 12290 22370 12302
rect 30718 12290 30770 12302
rect 28466 12238 28478 12290
rect 28530 12238 28542 12290
rect 29810 12238 29822 12290
rect 29874 12238 29886 12290
rect 22318 12226 22370 12238
rect 30718 12226 30770 12238
rect 31390 12290 31442 12302
rect 31390 12226 31442 12238
rect 33294 12290 33346 12302
rect 49534 12290 49586 12302
rect 56590 12290 56642 12302
rect 35074 12238 35086 12290
rect 35138 12238 35150 12290
rect 52658 12238 52670 12290
rect 52722 12238 52734 12290
rect 55122 12238 55134 12290
rect 55186 12238 55198 12290
rect 33294 12226 33346 12238
rect 49534 12226 49586 12238
rect 56590 12226 56642 12238
rect 2382 12178 2434 12190
rect 6302 12178 6354 12190
rect 3490 12126 3502 12178
rect 3554 12126 3566 12178
rect 2382 12114 2434 12126
rect 6302 12114 6354 12126
rect 6414 12178 6466 12190
rect 7198 12178 7250 12190
rect 8766 12178 8818 12190
rect 9550 12178 9602 12190
rect 13918 12178 13970 12190
rect 6738 12126 6750 12178
rect 6802 12126 6814 12178
rect 7522 12126 7534 12178
rect 7586 12126 7598 12178
rect 8978 12126 8990 12178
rect 9042 12126 9054 12178
rect 11666 12126 11678 12178
rect 11730 12126 11742 12178
rect 6414 12114 6466 12126
rect 7198 12114 7250 12126
rect 8766 12114 8818 12126
rect 9550 12114 9602 12126
rect 13918 12114 13970 12126
rect 14366 12178 14418 12190
rect 14366 12114 14418 12126
rect 16270 12178 16322 12190
rect 16270 12114 16322 12126
rect 16494 12178 16546 12190
rect 16494 12114 16546 12126
rect 16942 12178 16994 12190
rect 19182 12178 19234 12190
rect 17714 12126 17726 12178
rect 17778 12126 17790 12178
rect 16942 12114 16994 12126
rect 19182 12114 19234 12126
rect 21086 12178 21138 12190
rect 23214 12178 23266 12190
rect 30606 12178 30658 12190
rect 31502 12178 31554 12190
rect 21858 12126 21870 12178
rect 21922 12126 21934 12178
rect 23762 12126 23774 12178
rect 23826 12126 23838 12178
rect 27122 12126 27134 12178
rect 27186 12126 27198 12178
rect 27458 12126 27470 12178
rect 27522 12126 27534 12178
rect 28242 12126 28254 12178
rect 28306 12126 28318 12178
rect 29586 12126 29598 12178
rect 29650 12126 29662 12178
rect 30930 12126 30942 12178
rect 30994 12126 31006 12178
rect 21086 12114 21138 12126
rect 23214 12114 23266 12126
rect 30606 12114 30658 12126
rect 31502 12114 31554 12126
rect 33406 12178 33458 12190
rect 33406 12114 33458 12126
rect 33854 12178 33906 12190
rect 33854 12114 33906 12126
rect 33966 12178 34018 12190
rect 33966 12114 34018 12126
rect 34078 12178 34130 12190
rect 36430 12178 36482 12190
rect 37214 12178 37266 12190
rect 43598 12178 43650 12190
rect 47630 12178 47682 12190
rect 34962 12126 34974 12178
rect 35026 12126 35038 12178
rect 35970 12126 35982 12178
rect 36034 12126 36046 12178
rect 36642 12126 36654 12178
rect 36706 12126 36718 12178
rect 37986 12126 37998 12178
rect 38050 12126 38062 12178
rect 38658 12126 38670 12178
rect 38722 12126 38734 12178
rect 39554 12126 39566 12178
rect 39618 12126 39630 12178
rect 42018 12126 42030 12178
rect 42082 12126 42094 12178
rect 42578 12126 42590 12178
rect 42642 12126 42654 12178
rect 44034 12126 44046 12178
rect 44098 12126 44110 12178
rect 44594 12126 44606 12178
rect 44658 12126 44670 12178
rect 45154 12126 45166 12178
rect 45218 12126 45230 12178
rect 34078 12114 34130 12126
rect 36430 12114 36482 12126
rect 37214 12114 37266 12126
rect 43598 12114 43650 12126
rect 47630 12114 47682 12126
rect 48078 12178 48130 12190
rect 48078 12114 48130 12126
rect 49982 12178 50034 12190
rect 49982 12114 50034 12126
rect 50206 12178 50258 12190
rect 50206 12114 50258 12126
rect 50654 12178 50706 12190
rect 50654 12114 50706 12126
rect 51438 12178 51490 12190
rect 51874 12126 51886 12178
rect 51938 12126 51950 12178
rect 53778 12126 53790 12178
rect 53842 12126 53854 12178
rect 55682 12126 55694 12178
rect 55746 12126 55758 12178
rect 57026 12126 57038 12178
rect 57090 12126 57102 12178
rect 51438 12114 51490 12126
rect 5182 12066 5234 12078
rect 3826 12014 3838 12066
rect 3890 12014 3902 12066
rect 5182 12002 5234 12014
rect 7982 12066 8034 12078
rect 12350 12066 12402 12078
rect 23326 12066 23378 12078
rect 47070 12066 47122 12078
rect 11554 12014 11566 12066
rect 11618 12014 11630 12066
rect 15810 12014 15822 12066
rect 15874 12014 15886 12066
rect 21410 12014 21422 12066
rect 21474 12014 21486 12066
rect 28130 12014 28142 12066
rect 28194 12014 28206 12066
rect 39778 12014 39790 12066
rect 39842 12014 39854 12066
rect 42466 12014 42478 12066
rect 42530 12014 42542 12066
rect 45042 12014 45054 12066
rect 45106 12014 45118 12066
rect 49634 12014 49646 12066
rect 49698 12014 49710 12066
rect 50978 12014 50990 12066
rect 51042 12014 51054 12066
rect 57362 12014 57374 12066
rect 57426 12014 57438 12066
rect 7982 12002 8034 12014
rect 12350 12002 12402 12014
rect 23326 12002 23378 12014
rect 47070 12002 47122 12014
rect 13806 11954 13858 11966
rect 13806 11890 13858 11902
rect 14254 11954 14306 11966
rect 14254 11890 14306 11902
rect 26798 11954 26850 11966
rect 49310 11954 49362 11966
rect 34514 11902 34526 11954
rect 34578 11902 34590 11954
rect 40002 11902 40014 11954
rect 40066 11902 40078 11954
rect 42914 11902 42926 11954
rect 42978 11902 42990 11954
rect 45266 11902 45278 11954
rect 45330 11902 45342 11954
rect 26798 11890 26850 11902
rect 49310 11890 49362 11902
rect 1344 11786 58576 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 58576 11786
rect 1344 11700 58576 11734
rect 16382 11618 16434 11630
rect 35646 11618 35698 11630
rect 6290 11566 6302 11618
rect 6354 11566 6366 11618
rect 14466 11566 14478 11618
rect 14530 11566 14542 11618
rect 18722 11566 18734 11618
rect 18786 11566 18798 11618
rect 27458 11566 27470 11618
rect 27522 11566 27534 11618
rect 16382 11554 16434 11566
rect 35646 11554 35698 11566
rect 35982 11618 36034 11630
rect 35982 11554 36034 11566
rect 39566 11618 39618 11630
rect 39566 11554 39618 11566
rect 42254 11618 42306 11630
rect 53554 11566 53566 11618
rect 53618 11566 53630 11618
rect 42254 11554 42306 11566
rect 4622 11506 4674 11518
rect 9214 11506 9266 11518
rect 4946 11454 4958 11506
rect 5010 11454 5022 11506
rect 4622 11442 4674 11454
rect 9214 11442 9266 11454
rect 11902 11506 11954 11518
rect 15934 11506 15986 11518
rect 14354 11454 14366 11506
rect 14418 11454 14430 11506
rect 11902 11442 11954 11454
rect 15934 11442 15986 11454
rect 21534 11506 21586 11518
rect 21534 11442 21586 11454
rect 26798 11506 26850 11518
rect 26798 11442 26850 11454
rect 33182 11506 33234 11518
rect 33182 11442 33234 11454
rect 38446 11506 38498 11518
rect 38446 11442 38498 11454
rect 40686 11506 40738 11518
rect 47630 11506 47682 11518
rect 41570 11454 41582 11506
rect 41634 11454 41646 11506
rect 55570 11454 55582 11506
rect 55634 11454 55646 11506
rect 40686 11442 40738 11454
rect 47630 11442 47682 11454
rect 3726 11394 3778 11406
rect 12798 11394 12850 11406
rect 15486 11394 15538 11406
rect 2818 11342 2830 11394
rect 2882 11342 2894 11394
rect 5618 11342 5630 11394
rect 5682 11342 5694 11394
rect 6402 11342 6414 11394
rect 6466 11342 6478 11394
rect 6850 11342 6862 11394
rect 6914 11342 6926 11394
rect 9986 11342 9998 11394
rect 10050 11342 10062 11394
rect 10882 11342 10894 11394
rect 10946 11342 10958 11394
rect 12562 11342 12574 11394
rect 12626 11342 12638 11394
rect 14018 11342 14030 11394
rect 14082 11342 14094 11394
rect 3726 11330 3778 11342
rect 12798 11330 12850 11342
rect 15486 11330 15538 11342
rect 15710 11394 15762 11406
rect 27134 11394 27186 11406
rect 33294 11394 33346 11406
rect 35870 11394 35922 11406
rect 17154 11342 17166 11394
rect 17218 11342 17230 11394
rect 17714 11342 17726 11394
rect 17778 11342 17790 11394
rect 18498 11342 18510 11394
rect 18562 11342 18574 11394
rect 19170 11342 19182 11394
rect 19234 11342 19246 11394
rect 20290 11342 20302 11394
rect 20354 11342 20366 11394
rect 22866 11342 22878 11394
rect 22930 11342 22942 11394
rect 25442 11342 25454 11394
rect 25506 11342 25518 11394
rect 27794 11342 27806 11394
rect 27858 11342 27870 11394
rect 28578 11342 28590 11394
rect 28642 11342 28654 11394
rect 33954 11342 33966 11394
rect 34018 11342 34030 11394
rect 35074 11342 35086 11394
rect 35138 11342 35150 11394
rect 35410 11342 35422 11394
rect 35474 11342 35486 11394
rect 15710 11330 15762 11342
rect 27134 11330 27186 11342
rect 33294 11330 33346 11342
rect 35870 11330 35922 11342
rect 37550 11394 37602 11406
rect 39902 11394 39954 11406
rect 37874 11342 37886 11394
rect 37938 11342 37950 11394
rect 37550 11330 37602 11342
rect 39902 11330 39954 11342
rect 40238 11394 40290 11406
rect 49870 11394 49922 11406
rect 41346 11342 41358 11394
rect 41410 11342 41422 11394
rect 42018 11342 42030 11394
rect 42082 11342 42094 11394
rect 45826 11342 45838 11394
rect 45890 11342 45902 11394
rect 40238 11330 40290 11342
rect 49870 11330 49922 11342
rect 50430 11394 50482 11406
rect 50430 11330 50482 11342
rect 51886 11394 51938 11406
rect 53566 11394 53618 11406
rect 53330 11342 53342 11394
rect 53394 11342 53406 11394
rect 51886 11330 51938 11342
rect 53566 11330 53618 11342
rect 1710 11282 1762 11294
rect 1710 11218 1762 11230
rect 3390 11282 3442 11294
rect 11342 11282 11394 11294
rect 4274 11230 4286 11282
rect 4338 11230 4350 11282
rect 5730 11230 5742 11282
rect 5794 11230 5806 11282
rect 9762 11230 9774 11282
rect 9826 11230 9838 11282
rect 3390 11218 3442 11230
rect 11342 11218 11394 11230
rect 11454 11282 11506 11294
rect 29038 11282 29090 11294
rect 16818 11230 16830 11282
rect 16882 11230 16894 11282
rect 21634 11230 21646 11282
rect 21698 11230 21710 11282
rect 25106 11230 25118 11282
rect 25170 11230 25182 11282
rect 26562 11230 26574 11282
rect 26626 11230 26638 11282
rect 27346 11230 27358 11282
rect 27410 11230 27422 11282
rect 11454 11218 11506 11230
rect 29038 11218 29090 11230
rect 29262 11282 29314 11294
rect 29262 11218 29314 11230
rect 29374 11282 29426 11294
rect 33630 11282 33682 11294
rect 38782 11282 38834 11294
rect 30930 11230 30942 11282
rect 30994 11230 31006 11282
rect 34178 11230 34190 11282
rect 34242 11230 34254 11282
rect 29374 11218 29426 11230
rect 33630 11218 33682 11230
rect 38782 11218 38834 11230
rect 39118 11282 39170 11294
rect 39118 11218 39170 11230
rect 39566 11282 39618 11294
rect 39566 11218 39618 11230
rect 39678 11282 39730 11294
rect 39678 11218 39730 11230
rect 40574 11282 40626 11294
rect 40574 11218 40626 11230
rect 43262 11282 43314 11294
rect 43262 11218 43314 11230
rect 43598 11282 43650 11294
rect 47966 11282 48018 11294
rect 45602 11230 45614 11282
rect 45666 11230 45678 11282
rect 43598 11218 43650 11230
rect 47966 11218 48018 11230
rect 50318 11282 50370 11294
rect 50318 11218 50370 11230
rect 52222 11282 52274 11294
rect 52222 11218 52274 11230
rect 55134 11282 55186 11294
rect 55794 11230 55806 11282
rect 55858 11230 55870 11282
rect 57474 11230 57486 11282
rect 57538 11230 57550 11282
rect 55134 11218 55186 11230
rect 2046 11170 2098 11182
rect 3502 11170 3554 11182
rect 3042 11118 3054 11170
rect 3106 11118 3118 11170
rect 2046 11106 2098 11118
rect 3502 11106 3554 11118
rect 3950 11170 4002 11182
rect 3950 11106 4002 11118
rect 4846 11170 4898 11182
rect 11118 11170 11170 11182
rect 29822 11170 29874 11182
rect 10770 11118 10782 11170
rect 10834 11118 10846 11170
rect 17602 11118 17614 11170
rect 17666 11118 17678 11170
rect 23202 11118 23214 11170
rect 23266 11118 23278 11170
rect 4846 11106 4898 11118
rect 11118 11106 11170 11118
rect 29822 11106 29874 11118
rect 30270 11170 30322 11182
rect 30270 11106 30322 11118
rect 31278 11170 31330 11182
rect 31278 11106 31330 11118
rect 33518 11170 33570 11182
rect 40126 11170 40178 11182
rect 34962 11118 34974 11170
rect 35026 11118 35038 11170
rect 33518 11106 33570 11118
rect 40126 11106 40178 11118
rect 43374 11170 43426 11182
rect 43374 11106 43426 11118
rect 45390 11170 45442 11182
rect 45390 11106 45442 11118
rect 48078 11170 48130 11182
rect 48078 11106 48130 11118
rect 48302 11170 48354 11182
rect 48302 11106 48354 11118
rect 50206 11170 50258 11182
rect 50206 11106 50258 11118
rect 51662 11170 51714 11182
rect 51662 11106 51714 11118
rect 51998 11170 52050 11182
rect 51998 11106 52050 11118
rect 54574 11170 54626 11182
rect 54574 11106 54626 11118
rect 54686 11170 54738 11182
rect 54686 11106 54738 11118
rect 54910 11170 54962 11182
rect 57362 11118 57374 11170
rect 57426 11118 57438 11170
rect 54910 11106 54962 11118
rect 1344 11002 58576 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 50558 11002
rect 50610 10950 50662 11002
rect 50714 10950 50766 11002
rect 50818 10950 58576 11002
rect 1344 10916 58576 10950
rect 1822 10834 1874 10846
rect 3502 10834 3554 10846
rect 13918 10834 13970 10846
rect 3154 10782 3166 10834
rect 3218 10782 3230 10834
rect 3826 10782 3838 10834
rect 3890 10782 3902 10834
rect 1822 10770 1874 10782
rect 3502 10770 3554 10782
rect 13918 10770 13970 10782
rect 14478 10834 14530 10846
rect 14478 10770 14530 10782
rect 16382 10834 16434 10846
rect 16382 10770 16434 10782
rect 20414 10834 20466 10846
rect 20414 10770 20466 10782
rect 23550 10834 23602 10846
rect 28254 10834 28306 10846
rect 28018 10782 28030 10834
rect 28082 10782 28094 10834
rect 23550 10770 23602 10782
rect 28254 10770 28306 10782
rect 28478 10834 28530 10846
rect 28478 10770 28530 10782
rect 29598 10834 29650 10846
rect 36654 10834 36706 10846
rect 34178 10782 34190 10834
rect 34242 10782 34254 10834
rect 29598 10770 29650 10782
rect 36654 10770 36706 10782
rect 37886 10834 37938 10846
rect 37886 10770 37938 10782
rect 38110 10834 38162 10846
rect 41806 10834 41858 10846
rect 56702 10834 56754 10846
rect 39890 10782 39902 10834
rect 39954 10782 39966 10834
rect 53218 10782 53230 10834
rect 53282 10782 53294 10834
rect 38110 10770 38162 10782
rect 41806 10770 41858 10782
rect 56702 10770 56754 10782
rect 7758 10722 7810 10734
rect 2482 10670 2494 10722
rect 2546 10670 2558 10722
rect 4498 10670 4510 10722
rect 4562 10670 4574 10722
rect 5058 10670 5070 10722
rect 5122 10670 5134 10722
rect 7758 10658 7810 10670
rect 9662 10722 9714 10734
rect 19966 10722 20018 10734
rect 32510 10722 32562 10734
rect 35086 10722 35138 10734
rect 11106 10670 11118 10722
rect 11170 10670 11182 10722
rect 27122 10670 27134 10722
rect 27186 10670 27198 10722
rect 30594 10670 30606 10722
rect 30658 10670 30670 10722
rect 33954 10670 33966 10722
rect 34018 10670 34030 10722
rect 34514 10670 34526 10722
rect 34578 10670 34590 10722
rect 9662 10658 9714 10670
rect 19966 10658 20018 10670
rect 32510 10658 32562 10670
rect 35086 10658 35138 10670
rect 36766 10722 36818 10734
rect 36766 10658 36818 10670
rect 38222 10722 38274 10734
rect 41022 10722 41074 10734
rect 39106 10670 39118 10722
rect 39170 10670 39182 10722
rect 38222 10658 38274 10670
rect 41022 10658 41074 10670
rect 41582 10722 41634 10734
rect 41582 10658 41634 10670
rect 44494 10722 44546 10734
rect 44494 10658 44546 10670
rect 47742 10722 47794 10734
rect 47742 10658 47794 10670
rect 48750 10722 48802 10734
rect 48750 10658 48802 10670
rect 51102 10722 51154 10734
rect 52322 10670 52334 10722
rect 52386 10670 52398 10722
rect 55682 10670 55694 10722
rect 55746 10670 55758 10722
rect 51102 10658 51154 10670
rect 2830 10610 2882 10622
rect 7982 10610 8034 10622
rect 2258 10558 2270 10610
rect 2322 10558 2334 10610
rect 4274 10558 4286 10610
rect 4338 10558 4350 10610
rect 5282 10558 5294 10610
rect 5346 10558 5358 10610
rect 5842 10558 5854 10610
rect 5906 10558 5918 10610
rect 6402 10558 6414 10610
rect 6466 10558 6478 10610
rect 2830 10546 2882 10558
rect 7982 10546 8034 10558
rect 9774 10610 9826 10622
rect 9774 10546 9826 10558
rect 9886 10610 9938 10622
rect 14590 10610 14642 10622
rect 27470 10610 27522 10622
rect 11218 10558 11230 10610
rect 11282 10558 11294 10610
rect 12450 10558 12462 10610
rect 12514 10558 12526 10610
rect 17826 10558 17838 10610
rect 17890 10558 17902 10610
rect 19170 10558 19182 10610
rect 19234 10558 19246 10610
rect 22306 10558 22318 10610
rect 22370 10558 22382 10610
rect 25666 10558 25678 10610
rect 25730 10558 25742 10610
rect 26450 10558 26462 10610
rect 26514 10558 26526 10610
rect 9886 10546 9938 10558
rect 14590 10546 14642 10558
rect 27470 10546 27522 10558
rect 28590 10610 28642 10622
rect 28590 10546 28642 10558
rect 29934 10610 29986 10622
rect 38782 10610 38834 10622
rect 40238 10610 40290 10622
rect 31154 10558 31166 10610
rect 31218 10558 31230 10610
rect 32050 10558 32062 10610
rect 32114 10558 32126 10610
rect 33618 10558 33630 10610
rect 33682 10558 33694 10610
rect 35970 10558 35982 10610
rect 36034 10558 36046 10610
rect 39330 10558 39342 10610
rect 39394 10558 39406 10610
rect 29934 10546 29986 10558
rect 38782 10546 38834 10558
rect 40238 10546 40290 10558
rect 40910 10610 40962 10622
rect 40910 10546 40962 10558
rect 41246 10610 41298 10622
rect 41246 10546 41298 10558
rect 41470 10610 41522 10622
rect 47518 10610 47570 10622
rect 43586 10558 43598 10610
rect 43650 10558 43662 10610
rect 46050 10558 46062 10610
rect 46114 10558 46126 10610
rect 41470 10546 41522 10558
rect 47518 10546 47570 10558
rect 47966 10610 48018 10622
rect 47966 10546 48018 10558
rect 48190 10610 48242 10622
rect 53678 10610 53730 10622
rect 49186 10558 49198 10610
rect 49250 10558 49262 10610
rect 51538 10558 51550 10610
rect 51602 10558 51614 10610
rect 52210 10558 52222 10610
rect 52274 10558 52286 10610
rect 53330 10558 53342 10610
rect 53394 10558 53406 10610
rect 48190 10546 48242 10558
rect 53678 10546 53730 10558
rect 53902 10610 53954 10622
rect 56478 10610 56530 10622
rect 54562 10558 54574 10610
rect 54626 10558 54638 10610
rect 55570 10558 55582 10610
rect 55634 10558 55646 10610
rect 55906 10558 55918 10610
rect 55970 10558 55982 10610
rect 53902 10546 53954 10558
rect 56478 10546 56530 10558
rect 56814 10610 56866 10622
rect 56814 10546 56866 10558
rect 57038 10610 57090 10622
rect 57038 10546 57090 10558
rect 14926 10498 14978 10510
rect 27694 10498 27746 10510
rect 8978 10446 8990 10498
rect 9042 10446 9054 10498
rect 11890 10446 11902 10498
rect 11954 10446 11966 10498
rect 14018 10446 14030 10498
rect 14082 10446 14094 10498
rect 16482 10446 16494 10498
rect 16546 10446 16558 10498
rect 17714 10446 17726 10498
rect 17778 10446 17790 10498
rect 22754 10446 22766 10498
rect 22818 10446 22830 10498
rect 26338 10446 26350 10498
rect 26402 10446 26414 10498
rect 14926 10434 14978 10446
rect 27694 10434 27746 10446
rect 29150 10498 29202 10510
rect 43038 10498 43090 10510
rect 45726 10498 45778 10510
rect 35858 10446 35870 10498
rect 35922 10446 35934 10498
rect 43474 10446 43486 10498
rect 43538 10446 43550 10498
rect 46386 10446 46398 10498
rect 46450 10446 46462 10498
rect 49634 10446 49646 10498
rect 49698 10446 49710 10498
rect 54226 10446 54238 10498
rect 54290 10446 54302 10498
rect 29150 10434 29202 10446
rect 43038 10434 43090 10446
rect 45726 10434 45778 10446
rect 8206 10386 8258 10398
rect 6178 10334 6190 10386
rect 6242 10334 6254 10386
rect 8206 10322 8258 10334
rect 8430 10386 8482 10398
rect 13694 10386 13746 10398
rect 10322 10334 10334 10386
rect 10386 10334 10398 10386
rect 8430 10322 8482 10334
rect 13694 10322 13746 10334
rect 14478 10386 14530 10398
rect 14478 10322 14530 10334
rect 15038 10386 15090 10398
rect 15038 10322 15090 10334
rect 16158 10386 16210 10398
rect 16158 10322 16210 10334
rect 36542 10386 36594 10398
rect 36542 10322 36594 10334
rect 44382 10386 44434 10398
rect 44382 10322 44434 10334
rect 1344 10218 58576 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 58576 10218
rect 1344 10132 58576 10166
rect 11790 10050 11842 10062
rect 11790 9986 11842 9998
rect 12126 10050 12178 10062
rect 12126 9986 12178 9998
rect 26462 10050 26514 10062
rect 26462 9986 26514 9998
rect 30606 10050 30658 10062
rect 30606 9986 30658 9998
rect 31166 10050 31218 10062
rect 31166 9986 31218 9998
rect 55022 10050 55074 10062
rect 57474 9998 57486 10050
rect 57538 9998 57550 10050
rect 55022 9986 55074 9998
rect 6750 9938 6802 9950
rect 12350 9938 12402 9950
rect 23326 9938 23378 9950
rect 4946 9886 4958 9938
rect 5010 9886 5022 9938
rect 9538 9886 9550 9938
rect 9602 9886 9614 9938
rect 14354 9886 14366 9938
rect 14418 9886 14430 9938
rect 15026 9886 15038 9938
rect 15090 9886 15102 9938
rect 6750 9874 6802 9886
rect 12350 9874 12402 9886
rect 23326 9874 23378 9886
rect 25566 9938 25618 9950
rect 25566 9874 25618 9886
rect 37102 9938 37154 9950
rect 42590 9938 42642 9950
rect 44046 9938 44098 9950
rect 38322 9886 38334 9938
rect 38386 9886 38398 9938
rect 43026 9886 43038 9938
rect 43090 9886 43102 9938
rect 37102 9874 37154 9886
rect 42590 9874 42642 9886
rect 44046 9874 44098 9886
rect 45278 9938 45330 9950
rect 45278 9874 45330 9886
rect 50430 9938 50482 9950
rect 54126 9938 54178 9950
rect 53330 9886 53342 9938
rect 53394 9886 53406 9938
rect 55570 9886 55582 9938
rect 55634 9886 55646 9938
rect 50430 9874 50482 9886
rect 54126 9874 54178 9886
rect 1710 9826 1762 9838
rect 1710 9762 1762 9774
rect 3278 9826 3330 9838
rect 8206 9826 8258 9838
rect 17614 9826 17666 9838
rect 20414 9826 20466 9838
rect 4162 9774 4174 9826
rect 4226 9774 4238 9826
rect 4834 9774 4846 9826
rect 4898 9774 4910 9826
rect 6290 9774 6302 9826
rect 6354 9774 6366 9826
rect 6962 9774 6974 9826
rect 7026 9774 7038 9826
rect 8418 9774 8430 9826
rect 8482 9774 8494 9826
rect 9314 9774 9326 9826
rect 9378 9774 9390 9826
rect 10322 9774 10334 9826
rect 10386 9774 10398 9826
rect 13794 9774 13806 9826
rect 13858 9774 13870 9826
rect 14018 9774 14030 9826
rect 14082 9774 14094 9826
rect 15138 9774 15150 9826
rect 15202 9774 15214 9826
rect 19058 9774 19070 9826
rect 19122 9774 19134 9826
rect 19730 9774 19742 9826
rect 19794 9774 19806 9826
rect 3278 9762 3330 9774
rect 8206 9762 8258 9774
rect 17614 9762 17666 9774
rect 20414 9762 20466 9774
rect 21422 9826 21474 9838
rect 23774 9826 23826 9838
rect 21522 9774 21534 9826
rect 21586 9774 21598 9826
rect 21422 9762 21474 9774
rect 23774 9762 23826 9774
rect 25790 9826 25842 9838
rect 25790 9762 25842 9774
rect 26014 9826 26066 9838
rect 29710 9826 29762 9838
rect 29250 9774 29262 9826
rect 29314 9774 29326 9826
rect 26014 9762 26066 9774
rect 29710 9762 29762 9774
rect 32062 9826 32114 9838
rect 32062 9762 32114 9774
rect 35646 9826 35698 9838
rect 35646 9762 35698 9774
rect 35982 9826 36034 9838
rect 35982 9762 36034 9774
rect 36542 9826 36594 9838
rect 37886 9826 37938 9838
rect 37650 9774 37662 9826
rect 37714 9774 37726 9826
rect 36542 9762 36594 9774
rect 37886 9762 37938 9774
rect 38446 9826 38498 9838
rect 38446 9762 38498 9774
rect 38670 9826 38722 9838
rect 47182 9826 47234 9838
rect 50542 9826 50594 9838
rect 51774 9826 51826 9838
rect 39890 9774 39902 9826
rect 39954 9774 39966 9826
rect 40786 9774 40798 9826
rect 40850 9774 40862 9826
rect 43138 9774 43150 9826
rect 43202 9774 43214 9826
rect 44258 9774 44270 9826
rect 44322 9774 44334 9826
rect 48514 9774 48526 9826
rect 48578 9774 48590 9826
rect 50978 9774 50990 9826
rect 51042 9774 51054 9826
rect 38670 9762 38722 9774
rect 47182 9762 47234 9774
rect 50542 9762 50594 9774
rect 51774 9762 51826 9774
rect 52110 9826 52162 9838
rect 54350 9826 54402 9838
rect 52658 9774 52670 9826
rect 52722 9774 52734 9826
rect 53666 9774 53678 9826
rect 53730 9774 53742 9826
rect 52110 9762 52162 9774
rect 54350 9762 54402 9774
rect 54574 9826 54626 9838
rect 56018 9774 56030 9826
rect 56082 9774 56094 9826
rect 57138 9774 57150 9826
rect 57202 9774 57214 9826
rect 54574 9762 54626 9774
rect 2046 9714 2098 9726
rect 2046 9650 2098 9662
rect 2718 9714 2770 9726
rect 2718 9650 2770 9662
rect 3838 9714 3890 9726
rect 14814 9714 14866 9726
rect 4946 9662 4958 9714
rect 5010 9662 5022 9714
rect 6178 9662 6190 9714
rect 6242 9662 6254 9714
rect 6738 9662 6750 9714
rect 6802 9662 6814 9714
rect 9650 9662 9662 9714
rect 9714 9662 9726 9714
rect 10434 9662 10446 9714
rect 10498 9662 10510 9714
rect 10994 9662 11006 9714
rect 11058 9662 11070 9714
rect 3838 9650 3890 9662
rect 14814 9650 14866 9662
rect 17726 9714 17778 9726
rect 23214 9714 23266 9726
rect 18722 9662 18734 9714
rect 18786 9662 18798 9714
rect 17726 9650 17778 9662
rect 23214 9650 23266 9662
rect 23550 9714 23602 9726
rect 30718 9714 30770 9726
rect 28578 9662 28590 9714
rect 28642 9662 28654 9714
rect 23550 9650 23602 9662
rect 30718 9650 30770 9662
rect 31054 9714 31106 9726
rect 31054 9650 31106 9662
rect 31726 9714 31778 9726
rect 31726 9650 31778 9662
rect 31838 9714 31890 9726
rect 31838 9650 31890 9662
rect 34750 9714 34802 9726
rect 34750 9650 34802 9662
rect 34974 9714 35026 9726
rect 34974 9650 35026 9662
rect 35310 9714 35362 9726
rect 35310 9650 35362 9662
rect 36206 9714 36258 9726
rect 36206 9650 36258 9662
rect 36318 9714 36370 9726
rect 36318 9650 36370 9662
rect 38894 9714 38946 9726
rect 43934 9714 43986 9726
rect 40114 9662 40126 9714
rect 40178 9662 40190 9714
rect 41682 9662 41694 9714
rect 41746 9662 41758 9714
rect 38894 9650 38946 9662
rect 43934 9650 43986 9662
rect 45614 9714 45666 9726
rect 45614 9650 45666 9662
rect 45726 9714 45778 9726
rect 45726 9650 45778 9662
rect 46846 9714 46898 9726
rect 51886 9714 51938 9726
rect 48178 9662 48190 9714
rect 48242 9662 48254 9714
rect 49858 9662 49870 9714
rect 49922 9662 49934 9714
rect 52770 9662 52782 9714
rect 52834 9662 52846 9714
rect 46846 9650 46898 9662
rect 51886 9650 51938 9662
rect 17950 9602 18002 9614
rect 11106 9550 11118 9602
rect 11170 9550 11182 9602
rect 17950 9538 18002 9550
rect 22766 9602 22818 9614
rect 22766 9538 22818 9550
rect 27918 9602 27970 9614
rect 27918 9538 27970 9550
rect 28254 9602 28306 9614
rect 28254 9538 28306 9550
rect 30606 9602 30658 9614
rect 30606 9538 30658 9550
rect 31166 9602 31218 9614
rect 31166 9538 31218 9550
rect 34414 9602 34466 9614
rect 34414 9538 34466 9550
rect 35086 9602 35138 9614
rect 35086 9538 35138 9550
rect 35758 9602 35810 9614
rect 35758 9538 35810 9550
rect 38334 9602 38386 9614
rect 38334 9538 38386 9550
rect 39342 9602 39394 9614
rect 41358 9602 41410 9614
rect 40898 9550 40910 9602
rect 40962 9550 40974 9602
rect 39342 9538 39394 9550
rect 41358 9538 41410 9550
rect 45950 9602 46002 9614
rect 45950 9538 46002 9550
rect 46174 9602 46226 9614
rect 46958 9602 47010 9614
rect 46498 9550 46510 9602
rect 46562 9550 46574 9602
rect 49746 9550 49758 9602
rect 49810 9550 49822 9602
rect 46174 9538 46226 9550
rect 46958 9538 47010 9550
rect 1344 9434 58576 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 50558 9434
rect 50610 9382 50662 9434
rect 50714 9382 50766 9434
rect 50818 9382 58576 9434
rect 1344 9348 58576 9382
rect 3166 9266 3218 9278
rect 2706 9214 2718 9266
rect 2770 9214 2782 9266
rect 3166 9202 3218 9214
rect 5406 9266 5458 9278
rect 8654 9266 8706 9278
rect 20974 9266 21026 9278
rect 6626 9214 6638 9266
rect 6690 9214 6702 9266
rect 7298 9214 7310 9266
rect 7362 9214 7374 9266
rect 9874 9214 9886 9266
rect 9938 9214 9950 9266
rect 5406 9202 5458 9214
rect 8654 9202 8706 9214
rect 14702 9210 14754 9222
rect 1710 9154 1762 9166
rect 1710 9090 1762 9102
rect 2046 9154 2098 9166
rect 2046 9090 2098 9102
rect 4286 9154 4338 9166
rect 5294 9154 5346 9166
rect 4498 9102 4510 9154
rect 4562 9102 4574 9154
rect 4286 9090 4338 9102
rect 5294 9090 5346 9102
rect 7758 9154 7810 9166
rect 13918 9154 13970 9166
rect 11330 9102 11342 9154
rect 11394 9102 11406 9154
rect 12226 9102 12238 9154
rect 12290 9102 12302 9154
rect 7758 9090 7810 9102
rect 13918 9090 13970 9102
rect 14590 9154 14642 9166
rect 20974 9202 21026 9214
rect 22318 9266 22370 9278
rect 35198 9266 35250 9278
rect 34738 9214 34750 9266
rect 34802 9214 34814 9266
rect 22318 9202 22370 9214
rect 35198 9202 35250 9214
rect 35534 9266 35586 9278
rect 38894 9266 38946 9278
rect 36866 9214 36878 9266
rect 36930 9214 36942 9266
rect 38434 9214 38446 9266
rect 38498 9214 38510 9266
rect 35534 9202 35586 9214
rect 38894 9202 38946 9214
rect 40238 9266 40290 9278
rect 40238 9202 40290 9214
rect 40462 9266 40514 9278
rect 40462 9202 40514 9214
rect 47518 9266 47570 9278
rect 47518 9202 47570 9214
rect 48078 9266 48130 9278
rect 48078 9202 48130 9214
rect 51774 9266 51826 9278
rect 51774 9202 51826 9214
rect 52334 9266 52386 9278
rect 52334 9202 52386 9214
rect 53454 9266 53506 9278
rect 53454 9202 53506 9214
rect 53566 9266 53618 9278
rect 53566 9202 53618 9214
rect 54238 9266 54290 9278
rect 54238 9202 54290 9214
rect 55694 9266 55746 9278
rect 55694 9202 55746 9214
rect 14702 9146 14754 9158
rect 20862 9154 20914 9166
rect 15474 9102 15486 9154
rect 15538 9102 15550 9154
rect 19842 9102 19854 9154
rect 19906 9102 19918 9154
rect 14590 9090 14642 9102
rect 20862 9090 20914 9102
rect 21198 9154 21250 9166
rect 21198 9090 21250 9102
rect 21982 9154 22034 9166
rect 21982 9090 22034 9102
rect 22094 9154 22146 9166
rect 22094 9090 22146 9102
rect 26350 9154 26402 9166
rect 26350 9090 26402 9102
rect 26798 9154 26850 9166
rect 26798 9090 26850 9102
rect 32286 9154 32338 9166
rect 32286 9090 32338 9102
rect 35310 9154 35362 9166
rect 35310 9090 35362 9102
rect 35982 9154 36034 9166
rect 35982 9090 36034 9102
rect 36542 9154 36594 9166
rect 36542 9090 36594 9102
rect 40126 9154 40178 9166
rect 40126 9090 40178 9102
rect 42926 9154 42978 9166
rect 42926 9090 42978 9102
rect 43038 9154 43090 9166
rect 43038 9090 43090 9102
rect 47182 9154 47234 9166
rect 47182 9090 47234 9102
rect 47294 9154 47346 9166
rect 47294 9090 47346 9102
rect 47854 9154 47906 9166
rect 47854 9090 47906 9102
rect 52894 9154 52946 9166
rect 52894 9090 52946 9102
rect 55918 9154 55970 9166
rect 55918 9090 55970 9102
rect 2382 9042 2434 9054
rect 2382 8978 2434 8990
rect 4174 9042 4226 9054
rect 5070 9042 5122 9054
rect 4610 8990 4622 9042
rect 4674 8990 4686 9042
rect 4174 8978 4226 8990
rect 5070 8978 5122 8990
rect 5630 9042 5682 9054
rect 14926 9042 14978 9054
rect 31390 9042 31442 9054
rect 35086 9042 35138 9054
rect 6402 8990 6414 9042
rect 6466 8990 6478 9042
rect 7074 8990 7086 9042
rect 7138 8990 7150 9042
rect 8082 8990 8094 9042
rect 8146 8990 8158 9042
rect 9650 8990 9662 9042
rect 9714 8990 9726 9042
rect 10210 8990 10222 9042
rect 10274 8990 10286 9042
rect 11106 8990 11118 9042
rect 11170 8990 11182 9042
rect 13234 8990 13246 9042
rect 13298 8990 13310 9042
rect 15138 8990 15150 9042
rect 15202 8990 15214 9042
rect 16258 8990 16270 9042
rect 16322 8990 16334 9042
rect 17938 8990 17950 9042
rect 18002 8990 18014 9042
rect 19282 8990 19294 9042
rect 19346 8990 19358 9042
rect 25890 8990 25902 9042
rect 25954 8990 25966 9042
rect 27570 8990 27582 9042
rect 27634 8990 27646 9042
rect 28578 8990 28590 9042
rect 28642 8990 28654 9042
rect 31602 8990 31614 9042
rect 31666 8990 31678 9042
rect 5630 8978 5682 8990
rect 14926 8978 14978 8990
rect 31390 8978 31442 8990
rect 35086 8978 35138 8990
rect 36094 9042 36146 9054
rect 39230 9042 39282 9054
rect 38210 8990 38222 9042
rect 38274 8990 38286 9042
rect 36094 8978 36146 8990
rect 39230 8978 39282 8990
rect 39790 9042 39842 9054
rect 39790 8978 39842 8990
rect 43598 9042 43650 9054
rect 47742 9042 47794 9054
rect 43810 8990 43822 9042
rect 43874 8990 43886 9042
rect 44258 8990 44270 9042
rect 44322 8990 44334 9042
rect 45154 8990 45166 9042
rect 45218 8990 45230 9042
rect 43598 8978 43650 8990
rect 47742 8978 47794 8990
rect 51662 9042 51714 9054
rect 51662 8978 51714 8990
rect 52782 9042 52834 9054
rect 52782 8978 52834 8990
rect 53118 9042 53170 9054
rect 53118 8978 53170 8990
rect 54014 9042 54066 9054
rect 54014 8978 54066 8990
rect 54126 9042 54178 9054
rect 56030 9042 56082 9054
rect 54562 8990 54574 9042
rect 54626 8990 54638 9042
rect 54126 8978 54178 8990
rect 56030 8978 56082 8990
rect 56590 9042 56642 9054
rect 56590 8978 56642 8990
rect 56702 9042 56754 9054
rect 57026 8990 57038 9042
rect 57090 8990 57102 9042
rect 56702 8978 56754 8990
rect 3614 8930 3666 8942
rect 11902 8930 11954 8942
rect 34190 8930 34242 8942
rect 7970 8878 7982 8930
rect 8034 8878 8046 8930
rect 10994 8878 11006 8930
rect 11058 8878 11070 8930
rect 15698 8878 15710 8930
rect 15762 8878 15774 8930
rect 20066 8878 20078 8930
rect 20130 8878 20142 8930
rect 25554 8878 25566 8930
rect 25618 8878 25630 8930
rect 29026 8878 29038 8930
rect 29090 8878 29102 8930
rect 3614 8866 3666 8878
rect 11902 8866 11954 8878
rect 34190 8866 34242 8878
rect 42478 8930 42530 8942
rect 42478 8866 42530 8878
rect 42590 8930 42642 8942
rect 51326 8930 51378 8942
rect 45378 8878 45390 8930
rect 45442 8878 45454 8930
rect 42590 8866 42642 8878
rect 51326 8866 51378 8878
rect 34414 8818 34466 8830
rect 34414 8754 34466 8766
rect 43038 8818 43090 8830
rect 51774 8818 51826 8830
rect 45266 8766 45278 8818
rect 45330 8766 45342 8818
rect 43038 8754 43090 8766
rect 51774 8754 51826 8766
rect 53678 8818 53730 8830
rect 53678 8754 53730 8766
rect 1344 8650 58576 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 58576 8650
rect 1344 8564 58576 8598
rect 24670 8482 24722 8494
rect 24670 8418 24722 8430
rect 30382 8482 30434 8494
rect 30382 8418 30434 8430
rect 2494 8370 2546 8382
rect 14478 8370 14530 8382
rect 7970 8318 7982 8370
rect 8034 8318 8046 8370
rect 10210 8318 10222 8370
rect 10274 8318 10286 8370
rect 13570 8318 13582 8370
rect 13634 8318 13646 8370
rect 2494 8306 2546 8318
rect 14478 8306 14530 8318
rect 15038 8370 15090 8382
rect 25006 8370 25058 8382
rect 15362 8318 15374 8370
rect 15426 8318 15438 8370
rect 18162 8318 18174 8370
rect 18226 8318 18238 8370
rect 15038 8306 15090 8318
rect 25006 8306 25058 8318
rect 28142 8370 28194 8382
rect 49646 8370 49698 8382
rect 31938 8318 31950 8370
rect 32002 8318 32014 8370
rect 42130 8318 42142 8370
rect 42194 8318 42206 8370
rect 28142 8306 28194 8318
rect 49646 8306 49698 8318
rect 51214 8370 51266 8382
rect 51214 8306 51266 8318
rect 52110 8370 52162 8382
rect 52110 8306 52162 8318
rect 4398 8258 4450 8270
rect 4398 8194 4450 8206
rect 4734 8258 4786 8270
rect 4734 8194 4786 8206
rect 5742 8258 5794 8270
rect 6638 8258 6690 8270
rect 5954 8206 5966 8258
rect 6018 8206 6030 8258
rect 5742 8194 5794 8206
rect 6638 8194 6690 8206
rect 7310 8258 7362 8270
rect 19406 8258 19458 8270
rect 8306 8206 8318 8258
rect 8370 8206 8382 8258
rect 9426 8206 9438 8258
rect 9490 8206 9502 8258
rect 11106 8206 11118 8258
rect 11170 8206 11182 8258
rect 13794 8206 13806 8258
rect 13858 8206 13870 8258
rect 16818 8206 16830 8258
rect 16882 8206 16894 8258
rect 18834 8206 18846 8258
rect 18898 8206 18910 8258
rect 7310 8194 7362 8206
rect 19406 8194 19458 8206
rect 20190 8258 20242 8270
rect 25230 8258 25282 8270
rect 24658 8206 24670 8258
rect 24722 8206 24734 8258
rect 20190 8194 20242 8206
rect 25230 8194 25282 8206
rect 27470 8258 27522 8270
rect 27470 8194 27522 8206
rect 28702 8258 28754 8270
rect 34638 8258 34690 8270
rect 38782 8258 38834 8270
rect 31826 8206 31838 8258
rect 31890 8206 31902 8258
rect 32498 8206 32510 8258
rect 32562 8206 32574 8258
rect 33058 8206 33070 8258
rect 33122 8206 33134 8258
rect 35298 8206 35310 8258
rect 35362 8206 35374 8258
rect 28702 8194 28754 8206
rect 34638 8194 34690 8206
rect 38782 8194 38834 8206
rect 39118 8258 39170 8270
rect 39118 8194 39170 8206
rect 39902 8258 39954 8270
rect 50990 8258 51042 8270
rect 54238 8258 54290 8270
rect 40338 8206 40350 8258
rect 40402 8206 40414 8258
rect 43586 8206 43598 8258
rect 43650 8206 43662 8258
rect 46386 8206 46398 8258
rect 46450 8206 46462 8258
rect 52882 8206 52894 8258
rect 52946 8206 52958 8258
rect 53666 8206 53678 8258
rect 53730 8206 53742 8258
rect 54002 8206 54014 8258
rect 54066 8206 54078 8258
rect 39902 8194 39954 8206
rect 50990 8194 51042 8206
rect 54238 8194 54290 8206
rect 54462 8258 54514 8270
rect 54462 8194 54514 8206
rect 55918 8258 55970 8270
rect 56578 8206 56590 8258
rect 56642 8206 56654 8258
rect 57250 8206 57262 8258
rect 57314 8206 57326 8258
rect 55918 8194 55970 8206
rect 1710 8146 1762 8158
rect 1710 8082 1762 8094
rect 2942 8146 2994 8158
rect 2942 8082 2994 8094
rect 4510 8146 4562 8158
rect 4510 8082 4562 8094
rect 7086 8146 7138 8158
rect 19518 8146 19570 8158
rect 11442 8094 11454 8146
rect 11506 8094 11518 8146
rect 11666 8094 11678 8146
rect 11730 8094 11742 8146
rect 15810 8094 15822 8146
rect 15874 8094 15886 8146
rect 7086 8082 7138 8094
rect 19518 8082 19570 8094
rect 19854 8146 19906 8158
rect 19854 8082 19906 8094
rect 19966 8146 20018 8158
rect 19966 8082 20018 8094
rect 24334 8146 24386 8158
rect 24334 8082 24386 8094
rect 27134 8146 27186 8158
rect 27134 8082 27186 8094
rect 27246 8146 27298 8158
rect 27246 8082 27298 8094
rect 30494 8146 30546 8158
rect 33294 8146 33346 8158
rect 31154 8094 31166 8146
rect 31218 8094 31230 8146
rect 31602 8094 31614 8146
rect 31666 8094 31678 8146
rect 30494 8082 30546 8094
rect 33294 8082 33346 8094
rect 34078 8146 34130 8158
rect 34078 8082 34130 8094
rect 35534 8146 35586 8158
rect 35534 8082 35586 8094
rect 35870 8146 35922 8158
rect 35870 8082 35922 8094
rect 35982 8146 36034 8158
rect 35982 8082 36034 8094
rect 36990 8146 37042 8158
rect 36990 8082 37042 8094
rect 37774 8146 37826 8158
rect 37774 8082 37826 8094
rect 38894 8146 38946 8158
rect 38894 8082 38946 8094
rect 40798 8146 40850 8158
rect 53118 8146 53170 8158
rect 42578 8094 42590 8146
rect 42642 8094 42654 8146
rect 45938 8094 45950 8146
rect 46002 8094 46014 8146
rect 47506 8094 47518 8146
rect 47570 8094 47582 8146
rect 50194 8094 50206 8146
rect 50258 8094 50270 8146
rect 40798 8082 40850 8094
rect 53118 8082 53170 8094
rect 53230 8146 53282 8158
rect 53230 8082 53282 8094
rect 54574 8146 54626 8158
rect 57474 8094 57486 8146
rect 57538 8094 57550 8146
rect 54574 8082 54626 8094
rect 2046 8034 2098 8046
rect 2046 7970 2098 7982
rect 7422 8034 7474 8046
rect 7422 7970 7474 7982
rect 7534 8034 7586 8046
rect 26910 8034 26962 8046
rect 11890 7982 11902 8034
rect 11954 7982 11966 8034
rect 25554 7982 25566 8034
rect 25618 7982 25630 8034
rect 7534 7970 7586 7982
rect 26910 7970 26962 7982
rect 28030 8034 28082 8046
rect 28030 7970 28082 7982
rect 28254 8034 28306 8046
rect 28254 7970 28306 7982
rect 30382 8034 30434 8046
rect 30382 7970 30434 7982
rect 30830 8034 30882 8046
rect 30830 7970 30882 7982
rect 36206 8034 36258 8046
rect 36206 7970 36258 7982
rect 37102 8034 37154 8046
rect 37102 7970 37154 7982
rect 37326 8034 37378 8046
rect 37326 7970 37378 7982
rect 37886 8034 37938 8046
rect 37886 7970 37938 7982
rect 38110 8034 38162 8046
rect 38110 7970 38162 7982
rect 39454 8034 39506 8046
rect 39454 7970 39506 7982
rect 41246 8034 41298 8046
rect 49870 8034 49922 8046
rect 51774 8034 51826 8046
rect 43922 7982 43934 8034
rect 43986 7982 43998 8034
rect 47394 7982 47406 8034
rect 47458 7982 47470 8034
rect 50642 7982 50654 8034
rect 50706 7982 50718 8034
rect 41246 7970 41298 7982
rect 49870 7970 49922 7982
rect 51774 7970 51826 7982
rect 1344 7866 58576 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 50558 7866
rect 50610 7814 50662 7866
rect 50714 7814 50766 7866
rect 50818 7814 58576 7866
rect 1344 7780 58576 7814
rect 1822 7698 1874 7710
rect 1822 7634 1874 7646
rect 8878 7698 8930 7710
rect 26238 7698 26290 7710
rect 10098 7646 10110 7698
rect 10162 7646 10174 7698
rect 16482 7646 16494 7698
rect 16546 7646 16558 7698
rect 8878 7634 8930 7646
rect 26238 7634 26290 7646
rect 27246 7698 27298 7710
rect 33854 7698 33906 7710
rect 31378 7646 31390 7698
rect 31442 7646 31454 7698
rect 27246 7634 27298 7646
rect 33854 7634 33906 7646
rect 35310 7698 35362 7710
rect 41022 7698 41074 7710
rect 50654 7698 50706 7710
rect 37202 7695 37214 7698
rect 35310 7634 35362 7646
rect 37105 7649 37214 7695
rect 5406 7586 5458 7598
rect 5406 7522 5458 7534
rect 14702 7586 14754 7598
rect 14702 7522 14754 7534
rect 14814 7586 14866 7598
rect 14814 7522 14866 7534
rect 24670 7586 24722 7598
rect 24670 7522 24722 7534
rect 26462 7586 26514 7598
rect 26462 7522 26514 7534
rect 26910 7586 26962 7598
rect 26910 7522 26962 7534
rect 27022 7586 27074 7598
rect 27022 7522 27074 7534
rect 29822 7586 29874 7598
rect 29822 7522 29874 7534
rect 30606 7586 30658 7598
rect 36654 7586 36706 7598
rect 31714 7534 31726 7586
rect 31778 7534 31790 7586
rect 34290 7534 34302 7586
rect 34354 7534 34366 7586
rect 30606 7522 30658 7534
rect 36654 7522 36706 7534
rect 36766 7586 36818 7598
rect 36766 7522 36818 7534
rect 5630 7474 5682 7486
rect 5630 7410 5682 7422
rect 7982 7474 8034 7486
rect 7982 7410 8034 7422
rect 8430 7474 8482 7486
rect 8430 7410 8482 7422
rect 9550 7474 9602 7486
rect 9550 7410 9602 7422
rect 9774 7474 9826 7486
rect 23214 7474 23266 7486
rect 26574 7474 26626 7486
rect 30382 7474 30434 7486
rect 11890 7422 11902 7474
rect 11954 7422 11966 7474
rect 12562 7422 12574 7474
rect 12626 7422 12638 7474
rect 13794 7422 13806 7474
rect 13858 7422 13870 7474
rect 14466 7422 14478 7474
rect 14530 7422 14542 7474
rect 15922 7422 15934 7474
rect 15986 7422 15998 7474
rect 16146 7422 16158 7474
rect 16210 7422 16222 7474
rect 22866 7422 22878 7474
rect 22930 7422 22942 7474
rect 24210 7422 24222 7474
rect 24274 7422 24286 7474
rect 27682 7422 27694 7474
rect 27746 7422 27758 7474
rect 29026 7422 29038 7474
rect 29090 7422 29102 7474
rect 9774 7410 9826 7422
rect 23214 7410 23266 7422
rect 26574 7410 26626 7422
rect 30382 7410 30434 7422
rect 30718 7474 30770 7486
rect 32062 7474 32114 7486
rect 31154 7422 31166 7474
rect 31218 7422 31230 7474
rect 30718 7410 30770 7422
rect 32062 7410 32114 7422
rect 34638 7474 34690 7486
rect 35758 7474 35810 7486
rect 35074 7422 35086 7474
rect 35138 7422 35150 7474
rect 34638 7410 34690 7422
rect 35758 7410 35810 7422
rect 36318 7474 36370 7486
rect 36318 7410 36370 7422
rect 36990 7474 37042 7486
rect 36990 7410 37042 7422
rect 33182 7362 33234 7374
rect 15250 7310 15262 7362
rect 15314 7310 15326 7362
rect 15698 7310 15710 7362
rect 15762 7310 15774 7362
rect 27570 7310 27582 7362
rect 27634 7310 27646 7362
rect 33182 7298 33234 7310
rect 33630 7362 33682 7374
rect 33954 7310 33966 7362
rect 34018 7310 34030 7362
rect 33630 7298 33682 7310
rect 5966 7250 6018 7262
rect 5966 7186 6018 7198
rect 8206 7250 8258 7262
rect 37105 7250 37151 7649
rect 37202 7646 37214 7649
rect 37266 7646 37278 7698
rect 49298 7646 49310 7698
rect 49362 7646 49374 7698
rect 56690 7646 56702 7698
rect 56754 7646 56766 7698
rect 41022 7634 41074 7646
rect 50654 7634 50706 7646
rect 38894 7586 38946 7598
rect 41582 7586 41634 7598
rect 40114 7534 40126 7586
rect 40178 7534 40190 7586
rect 38894 7522 38946 7534
rect 41582 7522 41634 7534
rect 41694 7586 41746 7598
rect 41694 7522 41746 7534
rect 44606 7586 44658 7598
rect 44606 7522 44658 7534
rect 47630 7586 47682 7598
rect 47630 7522 47682 7534
rect 48750 7586 48802 7598
rect 51986 7534 51998 7586
rect 52050 7534 52062 7586
rect 53442 7534 53454 7586
rect 53506 7534 53518 7586
rect 55906 7534 55918 7586
rect 55970 7534 55982 7586
rect 57250 7534 57262 7586
rect 57314 7534 57326 7586
rect 48750 7522 48802 7534
rect 39230 7474 39282 7486
rect 40798 7474 40850 7486
rect 38098 7422 38110 7474
rect 38162 7422 38174 7474
rect 39890 7422 39902 7474
rect 39954 7422 39966 7474
rect 39230 7410 39282 7422
rect 40798 7410 40850 7422
rect 41134 7474 41186 7486
rect 41134 7410 41186 7422
rect 41358 7474 41410 7486
rect 47518 7474 47570 7486
rect 44146 7422 44158 7474
rect 44210 7422 44222 7474
rect 47170 7422 47182 7474
rect 47234 7422 47246 7474
rect 50194 7422 50206 7474
rect 50258 7422 50270 7474
rect 50418 7422 50430 7474
rect 50482 7422 50494 7474
rect 50866 7422 50878 7474
rect 50930 7422 50942 7474
rect 51650 7422 51662 7474
rect 51714 7422 51726 7474
rect 54674 7422 54686 7474
rect 54738 7422 54750 7474
rect 56578 7422 56590 7474
rect 56642 7422 56654 7474
rect 57138 7422 57150 7474
rect 57202 7422 57214 7474
rect 41358 7410 41410 7422
rect 47518 7410 47570 7422
rect 37550 7362 37602 7374
rect 50766 7362 50818 7374
rect 38322 7310 38334 7362
rect 38386 7310 38398 7362
rect 43698 7310 43710 7362
rect 43762 7310 43774 7362
rect 51538 7310 51550 7362
rect 51602 7310 51614 7362
rect 53330 7310 53342 7362
rect 53394 7310 53406 7362
rect 37550 7298 37602 7310
rect 50766 7298 50818 7310
rect 48974 7250 49026 7262
rect 14018 7198 14030 7250
rect 14082 7198 14094 7250
rect 37090 7198 37102 7250
rect 37154 7198 37166 7250
rect 8206 7186 8258 7198
rect 48974 7186 49026 7198
rect 1344 7082 58576 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 58576 7082
rect 1344 6996 58576 7030
rect 29262 6914 29314 6926
rect 24322 6862 24334 6914
rect 24386 6862 24398 6914
rect 29262 6850 29314 6862
rect 33406 6914 33458 6926
rect 33406 6850 33458 6862
rect 37886 6914 37938 6926
rect 37886 6850 37938 6862
rect 37438 6802 37490 6814
rect 51102 6802 51154 6814
rect 13570 6750 13582 6802
rect 13634 6750 13646 6802
rect 24658 6750 24670 6802
rect 24722 6750 24734 6802
rect 28242 6750 28254 6802
rect 28306 6750 28318 6802
rect 35746 6750 35758 6802
rect 35810 6750 35822 6802
rect 40898 6750 40910 6802
rect 40962 6750 40974 6802
rect 43138 6750 43150 6802
rect 43202 6750 43214 6802
rect 48962 6750 48974 6802
rect 49026 6750 49038 6802
rect 37438 6738 37490 6750
rect 51102 6738 51154 6750
rect 14702 6690 14754 6702
rect 13906 6638 13918 6690
rect 13970 6638 13982 6690
rect 14702 6626 14754 6638
rect 15038 6690 15090 6702
rect 27918 6690 27970 6702
rect 24434 6638 24446 6690
rect 24498 6638 24510 6690
rect 15038 6626 15090 6638
rect 27918 6626 27970 6638
rect 28366 6690 28418 6702
rect 28366 6626 28418 6638
rect 29150 6690 29202 6702
rect 29150 6626 29202 6638
rect 29374 6690 29426 6702
rect 29374 6626 29426 6638
rect 29598 6690 29650 6702
rect 29598 6626 29650 6638
rect 29822 6690 29874 6702
rect 29822 6626 29874 6638
rect 32174 6690 32226 6702
rect 32174 6626 32226 6638
rect 32510 6690 32562 6702
rect 36542 6690 36594 6702
rect 35858 6638 35870 6690
rect 35922 6638 35934 6690
rect 32510 6626 32562 6638
rect 36542 6626 36594 6638
rect 36990 6690 37042 6702
rect 36990 6626 37042 6638
rect 37214 6690 37266 6702
rect 39902 6690 39954 6702
rect 50878 6690 50930 6702
rect 38098 6638 38110 6690
rect 38162 6638 38174 6690
rect 39106 6638 39118 6690
rect 39170 6638 39182 6690
rect 41010 6638 41022 6690
rect 41074 6638 41086 6690
rect 42354 6638 42366 6690
rect 42418 6638 42430 6690
rect 47842 6638 47854 6690
rect 47906 6638 47918 6690
rect 48178 6638 48190 6690
rect 48242 6638 48254 6690
rect 49074 6638 49086 6690
rect 49138 6638 49150 6690
rect 37214 6626 37266 6638
rect 39902 6626 39954 6638
rect 50878 6626 50930 6638
rect 51438 6690 51490 6702
rect 52994 6638 53006 6690
rect 53058 6638 53070 6690
rect 53890 6638 53902 6690
rect 53954 6638 53966 6690
rect 51438 6626 51490 6638
rect 14814 6578 14866 6590
rect 32286 6578 32338 6590
rect 26114 6526 26126 6578
rect 26178 6526 26190 6578
rect 26786 6526 26798 6578
rect 26850 6526 26862 6578
rect 27458 6526 27470 6578
rect 27522 6526 27534 6578
rect 31826 6526 31838 6578
rect 31890 6526 31902 6578
rect 14814 6514 14866 6526
rect 32286 6514 32338 6526
rect 32734 6578 32786 6590
rect 32734 6514 32786 6526
rect 33294 6578 33346 6590
rect 35198 6578 35250 6590
rect 34402 6526 34414 6578
rect 34466 6526 34478 6578
rect 33294 6514 33346 6526
rect 35198 6514 35250 6526
rect 35422 6578 35474 6590
rect 35422 6514 35474 6526
rect 36206 6578 36258 6590
rect 49758 6578 49810 6590
rect 38210 6526 38222 6578
rect 38274 6526 38286 6578
rect 47394 6526 47406 6578
rect 47458 6526 47470 6578
rect 36206 6514 36258 6526
rect 49758 6514 49810 6526
rect 51326 6578 51378 6590
rect 53106 6526 53118 6578
rect 53170 6526 53182 6578
rect 51326 6514 51378 6526
rect 25790 6466 25842 6478
rect 25790 6402 25842 6414
rect 26462 6466 26514 6478
rect 26462 6402 26514 6414
rect 27134 6466 27186 6478
rect 27134 6402 27186 6414
rect 28030 6466 28082 6478
rect 28030 6402 28082 6414
rect 28254 6466 28306 6478
rect 28254 6402 28306 6414
rect 30942 6466 30994 6478
rect 30942 6402 30994 6414
rect 31502 6466 31554 6478
rect 31502 6402 31554 6414
rect 32846 6466 32898 6478
rect 32846 6402 32898 6414
rect 33070 6466 33122 6478
rect 33070 6402 33122 6414
rect 33406 6466 33458 6478
rect 33406 6402 33458 6414
rect 34078 6466 34130 6478
rect 34078 6402 34130 6414
rect 34862 6466 34914 6478
rect 34862 6402 34914 6414
rect 35646 6466 35698 6478
rect 35646 6402 35698 6414
rect 36318 6466 36370 6478
rect 39678 6466 39730 6478
rect 39106 6414 39118 6466
rect 39170 6414 39182 6466
rect 36318 6402 36370 6414
rect 39678 6402 39730 6414
rect 40238 6466 40290 6478
rect 40238 6402 40290 6414
rect 40462 6466 40514 6478
rect 40462 6402 40514 6414
rect 40574 6466 40626 6478
rect 40574 6402 40626 6414
rect 45502 6466 45554 6478
rect 50094 6466 50146 6478
rect 48290 6414 48302 6466
rect 48354 6414 48366 6466
rect 45502 6402 45554 6414
rect 50094 6402 50146 6414
rect 50206 6466 50258 6478
rect 50206 6402 50258 6414
rect 50318 6466 50370 6478
rect 50318 6402 50370 6414
rect 50542 6466 50594 6478
rect 54002 6414 54014 6466
rect 54066 6414 54078 6466
rect 50542 6402 50594 6414
rect 1344 6298 58576 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 50558 6298
rect 50610 6246 50662 6298
rect 50714 6246 50766 6298
rect 50818 6246 58576 6298
rect 1344 6212 58576 6246
rect 25342 6130 25394 6142
rect 25342 6066 25394 6078
rect 25566 6130 25618 6142
rect 25566 6066 25618 6078
rect 26798 6130 26850 6142
rect 26798 6066 26850 6078
rect 27022 6130 27074 6142
rect 27022 6066 27074 6078
rect 27358 6130 27410 6142
rect 27358 6066 27410 6078
rect 27582 6130 27634 6142
rect 27582 6066 27634 6078
rect 31166 6130 31218 6142
rect 31166 6066 31218 6078
rect 33742 6130 33794 6142
rect 33742 6066 33794 6078
rect 35422 6130 35474 6142
rect 40014 6130 40066 6142
rect 47742 6130 47794 6142
rect 53342 6130 53394 6142
rect 35858 6078 35870 6130
rect 35922 6078 35934 6130
rect 41906 6078 41918 6130
rect 41970 6078 41982 6130
rect 52546 6078 52558 6130
rect 52610 6078 52622 6130
rect 35422 6066 35474 6078
rect 40014 6066 40066 6078
rect 47742 6066 47794 6078
rect 53342 6066 53394 6078
rect 53566 6130 53618 6142
rect 53566 6066 53618 6078
rect 26686 6018 26738 6030
rect 26686 5954 26738 5966
rect 27246 6018 27298 6030
rect 27246 5954 27298 5966
rect 32174 6018 32226 6030
rect 32174 5954 32226 5966
rect 33070 6018 33122 6030
rect 40350 6018 40402 6030
rect 49198 6018 49250 6030
rect 37202 5966 37214 6018
rect 37266 5966 37278 6018
rect 37538 5966 37550 6018
rect 37602 5966 37614 6018
rect 41010 5966 41022 6018
rect 41074 5966 41086 6018
rect 45266 5966 45278 6018
rect 45330 5966 45342 6018
rect 33070 5954 33122 5966
rect 40350 5954 40402 5966
rect 49198 5954 49250 5966
rect 49646 6018 49698 6030
rect 49646 5954 49698 5966
rect 53230 6018 53282 6030
rect 53230 5954 53282 5966
rect 25678 5906 25730 5918
rect 31502 5906 31554 5918
rect 29922 5854 29934 5906
rect 29986 5854 29998 5906
rect 25678 5842 25730 5854
rect 31502 5842 31554 5854
rect 31838 5906 31890 5918
rect 34078 5906 34130 5918
rect 33282 5854 33294 5906
rect 33346 5854 33358 5906
rect 31838 5842 31890 5854
rect 34078 5842 34130 5854
rect 34526 5906 34578 5918
rect 34526 5842 34578 5854
rect 34638 5906 34690 5918
rect 34638 5842 34690 5854
rect 34750 5906 34802 5918
rect 34750 5842 34802 5854
rect 35198 5906 35250 5918
rect 39790 5906 39842 5918
rect 36306 5854 36318 5906
rect 36370 5854 36382 5906
rect 36754 5854 36766 5906
rect 36818 5854 36830 5906
rect 37762 5854 37774 5906
rect 37826 5854 37838 5906
rect 35198 5842 35250 5854
rect 39790 5842 39842 5854
rect 40126 5906 40178 5918
rect 42366 5906 42418 5918
rect 40898 5854 40910 5906
rect 40962 5854 40974 5906
rect 41794 5854 41806 5906
rect 41858 5854 41870 5906
rect 40126 5842 40178 5854
rect 42366 5842 42418 5854
rect 42590 5906 42642 5918
rect 47182 5906 47234 5918
rect 51102 5906 51154 5918
rect 44370 5854 44382 5906
rect 44434 5854 44446 5906
rect 44818 5854 44830 5906
rect 44882 5854 44894 5906
rect 46274 5854 46286 5906
rect 46338 5854 46350 5906
rect 50418 5854 50430 5906
rect 50482 5854 50494 5906
rect 51426 5854 51438 5906
rect 51490 5854 51502 5906
rect 52770 5854 52782 5906
rect 52834 5854 52846 5906
rect 42590 5842 42642 5854
rect 47182 5842 47234 5854
rect 51102 5842 51154 5854
rect 30942 5794 30994 5806
rect 38222 5794 38274 5806
rect 37090 5742 37102 5794
rect 37154 5742 37166 5794
rect 30942 5730 30994 5742
rect 38222 5730 38274 5742
rect 38894 5794 38946 5806
rect 38894 5730 38946 5742
rect 43374 5794 43426 5806
rect 43374 5730 43426 5742
rect 43822 5794 43874 5806
rect 44930 5742 44942 5794
rect 44994 5742 45006 5794
rect 46498 5742 46510 5794
rect 46562 5742 46574 5794
rect 47842 5742 47854 5794
rect 47906 5742 47918 5794
rect 49298 5742 49310 5794
rect 49362 5742 49374 5794
rect 43822 5730 43874 5742
rect 28030 5682 28082 5694
rect 28030 5618 28082 5630
rect 38446 5682 38498 5694
rect 38446 5618 38498 5630
rect 38670 5682 38722 5694
rect 38670 5618 38722 5630
rect 39342 5682 39394 5694
rect 47518 5682 47570 5694
rect 42914 5630 42926 5682
rect 42978 5630 42990 5682
rect 39342 5618 39394 5630
rect 47518 5618 47570 5630
rect 48974 5682 49026 5694
rect 48974 5618 49026 5630
rect 1344 5514 58576 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 58576 5514
rect 1344 5428 58576 5462
rect 40910 5346 40962 5358
rect 44382 5346 44434 5358
rect 39666 5294 39678 5346
rect 39730 5294 39742 5346
rect 41234 5294 41246 5346
rect 41298 5294 41310 5346
rect 40910 5282 40962 5294
rect 44382 5282 44434 5294
rect 48078 5346 48130 5358
rect 48078 5282 48130 5294
rect 50318 5346 50370 5358
rect 50318 5282 50370 5294
rect 50766 5346 50818 5358
rect 50766 5282 50818 5294
rect 28702 5234 28754 5246
rect 28702 5170 28754 5182
rect 30606 5234 30658 5246
rect 30606 5170 30658 5182
rect 33518 5234 33570 5246
rect 33518 5170 33570 5182
rect 36430 5234 36482 5246
rect 40686 5234 40738 5246
rect 38882 5182 38894 5234
rect 38946 5182 38958 5234
rect 39330 5182 39342 5234
rect 39394 5182 39406 5234
rect 36430 5170 36482 5182
rect 40686 5170 40738 5182
rect 44942 5234 44994 5246
rect 48414 5234 48466 5246
rect 47058 5182 47070 5234
rect 47122 5182 47134 5234
rect 44942 5170 44994 5182
rect 48414 5170 48466 5182
rect 49870 5234 49922 5246
rect 49870 5170 49922 5182
rect 50094 5234 50146 5246
rect 50094 5170 50146 5182
rect 29822 5122 29874 5134
rect 29822 5058 29874 5070
rect 30942 5122 30994 5134
rect 32622 5122 32674 5134
rect 31938 5070 31950 5122
rect 32002 5070 32014 5122
rect 30942 5058 30994 5070
rect 32622 5058 32674 5070
rect 32846 5122 32898 5134
rect 36094 5122 36146 5134
rect 37662 5122 37714 5134
rect 43710 5122 43762 5134
rect 44718 5122 44770 5134
rect 33170 5070 33182 5122
rect 33234 5070 33246 5122
rect 33730 5070 33742 5122
rect 33794 5070 33806 5122
rect 34626 5070 34638 5122
rect 34690 5070 34702 5122
rect 34962 5070 34974 5122
rect 35026 5070 35038 5122
rect 35858 5070 35870 5122
rect 35922 5070 35934 5122
rect 37202 5070 37214 5122
rect 37266 5070 37278 5122
rect 38658 5070 38670 5122
rect 38722 5070 38734 5122
rect 39778 5070 39790 5122
rect 39842 5070 39854 5122
rect 44034 5070 44046 5122
rect 44098 5070 44110 5122
rect 32846 5058 32898 5070
rect 36094 5058 36146 5070
rect 37662 5058 37714 5070
rect 43710 5058 43762 5070
rect 44718 5058 44770 5070
rect 45166 5122 45218 5134
rect 45166 5058 45218 5070
rect 45390 5122 45442 5134
rect 45390 5058 45442 5070
rect 45726 5122 45778 5134
rect 48190 5122 48242 5134
rect 46946 5070 46958 5122
rect 47010 5070 47022 5122
rect 47506 5070 47518 5122
rect 47570 5070 47582 5122
rect 45726 5058 45778 5070
rect 48190 5058 48242 5070
rect 48526 5122 48578 5134
rect 48526 5058 48578 5070
rect 29374 5010 29426 5022
rect 29374 4946 29426 4958
rect 29486 5010 29538 5022
rect 29486 4946 29538 4958
rect 30158 5010 30210 5022
rect 32174 5010 32226 5022
rect 31266 4958 31278 5010
rect 31330 4958 31342 5010
rect 30158 4946 30210 4958
rect 32174 4946 32226 4958
rect 32734 5010 32786 5022
rect 32734 4946 32786 4958
rect 33966 5010 34018 5022
rect 44270 5010 44322 5022
rect 35186 4958 35198 5010
rect 35250 4958 35262 5010
rect 36306 4958 36318 5010
rect 36370 4958 36382 5010
rect 36978 4958 36990 5010
rect 37042 4958 37054 5010
rect 37986 4958 37998 5010
rect 38050 4958 38062 5010
rect 43138 4958 43150 5010
rect 43202 4958 43214 5010
rect 33966 4946 34018 4958
rect 44270 4946 44322 4958
rect 45950 5010 46002 5022
rect 45950 4946 46002 4958
rect 46062 5010 46114 5022
rect 46610 4958 46622 5010
rect 46674 4958 46686 5010
rect 46062 4946 46114 4958
rect 29150 4898 29202 4910
rect 29150 4834 29202 4846
rect 35422 4898 35474 4910
rect 35422 4834 35474 4846
rect 42030 4898 42082 4910
rect 42030 4834 42082 4846
rect 42254 4898 42306 4910
rect 42254 4834 42306 4846
rect 42366 4898 42418 4910
rect 42366 4834 42418 4846
rect 42478 4898 42530 4910
rect 42478 4834 42530 4846
rect 42814 4898 42866 4910
rect 42814 4834 42866 4846
rect 1344 4730 58576 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 50558 4730
rect 50610 4678 50662 4730
rect 50714 4678 50766 4730
rect 50818 4678 58576 4730
rect 1344 4644 58576 4678
rect 31390 4562 31442 4574
rect 32062 4562 32114 4574
rect 33406 4562 33458 4574
rect 31714 4510 31726 4562
rect 31778 4510 31790 4562
rect 32386 4510 32398 4562
rect 32450 4510 32462 4562
rect 33058 4510 33070 4562
rect 33122 4510 33134 4562
rect 31390 4498 31442 4510
rect 32062 4498 32114 4510
rect 33406 4498 33458 4510
rect 40910 4562 40962 4574
rect 40910 4498 40962 4510
rect 37202 4398 37214 4450
rect 37266 4398 37278 4450
rect 42130 4398 42142 4450
rect 42194 4398 42206 4450
rect 45714 4398 45726 4450
rect 45778 4398 45790 4450
rect 47954 4398 47966 4450
rect 48018 4398 48030 4450
rect 40014 4338 40066 4350
rect 30594 4286 30606 4338
rect 30658 4286 30670 4338
rect 33842 4286 33854 4338
rect 33906 4286 33918 4338
rect 36978 4286 36990 4338
rect 37042 4286 37054 4338
rect 37874 4286 37886 4338
rect 37938 4286 37950 4338
rect 39330 4286 39342 4338
rect 39394 4286 39406 4338
rect 42354 4286 42366 4338
rect 42418 4286 42430 4338
rect 44034 4286 44046 4338
rect 44098 4286 44110 4338
rect 44930 4286 44942 4338
rect 44994 4286 45006 4338
rect 45938 4286 45950 4338
rect 46002 4286 46014 4338
rect 47170 4286 47182 4338
rect 47234 4286 47246 4338
rect 40014 4274 40066 4286
rect 26910 4226 26962 4238
rect 26910 4162 26962 4174
rect 28254 4226 28306 4238
rect 28254 4162 28306 4174
rect 37438 4226 37490 4238
rect 37438 4162 37490 4174
rect 37550 4226 37602 4238
rect 44718 4226 44770 4238
rect 39106 4174 39118 4226
rect 39170 4174 39182 4226
rect 41346 4174 41358 4226
rect 41410 4174 41422 4226
rect 44146 4174 44158 4226
rect 44210 4174 44222 4226
rect 37550 4162 37602 4174
rect 44718 4162 44770 4174
rect 28702 4114 28754 4126
rect 28702 4050 28754 4062
rect 34862 4114 34914 4126
rect 34862 4050 34914 4062
rect 44606 4114 44658 4126
rect 44606 4050 44658 4062
rect 1344 3946 58576 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 58576 3946
rect 1344 3860 58576 3894
rect 35086 3778 35138 3790
rect 35086 3714 35138 3726
rect 40350 3778 40402 3790
rect 40350 3714 40402 3726
rect 42366 3778 42418 3790
rect 42366 3714 42418 3726
rect 42590 3778 42642 3790
rect 42590 3714 42642 3726
rect 43038 3778 43090 3790
rect 48178 3726 48190 3778
rect 48242 3726 48254 3778
rect 43038 3714 43090 3726
rect 29262 3666 29314 3678
rect 29262 3602 29314 3614
rect 36206 3666 36258 3678
rect 36206 3602 36258 3614
rect 39790 3666 39842 3678
rect 39790 3602 39842 3614
rect 42142 3666 42194 3678
rect 42142 3602 42194 3614
rect 25118 3554 25170 3566
rect 32510 3554 32562 3566
rect 40014 3554 40066 3566
rect 45614 3554 45666 3566
rect 26002 3502 26014 3554
rect 26066 3502 26078 3554
rect 31154 3502 31166 3554
rect 31218 3502 31230 3554
rect 32946 3502 32958 3554
rect 33010 3502 33022 3554
rect 33506 3502 33518 3554
rect 33570 3502 33582 3554
rect 34290 3502 34302 3554
rect 34354 3502 34366 3554
rect 34850 3502 34862 3554
rect 34914 3502 34926 3554
rect 38098 3502 38110 3554
rect 38162 3502 38174 3554
rect 39106 3502 39118 3554
rect 39170 3502 39182 3554
rect 40898 3502 40910 3554
rect 40962 3502 40974 3554
rect 41570 3502 41582 3554
rect 41634 3502 41646 3554
rect 43810 3502 43822 3554
rect 43874 3502 43886 3554
rect 45154 3502 45166 3554
rect 45218 3502 45230 3554
rect 25118 3490 25170 3502
rect 32510 3490 32562 3502
rect 40014 3490 40066 3502
rect 45614 3490 45666 3502
rect 45950 3554 46002 3566
rect 45950 3490 46002 3502
rect 46286 3554 46338 3566
rect 47630 3554 47682 3566
rect 47394 3502 47406 3554
rect 47458 3502 47470 3554
rect 46286 3490 46338 3502
rect 47630 3490 47682 3502
rect 47742 3554 47794 3566
rect 47742 3490 47794 3502
rect 14142 3442 14194 3454
rect 14142 3378 14194 3390
rect 14366 3442 14418 3454
rect 25566 3442 25618 3454
rect 14690 3390 14702 3442
rect 14754 3390 14766 3442
rect 14366 3378 14418 3390
rect 25566 3378 25618 3390
rect 25790 3442 25842 3454
rect 25790 3378 25842 3390
rect 26462 3442 26514 3454
rect 26462 3378 26514 3390
rect 26798 3442 26850 3454
rect 26798 3378 26850 3390
rect 27134 3442 27186 3454
rect 28366 3442 28418 3454
rect 27458 3390 27470 3442
rect 27522 3390 27534 3442
rect 27134 3378 27186 3390
rect 28366 3378 28418 3390
rect 28702 3442 28754 3454
rect 33742 3442 33794 3454
rect 32162 3390 32174 3442
rect 32226 3390 32238 3442
rect 33170 3390 33182 3442
rect 33234 3390 33246 3442
rect 28702 3378 28754 3390
rect 33742 3378 33794 3390
rect 35534 3442 35586 3454
rect 35534 3378 35586 3390
rect 38894 3442 38946 3454
rect 43598 3442 43650 3454
rect 44606 3442 44658 3454
rect 45726 3442 45778 3454
rect 40674 3390 40686 3442
rect 40738 3390 40750 3442
rect 41346 3390 41358 3442
rect 41410 3390 41422 3442
rect 44258 3390 44270 3442
rect 44322 3390 44334 3442
rect 44930 3390 44942 3442
rect 44994 3390 45006 3442
rect 38894 3378 38946 3390
rect 43598 3378 43650 3390
rect 44606 3378 44658 3390
rect 45726 3378 45778 3390
rect 46734 3442 46786 3454
rect 46734 3378 46786 3390
rect 21758 3330 21810 3342
rect 21758 3266 21810 3278
rect 1344 3162 58576 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 50558 3162
rect 50610 3110 50662 3162
rect 50714 3110 50766 3162
rect 50818 3110 58576 3162
rect 1344 3076 58576 3110
<< via1 >>
rect 27582 46958 27634 47010
rect 28254 46958 28306 47010
rect 30270 46622 30322 46674
rect 31054 46622 31106 46674
rect 31502 46622 31554 46674
rect 10110 46510 10162 46562
rect 10782 46510 10834 46562
rect 8766 46398 8818 46450
rect 9102 46398 9154 46450
rect 9438 46398 9490 46450
rect 42366 46398 42418 46450
rect 44942 46398 44994 46450
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 29374 46062 29426 46114
rect 9662 45950 9714 46002
rect 14478 45950 14530 46002
rect 16046 45950 16098 46002
rect 19182 45950 19234 46002
rect 26798 45950 26850 46002
rect 35086 45950 35138 46002
rect 44606 45950 44658 46002
rect 49982 45950 50034 46002
rect 53790 45950 53842 46002
rect 8766 45838 8818 45890
rect 9998 45838 10050 45890
rect 10782 45838 10834 45890
rect 11902 45838 11954 45890
rect 12350 45838 12402 45890
rect 13134 45838 13186 45890
rect 13806 45838 13858 45890
rect 16494 45838 16546 45890
rect 17054 45838 17106 45890
rect 17726 45838 17778 45890
rect 18622 45838 18674 45890
rect 21086 45838 21138 45890
rect 27134 45838 27186 45890
rect 27582 45838 27634 45890
rect 28366 45838 28418 45890
rect 31502 45838 31554 45890
rect 36542 45838 36594 45890
rect 37214 45838 37266 45890
rect 38110 45838 38162 45890
rect 38670 45838 38722 45890
rect 40014 45838 40066 45890
rect 40462 45838 40514 45890
rect 41358 45838 41410 45890
rect 41806 45838 41858 45890
rect 42254 45838 42306 45890
rect 42814 45838 42866 45890
rect 43598 45838 43650 45890
rect 45054 45838 45106 45890
rect 45502 45838 45554 45890
rect 50094 45838 50146 45890
rect 51438 45838 51490 45890
rect 52110 45838 52162 45890
rect 52782 45838 52834 45890
rect 54238 45838 54290 45890
rect 8206 45726 8258 45778
rect 11566 45726 11618 45778
rect 12574 45726 12626 45778
rect 13246 45726 13298 45778
rect 13470 45726 13522 45778
rect 15374 45726 15426 45778
rect 20750 45726 20802 45778
rect 21310 45726 21362 45778
rect 35534 45726 35586 45778
rect 42366 45726 42418 45778
rect 42590 45726 42642 45778
rect 46062 45726 46114 45778
rect 46734 45726 46786 45778
rect 47406 45726 47458 45778
rect 47742 45726 47794 45778
rect 49646 45726 49698 45778
rect 53342 45726 53394 45778
rect 8430 45614 8482 45666
rect 10222 45614 10274 45666
rect 10558 45614 10610 45666
rect 14142 45614 14194 45666
rect 15038 45614 15090 45666
rect 17390 45614 17442 45666
rect 18062 45614 18114 45666
rect 18398 45614 18450 45666
rect 21086 45614 21138 45666
rect 27806 45614 27858 45666
rect 31278 45614 31330 45666
rect 36878 45614 36930 45666
rect 37550 45614 37602 45666
rect 37886 45614 37938 45666
rect 38894 45614 38946 45666
rect 39790 45614 39842 45666
rect 40798 45614 40850 45666
rect 43150 45614 43202 45666
rect 44158 45614 44210 45666
rect 46398 45614 46450 45666
rect 48078 45614 48130 45666
rect 48414 45614 48466 45666
rect 48750 45614 48802 45666
rect 49086 45614 49138 45666
rect 51214 45614 51266 45666
rect 51886 45614 51938 45666
rect 52558 45614 52610 45666
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 50558 45446 50610 45498
rect 50662 45446 50714 45498
rect 50766 45446 50818 45498
rect 9102 45278 9154 45330
rect 10446 45278 10498 45330
rect 14814 45278 14866 45330
rect 21086 45278 21138 45330
rect 21870 45278 21922 45330
rect 30046 45278 30098 45330
rect 31054 45278 31106 45330
rect 52222 45278 52274 45330
rect 9886 45166 9938 45218
rect 11566 45166 11618 45218
rect 12238 45166 12290 45218
rect 13918 45166 13970 45218
rect 14142 45166 14194 45218
rect 16606 45166 16658 45218
rect 17726 45166 17778 45218
rect 22542 45166 22594 45218
rect 30382 45166 30434 45218
rect 40238 45166 40290 45218
rect 42254 45166 42306 45218
rect 43038 45166 43090 45218
rect 43822 45166 43874 45218
rect 44718 45166 44770 45218
rect 50990 45166 51042 45218
rect 53230 45166 53282 45218
rect 9662 45054 9714 45106
rect 10222 45054 10274 45106
rect 11118 45054 11170 45106
rect 12126 45054 12178 45106
rect 12686 45054 12738 45106
rect 13358 45054 13410 45106
rect 14366 45054 14418 45106
rect 15374 45054 15426 45106
rect 15598 45054 15650 45106
rect 16830 45054 16882 45106
rect 18174 45054 18226 45106
rect 18958 45054 19010 45106
rect 20190 45054 20242 45106
rect 21758 45054 21810 45106
rect 21982 45054 22034 45106
rect 22430 45054 22482 45106
rect 22766 45054 22818 45106
rect 29262 45054 29314 45106
rect 36654 45054 36706 45106
rect 38222 45054 38274 45106
rect 39566 45054 39618 45106
rect 40350 45054 40402 45106
rect 41022 45054 41074 45106
rect 42030 45054 42082 45106
rect 42926 45054 42978 45106
rect 44158 45054 44210 45106
rect 45390 45054 45442 45106
rect 46286 45054 46338 45106
rect 47630 45054 47682 45106
rect 49870 45054 49922 45106
rect 51998 45054 52050 45106
rect 11566 44942 11618 44994
rect 13806 44942 13858 44994
rect 15710 44942 15762 44994
rect 19630 44942 19682 44994
rect 19966 44942 20018 44994
rect 20638 44942 20690 44994
rect 21310 44942 21362 44994
rect 21534 44942 21586 44994
rect 27358 44942 27410 44994
rect 34750 44942 34802 44994
rect 37438 44942 37490 44994
rect 39118 44942 39170 44994
rect 41358 44942 41410 44994
rect 43374 44942 43426 44994
rect 45278 44942 45330 44994
rect 49086 44942 49138 44994
rect 51550 44942 51602 44994
rect 52110 44942 52162 44994
rect 52782 44942 52834 44994
rect 11902 44830 11954 44882
rect 16494 44830 16546 44882
rect 20414 44830 20466 44882
rect 40238 44830 40290 44882
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 16270 44494 16322 44546
rect 36318 44494 36370 44546
rect 52894 44494 52946 44546
rect 10558 44382 10610 44434
rect 12126 44382 12178 44434
rect 15598 44382 15650 44434
rect 28702 44382 28754 44434
rect 30046 44382 30098 44434
rect 30382 44382 30434 44434
rect 32510 44382 32562 44434
rect 37214 44382 37266 44434
rect 44382 44382 44434 44434
rect 44942 44382 44994 44434
rect 49982 44382 50034 44434
rect 50878 44382 50930 44434
rect 52670 44382 52722 44434
rect 9662 44270 9714 44322
rect 9886 44270 9938 44322
rect 10110 44270 10162 44322
rect 11454 44270 11506 44322
rect 12462 44270 12514 44322
rect 13806 44270 13858 44322
rect 16382 44270 16434 44322
rect 17054 44270 17106 44322
rect 17502 44270 17554 44322
rect 18958 44270 19010 44322
rect 19742 44270 19794 44322
rect 20414 44270 20466 44322
rect 21310 44270 21362 44322
rect 22094 44270 22146 44322
rect 23214 44270 23266 44322
rect 29374 44270 29426 44322
rect 33518 44270 33570 44322
rect 34078 44270 34130 44322
rect 36206 44270 36258 44322
rect 38894 44270 38946 44322
rect 39118 44270 39170 44322
rect 39678 44270 39730 44322
rect 40350 44270 40402 44322
rect 41470 44270 41522 44322
rect 44270 44270 44322 44322
rect 46286 44270 46338 44322
rect 47294 44270 47346 44322
rect 48862 44270 48914 44322
rect 49086 44270 49138 44322
rect 50206 44270 50258 44322
rect 50654 44270 50706 44322
rect 1710 44158 1762 44210
rect 7982 44158 8034 44210
rect 9774 44158 9826 44210
rect 11790 44158 11842 44210
rect 12126 44158 12178 44210
rect 15262 44158 15314 44210
rect 15486 44158 15538 44210
rect 17614 44158 17666 44210
rect 17838 44158 17890 44210
rect 19294 44158 19346 44210
rect 20750 44158 20802 44210
rect 22766 44158 22818 44210
rect 32174 44158 32226 44210
rect 33630 44158 33682 44210
rect 36318 44158 36370 44210
rect 37550 44158 37602 44210
rect 37662 44158 37714 44210
rect 39342 44158 39394 44210
rect 40686 44158 40738 44210
rect 41918 44158 41970 44210
rect 42814 44158 42866 44210
rect 45838 44158 45890 44210
rect 48078 44158 48130 44210
rect 2046 44046 2098 44098
rect 2494 44046 2546 44098
rect 7646 44046 7698 44098
rect 8766 44046 8818 44098
rect 9102 44046 9154 44098
rect 13470 44046 13522 44098
rect 16270 44046 16322 44098
rect 16718 44046 16770 44098
rect 19742 44046 19794 44098
rect 21646 44046 21698 44098
rect 22206 44046 22258 44098
rect 29150 44046 29202 44098
rect 37326 44046 37378 44098
rect 40014 44046 40066 44098
rect 51886 44046 51938 44098
rect 53230 44046 53282 44098
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 50558 43878 50610 43930
rect 50662 43878 50714 43930
rect 50766 43878 50818 43930
rect 7086 43710 7138 43762
rect 9886 43710 9938 43762
rect 13246 43710 13298 43762
rect 39342 43710 39394 43762
rect 46286 43710 46338 43762
rect 10222 43598 10274 43650
rect 10670 43598 10722 43650
rect 14366 43598 14418 43650
rect 34414 43598 34466 43650
rect 37774 43598 37826 43650
rect 38110 43598 38162 43650
rect 38446 43598 38498 43650
rect 39566 43598 39618 43650
rect 40126 43598 40178 43650
rect 41022 43598 41074 43650
rect 42030 43598 42082 43650
rect 42926 43598 42978 43650
rect 44158 43598 44210 43650
rect 46062 43598 46114 43650
rect 47294 43598 47346 43650
rect 47630 43598 47682 43650
rect 48862 43598 48914 43650
rect 49086 43598 49138 43650
rect 7198 43486 7250 43538
rect 7870 43486 7922 43538
rect 10558 43486 10610 43538
rect 11342 43486 11394 43538
rect 11790 43486 11842 43538
rect 12798 43486 12850 43538
rect 13470 43486 13522 43538
rect 15598 43486 15650 43538
rect 17838 43486 17890 43538
rect 20526 43486 20578 43538
rect 20750 43486 20802 43538
rect 22206 43486 22258 43538
rect 23438 43486 23490 43538
rect 35870 43486 35922 43538
rect 37214 43486 37266 43538
rect 38782 43486 38834 43538
rect 39678 43486 39730 43538
rect 40014 43486 40066 43538
rect 41358 43486 41410 43538
rect 41806 43486 41858 43538
rect 42590 43486 42642 43538
rect 45614 43486 45666 43538
rect 46510 43486 46562 43538
rect 46958 43486 47010 43538
rect 47966 43486 48018 43538
rect 48750 43486 48802 43538
rect 49310 43486 49362 43538
rect 49534 43486 49586 43538
rect 49758 43486 49810 43538
rect 51214 43486 51266 43538
rect 51550 43486 51602 43538
rect 53006 43486 53058 43538
rect 53342 43486 53394 43538
rect 53566 43486 53618 43538
rect 2158 43374 2210 43426
rect 8206 43374 8258 43426
rect 8542 43374 8594 43426
rect 13358 43374 13410 43426
rect 14142 43374 14194 43426
rect 16270 43374 16322 43426
rect 17502 43374 17554 43426
rect 21870 43374 21922 43426
rect 22654 43374 22706 43426
rect 23662 43374 23714 43426
rect 34302 43374 34354 43426
rect 35086 43374 35138 43426
rect 37102 43374 37154 43426
rect 45390 43374 45442 43426
rect 47182 43374 47234 43426
rect 47742 43374 47794 43426
rect 51662 43374 51714 43426
rect 7086 43262 7138 43314
rect 11342 43262 11394 43314
rect 20974 43262 21026 43314
rect 21422 43262 21474 43314
rect 23998 43262 24050 43314
rect 34638 43262 34690 43314
rect 40126 43262 40178 43314
rect 50206 43262 50258 43314
rect 53902 43262 53954 43314
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 8206 42926 8258 42978
rect 15038 42926 15090 42978
rect 15262 42926 15314 42978
rect 34414 42926 34466 42978
rect 34750 42926 34802 42978
rect 37102 42926 37154 42978
rect 41134 42926 41186 42978
rect 45390 42926 45442 42978
rect 51326 42926 51378 42978
rect 7982 42814 8034 42866
rect 11454 42814 11506 42866
rect 14814 42814 14866 42866
rect 33518 42814 33570 42866
rect 40686 42814 40738 42866
rect 47070 42814 47122 42866
rect 49198 42814 49250 42866
rect 50094 42814 50146 42866
rect 52894 42814 52946 42866
rect 1822 42702 1874 42754
rect 7646 42702 7698 42754
rect 8878 42702 8930 42754
rect 10110 42702 10162 42754
rect 10558 42702 10610 42754
rect 11118 42702 11170 42754
rect 12126 42702 12178 42754
rect 13918 42702 13970 42754
rect 15710 42702 15762 42754
rect 16158 42702 16210 42754
rect 19182 42702 19234 42754
rect 19518 42702 19570 42754
rect 23326 42702 23378 42754
rect 23662 42702 23714 42754
rect 31950 42702 32002 42754
rect 33630 42702 33682 42754
rect 34190 42702 34242 42754
rect 34974 42702 35026 42754
rect 37214 42702 37266 42754
rect 37550 42702 37602 42754
rect 39006 42702 39058 42754
rect 41022 42702 41074 42754
rect 41806 42702 41858 42754
rect 42142 42702 42194 42754
rect 43038 42702 43090 42754
rect 44046 42702 44098 42754
rect 45054 42702 45106 42754
rect 46174 42702 46226 42754
rect 47854 42702 47906 42754
rect 48750 42702 48802 42754
rect 49534 42702 49586 42754
rect 54350 42702 54402 42754
rect 2382 42590 2434 42642
rect 7310 42590 7362 42642
rect 10894 42590 10946 42642
rect 13582 42590 13634 42642
rect 19630 42590 19682 42642
rect 22990 42590 23042 42642
rect 23438 42590 23490 42642
rect 30046 42590 30098 42642
rect 30158 42590 30210 42642
rect 31726 42590 31778 42642
rect 35310 42590 35362 42642
rect 39342 42590 39394 42642
rect 41918 42590 41970 42642
rect 42702 42590 42754 42642
rect 51550 42590 51602 42642
rect 53454 42590 53506 42642
rect 55694 42590 55746 42642
rect 2046 42478 2098 42530
rect 2718 42478 2770 42530
rect 3166 42478 3218 42530
rect 7534 42478 7586 42530
rect 8542 42478 8594 42530
rect 9214 42478 9266 42530
rect 11342 42478 11394 42530
rect 11454 42478 11506 42530
rect 11902 42478 11954 42530
rect 13694 42478 13746 42530
rect 16270 42478 16322 42530
rect 16382 42478 16434 42530
rect 16494 42478 16546 42530
rect 16606 42478 16658 42530
rect 22654 42478 22706 42530
rect 22878 42478 22930 42530
rect 30382 42478 30434 42530
rect 30718 42478 30770 42530
rect 35198 42478 35250 42530
rect 37102 42478 37154 42530
rect 37662 42478 37714 42530
rect 37886 42478 37938 42530
rect 39230 42478 39282 42530
rect 39902 42478 39954 42530
rect 40238 42478 40290 42530
rect 41134 42478 41186 42530
rect 42366 42478 42418 42530
rect 43374 42478 43426 42530
rect 43710 42478 43762 42530
rect 45278 42478 45330 42530
rect 45838 42478 45890 42530
rect 51438 42478 51490 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 50558 42310 50610 42362
rect 50662 42310 50714 42362
rect 50766 42310 50818 42362
rect 4398 42142 4450 42194
rect 9774 42142 9826 42194
rect 10558 42142 10610 42194
rect 14030 42142 14082 42194
rect 14590 42142 14642 42194
rect 30046 42142 30098 42194
rect 30494 42142 30546 42194
rect 44606 42142 44658 42194
rect 44830 42142 44882 42194
rect 50766 42142 50818 42194
rect 2046 42030 2098 42082
rect 2718 42030 2770 42082
rect 7646 42030 7698 42082
rect 11454 42030 11506 42082
rect 12686 42030 12738 42082
rect 13470 42030 13522 42082
rect 14478 42030 14530 42082
rect 15374 42030 15426 42082
rect 19070 42030 19122 42082
rect 29710 42030 29762 42082
rect 37550 42030 37602 42082
rect 39454 42030 39506 42082
rect 41358 42030 41410 42082
rect 41470 42030 41522 42082
rect 42254 42030 42306 42082
rect 43374 42030 43426 42082
rect 44158 42030 44210 42082
rect 47070 42030 47122 42082
rect 47966 42030 48018 42082
rect 48078 42030 48130 42082
rect 49198 42030 49250 42082
rect 49758 42030 49810 42082
rect 1710 41918 1762 41970
rect 2382 41918 2434 41970
rect 3614 41918 3666 41970
rect 4510 41918 4562 41970
rect 7422 41918 7474 41970
rect 9550 41918 9602 41970
rect 9998 41918 10050 41970
rect 10222 41918 10274 41970
rect 11678 41918 11730 41970
rect 12462 41918 12514 41970
rect 13358 41918 13410 41970
rect 14030 41918 14082 41970
rect 14814 41918 14866 41970
rect 15598 41918 15650 41970
rect 16158 41918 16210 41970
rect 16718 41918 16770 41970
rect 19966 41918 20018 41970
rect 20638 41918 20690 41970
rect 22206 41918 22258 41970
rect 22654 41918 22706 41970
rect 23326 41918 23378 41970
rect 23662 41918 23714 41970
rect 30270 41918 30322 41970
rect 30606 41918 30658 41970
rect 33182 41918 33234 41970
rect 33406 41918 33458 41970
rect 37438 41918 37490 41970
rect 37662 41918 37714 41970
rect 38558 41918 38610 41970
rect 39678 41918 39730 41970
rect 40350 41918 40402 41970
rect 41694 41918 41746 41970
rect 42030 41918 42082 41970
rect 42702 41918 42754 41970
rect 43150 41918 43202 41970
rect 43822 41918 43874 41970
rect 44494 41918 44546 41970
rect 45614 41918 45666 41970
rect 45838 41918 45890 41970
rect 46622 41918 46674 41970
rect 48302 41918 48354 41970
rect 48862 41918 48914 41970
rect 49982 41918 50034 41970
rect 50654 41918 50706 41970
rect 52446 41918 52498 41970
rect 53006 41918 53058 41970
rect 53342 41918 53394 41970
rect 53566 41918 53618 41970
rect 53790 41918 53842 41970
rect 54686 41918 54738 41970
rect 55134 41918 55186 41970
rect 3166 41806 3218 41858
rect 9886 41806 9938 41858
rect 11118 41806 11170 41858
rect 18622 41806 18674 41858
rect 21982 41806 22034 41858
rect 23438 41806 23490 41858
rect 31054 41806 31106 41858
rect 34078 41806 34130 41858
rect 43486 41806 43538 41858
rect 45054 41806 45106 41858
rect 46510 41806 46562 41858
rect 4398 41694 4450 41746
rect 16942 41694 16994 41746
rect 42478 41694 42530 41746
rect 45278 41694 45330 41746
rect 52670 41694 52722 41746
rect 54014 41694 54066 41746
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 10334 41358 10386 41410
rect 32958 41358 33010 41410
rect 38558 41358 38610 41410
rect 44158 41358 44210 41410
rect 45726 41358 45778 41410
rect 45950 41358 46002 41410
rect 50318 41358 50370 41410
rect 51550 41358 51602 41410
rect 53006 41358 53058 41410
rect 10670 41246 10722 41298
rect 13582 41246 13634 41298
rect 18062 41246 18114 41298
rect 23214 41246 23266 41298
rect 37662 41246 37714 41298
rect 42590 41246 42642 41298
rect 43150 41246 43202 41298
rect 44942 41246 44994 41298
rect 45502 41246 45554 41298
rect 47518 41246 47570 41298
rect 48078 41246 48130 41298
rect 51326 41246 51378 41298
rect 54238 41246 54290 41298
rect 2270 41134 2322 41186
rect 2606 41134 2658 41186
rect 3390 41134 3442 41186
rect 4846 41134 4898 41186
rect 5966 41134 6018 41186
rect 6414 41134 6466 41186
rect 6974 41134 7026 41186
rect 7310 41134 7362 41186
rect 8318 41134 8370 41186
rect 8878 41134 8930 41186
rect 8990 41134 9042 41186
rect 9438 41134 9490 41186
rect 12910 41134 12962 41186
rect 15038 41134 15090 41186
rect 17390 41134 17442 41186
rect 18510 41134 18562 41186
rect 19518 41134 19570 41186
rect 19630 41134 19682 41186
rect 19966 41134 20018 41186
rect 21422 41134 21474 41186
rect 21646 41134 21698 41186
rect 23102 41134 23154 41186
rect 30046 41134 30098 41186
rect 32174 41134 32226 41186
rect 32510 41134 32562 41186
rect 36206 41134 36258 41186
rect 37326 41134 37378 41186
rect 37774 41134 37826 41186
rect 38334 41134 38386 41186
rect 39006 41134 39058 41186
rect 39790 41134 39842 41186
rect 40462 41134 40514 41186
rect 40798 41134 40850 41186
rect 42142 41134 42194 41186
rect 42254 41134 42306 41186
rect 42478 41134 42530 41186
rect 43598 41134 43650 41186
rect 43934 41134 43986 41186
rect 47070 41134 47122 41186
rect 48750 41134 48802 41186
rect 49310 41134 49362 41186
rect 49646 41134 49698 41186
rect 50094 41134 50146 41186
rect 51774 41134 51826 41186
rect 52670 41134 52722 41186
rect 55694 41134 55746 41186
rect 4062 41022 4114 41074
rect 5070 41022 5122 41074
rect 7198 41022 7250 41074
rect 9214 41022 9266 41074
rect 9774 41022 9826 41074
rect 10110 41022 10162 41074
rect 12574 41022 12626 41074
rect 13806 41022 13858 41074
rect 16382 41022 16434 41074
rect 18398 41022 18450 41074
rect 19182 41022 19234 41074
rect 19294 41022 19346 41074
rect 22318 41022 22370 41074
rect 23998 41022 24050 41074
rect 29822 41022 29874 41074
rect 31166 41022 31218 41074
rect 32398 41022 32450 41074
rect 37550 41022 37602 41074
rect 38558 41022 38610 41074
rect 41694 41022 41746 41074
rect 46622 41022 46674 41074
rect 49422 41022 49474 41074
rect 50654 41022 50706 41074
rect 54462 41022 54514 41074
rect 5630 40910 5682 40962
rect 6638 40910 6690 40962
rect 7982 40910 8034 40962
rect 12798 40910 12850 40962
rect 16718 40910 16770 40962
rect 17054 40910 17106 40962
rect 19854 40910 19906 40962
rect 31278 40910 31330 40962
rect 33406 40910 33458 40962
rect 36430 40910 36482 40962
rect 37886 40910 37938 40962
rect 40126 40910 40178 40962
rect 41134 40910 41186 40962
rect 41358 40910 41410 40962
rect 41582 40910 41634 40962
rect 42590 40910 42642 40962
rect 46398 40910 46450 40962
rect 48862 40910 48914 40962
rect 49086 40910 49138 40962
rect 52222 40910 52274 40962
rect 52894 40910 52946 40962
rect 56030 40910 56082 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 50558 40742 50610 40794
rect 50662 40742 50714 40794
rect 50766 40742 50818 40794
rect 4510 40574 4562 40626
rect 4958 40574 5010 40626
rect 5294 40574 5346 40626
rect 5854 40574 5906 40626
rect 10670 40574 10722 40626
rect 18846 40574 18898 40626
rect 22766 40574 22818 40626
rect 28478 40574 28530 40626
rect 36318 40574 36370 40626
rect 37326 40574 37378 40626
rect 37998 40574 38050 40626
rect 43710 40574 43762 40626
rect 44158 40574 44210 40626
rect 44718 40574 44770 40626
rect 45390 40574 45442 40626
rect 45950 40574 46002 40626
rect 3502 40462 3554 40514
rect 5518 40462 5570 40514
rect 6190 40462 6242 40514
rect 7086 40462 7138 40514
rect 7870 40462 7922 40514
rect 7982 40462 8034 40514
rect 12238 40462 12290 40514
rect 13134 40462 13186 40514
rect 13246 40462 13298 40514
rect 13358 40462 13410 40514
rect 18398 40462 18450 40514
rect 19518 40462 19570 40514
rect 19630 40462 19682 40514
rect 19854 40462 19906 40514
rect 21534 40462 21586 40514
rect 23550 40462 23602 40514
rect 23662 40462 23714 40514
rect 28702 40462 28754 40514
rect 28814 40462 28866 40514
rect 31838 40462 31890 40514
rect 35086 40462 35138 40514
rect 36542 40462 36594 40514
rect 36654 40462 36706 40514
rect 36990 40462 37042 40514
rect 37662 40462 37714 40514
rect 41246 40462 41298 40514
rect 42814 40462 42866 40514
rect 43038 40462 43090 40514
rect 46286 40462 46338 40514
rect 47182 40462 47234 40514
rect 51662 40462 51714 40514
rect 2606 40350 2658 40402
rect 2942 40350 2994 40402
rect 3278 40350 3330 40402
rect 3614 40350 3666 40402
rect 5070 40350 5122 40402
rect 7310 40350 7362 40402
rect 7646 40350 7698 40402
rect 11118 40350 11170 40402
rect 11566 40350 11618 40402
rect 11902 40350 11954 40402
rect 12686 40350 12738 40402
rect 13806 40350 13858 40402
rect 14142 40350 14194 40402
rect 14590 40350 14642 40402
rect 14702 40350 14754 40402
rect 17390 40350 17442 40402
rect 17950 40350 18002 40402
rect 19070 40350 19122 40402
rect 20190 40350 20242 40402
rect 22430 40350 22482 40402
rect 23326 40350 23378 40402
rect 29038 40350 29090 40402
rect 29822 40350 29874 40402
rect 30158 40350 30210 40402
rect 30382 40350 30434 40402
rect 31390 40350 31442 40402
rect 31502 40350 31554 40402
rect 33070 40350 33122 40402
rect 33966 40350 34018 40402
rect 35758 40350 35810 40402
rect 41022 40350 41074 40402
rect 43262 40350 43314 40402
rect 44606 40350 44658 40402
rect 44942 40350 44994 40402
rect 46622 40350 46674 40402
rect 46846 40350 46898 40402
rect 47406 40350 47458 40402
rect 49534 40350 49586 40402
rect 50206 40350 50258 40402
rect 51998 40350 52050 40402
rect 52894 40350 52946 40402
rect 54910 40350 54962 40402
rect 2046 40238 2098 40290
rect 4062 40238 4114 40290
rect 5182 40238 5234 40290
rect 10222 40238 10274 40290
rect 14366 40238 14418 40290
rect 18398 40238 18450 40290
rect 20974 40238 21026 40290
rect 31726 40238 31778 40290
rect 33854 40238 33906 40290
rect 35870 40238 35922 40290
rect 42702 40238 42754 40290
rect 44046 40238 44098 40290
rect 49310 40238 49362 40290
rect 55134 40238 55186 40290
rect 55582 40238 55634 40290
rect 12574 40126 12626 40178
rect 43934 40126 43986 40178
rect 54238 40126 54290 40178
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 13918 39790 13970 39842
rect 14366 39790 14418 39842
rect 32286 39790 32338 39842
rect 32846 39790 32898 39842
rect 33854 39790 33906 39842
rect 35870 39790 35922 39842
rect 49870 39790 49922 39842
rect 5742 39678 5794 39730
rect 6526 39678 6578 39730
rect 12686 39678 12738 39730
rect 14702 39678 14754 39730
rect 22542 39678 22594 39730
rect 23438 39678 23490 39730
rect 29486 39678 29538 39730
rect 32062 39678 32114 39730
rect 34078 39678 34130 39730
rect 40686 39678 40738 39730
rect 43710 39678 43762 39730
rect 49646 39678 49698 39730
rect 51550 39678 51602 39730
rect 54238 39678 54290 39730
rect 2270 39566 2322 39618
rect 3838 39566 3890 39618
rect 4398 39566 4450 39618
rect 5070 39566 5122 39618
rect 5182 39566 5234 39618
rect 5518 39566 5570 39618
rect 6302 39566 6354 39618
rect 8654 39566 8706 39618
rect 9662 39566 9714 39618
rect 11566 39566 11618 39618
rect 18286 39566 18338 39618
rect 19070 39566 19122 39618
rect 22766 39566 22818 39618
rect 23102 39566 23154 39618
rect 28702 39566 28754 39618
rect 29374 39566 29426 39618
rect 31054 39566 31106 39618
rect 31950 39566 32002 39618
rect 32622 39566 32674 39618
rect 35982 39566 36034 39618
rect 36430 39566 36482 39618
rect 37438 39566 37490 39618
rect 39566 39566 39618 39618
rect 39678 39566 39730 39618
rect 40350 39566 40402 39618
rect 42478 39566 42530 39618
rect 43598 39566 43650 39618
rect 46286 39566 46338 39618
rect 46958 39566 47010 39618
rect 51102 39566 51154 39618
rect 51438 39566 51490 39618
rect 54014 39566 54066 39618
rect 55358 39566 55410 39618
rect 2942 39454 2994 39506
rect 3054 39454 3106 39506
rect 4846 39454 4898 39506
rect 11118 39454 11170 39506
rect 12014 39454 12066 39506
rect 14030 39454 14082 39506
rect 14590 39454 14642 39506
rect 18622 39454 18674 39506
rect 18958 39454 19010 39506
rect 21870 39454 21922 39506
rect 21982 39454 22034 39506
rect 28366 39454 28418 39506
rect 28478 39454 28530 39506
rect 31502 39454 31554 39506
rect 35870 39454 35922 39506
rect 37326 39454 37378 39506
rect 39790 39454 39842 39506
rect 41134 39454 41186 39506
rect 43150 39454 43202 39506
rect 46622 39454 46674 39506
rect 51774 39454 51826 39506
rect 54574 39454 54626 39506
rect 1710 39342 1762 39394
rect 2718 39342 2770 39394
rect 8318 39342 8370 39394
rect 13918 39342 13970 39394
rect 17950 39342 18002 39394
rect 18174 39342 18226 39394
rect 18846 39342 18898 39394
rect 22206 39342 22258 39394
rect 28142 39342 28194 39394
rect 33182 39342 33234 39394
rect 33518 39342 33570 39394
rect 37102 39342 37154 39394
rect 39118 39342 39170 39394
rect 41470 39342 41522 39394
rect 42254 39342 42306 39394
rect 42814 39342 42866 39394
rect 43374 39342 43426 39394
rect 43710 39342 43762 39394
rect 45950 39342 46002 39394
rect 46734 39342 46786 39394
rect 47294 39342 47346 39394
rect 50206 39342 50258 39394
rect 55470 39342 55522 39394
rect 55694 39342 55746 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 50558 39174 50610 39226
rect 50662 39174 50714 39226
rect 50766 39174 50818 39226
rect 2046 39006 2098 39058
rect 2718 39006 2770 39058
rect 3054 39006 3106 39058
rect 3726 39006 3778 39058
rect 4734 39006 4786 39058
rect 5854 39006 5906 39058
rect 6974 39006 7026 39058
rect 8430 39006 8482 39058
rect 8766 39006 8818 39058
rect 10782 39006 10834 39058
rect 11006 39006 11058 39058
rect 13246 39006 13298 39058
rect 13470 39006 13522 39058
rect 16830 39006 16882 39058
rect 28702 39006 28754 39058
rect 30382 39006 30434 39058
rect 42926 39006 42978 39058
rect 44830 39006 44882 39058
rect 45166 39006 45218 39058
rect 51102 39006 51154 39058
rect 4622 38894 4674 38946
rect 6414 38894 6466 38946
rect 6526 38894 6578 38946
rect 6862 38894 6914 38946
rect 10110 38894 10162 38946
rect 10222 38894 10274 38946
rect 10558 38894 10610 38946
rect 14142 38894 14194 38946
rect 17950 38894 18002 38946
rect 18622 38894 18674 38946
rect 21982 38894 22034 38946
rect 23662 38894 23714 38946
rect 25454 38894 25506 38946
rect 29038 38894 29090 38946
rect 29374 38894 29426 38946
rect 29822 38894 29874 38946
rect 29934 38894 29986 38946
rect 31502 38894 31554 38946
rect 37102 38894 37154 38946
rect 38446 38894 38498 38946
rect 39678 38894 39730 38946
rect 41022 38894 41074 38946
rect 42254 38894 42306 38946
rect 45502 38894 45554 38946
rect 46734 38894 46786 38946
rect 47070 38894 47122 38946
rect 51550 38894 51602 38946
rect 1822 38782 1874 38834
rect 4286 38782 4338 38834
rect 5742 38782 5794 38834
rect 6078 38782 6130 38834
rect 11230 38782 11282 38834
rect 12014 38782 12066 38834
rect 12238 38782 12290 38834
rect 12798 38782 12850 38834
rect 15374 38782 15426 38834
rect 16606 38782 16658 38834
rect 17726 38782 17778 38834
rect 19854 38782 19906 38834
rect 20526 38782 20578 38834
rect 20862 38782 20914 38834
rect 21870 38782 21922 38834
rect 22318 38782 22370 38834
rect 22542 38782 22594 38834
rect 22766 38782 22818 38834
rect 23214 38782 23266 38834
rect 23438 38782 23490 38834
rect 31838 38782 31890 38834
rect 35086 38782 35138 38834
rect 35198 38782 35250 38834
rect 38670 38782 38722 38834
rect 39006 38782 39058 38834
rect 39902 38782 39954 38834
rect 40910 38782 40962 38834
rect 41918 38782 41970 38834
rect 43150 38782 43202 38834
rect 45838 38782 45890 38834
rect 46062 38782 46114 38834
rect 49198 38782 49250 38834
rect 50094 38782 50146 38834
rect 50318 38782 50370 38834
rect 51774 38782 51826 38834
rect 52222 38782 52274 38834
rect 53790 38782 53842 38834
rect 55134 38782 55186 38834
rect 10894 38670 10946 38722
rect 11902 38670 11954 38722
rect 13358 38670 13410 38722
rect 13918 38670 13970 38722
rect 16046 38670 16098 38722
rect 18398 38670 18450 38722
rect 21534 38670 21586 38722
rect 23550 38670 23602 38722
rect 25230 38670 25282 38722
rect 31614 38670 31666 38722
rect 31950 38670 32002 38722
rect 34750 38670 34802 38722
rect 36542 38670 36594 38722
rect 39454 38670 39506 38722
rect 41470 38670 41522 38722
rect 46398 38670 46450 38722
rect 48750 38670 48802 38722
rect 49534 38670 49586 38722
rect 51438 38670 51490 38722
rect 54014 38670 54066 38722
rect 57822 38670 57874 38722
rect 58270 38670 58322 38722
rect 4734 38558 4786 38610
rect 6414 38558 6466 38610
rect 6974 38558 7026 38610
rect 10110 38558 10162 38610
rect 25566 38558 25618 38610
rect 29822 38558 29874 38610
rect 34526 38558 34578 38610
rect 50654 38558 50706 38610
rect 52446 38558 52498 38610
rect 55806 38558 55858 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 14366 38222 14418 38274
rect 14590 38222 14642 38274
rect 24334 38222 24386 38274
rect 39678 38222 39730 38274
rect 41806 38222 41858 38274
rect 50542 38222 50594 38274
rect 54910 38222 54962 38274
rect 1822 38110 1874 38162
rect 2270 38110 2322 38162
rect 6078 38110 6130 38162
rect 8878 38110 8930 38162
rect 11118 38110 11170 38162
rect 14142 38110 14194 38162
rect 18510 38110 18562 38162
rect 21870 38110 21922 38162
rect 21982 38110 22034 38162
rect 25566 38110 25618 38162
rect 29598 38110 29650 38162
rect 30158 38110 30210 38162
rect 45950 38110 46002 38162
rect 51214 38110 51266 38162
rect 54686 38110 54738 38162
rect 2158 37998 2210 38050
rect 3390 37998 3442 38050
rect 3838 37998 3890 38050
rect 4734 37998 4786 38050
rect 7646 37998 7698 38050
rect 8206 37998 8258 38050
rect 8766 37998 8818 38050
rect 9662 37998 9714 38050
rect 9998 37998 10050 38050
rect 10334 37998 10386 38050
rect 10894 37998 10946 38050
rect 16718 37998 16770 38050
rect 17166 37998 17218 38050
rect 18734 37998 18786 38050
rect 22206 37998 22258 38050
rect 23886 37998 23938 38050
rect 24110 37998 24162 38050
rect 25006 37998 25058 38050
rect 28254 37998 28306 38050
rect 29822 37998 29874 38050
rect 32734 37998 32786 38050
rect 33630 37998 33682 38050
rect 33966 37998 34018 38050
rect 34862 37998 34914 38050
rect 35086 37998 35138 38050
rect 35534 37998 35586 38050
rect 39118 37998 39170 38050
rect 39342 37998 39394 38050
rect 40238 37998 40290 38050
rect 41134 37998 41186 38050
rect 41582 37998 41634 38050
rect 43598 37998 43650 38050
rect 46622 37998 46674 38050
rect 48526 37998 48578 38050
rect 51438 37998 51490 38050
rect 53230 37998 53282 38050
rect 54238 37998 54290 38050
rect 58046 37998 58098 38050
rect 3950 37886 4002 37938
rect 5070 37886 5122 37938
rect 6414 37886 6466 37938
rect 11566 37886 11618 37938
rect 16270 37886 16322 37938
rect 19406 37886 19458 37938
rect 24446 37886 24498 37938
rect 25902 37886 25954 37938
rect 33294 37886 33346 37938
rect 34302 37886 34354 37938
rect 39566 37886 39618 37938
rect 41246 37886 41298 37938
rect 42478 37886 42530 37938
rect 42702 37886 42754 37938
rect 44158 37886 44210 37938
rect 46286 37886 46338 37938
rect 46398 37886 46450 37938
rect 47070 37886 47122 37938
rect 47406 37886 47458 37938
rect 48302 37886 48354 37938
rect 49646 37886 49698 37938
rect 54014 37886 54066 37938
rect 55806 37886 55858 37938
rect 55918 37886 55970 37938
rect 57486 37886 57538 37938
rect 57822 37886 57874 37938
rect 2382 37774 2434 37826
rect 2606 37774 2658 37826
rect 10110 37774 10162 37826
rect 15038 37774 15090 37826
rect 17390 37774 17442 37826
rect 17502 37774 17554 37826
rect 28590 37774 28642 37826
rect 33182 37774 33234 37826
rect 33406 37774 33458 37826
rect 33854 37774 33906 37826
rect 34974 37774 35026 37826
rect 40350 37774 40402 37826
rect 42142 37774 42194 37826
rect 42590 37774 42642 37826
rect 43262 37774 43314 37826
rect 43822 37774 43874 37826
rect 44046 37774 44098 37826
rect 44942 37774 44994 37826
rect 47182 37774 47234 37826
rect 49534 37774 49586 37826
rect 50318 37774 50370 37826
rect 50430 37774 50482 37826
rect 51774 37774 51826 37826
rect 53454 37774 53506 37826
rect 55246 37774 55298 37826
rect 56142 37774 56194 37826
rect 56926 37774 56978 37826
rect 57150 37774 57202 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 50558 37606 50610 37658
rect 50662 37606 50714 37658
rect 50766 37606 50818 37658
rect 2270 37438 2322 37490
rect 6078 37438 6130 37490
rect 6750 37438 6802 37490
rect 7086 37438 7138 37490
rect 8542 37438 8594 37490
rect 2830 37326 2882 37378
rect 2942 37326 2994 37378
rect 3054 37326 3106 37378
rect 6414 37326 6466 37378
rect 8766 37326 8818 37378
rect 8878 37326 8930 37378
rect 9102 37326 9154 37378
rect 9662 37326 9714 37378
rect 9774 37382 9826 37434
rect 13470 37438 13522 37490
rect 14478 37438 14530 37490
rect 16494 37438 16546 37490
rect 20078 37438 20130 37490
rect 29598 37438 29650 37490
rect 29822 37438 29874 37490
rect 30494 37438 30546 37490
rect 30942 37438 30994 37490
rect 32062 37438 32114 37490
rect 34414 37438 34466 37490
rect 39790 37438 39842 37490
rect 40462 37438 40514 37490
rect 43486 37438 43538 37490
rect 43934 37438 43986 37490
rect 57822 37438 57874 37490
rect 12462 37326 12514 37378
rect 14590 37326 14642 37378
rect 19966 37326 20018 37378
rect 25902 37326 25954 37378
rect 28478 37326 28530 37378
rect 28814 37326 28866 37378
rect 29262 37326 29314 37378
rect 29374 37326 29426 37378
rect 29934 37326 29986 37378
rect 32398 37326 32450 37378
rect 32510 37326 32562 37378
rect 33630 37326 33682 37378
rect 35534 37326 35586 37378
rect 40126 37326 40178 37378
rect 40238 37326 40290 37378
rect 41470 37326 41522 37378
rect 43374 37326 43426 37378
rect 44270 37326 44322 37378
rect 52222 37326 52274 37378
rect 56590 37326 56642 37378
rect 4174 37214 4226 37266
rect 4398 37214 4450 37266
rect 10334 37214 10386 37266
rect 11678 37214 11730 37266
rect 14030 37214 14082 37266
rect 14254 37214 14306 37266
rect 16158 37214 16210 37266
rect 16270 37214 16322 37266
rect 16606 37214 16658 37266
rect 17502 37214 17554 37266
rect 18398 37214 18450 37266
rect 19070 37214 19122 37266
rect 19294 37214 19346 37266
rect 19518 37214 19570 37266
rect 20302 37214 20354 37266
rect 23326 37214 23378 37266
rect 23550 37214 23602 37266
rect 25230 37214 25282 37266
rect 25790 37214 25842 37266
rect 33406 37214 33458 37266
rect 34302 37214 34354 37266
rect 34526 37214 34578 37266
rect 36318 37214 36370 37266
rect 37326 37214 37378 37266
rect 41806 37214 41858 37266
rect 42366 37214 42418 37266
rect 43710 37214 43762 37266
rect 45054 37214 45106 37266
rect 46734 37214 46786 37266
rect 49198 37214 49250 37266
rect 49534 37214 49586 37266
rect 50654 37214 50706 37266
rect 51102 37214 51154 37266
rect 52446 37214 52498 37266
rect 53230 37214 53282 37266
rect 55134 37214 55186 37266
rect 55358 37214 55410 37266
rect 56814 37214 56866 37266
rect 57150 37214 57202 37266
rect 58158 37214 58210 37266
rect 1822 37102 1874 37154
rect 8654 37102 8706 37154
rect 10222 37102 10274 37154
rect 16382 37102 16434 37154
rect 17950 37102 18002 37154
rect 19182 37102 19234 37154
rect 26014 37102 26066 37154
rect 37774 37102 37826 37154
rect 41694 37102 41746 37154
rect 44718 37102 44770 37154
rect 45614 37102 45666 37154
rect 47070 37102 47122 37154
rect 50430 37102 50482 37154
rect 54238 37102 54290 37154
rect 56702 37102 56754 37154
rect 3502 36990 3554 37042
rect 3838 36990 3890 37042
rect 9662 36990 9714 37042
rect 18398 36990 18450 37042
rect 23998 36990 24050 37042
rect 29262 36990 29314 37042
rect 32398 36990 32450 37042
rect 33070 36990 33122 37042
rect 34078 36990 34130 37042
rect 46398 36990 46450 37042
rect 50318 36990 50370 37042
rect 55022 36990 55074 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 10334 36654 10386 36706
rect 23438 36654 23490 36706
rect 24558 36654 24610 36706
rect 33742 36654 33794 36706
rect 53006 36654 53058 36706
rect 54462 36654 54514 36706
rect 3838 36542 3890 36594
rect 4398 36542 4450 36594
rect 8878 36542 8930 36594
rect 18622 36542 18674 36594
rect 20750 36542 20802 36594
rect 21310 36542 21362 36594
rect 23214 36542 23266 36594
rect 25342 36542 25394 36594
rect 29486 36542 29538 36594
rect 41470 36542 41522 36594
rect 53230 36542 53282 36594
rect 57038 36542 57090 36594
rect 2830 36430 2882 36482
rect 3502 36430 3554 36482
rect 4174 36430 4226 36482
rect 7422 36430 7474 36482
rect 8318 36430 8370 36482
rect 8654 36430 8706 36482
rect 9438 36430 9490 36482
rect 10222 36430 10274 36482
rect 12238 36430 12290 36482
rect 12350 36430 12402 36482
rect 12462 36430 12514 36482
rect 14254 36430 14306 36482
rect 15150 36430 15202 36482
rect 17950 36430 18002 36482
rect 20190 36430 20242 36482
rect 21534 36430 21586 36482
rect 21758 36430 21810 36482
rect 22206 36430 22258 36482
rect 22654 36430 22706 36482
rect 24334 36430 24386 36482
rect 24782 36430 24834 36482
rect 25790 36430 25842 36482
rect 29374 36430 29426 36482
rect 30830 36430 30882 36482
rect 32398 36430 32450 36482
rect 32734 36430 32786 36482
rect 33518 36430 33570 36482
rect 36430 36430 36482 36482
rect 37102 36430 37154 36482
rect 37662 36430 37714 36482
rect 38334 36430 38386 36482
rect 38446 36430 38498 36482
rect 39006 36430 39058 36482
rect 40686 36430 40738 36482
rect 41582 36430 41634 36482
rect 41918 36430 41970 36482
rect 44046 36430 44098 36482
rect 44382 36430 44434 36482
rect 44830 36430 44882 36482
rect 45726 36430 45778 36482
rect 46286 36430 46338 36482
rect 46622 36430 46674 36482
rect 47070 36430 47122 36482
rect 50318 36430 50370 36482
rect 51438 36430 51490 36482
rect 51886 36430 51938 36482
rect 54574 36430 54626 36482
rect 1710 36318 1762 36370
rect 2718 36318 2770 36370
rect 8766 36318 8818 36370
rect 9662 36318 9714 36370
rect 9774 36318 9826 36370
rect 10334 36318 10386 36370
rect 14030 36318 14082 36370
rect 16494 36318 16546 36370
rect 18062 36318 18114 36370
rect 18286 36318 18338 36370
rect 18958 36318 19010 36370
rect 23774 36318 23826 36370
rect 23998 36318 24050 36370
rect 24334 36318 24386 36370
rect 26238 36318 26290 36370
rect 30270 36318 30322 36370
rect 36990 36318 37042 36370
rect 40574 36318 40626 36370
rect 41134 36318 41186 36370
rect 42030 36318 42082 36370
rect 43486 36318 43538 36370
rect 43598 36318 43650 36370
rect 45278 36318 45330 36370
rect 48302 36318 48354 36370
rect 51214 36318 51266 36370
rect 54462 36318 54514 36370
rect 56478 36318 56530 36370
rect 58158 36318 58210 36370
rect 2046 36206 2098 36258
rect 2494 36206 2546 36258
rect 7086 36206 7138 36258
rect 7310 36206 7362 36258
rect 10894 36206 10946 36258
rect 12910 36206 12962 36258
rect 22318 36206 22370 36258
rect 22542 36206 22594 36258
rect 24446 36206 24498 36258
rect 31054 36206 31106 36258
rect 36094 36206 36146 36258
rect 38558 36206 38610 36258
rect 40350 36206 40402 36258
rect 41358 36206 41410 36258
rect 42254 36206 42306 36258
rect 43262 36206 43314 36258
rect 44158 36206 44210 36258
rect 45838 36206 45890 36258
rect 46398 36206 46450 36258
rect 47406 36206 47458 36258
rect 48414 36206 48466 36258
rect 48526 36206 48578 36258
rect 49982 36206 50034 36258
rect 51998 36206 52050 36258
rect 52670 36206 52722 36258
rect 55694 36206 55746 36258
rect 57822 36206 57874 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 50558 36038 50610 36090
rect 50662 36038 50714 36090
rect 50766 36038 50818 36090
rect 4734 35870 4786 35922
rect 13918 35870 13970 35922
rect 17502 35870 17554 35922
rect 20638 35870 20690 35922
rect 23438 35870 23490 35922
rect 24558 35870 24610 35922
rect 28254 35870 28306 35922
rect 28478 35870 28530 35922
rect 33742 35870 33794 35922
rect 37886 35870 37938 35922
rect 44606 35870 44658 35922
rect 49086 35870 49138 35922
rect 50766 35870 50818 35922
rect 50990 35870 51042 35922
rect 51326 35870 51378 35922
rect 2494 35758 2546 35810
rect 4958 35758 5010 35810
rect 6078 35758 6130 35810
rect 8206 35758 8258 35810
rect 13022 35758 13074 35810
rect 16606 35758 16658 35810
rect 17614 35758 17666 35810
rect 22542 35758 22594 35810
rect 28926 35758 28978 35810
rect 29822 35758 29874 35810
rect 31838 35758 31890 35810
rect 34190 35758 34242 35810
rect 35422 35758 35474 35810
rect 36318 35758 36370 35810
rect 36542 35758 36594 35810
rect 37326 35758 37378 35810
rect 41246 35758 41298 35810
rect 42478 35758 42530 35810
rect 42590 35758 42642 35810
rect 44942 35758 44994 35810
rect 45278 35758 45330 35810
rect 45390 35758 45442 35810
rect 49310 35758 49362 35810
rect 49646 35758 49698 35810
rect 57822 35758 57874 35810
rect 2606 35646 2658 35698
rect 3614 35646 3666 35698
rect 4398 35646 4450 35698
rect 6414 35646 6466 35698
rect 6638 35646 6690 35698
rect 7310 35646 7362 35698
rect 13246 35646 13298 35698
rect 14142 35646 14194 35698
rect 14478 35646 14530 35698
rect 14702 35646 14754 35698
rect 16270 35646 16322 35698
rect 17390 35646 17442 35698
rect 17950 35646 18002 35698
rect 18622 35646 18674 35698
rect 19518 35646 19570 35698
rect 20190 35646 20242 35698
rect 20526 35646 20578 35698
rect 20862 35646 20914 35698
rect 21758 35646 21810 35698
rect 22094 35646 22146 35698
rect 23550 35646 23602 35698
rect 24446 35646 24498 35698
rect 24782 35646 24834 35698
rect 25342 35646 25394 35698
rect 26126 35646 26178 35698
rect 28590 35646 28642 35698
rect 29262 35646 29314 35698
rect 29710 35646 29762 35698
rect 30046 35646 30098 35698
rect 30494 35646 30546 35698
rect 31166 35646 31218 35698
rect 31614 35646 31666 35698
rect 31950 35646 32002 35698
rect 33630 35646 33682 35698
rect 33966 35646 34018 35698
rect 35086 35646 35138 35698
rect 36878 35646 36930 35698
rect 37102 35646 37154 35698
rect 37438 35646 37490 35698
rect 38110 35646 38162 35698
rect 38446 35646 38498 35698
rect 38782 35646 38834 35698
rect 39230 35646 39282 35698
rect 40126 35646 40178 35698
rect 40910 35646 40962 35698
rect 43262 35646 43314 35698
rect 43934 35646 43986 35698
rect 45614 35646 45666 35698
rect 47406 35646 47458 35698
rect 47630 35646 47682 35698
rect 47854 35646 47906 35698
rect 48638 35646 48690 35698
rect 49982 35646 50034 35698
rect 50654 35646 50706 35698
rect 51214 35646 51266 35698
rect 51550 35646 51602 35698
rect 51998 35646 52050 35698
rect 52222 35646 52274 35698
rect 53678 35646 53730 35698
rect 57150 35646 57202 35698
rect 58158 35646 58210 35698
rect 4174 35534 4226 35586
rect 4958 35534 5010 35586
rect 7422 35534 7474 35586
rect 14926 35534 14978 35586
rect 19294 35534 19346 35586
rect 21982 35534 22034 35586
rect 23998 35534 24050 35586
rect 26014 35534 26066 35586
rect 32398 35534 32450 35586
rect 34414 35534 34466 35586
rect 38334 35534 38386 35586
rect 40014 35534 40066 35586
rect 41134 35534 41186 35586
rect 43150 35534 43202 35586
rect 45950 35534 46002 35586
rect 49198 35534 49250 35586
rect 52670 35534 52722 35586
rect 53454 35534 53506 35586
rect 57598 35534 57650 35586
rect 15038 35422 15090 35474
rect 23438 35422 23490 35474
rect 25566 35422 25618 35474
rect 31278 35422 31330 35474
rect 34750 35422 34802 35474
rect 35086 35422 35138 35474
rect 36654 35422 36706 35474
rect 43486 35422 43538 35474
rect 48302 35422 48354 35474
rect 52334 35422 52386 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 3166 35086 3218 35138
rect 9774 35086 9826 35138
rect 33406 35086 33458 35138
rect 53006 35086 53058 35138
rect 4510 34974 4562 35026
rect 8430 34974 8482 35026
rect 9214 34974 9266 35026
rect 11566 34974 11618 35026
rect 17838 34974 17890 35026
rect 22766 34974 22818 35026
rect 25230 34974 25282 35026
rect 30382 34974 30434 35026
rect 33630 34974 33682 35026
rect 34974 34974 35026 35026
rect 37102 34974 37154 35026
rect 39566 34974 39618 35026
rect 40014 34974 40066 35026
rect 47518 34974 47570 35026
rect 50990 34974 51042 35026
rect 53566 34974 53618 35026
rect 3054 34862 3106 34914
rect 4174 34862 4226 34914
rect 5070 34862 5122 34914
rect 7086 34862 7138 34914
rect 8766 34862 8818 34914
rect 10670 34862 10722 34914
rect 11118 34862 11170 34914
rect 14030 34862 14082 34914
rect 14366 34862 14418 34914
rect 17390 34862 17442 34914
rect 17950 34862 18002 34914
rect 18846 34862 18898 34914
rect 19742 34862 19794 34914
rect 22430 34862 22482 34914
rect 23438 34862 23490 34914
rect 23774 34862 23826 34914
rect 24334 34862 24386 34914
rect 25342 34862 25394 34914
rect 26014 34862 26066 34914
rect 26350 34862 26402 34914
rect 26686 34862 26738 34914
rect 26910 34862 26962 34914
rect 29150 34862 29202 34914
rect 29374 34862 29426 34914
rect 29710 34862 29762 34914
rect 31278 34862 31330 34914
rect 31502 34862 31554 34914
rect 31838 34862 31890 34914
rect 32398 34862 32450 34914
rect 32734 34862 32786 34914
rect 33182 34862 33234 34914
rect 34414 34862 34466 34914
rect 35310 34862 35362 34914
rect 36094 34862 36146 34914
rect 37662 34862 37714 34914
rect 37998 34862 38050 34914
rect 40126 34862 40178 34914
rect 41358 34862 41410 34914
rect 43262 34862 43314 34914
rect 43598 34862 43650 34914
rect 45278 34862 45330 34914
rect 48974 34862 49026 34914
rect 55022 34862 55074 34914
rect 2830 34750 2882 34802
rect 3278 34750 3330 34802
rect 6190 34750 6242 34802
rect 6862 34750 6914 34802
rect 9886 34750 9938 34802
rect 18286 34750 18338 34802
rect 19518 34750 19570 34802
rect 20078 34750 20130 34802
rect 22654 34750 22706 34802
rect 23886 34750 23938 34802
rect 32286 34750 32338 34802
rect 33742 34750 33794 34802
rect 34526 34750 34578 34802
rect 35982 34750 36034 34802
rect 37438 34750 37490 34802
rect 47742 34750 47794 34802
rect 50318 34750 50370 34802
rect 53006 34750 53058 34802
rect 53118 34750 53170 34802
rect 53790 34750 53842 34802
rect 58158 34750 58210 34802
rect 6526 34638 6578 34690
rect 9774 34638 9826 34690
rect 14254 34638 14306 34690
rect 18958 34638 19010 34690
rect 19182 34638 19234 34690
rect 19630 34638 19682 34690
rect 22094 34638 22146 34690
rect 26574 34638 26626 34690
rect 29486 34638 29538 34690
rect 29598 34638 29650 34690
rect 31502 34638 31554 34690
rect 32174 34638 32226 34690
rect 35758 34638 35810 34690
rect 37326 34638 37378 34690
rect 38334 34638 38386 34690
rect 41134 34638 41186 34690
rect 41246 34638 41298 34690
rect 41582 34638 41634 34690
rect 43374 34638 43426 34690
rect 45054 34638 45106 34690
rect 55358 34638 55410 34690
rect 57598 34638 57650 34690
rect 57822 34638 57874 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 50558 34470 50610 34522
rect 50662 34470 50714 34522
rect 50766 34470 50818 34522
rect 2046 34302 2098 34354
rect 6862 34302 6914 34354
rect 7198 34302 7250 34354
rect 8094 34302 8146 34354
rect 9774 34302 9826 34354
rect 11230 34302 11282 34354
rect 21646 34302 21698 34354
rect 22990 34302 23042 34354
rect 25454 34302 25506 34354
rect 27918 34302 27970 34354
rect 29598 34302 29650 34354
rect 31502 34302 31554 34354
rect 34302 34302 34354 34354
rect 34862 34302 34914 34354
rect 35982 34302 36034 34354
rect 38782 34302 38834 34354
rect 42254 34302 42306 34354
rect 43262 34302 43314 34354
rect 47742 34302 47794 34354
rect 50766 34302 50818 34354
rect 4174 34190 4226 34242
rect 8542 34190 8594 34242
rect 8654 34190 8706 34242
rect 9886 34190 9938 34242
rect 10670 34190 10722 34242
rect 11678 34190 11730 34242
rect 11790 34190 11842 34242
rect 16606 34190 16658 34242
rect 18398 34190 18450 34242
rect 19182 34190 19234 34242
rect 21534 34190 21586 34242
rect 22318 34190 22370 34242
rect 22430 34190 22482 34242
rect 26126 34190 26178 34242
rect 27694 34190 27746 34242
rect 28814 34190 28866 34242
rect 28926 34190 28978 34242
rect 29486 34190 29538 34242
rect 31054 34190 31106 34242
rect 33742 34190 33794 34242
rect 36206 34190 36258 34242
rect 36318 34190 36370 34242
rect 37326 34190 37378 34242
rect 39006 34190 39058 34242
rect 40014 34190 40066 34242
rect 42590 34190 42642 34242
rect 45166 34190 45218 34242
rect 45502 34190 45554 34242
rect 45726 34190 45778 34242
rect 45838 34190 45890 34242
rect 47518 34190 47570 34242
rect 47966 34190 48018 34242
rect 48078 34190 48130 34242
rect 48974 34190 49026 34242
rect 49198 34190 49250 34242
rect 51774 34190 51826 34242
rect 53342 34190 53394 34242
rect 57822 34190 57874 34242
rect 1710 34078 1762 34130
rect 4398 34078 4450 34130
rect 5070 34078 5122 34130
rect 5854 34078 5906 34130
rect 8766 34078 8818 34130
rect 9550 34078 9602 34130
rect 10558 34078 10610 34130
rect 11118 34078 11170 34130
rect 12014 34078 12066 34130
rect 12686 34078 12738 34130
rect 13134 34078 13186 34130
rect 13582 34078 13634 34130
rect 13918 34078 13970 34130
rect 14366 34078 14418 34130
rect 14702 34078 14754 34130
rect 16718 34078 16770 34130
rect 17950 34078 18002 34130
rect 20302 34078 20354 34130
rect 21422 34078 21474 34130
rect 21982 34078 22034 34130
rect 23438 34078 23490 34130
rect 23662 34078 23714 34130
rect 24334 34078 24386 34130
rect 25230 34078 25282 34130
rect 25902 34078 25954 34130
rect 26350 34078 26402 34130
rect 27470 34078 27522 34130
rect 28590 34078 28642 34130
rect 29150 34078 29202 34130
rect 29822 34078 29874 34130
rect 30382 34078 30434 34130
rect 30830 34078 30882 34130
rect 31390 34078 31442 34130
rect 31614 34078 31666 34130
rect 32062 34078 32114 34130
rect 33966 34078 34018 34130
rect 34638 34078 34690 34130
rect 36542 34078 36594 34130
rect 36878 34078 36930 34130
rect 37102 34078 37154 34130
rect 37886 34078 37938 34130
rect 38446 34078 38498 34130
rect 40350 34078 40402 34130
rect 40910 34078 40962 34130
rect 41134 34078 41186 34130
rect 41358 34078 41410 34130
rect 41806 34078 41858 34130
rect 42030 34078 42082 34130
rect 42254 34078 42306 34130
rect 43038 34078 43090 34130
rect 43150 34078 43202 34130
rect 43598 34078 43650 34130
rect 45054 34078 45106 34130
rect 48750 34078 48802 34130
rect 49310 34078 49362 34130
rect 49758 34078 49810 34130
rect 50654 34078 50706 34130
rect 51662 34078 51714 34130
rect 53790 34078 53842 34130
rect 54238 34078 54290 34130
rect 55694 34078 55746 34130
rect 58158 34078 58210 34130
rect 2494 33966 2546 34018
rect 4510 33966 4562 34018
rect 6302 33966 6354 34018
rect 14926 33966 14978 34018
rect 17502 33966 17554 34018
rect 18846 33966 18898 34018
rect 20974 33966 21026 34018
rect 25342 33966 25394 34018
rect 30606 33966 30658 34018
rect 34750 33966 34802 34018
rect 37214 33966 37266 34018
rect 37662 33966 37714 34018
rect 40126 33966 40178 34018
rect 57598 33966 57650 34018
rect 16606 33854 16658 33906
rect 22318 33854 22370 33906
rect 26686 33854 26738 33906
rect 28030 33854 28082 33906
rect 28142 33854 28194 33906
rect 38222 33854 38274 33906
rect 38670 33854 38722 33906
rect 45166 33854 45218 33906
rect 47406 33854 47458 33906
rect 54798 33854 54850 33906
rect 55246 33854 55298 33906
rect 55470 33854 55522 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 4062 33518 4114 33570
rect 15710 33518 15762 33570
rect 17390 33518 17442 33570
rect 27806 33518 27858 33570
rect 28254 33518 28306 33570
rect 28478 33518 28530 33570
rect 39566 33518 39618 33570
rect 41134 33518 41186 33570
rect 44158 33518 44210 33570
rect 5966 33406 6018 33458
rect 13582 33406 13634 33458
rect 16494 33406 16546 33458
rect 17838 33406 17890 33458
rect 31838 33406 31890 33458
rect 37102 33406 37154 33458
rect 39678 33406 39730 33458
rect 42814 33406 42866 33458
rect 45390 33406 45442 33458
rect 45838 33406 45890 33458
rect 48750 33406 48802 33458
rect 50318 33406 50370 33458
rect 53342 33406 53394 33458
rect 2382 33294 2434 33346
rect 2718 33294 2770 33346
rect 3726 33294 3778 33346
rect 6414 33294 6466 33346
rect 6974 33294 7026 33346
rect 7982 33294 8034 33346
rect 8990 33294 9042 33346
rect 10558 33294 10610 33346
rect 11006 33294 11058 33346
rect 14030 33294 14082 33346
rect 15038 33294 15090 33346
rect 16830 33294 16882 33346
rect 17278 33294 17330 33346
rect 17950 33294 18002 33346
rect 18846 33294 18898 33346
rect 19182 33294 19234 33346
rect 19406 33294 19458 33346
rect 22318 33294 22370 33346
rect 22542 33294 22594 33346
rect 24894 33294 24946 33346
rect 25454 33294 25506 33346
rect 32062 33294 32114 33346
rect 34302 33294 34354 33346
rect 34638 33294 34690 33346
rect 34974 33294 35026 33346
rect 35086 33294 35138 33346
rect 35534 33294 35586 33346
rect 35646 33294 35698 33346
rect 35758 33294 35810 33346
rect 38670 33294 38722 33346
rect 41022 33294 41074 33346
rect 42590 33294 42642 33346
rect 45278 33294 45330 33346
rect 47182 33294 47234 33346
rect 47406 33294 47458 33346
rect 47742 33294 47794 33346
rect 48190 33294 48242 33346
rect 48974 33294 49026 33346
rect 49982 33294 50034 33346
rect 50654 33294 50706 33346
rect 51774 33294 51826 33346
rect 51998 33294 52050 33346
rect 55246 33294 55298 33346
rect 55470 33294 55522 33346
rect 5966 33182 6018 33234
rect 8654 33182 8706 33234
rect 22766 33182 22818 33234
rect 25342 33182 25394 33234
rect 27694 33182 27746 33234
rect 27918 33182 27970 33234
rect 32846 33182 32898 33234
rect 32958 33182 33010 33234
rect 37326 33182 37378 33234
rect 44158 33182 44210 33234
rect 44270 33182 44322 33234
rect 48414 33182 48466 33234
rect 49870 33182 49922 33234
rect 50094 33182 50146 33234
rect 51102 33182 51154 33234
rect 52670 33182 52722 33234
rect 52782 33182 52834 33234
rect 55022 33182 55074 33234
rect 58158 33182 58210 33234
rect 7310 33070 7362 33122
rect 7422 33070 7474 33122
rect 7534 33070 7586 33122
rect 9662 33070 9714 33122
rect 9998 33070 10050 33122
rect 19070 33070 19122 33122
rect 25118 33070 25170 33122
rect 29374 33070 29426 33122
rect 30382 33070 30434 33122
rect 32398 33070 32450 33122
rect 32622 33070 32674 33122
rect 34750 33070 34802 33122
rect 39006 33070 39058 33122
rect 47518 33070 47570 33122
rect 48526 33070 48578 33122
rect 53006 33070 53058 33122
rect 55358 33070 55410 33122
rect 57598 33070 57650 33122
rect 57822 33070 57874 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 50558 32902 50610 32954
rect 50662 32902 50714 32954
rect 50766 32902 50818 32954
rect 3614 32734 3666 32786
rect 6190 32734 6242 32786
rect 7982 32734 8034 32786
rect 9662 32734 9714 32786
rect 18398 32734 18450 32786
rect 31054 32734 31106 32786
rect 37550 32734 37602 32786
rect 39678 32734 39730 32786
rect 46286 32734 46338 32786
rect 46734 32734 46786 32786
rect 49422 32734 49474 32786
rect 2382 32622 2434 32674
rect 3726 32622 3778 32674
rect 6078 32622 6130 32674
rect 7758 32622 7810 32674
rect 10334 32622 10386 32674
rect 10670 32622 10722 32674
rect 11118 32622 11170 32674
rect 13694 32622 13746 32674
rect 14926 32622 14978 32674
rect 15262 32622 15314 32674
rect 16382 32622 16434 32674
rect 17390 32622 17442 32674
rect 18286 32622 18338 32674
rect 20078 32622 20130 32674
rect 23214 32622 23266 32674
rect 26126 32622 26178 32674
rect 26910 32622 26962 32674
rect 28366 32622 28418 32674
rect 32062 32622 32114 32674
rect 42702 32622 42754 32674
rect 43262 32622 43314 32674
rect 48862 32622 48914 32674
rect 49534 32622 49586 32674
rect 57822 32622 57874 32674
rect 2606 32510 2658 32562
rect 6302 32510 6354 32562
rect 6750 32510 6802 32562
rect 7086 32510 7138 32562
rect 7422 32510 7474 32562
rect 9774 32510 9826 32562
rect 11230 32510 11282 32562
rect 15710 32510 15762 32562
rect 16270 32510 16322 32562
rect 17726 32510 17778 32562
rect 17838 32510 17890 32562
rect 19966 32510 20018 32562
rect 20302 32510 20354 32562
rect 22318 32510 22370 32562
rect 22542 32510 22594 32562
rect 24222 32510 24274 32562
rect 26238 32510 26290 32562
rect 26686 32510 26738 32562
rect 27582 32510 27634 32562
rect 28590 32510 28642 32562
rect 29822 32510 29874 32562
rect 30046 32510 30098 32562
rect 30718 32510 30770 32562
rect 32286 32510 32338 32562
rect 32622 32510 32674 32562
rect 33630 32510 33682 32562
rect 37662 32510 37714 32562
rect 37774 32510 37826 32562
rect 38222 32510 38274 32562
rect 38894 32510 38946 32562
rect 41470 32510 41522 32562
rect 42366 32510 42418 32562
rect 42926 32510 42978 32562
rect 43150 32510 43202 32562
rect 45390 32510 45442 32562
rect 45838 32510 45890 32562
rect 46398 32510 46450 32562
rect 46510 32510 46562 32562
rect 48750 32510 48802 32562
rect 50766 32510 50818 32562
rect 50990 32510 51042 32562
rect 51886 32510 51938 32562
rect 52894 32510 52946 32562
rect 58158 32510 58210 32562
rect 6974 32398 7026 32450
rect 7870 32398 7922 32450
rect 13134 32398 13186 32450
rect 16718 32398 16770 32450
rect 18062 32398 18114 32450
rect 22766 32398 22818 32450
rect 23326 32398 23378 32450
rect 23774 32398 23826 32450
rect 24670 32398 24722 32450
rect 26350 32398 26402 32450
rect 28702 32398 28754 32450
rect 31726 32398 31778 32450
rect 32062 32398 32114 32450
rect 33182 32398 33234 32450
rect 34078 32398 34130 32450
rect 39006 32398 39058 32450
rect 41582 32398 41634 32450
rect 43710 32398 43762 32450
rect 44382 32398 44434 32450
rect 51774 32398 51826 32450
rect 57150 32398 57202 32450
rect 57598 32398 57650 32450
rect 9662 32286 9714 32338
rect 11118 32286 11170 32338
rect 38558 32286 38610 32338
rect 48862 32286 48914 32338
rect 49422 32286 49474 32338
rect 50430 32286 50482 32338
rect 53566 32286 53618 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 25118 31950 25170 32002
rect 39790 31950 39842 32002
rect 48750 31950 48802 32002
rect 4174 31838 4226 31890
rect 6638 31838 6690 31890
rect 7198 31838 7250 31890
rect 11342 31838 11394 31890
rect 17390 31838 17442 31890
rect 19630 31838 19682 31890
rect 26126 31838 26178 31890
rect 33182 31838 33234 31890
rect 34526 31838 34578 31890
rect 34862 31838 34914 31890
rect 36094 31838 36146 31890
rect 36990 31838 37042 31890
rect 39230 31838 39282 31890
rect 40350 31838 40402 31890
rect 42366 31838 42418 31890
rect 46846 31838 46898 31890
rect 49310 31838 49362 31890
rect 3278 31726 3330 31778
rect 3614 31726 3666 31778
rect 3726 31726 3778 31778
rect 3950 31726 4002 31778
rect 5070 31726 5122 31778
rect 6078 31726 6130 31778
rect 6974 31726 7026 31778
rect 11118 31726 11170 31778
rect 11790 31726 11842 31778
rect 12126 31726 12178 31778
rect 12574 31726 12626 31778
rect 16718 31726 16770 31778
rect 17726 31726 17778 31778
rect 18174 31726 18226 31778
rect 18510 31726 18562 31778
rect 18846 31726 18898 31778
rect 19966 31726 20018 31778
rect 20190 31726 20242 31778
rect 24110 31726 24162 31778
rect 24894 31726 24946 31778
rect 25342 31726 25394 31778
rect 25678 31726 25730 31778
rect 26574 31726 26626 31778
rect 27806 31726 27858 31778
rect 28254 31726 28306 31778
rect 29374 31726 29426 31778
rect 30942 31726 30994 31778
rect 31390 31726 31442 31778
rect 31838 31726 31890 31778
rect 33518 31726 33570 31778
rect 35198 31726 35250 31778
rect 38110 31726 38162 31778
rect 38558 31726 38610 31778
rect 39454 31726 39506 31778
rect 42478 31726 42530 31778
rect 43710 31726 43762 31778
rect 45502 31726 45554 31778
rect 45838 31726 45890 31778
rect 47966 31726 48018 31778
rect 48638 31726 48690 31778
rect 49422 31726 49474 31778
rect 50766 31726 50818 31778
rect 54574 31726 54626 31778
rect 55134 31726 55186 31778
rect 4510 31614 4562 31666
rect 7870 31614 7922 31666
rect 7982 31614 8034 31666
rect 8654 31614 8706 31666
rect 11566 31614 11618 31666
rect 14142 31614 14194 31666
rect 14926 31614 14978 31666
rect 15038 31614 15090 31666
rect 15486 31614 15538 31666
rect 18622 31614 18674 31666
rect 19294 31614 19346 31666
rect 19518 31614 19570 31666
rect 20414 31614 20466 31666
rect 24446 31614 24498 31666
rect 26014 31614 26066 31666
rect 26350 31614 26402 31666
rect 29150 31614 29202 31666
rect 36206 31614 36258 31666
rect 36430 31614 36482 31666
rect 37102 31614 37154 31666
rect 37326 31614 37378 31666
rect 39678 31614 39730 31666
rect 39790 31614 39842 31666
rect 43374 31614 43426 31666
rect 44942 31614 44994 31666
rect 45166 31614 45218 31666
rect 45950 31614 46002 31666
rect 46286 31614 46338 31666
rect 51550 31614 51602 31666
rect 53342 31614 53394 31666
rect 53678 31614 53730 31666
rect 53902 31614 53954 31666
rect 54238 31614 54290 31666
rect 56926 31614 56978 31666
rect 57486 31614 57538 31666
rect 4286 31502 4338 31554
rect 4734 31502 4786 31554
rect 4958 31502 5010 31554
rect 6190 31502 6242 31554
rect 6414 31502 6466 31554
rect 7646 31502 7698 31554
rect 8318 31502 8370 31554
rect 8542 31502 8594 31554
rect 9550 31502 9602 31554
rect 9886 31502 9938 31554
rect 12014 31502 12066 31554
rect 13918 31502 13970 31554
rect 14030 31502 14082 31554
rect 14366 31502 14418 31554
rect 14702 31502 14754 31554
rect 16494 31502 16546 31554
rect 20078 31502 20130 31554
rect 24222 31502 24274 31554
rect 25454 31502 25506 31554
rect 30382 31502 30434 31554
rect 42590 31502 42642 31554
rect 43150 31502 43202 31554
rect 44158 31502 44210 31554
rect 44830 31502 44882 31554
rect 46062 31502 46114 31554
rect 53454 31502 53506 31554
rect 54798 31502 54850 31554
rect 55022 31502 55074 31554
rect 57150 31502 57202 31554
rect 57822 31502 57874 31554
rect 58158 31502 58210 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 50558 31334 50610 31386
rect 50662 31334 50714 31386
rect 50766 31334 50818 31386
rect 2718 31166 2770 31218
rect 10894 31166 10946 31218
rect 11230 31166 11282 31218
rect 15934 31166 15986 31218
rect 17614 31166 17666 31218
rect 23214 31166 23266 31218
rect 26238 31166 26290 31218
rect 27918 31166 27970 31218
rect 28926 31166 28978 31218
rect 30046 31166 30098 31218
rect 37214 31166 37266 31218
rect 38110 31166 38162 31218
rect 39790 31166 39842 31218
rect 2830 31054 2882 31106
rect 4622 31054 4674 31106
rect 7198 31054 7250 31106
rect 11678 31054 11730 31106
rect 11790 31054 11842 31106
rect 12350 31054 12402 31106
rect 12462 31054 12514 31106
rect 13918 31054 13970 31106
rect 15598 31054 15650 31106
rect 17390 31054 17442 31106
rect 20078 31054 20130 31106
rect 21982 31054 22034 31106
rect 22094 31054 22146 31106
rect 23550 31054 23602 31106
rect 24558 31054 24610 31106
rect 28478 31054 28530 31106
rect 32510 31054 32562 31106
rect 36990 31054 37042 31106
rect 43822 31054 43874 31106
rect 44606 31054 44658 31106
rect 46174 31054 46226 31106
rect 47966 31054 48018 31106
rect 49198 31054 49250 31106
rect 49422 31054 49474 31106
rect 50094 31054 50146 31106
rect 52446 31054 52498 31106
rect 57822 31054 57874 31106
rect 2494 30942 2546 30994
rect 3502 30942 3554 30994
rect 3726 30942 3778 30994
rect 4062 30942 4114 30994
rect 4286 30942 4338 30994
rect 5406 30942 5458 30994
rect 6302 30942 6354 30994
rect 6862 30942 6914 30994
rect 7982 30942 8034 30994
rect 8654 30942 8706 30994
rect 9550 30942 9602 30994
rect 9662 30942 9714 30994
rect 11454 30942 11506 30994
rect 13022 30942 13074 30994
rect 14702 30942 14754 30994
rect 16270 30942 16322 30994
rect 17838 30942 17890 30994
rect 17950 30942 18002 30994
rect 20974 30942 21026 30994
rect 22878 30942 22930 30994
rect 23326 30942 23378 30994
rect 25902 30942 25954 30994
rect 26910 30942 26962 30994
rect 28254 30942 28306 30994
rect 28926 30942 28978 30994
rect 29822 30942 29874 30994
rect 32286 30942 32338 30994
rect 36094 30942 36146 30994
rect 38446 30942 38498 30994
rect 38670 30942 38722 30994
rect 41358 30942 41410 30994
rect 42814 30942 42866 30994
rect 43150 30942 43202 30994
rect 45278 30942 45330 30994
rect 45838 30942 45890 30994
rect 46062 30942 46114 30994
rect 47294 30942 47346 30994
rect 48190 30942 48242 30994
rect 49310 30942 49362 30994
rect 50206 30942 50258 30994
rect 50430 30942 50482 30994
rect 50878 30942 50930 30994
rect 51550 30942 51602 30994
rect 52334 30942 52386 30994
rect 52894 30942 52946 30994
rect 54350 30942 54402 30994
rect 58158 30942 58210 30994
rect 3838 30830 3890 30882
rect 6190 30830 6242 30882
rect 8542 30830 8594 30882
rect 13134 30830 13186 30882
rect 14366 30830 14418 30882
rect 15262 30830 15314 30882
rect 17726 30830 17778 30882
rect 19518 30830 19570 30882
rect 21646 30830 21698 30882
rect 24334 30830 24386 30882
rect 24670 30830 24722 30882
rect 25678 30830 25730 30882
rect 26574 30830 26626 30882
rect 26686 30830 26738 30882
rect 30494 30830 30546 30882
rect 31838 30830 31890 30882
rect 35422 30830 35474 30882
rect 39342 30830 39394 30882
rect 47630 30830 47682 30882
rect 51102 30830 51154 30882
rect 51326 30830 51378 30882
rect 53902 30830 53954 30882
rect 57598 30830 57650 30882
rect 6862 30718 6914 30770
rect 8654 30718 8706 30770
rect 12350 30718 12402 30770
rect 16494 30718 16546 30770
rect 16830 30718 16882 30770
rect 22094 30718 22146 30770
rect 29038 30718 29090 30770
rect 29262 30718 29314 30770
rect 34862 30718 34914 30770
rect 35198 30718 35250 30770
rect 35758 30718 35810 30770
rect 36094 30718 36146 30770
rect 37326 30718 37378 30770
rect 46622 30718 46674 30770
rect 48750 30718 48802 30770
rect 50094 30718 50146 30770
rect 53566 30718 53618 30770
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 4510 30382 4562 30434
rect 4734 30382 4786 30434
rect 7086 30382 7138 30434
rect 8990 30382 9042 30434
rect 21422 30382 21474 30434
rect 24670 30382 24722 30434
rect 28590 30382 28642 30434
rect 30494 30382 30546 30434
rect 32398 30382 32450 30434
rect 38894 30382 38946 30434
rect 39902 30382 39954 30434
rect 44046 30382 44098 30434
rect 44830 30382 44882 30434
rect 45390 30382 45442 30434
rect 45614 30382 45666 30434
rect 46398 30382 46450 30434
rect 6078 30270 6130 30322
rect 9886 30270 9938 30322
rect 17614 30270 17666 30322
rect 20190 30270 20242 30322
rect 21758 30270 21810 30322
rect 23550 30270 23602 30322
rect 29710 30270 29762 30322
rect 29934 30270 29986 30322
rect 31614 30270 31666 30322
rect 39230 30270 39282 30322
rect 40126 30270 40178 30322
rect 42590 30270 42642 30322
rect 43374 30270 43426 30322
rect 43822 30270 43874 30322
rect 47854 30270 47906 30322
rect 2494 30158 2546 30210
rect 3502 30158 3554 30210
rect 4286 30158 4338 30210
rect 6302 30158 6354 30210
rect 6638 30158 6690 30210
rect 7198 30158 7250 30210
rect 7982 30158 8034 30210
rect 8654 30158 8706 30210
rect 9214 30158 9266 30210
rect 10334 30158 10386 30210
rect 12686 30158 12738 30210
rect 13022 30158 13074 30210
rect 13470 30158 13522 30210
rect 13806 30158 13858 30210
rect 13918 30158 13970 30210
rect 14366 30158 14418 30210
rect 16606 30158 16658 30210
rect 16942 30158 16994 30210
rect 17166 30158 17218 30210
rect 17390 30158 17442 30210
rect 19742 30158 19794 30210
rect 22094 30158 22146 30210
rect 22318 30158 22370 30210
rect 23102 30158 23154 30210
rect 23326 30158 23378 30210
rect 24110 30158 24162 30210
rect 24334 30158 24386 30210
rect 24894 30158 24946 30210
rect 25230 30158 25282 30210
rect 26126 30158 26178 30210
rect 27022 30158 27074 30210
rect 27806 30158 27858 30210
rect 29486 30158 29538 30210
rect 31278 30158 31330 30210
rect 32510 30158 32562 30210
rect 34078 30158 34130 30210
rect 35086 30158 35138 30210
rect 36206 30158 36258 30210
rect 36990 30158 37042 30210
rect 37662 30158 37714 30210
rect 38670 30158 38722 30210
rect 39790 30158 39842 30210
rect 41470 30158 41522 30210
rect 41918 30158 41970 30210
rect 42142 30158 42194 30210
rect 43710 30158 43762 30210
rect 44270 30158 44322 30210
rect 44942 30158 44994 30210
rect 46622 30158 46674 30210
rect 47630 30158 47682 30210
rect 55582 30158 55634 30210
rect 2382 30046 2434 30098
rect 4846 30046 4898 30098
rect 7086 30046 7138 30098
rect 10782 30046 10834 30098
rect 14590 30046 14642 30098
rect 17950 30046 18002 30098
rect 19294 30046 19346 30098
rect 25342 30046 25394 30098
rect 26350 30046 26402 30098
rect 26910 30046 26962 30098
rect 28478 30046 28530 30098
rect 30270 30046 30322 30098
rect 31502 30046 31554 30098
rect 31950 30046 32002 30098
rect 32174 30046 32226 30098
rect 35310 30046 35362 30098
rect 36094 30046 36146 30098
rect 37326 30046 37378 30098
rect 39118 30046 39170 30098
rect 39342 30046 39394 30098
rect 40238 30046 40290 30098
rect 41134 30046 41186 30098
rect 41246 30046 41298 30098
rect 42478 30046 42530 30098
rect 43038 30046 43090 30098
rect 43262 30046 43314 30098
rect 45166 30046 45218 30098
rect 47294 30046 47346 30098
rect 57262 30046 57314 30098
rect 3614 29934 3666 29986
rect 12798 29934 12850 29986
rect 13582 29934 13634 29986
rect 14254 29934 14306 29986
rect 17054 29934 17106 29986
rect 17726 29934 17778 29986
rect 21646 29934 21698 29986
rect 24222 29934 24274 29986
rect 25566 29934 25618 29986
rect 28254 29934 28306 29986
rect 29038 29934 29090 29986
rect 30830 29934 30882 29986
rect 32734 29934 32786 29986
rect 33742 29934 33794 29986
rect 35198 29934 35250 29986
rect 37214 29934 37266 29986
rect 37774 29934 37826 29986
rect 37886 29934 37938 29986
rect 38110 29934 38162 29986
rect 40910 29934 40962 29986
rect 41694 29934 41746 29986
rect 46062 29934 46114 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 50558 29766 50610 29818
rect 50662 29766 50714 29818
rect 50766 29766 50818 29818
rect 3838 29598 3890 29650
rect 11454 29598 11506 29650
rect 3166 29486 3218 29538
rect 3278 29486 3330 29538
rect 3390 29486 3442 29538
rect 4398 29486 4450 29538
rect 10670 29486 10722 29538
rect 14478 29486 14530 29538
rect 14590 29542 14642 29594
rect 15038 29598 15090 29650
rect 15598 29598 15650 29650
rect 15934 29598 15986 29650
rect 16606 29598 16658 29650
rect 16830 29598 16882 29650
rect 17614 29598 17666 29650
rect 22206 29598 22258 29650
rect 22542 29598 22594 29650
rect 27134 29598 27186 29650
rect 28142 29598 28194 29650
rect 30046 29598 30098 29650
rect 30382 29598 30434 29650
rect 32062 29598 32114 29650
rect 33518 29598 33570 29650
rect 35758 29598 35810 29650
rect 43822 29598 43874 29650
rect 43934 29598 43986 29650
rect 44718 29598 44770 29650
rect 45390 29598 45442 29650
rect 45950 29598 46002 29650
rect 57598 29598 57650 29650
rect 16046 29486 16098 29538
rect 21758 29486 21810 29538
rect 26798 29486 26850 29538
rect 28478 29486 28530 29538
rect 28702 29486 28754 29538
rect 31726 29486 31778 29538
rect 35310 29486 35362 29538
rect 35982 29486 36034 29538
rect 36766 29486 36818 29538
rect 37102 29486 37154 29538
rect 37326 29486 37378 29538
rect 45502 29486 45554 29538
rect 57822 29486 57874 29538
rect 58158 29486 58210 29538
rect 4174 29374 4226 29426
rect 5070 29374 5122 29426
rect 7310 29374 7362 29426
rect 7758 29374 7810 29426
rect 8430 29374 8482 29426
rect 10446 29374 10498 29426
rect 11342 29374 11394 29426
rect 15710 29374 15762 29426
rect 16382 29374 16434 29426
rect 17390 29374 17442 29426
rect 18062 29374 18114 29426
rect 18398 29374 18450 29426
rect 18622 29374 18674 29426
rect 18958 29374 19010 29426
rect 19294 29374 19346 29426
rect 19518 29374 19570 29426
rect 19966 29374 20018 29426
rect 21422 29374 21474 29426
rect 22430 29374 22482 29426
rect 22654 29374 22706 29426
rect 29150 29374 29202 29426
rect 29598 29374 29650 29426
rect 31390 29374 31442 29426
rect 32398 29374 32450 29426
rect 33070 29374 33122 29426
rect 33630 29374 33682 29426
rect 33854 29374 33906 29426
rect 34750 29374 34802 29426
rect 34862 29374 34914 29426
rect 34974 29374 35026 29426
rect 35646 29374 35698 29426
rect 36206 29374 36258 29426
rect 38670 29374 38722 29426
rect 39118 29374 39170 29426
rect 40910 29374 40962 29426
rect 41694 29374 41746 29426
rect 43038 29374 43090 29426
rect 43710 29374 43762 29426
rect 44270 29374 44322 29426
rect 44942 29374 44994 29426
rect 4734 29262 4786 29314
rect 7422 29262 7474 29314
rect 8542 29262 8594 29314
rect 13134 29262 13186 29314
rect 16718 29262 16770 29314
rect 17502 29262 17554 29314
rect 18510 29262 18562 29314
rect 19406 29262 19458 29314
rect 20638 29262 20690 29314
rect 21086 29262 21138 29314
rect 21646 29262 21698 29314
rect 28814 29262 28866 29314
rect 35198 29262 35250 29314
rect 36878 29262 36930 29314
rect 42926 29262 42978 29314
rect 8318 29150 8370 29202
rect 14478 29150 14530 29202
rect 33294 29150 33346 29202
rect 38446 29150 38498 29202
rect 44606 29150 44658 29202
rect 45390 29150 45442 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 8766 28814 8818 28866
rect 9102 28814 9154 28866
rect 15262 28814 15314 28866
rect 18174 28814 18226 28866
rect 21758 28814 21810 28866
rect 29486 28814 29538 28866
rect 30046 28814 30098 28866
rect 4174 28702 4226 28754
rect 4958 28702 5010 28754
rect 8430 28702 8482 28754
rect 10782 28702 10834 28754
rect 14142 28702 14194 28754
rect 15710 28702 15762 28754
rect 16382 28702 16434 28754
rect 18734 28702 18786 28754
rect 20190 28702 20242 28754
rect 21982 28702 22034 28754
rect 26798 28702 26850 28754
rect 29710 28702 29762 28754
rect 32286 28702 32338 28754
rect 39230 28702 39282 28754
rect 39678 28702 39730 28754
rect 43598 28702 43650 28754
rect 44158 28702 44210 28754
rect 44942 28702 44994 28754
rect 57934 28702 57986 28754
rect 4286 28590 4338 28642
rect 6974 28590 7026 28642
rect 7870 28590 7922 28642
rect 8766 28590 8818 28642
rect 10558 28590 10610 28642
rect 11230 28590 11282 28642
rect 12574 28590 12626 28642
rect 12798 28590 12850 28642
rect 13918 28590 13970 28642
rect 14366 28590 14418 28642
rect 14926 28590 14978 28642
rect 17726 28590 17778 28642
rect 20414 28590 20466 28642
rect 20750 28590 20802 28642
rect 22878 28590 22930 28642
rect 23998 28590 24050 28642
rect 27022 28590 27074 28642
rect 30382 28590 30434 28642
rect 30830 28590 30882 28642
rect 31054 28590 31106 28642
rect 32734 28590 32786 28642
rect 35310 28590 35362 28642
rect 37102 28590 37154 28642
rect 37662 28590 37714 28642
rect 38110 28590 38162 28642
rect 38894 28590 38946 28642
rect 55246 28590 55298 28642
rect 55582 28590 55634 28642
rect 6526 28478 6578 28530
rect 12014 28478 12066 28530
rect 12126 28478 12178 28530
rect 12350 28478 12402 28530
rect 12910 28478 12962 28530
rect 13582 28478 13634 28530
rect 17502 28478 17554 28530
rect 18062 28478 18114 28530
rect 20638 28478 20690 28530
rect 22542 28478 22594 28530
rect 24670 28478 24722 28530
rect 27246 28478 27298 28530
rect 27358 28478 27410 28530
rect 27806 28478 27858 28530
rect 30718 28478 30770 28530
rect 34526 28478 34578 28530
rect 35534 28478 35586 28530
rect 36094 28478 36146 28530
rect 36206 28478 36258 28530
rect 39006 28478 39058 28530
rect 11790 28366 11842 28418
rect 15150 28366 15202 28418
rect 16942 28366 16994 28418
rect 17278 28366 17330 28418
rect 17614 28366 17666 28418
rect 18174 28366 18226 28418
rect 21422 28366 21474 28418
rect 22318 28366 22370 28418
rect 22430 28366 22482 28418
rect 29150 28366 29202 28418
rect 30158 28366 30210 28418
rect 34302 28366 34354 28418
rect 34414 28366 34466 28418
rect 34750 28366 34802 28418
rect 36430 28366 36482 28418
rect 38446 28366 38498 28418
rect 38670 28366 38722 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 50558 28198 50610 28250
rect 50662 28198 50714 28250
rect 50766 28198 50818 28250
rect 7422 28030 7474 28082
rect 10894 28030 10946 28082
rect 16270 28030 16322 28082
rect 17502 28030 17554 28082
rect 20750 28030 20802 28082
rect 21422 28030 21474 28082
rect 25342 28030 25394 28082
rect 25454 28030 25506 28082
rect 25678 28030 25730 28082
rect 27246 28030 27298 28082
rect 30942 28030 30994 28082
rect 33182 28030 33234 28082
rect 33294 28030 33346 28082
rect 34078 28030 34130 28082
rect 38110 28030 38162 28082
rect 38334 28030 38386 28082
rect 38446 28030 38498 28082
rect 41022 28030 41074 28082
rect 43038 28030 43090 28082
rect 43262 28030 43314 28082
rect 45502 28030 45554 28082
rect 46062 28030 46114 28082
rect 12574 27918 12626 27970
rect 13918 27918 13970 27970
rect 15822 27918 15874 27970
rect 18062 27918 18114 27970
rect 18958 27918 19010 27970
rect 21646 27918 21698 27970
rect 29934 27918 29986 27970
rect 33070 27918 33122 27970
rect 33854 27918 33906 27970
rect 34190 27918 34242 27970
rect 35534 27918 35586 27970
rect 38670 27918 38722 27970
rect 38782 27918 38834 27970
rect 39230 27918 39282 27970
rect 39678 27918 39730 27970
rect 40798 27918 40850 27970
rect 44270 27918 44322 27970
rect 44718 27918 44770 27970
rect 44830 27918 44882 27970
rect 57822 27918 57874 27970
rect 6862 27806 6914 27858
rect 7086 27806 7138 27858
rect 8094 27806 8146 27858
rect 8990 27806 9042 27858
rect 10334 27806 10386 27858
rect 10558 27806 10610 27858
rect 12798 27806 12850 27858
rect 14926 27806 14978 27858
rect 15598 27806 15650 27858
rect 17950 27806 18002 27858
rect 18510 27806 18562 27858
rect 18734 27806 18786 27858
rect 18846 27806 18898 27858
rect 19406 27806 19458 27858
rect 22542 27806 22594 27858
rect 25230 27806 25282 27858
rect 28366 27806 28418 27858
rect 28926 27806 28978 27858
rect 30158 27806 30210 27858
rect 30606 27806 30658 27858
rect 33742 27806 33794 27858
rect 34750 27806 34802 27858
rect 37998 27806 38050 27858
rect 39566 27806 39618 27858
rect 39902 27806 39954 27858
rect 41134 27806 41186 27858
rect 42702 27806 42754 27858
rect 42926 27806 42978 27858
rect 43822 27806 43874 27858
rect 44046 27806 44098 27858
rect 45054 27806 45106 27858
rect 58158 27806 58210 27858
rect 8430 27694 8482 27746
rect 14142 27694 14194 27746
rect 18286 27694 18338 27746
rect 20638 27694 20690 27746
rect 21534 27694 21586 27746
rect 22318 27694 22370 27746
rect 31502 27694 31554 27746
rect 37662 27694 37714 27746
rect 41582 27694 41634 27746
rect 44382 27694 44434 27746
rect 57598 27694 57650 27746
rect 20974 27582 21026 27634
rect 22990 27582 23042 27634
rect 43374 27582 43426 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 16270 27246 16322 27298
rect 43598 27246 43650 27298
rect 43822 27246 43874 27298
rect 43934 27246 43986 27298
rect 1934 27134 1986 27186
rect 13918 27134 13970 27186
rect 14254 27134 14306 27186
rect 16606 27134 16658 27186
rect 17950 27134 18002 27186
rect 21534 27134 21586 27186
rect 27134 27134 27186 27186
rect 28030 27134 28082 27186
rect 29262 27134 29314 27186
rect 30158 27134 30210 27186
rect 32398 27134 32450 27186
rect 34526 27134 34578 27186
rect 40014 27134 40066 27186
rect 42142 27134 42194 27186
rect 45950 27134 46002 27186
rect 46510 27134 46562 27186
rect 47070 27134 47122 27186
rect 47518 27134 47570 27186
rect 57934 27134 57986 27186
rect 4286 27022 4338 27074
rect 14702 27022 14754 27074
rect 15150 27022 15202 27074
rect 17054 27022 17106 27074
rect 18174 27022 18226 27074
rect 18622 27022 18674 27074
rect 19294 27022 19346 27074
rect 19854 27022 19906 27074
rect 20190 27022 20242 27074
rect 20750 27022 20802 27074
rect 21870 27022 21922 27074
rect 24222 27022 24274 27074
rect 28590 27022 28642 27074
rect 29598 27022 29650 27074
rect 30494 27022 30546 27074
rect 31054 27022 31106 27074
rect 31614 27022 31666 27074
rect 39230 27022 39282 27074
rect 45502 27022 45554 27074
rect 45726 27022 45778 27074
rect 55582 27022 55634 27074
rect 12014 26910 12066 26962
rect 12350 26910 12402 26962
rect 14478 26910 14530 26962
rect 16494 26910 16546 26962
rect 12238 26798 12290 26850
rect 17166 26854 17218 26906
rect 17390 26910 17442 26962
rect 17614 26910 17666 26962
rect 21646 26910 21698 26962
rect 22878 26910 22930 26962
rect 23102 26910 23154 26962
rect 23214 26910 23266 26962
rect 23774 26910 23826 26962
rect 25006 26910 25058 26962
rect 27358 26910 27410 26962
rect 27582 26910 27634 26962
rect 37438 26910 37490 26962
rect 42590 26910 42642 26962
rect 23438 26798 23490 26850
rect 27694 26854 27746 26906
rect 35086 26798 35138 26850
rect 37774 26798 37826 26850
rect 38222 26798 38274 26850
rect 43038 26798 43090 26850
rect 43934 26798 43986 26850
rect 44718 26798 44770 26850
rect 46398 26798 46450 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 50558 26630 50610 26682
rect 50662 26630 50714 26682
rect 50766 26630 50818 26682
rect 23774 26462 23826 26514
rect 28926 26462 28978 26514
rect 29150 26462 29202 26514
rect 34862 26462 34914 26514
rect 37102 26462 37154 26514
rect 38446 26462 38498 26514
rect 44942 26462 44994 26514
rect 49086 26462 49138 26514
rect 57598 26462 57650 26514
rect 11678 26350 11730 26402
rect 16270 26350 16322 26402
rect 16830 26350 16882 26402
rect 17726 26350 17778 26402
rect 27918 26350 27970 26402
rect 28366 26350 28418 26402
rect 28590 26350 28642 26402
rect 29262 26350 29314 26402
rect 29486 26350 29538 26402
rect 30382 26350 30434 26402
rect 31054 26350 31106 26402
rect 40126 26350 40178 26402
rect 44382 26350 44434 26402
rect 57822 26350 57874 26402
rect 58158 26350 58210 26402
rect 4286 26238 4338 26290
rect 12462 26238 12514 26290
rect 15710 26238 15762 26290
rect 16046 26238 16098 26290
rect 16382 26238 16434 26290
rect 18286 26238 18338 26290
rect 18622 26238 18674 26290
rect 19742 26238 19794 26290
rect 19966 26238 20018 26290
rect 23102 26238 23154 26290
rect 23550 26238 23602 26290
rect 24110 26238 24162 26290
rect 26126 26238 26178 26290
rect 26350 26238 26402 26290
rect 26686 26238 26738 26290
rect 27694 26238 27746 26290
rect 28254 26238 28306 26290
rect 30718 26238 30770 26290
rect 31166 26238 31218 26290
rect 32062 26238 32114 26290
rect 34638 26238 34690 26290
rect 35198 26238 35250 26290
rect 39006 26238 39058 26290
rect 39566 26238 39618 26290
rect 39902 26238 39954 26290
rect 41022 26238 41074 26290
rect 44158 26238 44210 26290
rect 44494 26238 44546 26290
rect 45390 26238 45442 26290
rect 48862 26238 48914 26290
rect 1934 26126 1986 26178
rect 9550 26126 9602 26178
rect 12910 26126 12962 26178
rect 15038 26126 15090 26178
rect 18734 26126 18786 26178
rect 20302 26126 20354 26178
rect 22430 26126 22482 26178
rect 23662 26126 23714 26178
rect 29710 26126 29762 26178
rect 30270 26126 30322 26178
rect 33406 26126 33458 26178
rect 34750 26126 34802 26178
rect 36766 26126 36818 26178
rect 39790 26126 39842 26178
rect 41694 26126 41746 26178
rect 43822 26126 43874 26178
rect 46062 26126 46114 26178
rect 48190 26126 48242 26178
rect 25678 26014 25730 26066
rect 32958 26014 33010 26066
rect 33406 26014 33458 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 12126 25678 12178 25730
rect 13582 25678 13634 25730
rect 37102 25678 37154 25730
rect 42030 25678 42082 25730
rect 1934 25566 1986 25618
rect 8654 25566 8706 25618
rect 14142 25566 14194 25618
rect 17390 25566 17442 25618
rect 19630 25566 19682 25618
rect 21870 25566 21922 25618
rect 27918 25566 27970 25618
rect 30046 25566 30098 25618
rect 30494 25566 30546 25618
rect 31390 25566 31442 25618
rect 31950 25566 32002 25618
rect 34302 25566 34354 25618
rect 36430 25566 36482 25618
rect 40798 25566 40850 25618
rect 41470 25566 41522 25618
rect 45054 25566 45106 25618
rect 45502 25566 45554 25618
rect 57934 25566 57986 25618
rect 4286 25454 4338 25506
rect 11566 25454 11618 25506
rect 12798 25454 12850 25506
rect 13694 25454 13746 25506
rect 14926 25454 14978 25506
rect 15262 25454 15314 25506
rect 17278 25454 17330 25506
rect 18286 25454 18338 25506
rect 18622 25454 18674 25506
rect 18734 25454 18786 25506
rect 19742 25454 19794 25506
rect 26574 25454 26626 25506
rect 29374 25454 29426 25506
rect 32510 25454 32562 25506
rect 32958 25454 33010 25506
rect 33630 25454 33682 25506
rect 38110 25454 38162 25506
rect 39006 25454 39058 25506
rect 40014 25454 40066 25506
rect 40350 25454 40402 25506
rect 41358 25454 41410 25506
rect 41918 25454 41970 25506
rect 42366 25454 42418 25506
rect 42702 25454 42754 25506
rect 44270 25454 44322 25506
rect 46286 25454 46338 25506
rect 55582 25454 55634 25506
rect 10782 25342 10834 25394
rect 12238 25342 12290 25394
rect 12462 25342 12514 25394
rect 12686 25342 12738 25394
rect 13582 25342 13634 25394
rect 17166 25342 17218 25394
rect 20078 25342 20130 25394
rect 20190 25342 20242 25394
rect 28254 25342 28306 25394
rect 32734 25342 32786 25394
rect 37102 25342 37154 25394
rect 38782 25342 38834 25394
rect 39454 25342 39506 25394
rect 12126 25230 12178 25282
rect 15150 25230 15202 25282
rect 16606 25230 16658 25282
rect 20414 25230 20466 25282
rect 26574 25230 26626 25282
rect 26798 25230 26850 25282
rect 27022 25230 27074 25282
rect 28590 25230 28642 25282
rect 29150 25230 29202 25282
rect 30942 25230 30994 25282
rect 31838 25230 31890 25282
rect 32062 25230 32114 25282
rect 37214 25286 37266 25338
rect 39790 25342 39842 25394
rect 41582 25342 41634 25394
rect 42030 25342 42082 25394
rect 42590 25342 42642 25394
rect 43038 25342 43090 25394
rect 43374 25342 43426 25394
rect 44158 25342 44210 25394
rect 45838 25342 45890 25394
rect 37774 25230 37826 25282
rect 40238 25230 40290 25282
rect 41134 25230 41186 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 50558 25062 50610 25114
rect 50662 25062 50714 25114
rect 50766 25062 50818 25114
rect 4734 24894 4786 24946
rect 13134 24894 13186 24946
rect 23214 24894 23266 24946
rect 23326 24894 23378 24946
rect 24222 24894 24274 24946
rect 24446 24894 24498 24946
rect 24558 24894 24610 24946
rect 25902 24894 25954 24946
rect 26014 24894 26066 24946
rect 30046 24894 30098 24946
rect 33182 24894 33234 24946
rect 33518 24894 33570 24946
rect 38894 24894 38946 24946
rect 41358 24894 41410 24946
rect 41582 24894 41634 24946
rect 44270 24894 44322 24946
rect 47854 24894 47906 24946
rect 18846 24782 18898 24834
rect 18958 24782 19010 24834
rect 20302 24782 20354 24834
rect 20526 24782 20578 24834
rect 20638 24782 20690 24834
rect 21086 24782 21138 24834
rect 22654 24782 22706 24834
rect 22766 24782 22818 24834
rect 26910 24782 26962 24834
rect 28030 24782 28082 24834
rect 28814 24782 28866 24834
rect 31726 24782 31778 24834
rect 32062 24782 32114 24834
rect 37550 24782 37602 24834
rect 39230 24782 39282 24834
rect 41806 24782 41858 24834
rect 43934 24782 43986 24834
rect 46398 24782 46450 24834
rect 47518 24782 47570 24834
rect 4286 24670 4338 24722
rect 11902 24670 11954 24722
rect 14590 24670 14642 24722
rect 15262 24670 15314 24722
rect 15710 24670 15762 24722
rect 18622 24670 18674 24722
rect 19294 24670 19346 24722
rect 19854 24670 19906 24722
rect 21534 24670 21586 24722
rect 22990 24670 23042 24722
rect 23438 24670 23490 24722
rect 23774 24670 23826 24722
rect 24670 24670 24722 24722
rect 25790 24670 25842 24722
rect 26462 24670 26514 24722
rect 27134 24670 27186 24722
rect 27358 24670 27410 24722
rect 27918 24670 27970 24722
rect 28590 24670 28642 24722
rect 29486 24670 29538 24722
rect 30718 24670 30770 24722
rect 31278 24670 31330 24722
rect 31838 24670 31890 24722
rect 32398 24670 32450 24722
rect 33070 24670 33122 24722
rect 33294 24670 33346 24722
rect 34190 24670 34242 24722
rect 37662 24670 37714 24722
rect 40910 24670 40962 24722
rect 41134 24670 41186 24722
rect 41918 24670 41970 24722
rect 44494 24670 44546 24722
rect 46510 24670 46562 24722
rect 46958 24670 47010 24722
rect 53454 24670 53506 24722
rect 1934 24558 1986 24610
rect 5294 24558 5346 24610
rect 10334 24558 10386 24610
rect 12126 24558 12178 24610
rect 12574 24558 12626 24610
rect 14366 24558 14418 24610
rect 25342 24558 25394 24610
rect 34974 24558 35026 24610
rect 37102 24558 37154 24610
rect 38110 24558 38162 24610
rect 40462 24558 40514 24610
rect 42366 24558 42418 24610
rect 10558 24446 10610 24498
rect 10894 24446 10946 24498
rect 15598 24446 15650 24498
rect 27246 24446 27298 24498
rect 37550 24446 37602 24498
rect 41470 24446 41522 24498
rect 42254 24446 42306 24498
rect 55358 24446 55410 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 1934 24110 1986 24162
rect 29710 24110 29762 24162
rect 45726 24110 45778 24162
rect 57934 24110 57986 24162
rect 4958 23998 5010 24050
rect 10110 23998 10162 24050
rect 15262 23998 15314 24050
rect 16718 23998 16770 24050
rect 18510 23998 18562 24050
rect 20638 23998 20690 24050
rect 21310 23998 21362 24050
rect 23438 23998 23490 24050
rect 33406 23998 33458 24050
rect 33854 23998 33906 24050
rect 35646 23998 35698 24050
rect 46846 23998 46898 24050
rect 47294 23998 47346 24050
rect 55358 23998 55410 24050
rect 4286 23886 4338 23938
rect 6414 23886 6466 23938
rect 7870 23886 7922 23938
rect 8318 23886 8370 23938
rect 9998 23886 10050 23938
rect 14030 23886 14082 23938
rect 15150 23886 15202 23938
rect 16830 23886 16882 23938
rect 17838 23886 17890 23938
rect 24110 23886 24162 23938
rect 24446 23886 24498 23938
rect 24782 23886 24834 23938
rect 25118 23886 25170 23938
rect 25454 23886 25506 23938
rect 26350 23886 26402 23938
rect 27246 23886 27298 23938
rect 27806 23886 27858 23938
rect 29150 23886 29202 23938
rect 30046 23886 30098 23938
rect 31614 23886 31666 23938
rect 32174 23886 32226 23938
rect 33070 23886 33122 23938
rect 33742 23886 33794 23938
rect 33966 23886 34018 23938
rect 34526 23886 34578 23938
rect 35086 23886 35138 23938
rect 35534 23886 35586 23938
rect 35758 23886 35810 23938
rect 36206 23886 36258 23938
rect 38558 23886 38610 23938
rect 40238 23886 40290 23938
rect 45166 23886 45218 23938
rect 45614 23886 45666 23938
rect 55582 23886 55634 23938
rect 4622 23774 4674 23826
rect 5630 23774 5682 23826
rect 6638 23774 6690 23826
rect 6750 23774 6802 23826
rect 8542 23774 8594 23826
rect 10670 23774 10722 23826
rect 11006 23774 11058 23826
rect 14254 23774 14306 23826
rect 14366 23774 14418 23826
rect 24670 23774 24722 23826
rect 25678 23774 25730 23826
rect 26126 23774 26178 23826
rect 27022 23774 27074 23826
rect 32622 23774 32674 23826
rect 32958 23774 33010 23826
rect 34190 23774 34242 23826
rect 34974 23774 35026 23826
rect 41246 23774 41298 23826
rect 44942 23774 44994 23826
rect 46398 23774 46450 23826
rect 46622 23774 46674 23826
rect 46958 23774 47010 23826
rect 4846 23662 4898 23714
rect 5070 23662 5122 23714
rect 5742 23662 5794 23714
rect 5966 23662 6018 23714
rect 7198 23662 7250 23714
rect 11118 23662 11170 23714
rect 25342 23662 25394 23714
rect 28366 23662 28418 23714
rect 29374 23662 29426 23714
rect 29598 23662 29650 23714
rect 30270 23662 30322 23714
rect 30830 23662 30882 23714
rect 35198 23662 35250 23714
rect 45726 23662 45778 23714
rect 47406 23662 47458 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 50558 23494 50610 23546
rect 50662 23494 50714 23546
rect 50766 23494 50818 23546
rect 13806 23326 13858 23378
rect 24222 23326 24274 23378
rect 24782 23326 24834 23378
rect 25230 23326 25282 23378
rect 25566 23326 25618 23378
rect 31614 23326 31666 23378
rect 37662 23326 37714 23378
rect 38558 23326 38610 23378
rect 6974 23214 7026 23266
rect 7870 23214 7922 23266
rect 12014 23214 12066 23266
rect 16158 23214 16210 23266
rect 18062 23214 18114 23266
rect 21646 23214 21698 23266
rect 24446 23214 24498 23266
rect 24558 23214 24610 23266
rect 29822 23214 29874 23266
rect 31950 23214 32002 23266
rect 32398 23214 32450 23266
rect 42030 23214 42082 23266
rect 45390 23214 45442 23266
rect 4286 23102 4338 23154
rect 5182 23102 5234 23154
rect 6190 23102 6242 23154
rect 8318 23102 8370 23154
rect 8990 23102 9042 23154
rect 10782 23102 10834 23154
rect 11790 23102 11842 23154
rect 13470 23102 13522 23154
rect 14254 23102 14306 23154
rect 15262 23102 15314 23154
rect 15486 23102 15538 23154
rect 17950 23102 18002 23154
rect 18286 23102 18338 23154
rect 19182 23102 19234 23154
rect 21534 23102 21586 23154
rect 22430 23102 22482 23154
rect 22766 23102 22818 23154
rect 22990 23102 23042 23154
rect 26798 23102 26850 23154
rect 37886 23102 37938 23154
rect 38334 23102 38386 23154
rect 38670 23102 38722 23154
rect 39006 23102 39058 23154
rect 39454 23102 39506 23154
rect 39790 23102 39842 23154
rect 41246 23102 41298 23154
rect 44606 23102 44658 23154
rect 47966 23102 48018 23154
rect 53454 23102 53506 23154
rect 1934 22990 1986 23042
rect 4734 22990 4786 23042
rect 8542 22990 8594 23042
rect 11006 22990 11058 23042
rect 18510 22990 18562 23042
rect 22206 22990 22258 23042
rect 22654 22990 22706 23042
rect 23662 22990 23714 23042
rect 39678 22990 39730 23042
rect 44158 22990 44210 23042
rect 47518 22990 47570 23042
rect 11118 22878 11170 22930
rect 14254 22878 14306 22930
rect 14590 22878 14642 22930
rect 18622 22878 18674 22930
rect 19294 22878 19346 22930
rect 38110 22878 38162 22930
rect 39230 22878 39282 22930
rect 55358 22878 55410 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 3054 22542 3106 22594
rect 3390 22542 3442 22594
rect 8990 22542 9042 22594
rect 12014 22542 12066 22594
rect 22094 22542 22146 22594
rect 37102 22542 37154 22594
rect 37550 22542 37602 22594
rect 38334 22542 38386 22594
rect 39790 22542 39842 22594
rect 57934 22542 57986 22594
rect 4510 22430 4562 22482
rect 4846 22430 4898 22482
rect 5966 22430 6018 22482
rect 8094 22430 8146 22482
rect 9886 22430 9938 22482
rect 12126 22430 12178 22482
rect 13582 22430 13634 22482
rect 15262 22430 15314 22482
rect 15710 22430 15762 22482
rect 16606 22430 16658 22482
rect 19070 22430 19122 22482
rect 24894 22430 24946 22482
rect 25678 22430 25730 22482
rect 29374 22430 29426 22482
rect 33518 22430 33570 22482
rect 36990 22430 37042 22482
rect 42590 22430 42642 22482
rect 43038 22430 43090 22482
rect 47630 22430 47682 22482
rect 49758 22430 49810 22482
rect 55022 22430 55074 22482
rect 2270 22318 2322 22370
rect 2830 22318 2882 22370
rect 4062 22318 4114 22370
rect 4958 22318 5010 22370
rect 7422 22318 7474 22370
rect 8430 22318 8482 22370
rect 8654 22318 8706 22370
rect 8878 22318 8930 22370
rect 11342 22318 11394 22370
rect 11566 22318 11618 22370
rect 12574 22318 12626 22370
rect 14030 22318 14082 22370
rect 14478 22318 14530 22370
rect 15934 22318 15986 22370
rect 18174 22318 18226 22370
rect 18398 22318 18450 22370
rect 21422 22318 21474 22370
rect 21646 22318 21698 22370
rect 23102 22318 23154 22370
rect 23438 22318 23490 22370
rect 24110 22318 24162 22370
rect 26798 22318 26850 22370
rect 27246 22318 27298 22370
rect 28254 22318 28306 22370
rect 29598 22318 29650 22370
rect 35422 22318 35474 22370
rect 37214 22318 37266 22370
rect 37774 22318 37826 22370
rect 39230 22318 39282 22370
rect 39566 22318 39618 22370
rect 40238 22318 40290 22370
rect 40910 22318 40962 22370
rect 42142 22318 42194 22370
rect 42478 22318 42530 22370
rect 42702 22318 42754 22370
rect 44046 22318 44098 22370
rect 46062 22318 46114 22370
rect 46398 22318 46450 22370
rect 46846 22318 46898 22370
rect 52670 22318 52722 22370
rect 55582 22318 55634 22370
rect 2494 22206 2546 22258
rect 6526 22206 6578 22258
rect 9550 22206 9602 22258
rect 11006 22206 11058 22258
rect 14926 22206 14978 22258
rect 17726 22206 17778 22258
rect 25342 22206 25394 22258
rect 25790 22206 25842 22258
rect 26462 22206 26514 22258
rect 27470 22206 27522 22258
rect 35982 22206 36034 22258
rect 36094 22206 36146 22258
rect 38222 22206 38274 22258
rect 38894 22206 38946 22258
rect 40350 22206 40402 22258
rect 40574 22206 40626 22258
rect 41246 22206 41298 22258
rect 41470 22206 41522 22258
rect 41806 22206 41858 22258
rect 45166 22206 45218 22258
rect 45502 22206 45554 22258
rect 46286 22206 46338 22258
rect 9774 22094 9826 22146
rect 11118 22094 11170 22146
rect 15150 22094 15202 22146
rect 17390 22094 17442 22146
rect 17614 22094 17666 22146
rect 25566 22094 25618 22146
rect 28702 22094 28754 22146
rect 35198 22094 35250 22146
rect 35758 22094 35810 22146
rect 38334 22094 38386 22146
rect 39006 22094 39058 22146
rect 39454 22094 39506 22146
rect 40798 22094 40850 22146
rect 41694 22094 41746 22146
rect 43598 22094 43650 22146
rect 44270 22094 44322 22146
rect 44830 22094 44882 22146
rect 45838 22094 45890 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 50558 21926 50610 21978
rect 50662 21926 50714 21978
rect 50766 21926 50818 21978
rect 3950 21758 4002 21810
rect 4734 21758 4786 21810
rect 5070 21758 5122 21810
rect 8094 21758 8146 21810
rect 10222 21758 10274 21810
rect 22542 21758 22594 21810
rect 23886 21758 23938 21810
rect 24334 21758 24386 21810
rect 40014 21758 40066 21810
rect 2270 21646 2322 21698
rect 4062 21646 4114 21698
rect 7198 21646 7250 21698
rect 11230 21646 11282 21698
rect 13582 21646 13634 21698
rect 14590 21646 14642 21698
rect 16494 21646 16546 21698
rect 19518 21646 19570 21698
rect 20750 21646 20802 21698
rect 22430 21646 22482 21698
rect 23102 21646 23154 21698
rect 32062 21646 32114 21698
rect 32510 21646 32562 21698
rect 37102 21646 37154 21698
rect 39678 21646 39730 21698
rect 2718 21534 2770 21586
rect 3166 21534 3218 21586
rect 3614 21534 3666 21586
rect 4286 21534 4338 21586
rect 4622 21534 4674 21586
rect 4846 21534 4898 21586
rect 7086 21534 7138 21586
rect 7982 21534 8034 21586
rect 9886 21534 9938 21586
rect 10334 21534 10386 21586
rect 12350 21534 12402 21586
rect 14702 21534 14754 21586
rect 15150 21534 15202 21586
rect 15598 21534 15650 21586
rect 15822 21534 15874 21586
rect 17614 21534 17666 21586
rect 19182 21534 19234 21586
rect 21310 21534 21362 21586
rect 25342 21534 25394 21586
rect 28814 21534 28866 21586
rect 33070 21534 33122 21586
rect 36318 21534 36370 21586
rect 40238 21534 40290 21586
rect 40910 21534 40962 21586
rect 53454 21534 53506 21586
rect 2942 21422 2994 21474
rect 12462 21422 12514 21474
rect 17726 21422 17778 21474
rect 23214 21422 23266 21474
rect 24670 21422 24722 21474
rect 26014 21422 26066 21474
rect 28142 21422 28194 21474
rect 29486 21422 29538 21474
rect 31614 21422 31666 21474
rect 33854 21422 33906 21474
rect 35982 21422 36034 21474
rect 39230 21422 39282 21474
rect 43710 21422 43762 21474
rect 46622 21422 46674 21474
rect 10110 21310 10162 21362
rect 11006 21310 11058 21362
rect 11342 21310 11394 21362
rect 14926 21310 14978 21362
rect 23326 21310 23378 21362
rect 55358 21310 55410 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 3390 20974 3442 21026
rect 4958 20974 5010 21026
rect 12350 20974 12402 21026
rect 16158 20974 16210 21026
rect 17502 20974 17554 21026
rect 19182 20974 19234 21026
rect 27022 20974 27074 21026
rect 28142 20974 28194 21026
rect 28478 20974 28530 21026
rect 30046 20974 30098 21026
rect 33518 20974 33570 21026
rect 34078 20974 34130 21026
rect 37550 20974 37602 21026
rect 43822 20974 43874 21026
rect 44158 20974 44210 21026
rect 57934 20974 57986 21026
rect 3166 20862 3218 20914
rect 6750 20862 6802 20914
rect 8766 20862 8818 20914
rect 12238 20862 12290 20914
rect 13806 20862 13858 20914
rect 14366 20862 14418 20914
rect 15262 20862 15314 20914
rect 32062 20862 32114 20914
rect 33854 20862 33906 20914
rect 35982 20862 36034 20914
rect 36990 20862 37042 20914
rect 38334 20862 38386 20914
rect 39566 20862 39618 20914
rect 41694 20862 41746 20914
rect 45278 20862 45330 20914
rect 45838 20862 45890 20914
rect 49758 20862 49810 20914
rect 3614 20750 3666 20802
rect 4062 20750 4114 20802
rect 4398 20750 4450 20802
rect 4622 20750 4674 20802
rect 6302 20750 6354 20802
rect 6638 20750 6690 20802
rect 7982 20750 8034 20802
rect 8878 20750 8930 20802
rect 9886 20750 9938 20802
rect 10110 20750 10162 20802
rect 10670 20750 10722 20802
rect 11118 20750 11170 20802
rect 11566 20750 11618 20802
rect 12462 20750 12514 20802
rect 13582 20750 13634 20802
rect 14590 20750 14642 20802
rect 15598 20750 15650 20802
rect 15822 20750 15874 20802
rect 16046 20750 16098 20802
rect 17166 20750 17218 20802
rect 17390 20750 17442 20802
rect 18510 20750 18562 20802
rect 22430 20750 22482 20802
rect 23998 20750 24050 20802
rect 26014 20750 26066 20802
rect 27246 20750 27298 20802
rect 29822 20750 29874 20802
rect 30382 20750 30434 20802
rect 33294 20750 33346 20802
rect 33966 20750 34018 20802
rect 34414 20750 34466 20802
rect 34862 20750 34914 20802
rect 35422 20750 35474 20802
rect 35758 20750 35810 20802
rect 37214 20750 37266 20802
rect 37886 20750 37938 20802
rect 38782 20750 38834 20802
rect 42590 20750 42642 20802
rect 43150 20750 43202 20802
rect 44830 20750 44882 20802
rect 46846 20750 46898 20802
rect 55582 20750 55634 20802
rect 10222 20638 10274 20690
rect 13918 20638 13970 20690
rect 16830 20638 16882 20690
rect 19070 20638 19122 20690
rect 21198 20638 21250 20690
rect 21422 20638 21474 20690
rect 21534 20638 21586 20690
rect 22206 20638 22258 20690
rect 24110 20638 24162 20690
rect 25454 20638 25506 20690
rect 27582 20638 27634 20690
rect 27806 20638 27858 20690
rect 29038 20638 29090 20690
rect 29374 20638 29426 20690
rect 30606 20638 30658 20690
rect 30830 20638 30882 20690
rect 31166 20638 31218 20690
rect 38110 20638 38162 20690
rect 38446 20638 38498 20690
rect 42030 20638 42082 20690
rect 43038 20638 43090 20690
rect 47630 20638 47682 20690
rect 55358 20638 55410 20690
rect 16942 20526 16994 20578
rect 17502 20526 17554 20578
rect 18734 20526 18786 20578
rect 19182 20526 19234 20578
rect 26910 20526 26962 20578
rect 28254 20526 28306 20578
rect 29262 20526 29314 20578
rect 29710 20526 29762 20578
rect 31054 20526 31106 20578
rect 31614 20526 31666 20578
rect 34638 20526 34690 20578
rect 34750 20526 34802 20578
rect 34974 20526 35026 20578
rect 36542 20526 36594 20578
rect 46510 20526 46562 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 50558 20358 50610 20410
rect 50662 20358 50714 20410
rect 50766 20358 50818 20410
rect 12462 20190 12514 20242
rect 14590 20190 14642 20242
rect 25902 20190 25954 20242
rect 40462 20190 40514 20242
rect 47630 20190 47682 20242
rect 5182 20078 5234 20130
rect 5406 20078 5458 20130
rect 6526 20078 6578 20130
rect 8206 20078 8258 20130
rect 11118 20078 11170 20130
rect 14254 20078 14306 20130
rect 14478 20078 14530 20130
rect 15262 20078 15314 20130
rect 15374 20078 15426 20130
rect 17502 20078 17554 20130
rect 20414 20078 20466 20130
rect 22542 20078 22594 20130
rect 24558 20078 24610 20130
rect 25678 20078 25730 20130
rect 26238 20078 26290 20130
rect 27694 20078 27746 20130
rect 28478 20078 28530 20130
rect 29710 20078 29762 20130
rect 31726 20078 31778 20130
rect 34302 20078 34354 20130
rect 39454 20078 39506 20130
rect 40910 20078 40962 20130
rect 42030 20078 42082 20130
rect 45838 20078 45890 20130
rect 47070 20078 47122 20130
rect 48974 20078 49026 20130
rect 2718 19966 2770 20018
rect 3950 19966 4002 20018
rect 4734 19966 4786 20018
rect 5518 19966 5570 20018
rect 7758 19966 7810 20018
rect 11342 19966 11394 20018
rect 12014 19966 12066 20018
rect 14702 19966 14754 20018
rect 14926 19966 14978 20018
rect 17614 19966 17666 20018
rect 20190 19966 20242 20018
rect 20526 19966 20578 20018
rect 21310 19966 21362 20018
rect 22766 19966 22818 20018
rect 23662 19966 23714 20018
rect 26014 19966 26066 20018
rect 27246 19966 27298 20018
rect 29038 19966 29090 20018
rect 29934 19966 29986 20018
rect 30382 19966 30434 20018
rect 30606 19966 30658 20018
rect 32062 19966 32114 20018
rect 33182 19966 33234 20018
rect 34190 19966 34242 20018
rect 35646 19966 35698 20018
rect 39902 19966 39954 20018
rect 41246 19966 41298 20018
rect 46510 19966 46562 20018
rect 47966 19966 48018 20018
rect 48862 19966 48914 20018
rect 49982 19966 50034 20018
rect 53678 19966 53730 20018
rect 2830 19854 2882 19906
rect 6414 19854 6466 19906
rect 7422 19854 7474 19906
rect 13246 19854 13298 19906
rect 15934 19854 15986 19906
rect 21534 19854 21586 19906
rect 23214 19854 23266 19906
rect 27022 19854 27074 19906
rect 28814 19854 28866 19906
rect 30494 19854 30546 19906
rect 35198 19854 35250 19906
rect 36318 19854 36370 19906
rect 38446 19854 38498 19906
rect 38894 19854 38946 19906
rect 42926 19854 42978 19906
rect 43710 19854 43762 19906
rect 6750 19742 6802 19794
rect 15374 19742 15426 19794
rect 17502 19742 17554 19794
rect 24110 19742 24162 19794
rect 33518 19742 33570 19794
rect 49646 19742 49698 19794
rect 55358 19742 55410 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 2494 19406 2546 19458
rect 6638 19406 6690 19458
rect 8318 19406 8370 19458
rect 8654 19406 8706 19458
rect 8990 19406 9042 19458
rect 12126 19406 12178 19458
rect 22766 19406 22818 19458
rect 25790 19406 25842 19458
rect 57934 19406 57986 19458
rect 3614 19294 3666 19346
rect 8990 19294 9042 19346
rect 19294 19294 19346 19346
rect 21310 19294 21362 19346
rect 23438 19294 23490 19346
rect 25454 19294 25506 19346
rect 29150 19294 29202 19346
rect 31278 19294 31330 19346
rect 33406 19294 33458 19346
rect 38782 19294 38834 19346
rect 40238 19294 40290 19346
rect 42366 19294 42418 19346
rect 42814 19294 42866 19346
rect 44270 19294 44322 19346
rect 47742 19294 47794 19346
rect 53230 19294 53282 19346
rect 2830 19182 2882 19234
rect 3054 19182 3106 19234
rect 3726 19182 3778 19234
rect 4174 19182 4226 19234
rect 4510 19182 4562 19234
rect 6974 19182 7026 19234
rect 7198 19182 7250 19234
rect 9662 19182 9714 19234
rect 10670 19182 10722 19234
rect 11342 19182 11394 19234
rect 11566 19182 11618 19234
rect 12574 19182 12626 19234
rect 16942 19182 16994 19234
rect 17502 19182 17554 19234
rect 18174 19182 18226 19234
rect 19406 19182 19458 19234
rect 19742 19182 19794 19234
rect 21422 19182 21474 19234
rect 21758 19182 21810 19234
rect 26126 19182 26178 19234
rect 27022 19182 27074 19234
rect 28142 19182 28194 19234
rect 28254 19182 28306 19234
rect 30494 19182 30546 19234
rect 37438 19182 37490 19234
rect 38222 19182 38274 19234
rect 39454 19182 39506 19234
rect 44830 19182 44882 19234
rect 55582 19182 55634 19234
rect 1710 19070 1762 19122
rect 3390 19070 3442 19122
rect 4398 19070 4450 19122
rect 5630 19070 5682 19122
rect 8430 19070 8482 19122
rect 9998 19070 10050 19122
rect 11678 19070 11730 19122
rect 12238 19070 12290 19122
rect 12686 19070 12738 19122
rect 16270 19070 16322 19122
rect 18734 19070 18786 19122
rect 22878 19070 22930 19122
rect 23550 19070 23602 19122
rect 25230 19070 25282 19122
rect 25902 19070 25954 19122
rect 27246 19070 27298 19122
rect 27694 19070 27746 19122
rect 28478 19070 28530 19122
rect 28590 19070 28642 19122
rect 29486 19070 29538 19122
rect 29598 19070 29650 19122
rect 29710 19070 29762 19122
rect 36094 19070 36146 19122
rect 36430 19070 36482 19122
rect 37102 19070 37154 19122
rect 37998 19070 38050 19122
rect 45614 19070 45666 19122
rect 52782 19070 52834 19122
rect 2046 18958 2098 19010
rect 5070 18958 5122 19010
rect 5966 18958 6018 19010
rect 7534 18958 7586 19010
rect 7870 18958 7922 19010
rect 8318 18958 8370 19010
rect 9886 18958 9938 19010
rect 12126 18958 12178 19010
rect 15934 18958 15986 19010
rect 22766 18958 22818 19010
rect 29934 18958 29986 19010
rect 52670 18958 52722 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 50558 18790 50610 18842
rect 50662 18790 50714 18842
rect 50766 18790 50818 18842
rect 1822 18622 1874 18674
rect 4846 18622 4898 18674
rect 7310 18622 7362 18674
rect 13470 18622 13522 18674
rect 14254 18622 14306 18674
rect 16942 18622 16994 18674
rect 18174 18622 18226 18674
rect 18622 18622 18674 18674
rect 18846 18622 18898 18674
rect 19182 18622 19234 18674
rect 19406 18622 19458 18674
rect 19966 18622 20018 18674
rect 23662 18622 23714 18674
rect 24446 18622 24498 18674
rect 30606 18622 30658 18674
rect 37886 18622 37938 18674
rect 45166 18622 45218 18674
rect 2942 18510 2994 18562
rect 4174 18510 4226 18562
rect 4958 18510 5010 18562
rect 5630 18510 5682 18562
rect 5742 18510 5794 18562
rect 6190 18510 6242 18562
rect 6750 18510 6802 18562
rect 7534 18510 7586 18562
rect 9998 18510 10050 18562
rect 10110 18510 10162 18562
rect 11790 18510 11842 18562
rect 13358 18510 13410 18562
rect 16718 18510 16770 18562
rect 17838 18510 17890 18562
rect 17950 18510 18002 18562
rect 18510 18510 18562 18562
rect 19518 18510 19570 18562
rect 19854 18510 19906 18562
rect 23774 18510 23826 18562
rect 27918 18510 27970 18562
rect 28030 18510 28082 18562
rect 41134 18510 41186 18562
rect 45726 18510 45778 18562
rect 48750 18510 48802 18562
rect 2718 18398 2770 18450
rect 3054 18398 3106 18450
rect 4062 18398 4114 18450
rect 6526 18398 6578 18450
rect 6862 18398 6914 18450
rect 7646 18398 7698 18450
rect 10558 18398 10610 18450
rect 11118 18398 11170 18450
rect 11454 18398 11506 18450
rect 13918 18398 13970 18450
rect 15150 18398 15202 18450
rect 15598 18398 15650 18450
rect 16606 18398 16658 18450
rect 20190 18398 20242 18450
rect 20750 18398 20802 18450
rect 21310 18398 21362 18450
rect 22094 18398 22146 18450
rect 24334 18398 24386 18450
rect 24670 18398 24722 18450
rect 27134 18398 27186 18450
rect 28254 18398 28306 18450
rect 28590 18398 28642 18450
rect 30270 18398 30322 18450
rect 37326 18398 37378 18450
rect 37774 18398 37826 18450
rect 37998 18398 38050 18450
rect 41358 18398 41410 18450
rect 42142 18398 42194 18450
rect 44942 18398 44994 18450
rect 45950 18398 46002 18450
rect 46734 18398 46786 18450
rect 49086 18398 49138 18450
rect 51662 18398 51714 18450
rect 52110 18398 52162 18450
rect 53454 18398 53506 18450
rect 2270 18286 2322 18338
rect 8094 18286 8146 18338
rect 12350 18286 12402 18338
rect 15262 18286 15314 18338
rect 22542 18286 22594 18338
rect 27358 18286 27410 18338
rect 27470 18286 27522 18338
rect 38558 18286 38610 18338
rect 39006 18286 39058 18338
rect 46398 18286 46450 18338
rect 51998 18286 52050 18338
rect 1710 18174 1762 18226
rect 2270 18174 2322 18226
rect 5630 18174 5682 18226
rect 10110 18174 10162 18226
rect 10782 18174 10834 18226
rect 13470 18174 13522 18226
rect 23550 18174 23602 18226
rect 41806 18174 41858 18226
rect 51550 18174 51602 18226
rect 55358 18174 55410 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 3726 17838 3778 17890
rect 15262 17838 15314 17890
rect 16270 17838 16322 17890
rect 26574 17838 26626 17890
rect 50766 17838 50818 17890
rect 51102 17838 51154 17890
rect 51214 17838 51266 17890
rect 57934 17838 57986 17890
rect 5854 17726 5906 17778
rect 7870 17726 7922 17778
rect 10782 17726 10834 17778
rect 13582 17726 13634 17778
rect 27918 17726 27970 17778
rect 31950 17726 32002 17778
rect 35310 17726 35362 17778
rect 35758 17726 35810 17778
rect 39230 17726 39282 17778
rect 46958 17726 47010 17778
rect 48078 17726 48130 17778
rect 50206 17726 50258 17778
rect 51662 17726 51714 17778
rect 55022 17726 55074 17778
rect 2270 17614 2322 17666
rect 2606 17614 2658 17666
rect 3390 17614 3442 17666
rect 4398 17614 4450 17666
rect 7310 17614 7362 17666
rect 8318 17614 8370 17666
rect 10334 17614 10386 17666
rect 11118 17614 11170 17666
rect 13022 17614 13074 17666
rect 13694 17614 13746 17666
rect 15038 17614 15090 17666
rect 18622 17614 18674 17666
rect 18846 17614 18898 17666
rect 19518 17614 19570 17666
rect 21870 17614 21922 17666
rect 23214 17614 23266 17666
rect 25118 17614 25170 17666
rect 27022 17614 27074 17666
rect 27246 17614 27298 17666
rect 30718 17614 30770 17666
rect 31390 17614 31442 17666
rect 34862 17614 34914 17666
rect 36318 17614 36370 17666
rect 37214 17614 37266 17666
rect 37662 17614 37714 17666
rect 38334 17614 38386 17666
rect 39454 17614 39506 17666
rect 39790 17614 39842 17666
rect 40126 17614 40178 17666
rect 40350 17614 40402 17666
rect 45278 17614 45330 17666
rect 45950 17614 46002 17666
rect 47294 17614 47346 17666
rect 50878 17614 50930 17666
rect 52222 17614 52274 17666
rect 52670 17614 52722 17666
rect 55582 17614 55634 17666
rect 4734 17502 4786 17554
rect 6190 17502 6242 17554
rect 9886 17502 9938 17554
rect 9998 17502 10050 17554
rect 11454 17502 11506 17554
rect 11678 17502 11730 17554
rect 11902 17502 11954 17554
rect 12014 17502 12066 17554
rect 12686 17502 12738 17554
rect 16382 17502 16434 17554
rect 20638 17502 20690 17554
rect 22094 17502 22146 17554
rect 24782 17502 24834 17554
rect 26462 17502 26514 17554
rect 29934 17502 29986 17554
rect 30382 17502 30434 17554
rect 31502 17502 31554 17554
rect 34078 17502 34130 17554
rect 37998 17502 38050 17554
rect 40574 17502 40626 17554
rect 43822 17502 43874 17554
rect 44942 17502 44994 17554
rect 45838 17502 45890 17554
rect 51550 17502 51602 17554
rect 8654 17390 8706 17442
rect 10222 17390 10274 17442
rect 10670 17390 10722 17442
rect 10894 17390 10946 17442
rect 11342 17390 11394 17442
rect 12798 17390 12850 17442
rect 16270 17390 16322 17442
rect 18286 17390 18338 17442
rect 25566 17390 25618 17442
rect 29598 17390 29650 17442
rect 36094 17390 36146 17442
rect 36990 17390 37042 17442
rect 38670 17390 38722 17442
rect 39118 17390 39170 17442
rect 39342 17390 39394 17442
rect 40686 17390 40738 17442
rect 40798 17390 40850 17442
rect 42142 17390 42194 17442
rect 43486 17390 43538 17442
rect 51774 17390 51826 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 50558 17222 50610 17274
rect 50662 17222 50714 17274
rect 50766 17222 50818 17274
rect 1710 17054 1762 17106
rect 2046 17054 2098 17106
rect 3950 17054 4002 17106
rect 5182 17054 5234 17106
rect 5854 17054 5906 17106
rect 6974 17054 7026 17106
rect 14702 17054 14754 17106
rect 26574 17054 26626 17106
rect 26798 17054 26850 17106
rect 33518 17054 33570 17106
rect 36430 17054 36482 17106
rect 36990 17054 37042 17106
rect 38110 17054 38162 17106
rect 39678 17054 39730 17106
rect 41806 17054 41858 17106
rect 45614 17054 45666 17106
rect 49982 17054 50034 17106
rect 3614 16942 3666 16994
rect 6078 16942 6130 16994
rect 8318 16942 8370 16994
rect 9774 16942 9826 16994
rect 10110 16942 10162 16994
rect 12014 16942 12066 16994
rect 15038 16942 15090 16994
rect 15374 16942 15426 16994
rect 17726 16942 17778 16994
rect 17838 16942 17890 16994
rect 18510 16942 18562 16994
rect 19070 16942 19122 16994
rect 20974 16942 21026 16994
rect 23214 16942 23266 16994
rect 24670 16942 24722 16994
rect 26014 16942 26066 16994
rect 29150 16942 29202 16994
rect 32062 16942 32114 16994
rect 35086 16942 35138 16994
rect 35758 16942 35810 16994
rect 43038 16942 43090 16994
rect 49086 16942 49138 16994
rect 50654 16942 50706 16994
rect 52222 16942 52274 16994
rect 2942 16830 2994 16882
rect 3390 16830 3442 16882
rect 4510 16830 4562 16882
rect 4958 16830 5010 16882
rect 5070 16830 5122 16882
rect 5518 16830 5570 16882
rect 6190 16830 6242 16882
rect 7310 16830 7362 16882
rect 7982 16830 8034 16882
rect 9102 16830 9154 16882
rect 9550 16830 9602 16882
rect 12238 16830 12290 16882
rect 14030 16830 14082 16882
rect 14366 16830 14418 16882
rect 18286 16830 18338 16882
rect 21982 16830 22034 16882
rect 23102 16830 23154 16882
rect 23998 16830 24050 16882
rect 26462 16830 26514 16882
rect 28478 16830 28530 16882
rect 33294 16830 33346 16882
rect 34078 16830 34130 16882
rect 35198 16830 35250 16882
rect 36206 16830 36258 16882
rect 36542 16830 36594 16882
rect 37438 16830 37490 16882
rect 39454 16830 39506 16882
rect 39902 16830 39954 16882
rect 40014 16830 40066 16882
rect 41358 16830 41410 16882
rect 41582 16830 41634 16882
rect 42254 16830 42306 16882
rect 48862 16830 48914 16882
rect 51326 16830 51378 16882
rect 51998 16830 52050 16882
rect 53566 16830 53618 16882
rect 7870 16718 7922 16770
rect 9998 16718 10050 16770
rect 16046 16718 16098 16770
rect 18174 16718 18226 16770
rect 23774 16718 23826 16770
rect 31278 16718 31330 16770
rect 34414 16718 34466 16770
rect 39790 16718 39842 16770
rect 41694 16718 41746 16770
rect 45166 16718 45218 16770
rect 16270 16606 16322 16658
rect 16494 16606 16546 16658
rect 16942 16606 16994 16658
rect 17726 16606 17778 16658
rect 25790 16606 25842 16658
rect 26126 16606 26178 16658
rect 31838 16606 31890 16658
rect 32174 16606 32226 16658
rect 40910 16606 40962 16658
rect 41134 16606 41186 16658
rect 49646 16606 49698 16658
rect 55358 16606 55410 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 7982 16270 8034 16322
rect 9550 16270 9602 16322
rect 9886 16270 9938 16322
rect 15710 16270 15762 16322
rect 16270 16270 16322 16322
rect 17614 16270 17666 16322
rect 20638 16270 20690 16322
rect 26910 16270 26962 16322
rect 31614 16270 31666 16322
rect 32510 16270 32562 16322
rect 40798 16270 40850 16322
rect 51998 16270 52050 16322
rect 52782 16270 52834 16322
rect 57934 16270 57986 16322
rect 2830 16158 2882 16210
rect 6750 16158 6802 16210
rect 10446 16158 10498 16210
rect 14814 16158 14866 16210
rect 16830 16158 16882 16210
rect 26238 16158 26290 16210
rect 30158 16158 30210 16210
rect 31166 16158 31218 16210
rect 32958 16158 33010 16210
rect 34190 16158 34242 16210
rect 34526 16158 34578 16210
rect 35198 16158 35250 16210
rect 41358 16158 41410 16210
rect 42590 16158 42642 16210
rect 46510 16158 46562 16210
rect 48638 16158 48690 16210
rect 1710 16046 1762 16098
rect 3390 16046 3442 16098
rect 4622 16046 4674 16098
rect 6190 16046 6242 16098
rect 7310 16046 7362 16098
rect 7870 16046 7922 16098
rect 9214 16046 9266 16098
rect 9550 16046 9602 16098
rect 10222 16046 10274 16098
rect 11790 16046 11842 16098
rect 12686 16046 12738 16098
rect 13806 16046 13858 16098
rect 14590 16046 14642 16098
rect 16718 16046 16770 16098
rect 17726 16046 17778 16098
rect 18174 16046 18226 16098
rect 19182 16046 19234 16098
rect 20526 16046 20578 16098
rect 22430 16046 22482 16098
rect 24110 16046 24162 16098
rect 25006 16046 25058 16098
rect 26350 16046 26402 16098
rect 29822 16046 29874 16098
rect 31390 16046 31442 16098
rect 31950 16046 32002 16098
rect 32286 16046 32338 16098
rect 32846 16046 32898 16098
rect 33182 16046 33234 16098
rect 34750 16046 34802 16098
rect 34974 16046 35026 16098
rect 35422 16046 35474 16098
rect 39118 16046 39170 16098
rect 39454 16046 39506 16098
rect 39566 16046 39618 16098
rect 39902 16046 39954 16098
rect 40350 16046 40402 16098
rect 40574 16046 40626 16098
rect 41134 16046 41186 16098
rect 42142 16046 42194 16098
rect 42478 16046 42530 16098
rect 42702 16046 42754 16098
rect 47070 16046 47122 16098
rect 52894 16046 52946 16098
rect 53118 16046 53170 16098
rect 55582 16046 55634 16098
rect 2046 15934 2098 15986
rect 2942 15934 2994 15986
rect 4062 15934 4114 15986
rect 4174 15934 4226 15986
rect 6302 15934 6354 15986
rect 8094 15934 8146 15986
rect 12014 15934 12066 15986
rect 14478 15934 14530 15986
rect 15262 15934 15314 15986
rect 22766 15934 22818 15986
rect 23998 15934 24050 15986
rect 25678 15934 25730 15986
rect 30046 15934 30098 15986
rect 30382 15934 30434 15986
rect 30606 15934 30658 15986
rect 33854 15934 33906 15986
rect 35198 15934 35250 15986
rect 38782 15934 38834 15986
rect 39790 15934 39842 15986
rect 41470 15934 41522 15986
rect 45278 15934 45330 15986
rect 48078 15934 48130 15986
rect 51662 15934 51714 15986
rect 55358 15934 55410 15986
rect 2718 15822 2770 15874
rect 3614 15822 3666 15874
rect 3838 15822 3890 15874
rect 12798 15822 12850 15874
rect 13022 15822 13074 15874
rect 15374 15822 15426 15874
rect 15598 15822 15650 15874
rect 15934 15822 15986 15874
rect 22542 15822 22594 15874
rect 23102 15822 23154 15874
rect 29150 15822 29202 15874
rect 29262 15822 29314 15874
rect 29374 15822 29426 15874
rect 32958 15822 33010 15874
rect 34078 15822 34130 15874
rect 38894 15822 38946 15874
rect 41246 15822 41298 15874
rect 45054 15822 45106 15874
rect 45166 15822 45218 15874
rect 51886 15822 51938 15874
rect 54238 15822 54290 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 50558 15654 50610 15706
rect 50662 15654 50714 15706
rect 50766 15654 50818 15706
rect 4846 15486 4898 15538
rect 4958 15486 5010 15538
rect 5518 15486 5570 15538
rect 5742 15486 5794 15538
rect 5966 15486 6018 15538
rect 6526 15486 6578 15538
rect 7310 15486 7362 15538
rect 8094 15486 8146 15538
rect 8878 15486 8930 15538
rect 9886 15486 9938 15538
rect 12462 15486 12514 15538
rect 16158 15486 16210 15538
rect 18398 15486 18450 15538
rect 23886 15486 23938 15538
rect 25902 15486 25954 15538
rect 26126 15486 26178 15538
rect 34526 15486 34578 15538
rect 37550 15486 37602 15538
rect 38558 15486 38610 15538
rect 40126 15486 40178 15538
rect 42142 15486 42194 15538
rect 47182 15486 47234 15538
rect 51998 15486 52050 15538
rect 6190 15374 6242 15426
rect 15598 15374 15650 15426
rect 17614 15374 17666 15426
rect 23662 15374 23714 15426
rect 23998 15374 24050 15426
rect 29038 15374 29090 15426
rect 30158 15374 30210 15426
rect 30942 15374 30994 15426
rect 33294 15374 33346 15426
rect 35982 15374 36034 15426
rect 40238 15374 40290 15426
rect 41134 15374 41186 15426
rect 42478 15374 42530 15426
rect 43710 15374 43762 15426
rect 46398 15374 46450 15426
rect 48750 15374 48802 15426
rect 2158 15262 2210 15314
rect 2606 15262 2658 15314
rect 3390 15262 3442 15314
rect 4510 15262 4562 15314
rect 4734 15262 4786 15314
rect 5182 15262 5234 15314
rect 5518 15262 5570 15314
rect 6750 15262 6802 15314
rect 7534 15262 7586 15314
rect 7870 15262 7922 15314
rect 8206 15262 8258 15314
rect 8542 15262 8594 15314
rect 9662 15262 9714 15314
rect 12126 15262 12178 15314
rect 13134 15262 13186 15314
rect 13694 15262 13746 15314
rect 15150 15262 15202 15314
rect 15486 15262 15538 15314
rect 15822 15262 15874 15314
rect 16494 15262 16546 15314
rect 16718 15262 16770 15314
rect 17838 15262 17890 15314
rect 18510 15262 18562 15314
rect 19182 15262 19234 15314
rect 20638 15262 20690 15314
rect 21310 15262 21362 15314
rect 22206 15262 22258 15314
rect 22430 15262 22482 15314
rect 23102 15262 23154 15314
rect 23438 15262 23490 15314
rect 25678 15262 25730 15314
rect 28590 15262 28642 15314
rect 29486 15262 29538 15314
rect 30494 15262 30546 15314
rect 31502 15262 31554 15314
rect 32062 15262 32114 15314
rect 33518 15262 33570 15314
rect 34190 15262 34242 15314
rect 35086 15262 35138 15314
rect 36318 15262 36370 15314
rect 36990 15262 37042 15314
rect 39006 15262 39058 15314
rect 39118 15262 39170 15314
rect 39342 15262 39394 15314
rect 39678 15262 39730 15314
rect 39902 15262 39954 15314
rect 41358 15262 41410 15314
rect 41582 15262 41634 15314
rect 41806 15262 41858 15314
rect 42030 15262 42082 15314
rect 42254 15262 42306 15314
rect 44382 15262 44434 15314
rect 45390 15262 45442 15314
rect 46174 15262 46226 15314
rect 46510 15262 46562 15314
rect 47070 15262 47122 15314
rect 47406 15262 47458 15314
rect 47966 15262 48018 15314
rect 49198 15262 49250 15314
rect 50878 15262 50930 15314
rect 53118 15262 53170 15314
rect 53454 15262 53506 15314
rect 14702 15150 14754 15202
rect 19294 15150 19346 15202
rect 25790 15150 25842 15202
rect 28142 15150 28194 15202
rect 30046 15150 30098 15202
rect 31614 15150 31666 15202
rect 33182 15150 33234 15202
rect 45278 15150 45330 15202
rect 47630 15150 47682 15202
rect 50990 15150 51042 15202
rect 52670 15150 52722 15202
rect 52894 15150 52946 15202
rect 3502 15038 3554 15090
rect 34862 15038 34914 15090
rect 47966 15038 48018 15090
rect 52446 15038 52498 15090
rect 55358 15038 55410 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 2942 14702 2994 14754
rect 7198 14702 7250 14754
rect 12798 14702 12850 14754
rect 26238 14702 26290 14754
rect 29486 14702 29538 14754
rect 31614 14702 31666 14754
rect 32174 14702 32226 14754
rect 42030 14702 42082 14754
rect 53006 14702 53058 14754
rect 57934 14702 57986 14754
rect 1822 14590 1874 14642
rect 3054 14590 3106 14642
rect 15710 14590 15762 14642
rect 18398 14590 18450 14642
rect 19070 14590 19122 14642
rect 22206 14590 22258 14642
rect 25678 14590 25730 14642
rect 27918 14590 27970 14642
rect 33518 14590 33570 14642
rect 34414 14590 34466 14642
rect 37774 14590 37826 14642
rect 41470 14590 41522 14642
rect 46062 14590 46114 14642
rect 48414 14590 48466 14642
rect 54126 14590 54178 14642
rect 54910 14590 54962 14642
rect 2606 14478 2658 14530
rect 3502 14478 3554 14530
rect 3838 14478 3890 14530
rect 6302 14478 6354 14530
rect 10110 14478 10162 14530
rect 10558 14478 10610 14530
rect 12126 14478 12178 14530
rect 14702 14478 14754 14530
rect 17390 14478 17442 14530
rect 19294 14478 19346 14530
rect 23550 14478 23602 14530
rect 24222 14478 24274 14530
rect 25006 14478 25058 14530
rect 25454 14478 25506 14530
rect 27022 14478 27074 14530
rect 27582 14478 27634 14530
rect 29486 14478 29538 14530
rect 30158 14478 30210 14530
rect 30830 14478 30882 14530
rect 31502 14478 31554 14530
rect 33182 14478 33234 14530
rect 35982 14478 36034 14530
rect 36206 14478 36258 14530
rect 36878 14478 36930 14530
rect 37662 14478 37714 14530
rect 39230 14478 39282 14530
rect 40910 14478 40962 14530
rect 41358 14478 41410 14530
rect 45166 14478 45218 14530
rect 45614 14478 45666 14530
rect 47742 14478 47794 14530
rect 48526 14478 48578 14530
rect 50542 14478 50594 14530
rect 51326 14478 51378 14530
rect 51998 14478 52050 14530
rect 52894 14478 52946 14530
rect 53342 14478 53394 14530
rect 53790 14478 53842 14530
rect 55582 14478 55634 14530
rect 4622 14366 4674 14418
rect 4958 14366 5010 14418
rect 6638 14366 6690 14418
rect 7198 14366 7250 14418
rect 7310 14366 7362 14418
rect 11230 14366 11282 14418
rect 12238 14366 12290 14418
rect 3726 14254 3778 14306
rect 10894 14254 10946 14306
rect 12462 14254 12514 14306
rect 12686 14310 12738 14362
rect 12798 14366 12850 14418
rect 14478 14366 14530 14418
rect 14590 14366 14642 14418
rect 16158 14366 16210 14418
rect 19966 14366 20018 14418
rect 20302 14366 20354 14418
rect 21422 14366 21474 14418
rect 21758 14366 21810 14418
rect 22430 14366 22482 14418
rect 24670 14366 24722 14418
rect 28030 14366 28082 14418
rect 29150 14366 29202 14418
rect 29822 14366 29874 14418
rect 32174 14366 32226 14418
rect 32286 14366 32338 14418
rect 33854 14366 33906 14418
rect 35534 14366 35586 14418
rect 35646 14366 35698 14418
rect 36318 14366 36370 14418
rect 38334 14366 38386 14418
rect 39006 14366 39058 14418
rect 40574 14366 40626 14418
rect 46174 14366 46226 14418
rect 49198 14366 49250 14418
rect 50430 14366 50482 14418
rect 51774 14366 51826 14418
rect 54798 14366 54850 14418
rect 15150 14254 15202 14306
rect 20414 14254 20466 14306
rect 20638 14254 20690 14306
rect 21534 14254 21586 14306
rect 24782 14254 24834 14306
rect 28590 14254 28642 14306
rect 29934 14254 29986 14306
rect 35310 14254 35362 14306
rect 40686 14254 40738 14306
rect 51214 14254 51266 14306
rect 55022 14254 55074 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 50558 14086 50610 14138
rect 50662 14086 50714 14138
rect 50766 14086 50818 14138
rect 2046 13918 2098 13970
rect 2718 13918 2770 13970
rect 3166 13918 3218 13970
rect 3726 13918 3778 13970
rect 4734 13918 4786 13970
rect 6974 13918 7026 13970
rect 15150 13918 15202 13970
rect 21646 13918 21698 13970
rect 22542 13918 22594 13970
rect 25454 13918 25506 13970
rect 41246 13918 41298 13970
rect 48862 13918 48914 13970
rect 50318 13918 50370 13970
rect 51214 13918 51266 13970
rect 53902 13918 53954 13970
rect 55358 13918 55410 13970
rect 2382 13806 2434 13858
rect 6526 13806 6578 13858
rect 23102 13806 23154 13858
rect 28142 13806 28194 13858
rect 35646 13806 35698 13858
rect 38558 13806 38610 13858
rect 40238 13806 40290 13858
rect 41022 13806 41074 13858
rect 45054 13806 45106 13858
rect 47406 13806 47458 13858
rect 47854 13806 47906 13858
rect 49086 13806 49138 13858
rect 49758 13806 49810 13858
rect 53566 13806 53618 13858
rect 56590 13806 56642 13858
rect 1822 13694 1874 13746
rect 3950 13694 4002 13746
rect 4398 13694 4450 13746
rect 6302 13694 6354 13746
rect 6862 13694 6914 13746
rect 11342 13694 11394 13746
rect 12686 13694 12738 13746
rect 12910 13694 12962 13746
rect 14142 13694 14194 13746
rect 14814 13694 14866 13746
rect 15710 13694 15762 13746
rect 16158 13694 16210 13746
rect 16606 13694 16658 13746
rect 16942 13694 16994 13746
rect 18062 13694 18114 13746
rect 18734 13694 18786 13746
rect 19742 13694 19794 13746
rect 20078 13694 20130 13746
rect 22206 13694 22258 13746
rect 22318 13694 22370 13746
rect 22654 13694 22706 13746
rect 25118 13694 25170 13746
rect 25454 13694 25506 13746
rect 25678 13694 25730 13746
rect 27358 13694 27410 13746
rect 30942 13694 30994 13746
rect 35086 13694 35138 13746
rect 38894 13694 38946 13746
rect 39790 13694 39842 13746
rect 40910 13694 40962 13746
rect 44606 13694 44658 13746
rect 46958 13694 47010 13746
rect 47742 13694 47794 13746
rect 48078 13694 48130 13746
rect 48750 13694 48802 13746
rect 49982 13694 50034 13746
rect 50654 13694 50706 13746
rect 52894 13694 52946 13746
rect 53454 13694 53506 13746
rect 54238 13694 54290 13746
rect 57038 13694 57090 13746
rect 10670 13582 10722 13634
rect 13582 13582 13634 13634
rect 13918 13582 13970 13634
rect 18286 13582 18338 13634
rect 20862 13582 20914 13634
rect 27918 13582 27970 13634
rect 29710 13582 29762 13634
rect 30158 13582 30210 13634
rect 30606 13582 30658 13634
rect 34750 13582 34802 13634
rect 41582 13582 41634 13634
rect 43038 13582 43090 13634
rect 44270 13582 44322 13634
rect 46510 13582 46562 13634
rect 54462 13582 54514 13634
rect 57374 13582 57426 13634
rect 6974 13470 7026 13522
rect 10894 13470 10946 13522
rect 14478 13470 14530 13522
rect 17726 13470 17778 13522
rect 23326 13470 23378 13522
rect 23662 13470 23714 13522
rect 43262 13470 43314 13522
rect 43598 13470 43650 13522
rect 50878 13470 50930 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 3502 13134 3554 13186
rect 25902 13134 25954 13186
rect 31278 13134 31330 13186
rect 39790 13134 39842 13186
rect 46734 13134 46786 13186
rect 4062 13022 4114 13074
rect 15262 13022 15314 13074
rect 16830 13022 16882 13074
rect 18734 13022 18786 13074
rect 22318 13022 22370 13074
rect 23102 13022 23154 13074
rect 26574 13022 26626 13074
rect 33070 13022 33122 13074
rect 53006 13022 53058 13074
rect 56814 13022 56866 13074
rect 1710 12910 1762 12962
rect 6638 12910 6690 12962
rect 7422 12910 7474 12962
rect 8654 12910 8706 12962
rect 8878 12910 8930 12962
rect 9102 12910 9154 12962
rect 10446 12910 10498 12962
rect 11342 12910 11394 12962
rect 11790 12910 11842 12962
rect 15710 12910 15762 12962
rect 17390 12910 17442 12962
rect 20750 12910 20802 12962
rect 21758 12910 21810 12962
rect 23214 12910 23266 12962
rect 23662 12910 23714 12962
rect 25790 12910 25842 12962
rect 30494 12910 30546 12962
rect 31166 12910 31218 12962
rect 34638 12910 34690 12962
rect 38558 12910 38610 12962
rect 38782 12910 38834 12962
rect 42702 12910 42754 12962
rect 43710 12910 43762 12962
rect 45166 12910 45218 12962
rect 46286 12910 46338 12962
rect 47070 12910 47122 12962
rect 48638 12910 48690 12962
rect 49758 12910 49810 12962
rect 50430 12910 50482 12962
rect 50654 12910 50706 12962
rect 51886 12910 51938 12962
rect 52222 12910 52274 12962
rect 52670 12910 52722 12962
rect 53566 12910 53618 12962
rect 55582 12910 55634 12962
rect 56142 12910 56194 12962
rect 56366 12910 56418 12962
rect 56926 12910 56978 12962
rect 57262 12910 57314 12962
rect 2046 12798 2098 12850
rect 2382 12798 2434 12850
rect 3502 12798 3554 12850
rect 3614 12798 3666 12850
rect 4510 12798 4562 12850
rect 5966 12798 6018 12850
rect 6862 12798 6914 12850
rect 7086 12798 7138 12850
rect 9550 12798 9602 12850
rect 10110 12798 10162 12850
rect 10558 12798 10610 12850
rect 12126 12798 12178 12850
rect 15598 12798 15650 12850
rect 19070 12798 19122 12850
rect 20414 12798 20466 12850
rect 26910 12798 26962 12850
rect 28366 12798 28418 12850
rect 33518 12798 33570 12850
rect 39006 12798 39058 12850
rect 39118 12798 39170 12850
rect 39790 12798 39842 12850
rect 39902 12798 39954 12850
rect 41694 12798 41746 12850
rect 42478 12798 42530 12850
rect 44270 12798 44322 12850
rect 44830 12798 44882 12850
rect 46174 12798 46226 12850
rect 47294 12798 47346 12850
rect 47854 12798 47906 12850
rect 48302 12798 48354 12850
rect 51998 12798 52050 12850
rect 53118 12798 53170 12850
rect 55246 12798 55298 12850
rect 55806 12798 55858 12850
rect 56702 12798 56754 12850
rect 2718 12686 2770 12738
rect 4958 12686 5010 12738
rect 6302 12686 6354 12738
rect 7646 12686 7698 12738
rect 9774 12686 9826 12738
rect 11454 12686 11506 12738
rect 12014 12686 12066 12738
rect 14702 12686 14754 12738
rect 25902 12686 25954 12738
rect 28478 12686 28530 12738
rect 34750 12686 34802 12738
rect 38110 12686 38162 12738
rect 38222 12686 38274 12738
rect 38446 12686 38498 12738
rect 41358 12686 41410 12738
rect 41582 12686 41634 12738
rect 44942 12686 44994 12738
rect 48414 12686 48466 12738
rect 55358 12686 55410 12738
rect 56030 12686 56082 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 50558 12518 50610 12570
rect 50662 12518 50714 12570
rect 50766 12518 50818 12570
rect 1710 12350 1762 12402
rect 4622 12350 4674 12402
rect 8542 12350 8594 12402
rect 8654 12350 8706 12402
rect 9662 12350 9714 12402
rect 10446 12350 10498 12402
rect 10670 12350 10722 12402
rect 13806 12350 13858 12402
rect 15374 12350 15426 12402
rect 18510 12350 18562 12402
rect 19742 12350 19794 12402
rect 20862 12350 20914 12402
rect 23438 12350 23490 12402
rect 26910 12350 26962 12402
rect 30158 12350 30210 12402
rect 31166 12350 31218 12402
rect 31950 12350 32002 12402
rect 33070 12350 33122 12402
rect 35982 12350 36034 12402
rect 38222 12350 38274 12402
rect 38894 12350 38946 12402
rect 47294 12350 47346 12402
rect 47518 12350 47570 12402
rect 47966 12350 48018 12402
rect 50094 12350 50146 12402
rect 52110 12350 52162 12402
rect 2046 12238 2098 12290
rect 2718 12238 2770 12290
rect 5518 12238 5570 12290
rect 5854 12238 5906 12290
rect 6526 12238 6578 12290
rect 8318 12238 8370 12290
rect 9886 12238 9938 12290
rect 10334 12238 10386 12290
rect 16382 12238 16434 12290
rect 17950 12238 18002 12290
rect 18286 12238 18338 12290
rect 19518 12238 19570 12290
rect 19966 12238 20018 12290
rect 20078 12238 20130 12290
rect 20750 12238 20802 12290
rect 22318 12238 22370 12290
rect 28478 12238 28530 12290
rect 29822 12238 29874 12290
rect 30718 12238 30770 12290
rect 31390 12238 31442 12290
rect 33294 12238 33346 12290
rect 35086 12238 35138 12290
rect 49534 12238 49586 12290
rect 52670 12238 52722 12290
rect 55134 12238 55186 12290
rect 56590 12238 56642 12290
rect 2382 12126 2434 12178
rect 3502 12126 3554 12178
rect 6302 12126 6354 12178
rect 6414 12126 6466 12178
rect 6750 12126 6802 12178
rect 7198 12126 7250 12178
rect 7534 12126 7586 12178
rect 8766 12126 8818 12178
rect 8990 12126 9042 12178
rect 9550 12126 9602 12178
rect 11678 12126 11730 12178
rect 13918 12126 13970 12178
rect 14366 12126 14418 12178
rect 16270 12126 16322 12178
rect 16494 12126 16546 12178
rect 16942 12126 16994 12178
rect 17726 12126 17778 12178
rect 19182 12126 19234 12178
rect 21086 12126 21138 12178
rect 21870 12126 21922 12178
rect 23214 12126 23266 12178
rect 23774 12126 23826 12178
rect 27134 12126 27186 12178
rect 27470 12126 27522 12178
rect 28254 12126 28306 12178
rect 29598 12126 29650 12178
rect 30606 12126 30658 12178
rect 30942 12126 30994 12178
rect 31502 12126 31554 12178
rect 33406 12126 33458 12178
rect 33854 12126 33906 12178
rect 33966 12126 34018 12178
rect 34078 12126 34130 12178
rect 34974 12126 35026 12178
rect 35982 12126 36034 12178
rect 36430 12126 36482 12178
rect 36654 12126 36706 12178
rect 37214 12126 37266 12178
rect 37998 12126 38050 12178
rect 38670 12126 38722 12178
rect 39566 12126 39618 12178
rect 42030 12126 42082 12178
rect 42590 12126 42642 12178
rect 43598 12126 43650 12178
rect 44046 12126 44098 12178
rect 44606 12126 44658 12178
rect 45166 12126 45218 12178
rect 47630 12126 47682 12178
rect 48078 12126 48130 12178
rect 49982 12126 50034 12178
rect 50206 12126 50258 12178
rect 50654 12126 50706 12178
rect 51438 12126 51490 12178
rect 51886 12126 51938 12178
rect 53790 12126 53842 12178
rect 55694 12126 55746 12178
rect 57038 12126 57090 12178
rect 3838 12014 3890 12066
rect 5182 12014 5234 12066
rect 7982 12014 8034 12066
rect 11566 12014 11618 12066
rect 12350 12014 12402 12066
rect 15822 12014 15874 12066
rect 21422 12014 21474 12066
rect 23326 12014 23378 12066
rect 28142 12014 28194 12066
rect 39790 12014 39842 12066
rect 42478 12014 42530 12066
rect 45054 12014 45106 12066
rect 47070 12014 47122 12066
rect 49646 12014 49698 12066
rect 50990 12014 51042 12066
rect 57374 12014 57426 12066
rect 13806 11902 13858 11954
rect 14254 11902 14306 11954
rect 26798 11902 26850 11954
rect 34526 11902 34578 11954
rect 40014 11902 40066 11954
rect 42926 11902 42978 11954
rect 45278 11902 45330 11954
rect 49310 11902 49362 11954
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 6302 11566 6354 11618
rect 14478 11566 14530 11618
rect 16382 11566 16434 11618
rect 18734 11566 18786 11618
rect 27470 11566 27522 11618
rect 35646 11566 35698 11618
rect 35982 11566 36034 11618
rect 39566 11566 39618 11618
rect 42254 11566 42306 11618
rect 53566 11566 53618 11618
rect 4622 11454 4674 11506
rect 4958 11454 5010 11506
rect 9214 11454 9266 11506
rect 11902 11454 11954 11506
rect 14366 11454 14418 11506
rect 15934 11454 15986 11506
rect 21534 11454 21586 11506
rect 26798 11454 26850 11506
rect 33182 11454 33234 11506
rect 38446 11454 38498 11506
rect 40686 11454 40738 11506
rect 41582 11454 41634 11506
rect 47630 11454 47682 11506
rect 55582 11454 55634 11506
rect 2830 11342 2882 11394
rect 3726 11342 3778 11394
rect 5630 11342 5682 11394
rect 6414 11342 6466 11394
rect 6862 11342 6914 11394
rect 9998 11342 10050 11394
rect 10894 11342 10946 11394
rect 12574 11342 12626 11394
rect 12798 11342 12850 11394
rect 14030 11342 14082 11394
rect 15486 11342 15538 11394
rect 15710 11342 15762 11394
rect 17166 11342 17218 11394
rect 17726 11342 17778 11394
rect 18510 11342 18562 11394
rect 19182 11342 19234 11394
rect 20302 11342 20354 11394
rect 22878 11342 22930 11394
rect 25454 11342 25506 11394
rect 27134 11342 27186 11394
rect 27806 11342 27858 11394
rect 28590 11342 28642 11394
rect 33294 11342 33346 11394
rect 33966 11342 34018 11394
rect 35086 11342 35138 11394
rect 35422 11342 35474 11394
rect 35870 11342 35922 11394
rect 37550 11342 37602 11394
rect 37886 11342 37938 11394
rect 39902 11342 39954 11394
rect 40238 11342 40290 11394
rect 41358 11342 41410 11394
rect 42030 11342 42082 11394
rect 45838 11342 45890 11394
rect 49870 11342 49922 11394
rect 50430 11342 50482 11394
rect 51886 11342 51938 11394
rect 53342 11342 53394 11394
rect 53566 11342 53618 11394
rect 1710 11230 1762 11282
rect 3390 11230 3442 11282
rect 4286 11230 4338 11282
rect 5742 11230 5794 11282
rect 9774 11230 9826 11282
rect 11342 11230 11394 11282
rect 11454 11230 11506 11282
rect 16830 11230 16882 11282
rect 21646 11230 21698 11282
rect 25118 11230 25170 11282
rect 26574 11230 26626 11282
rect 27358 11230 27410 11282
rect 29038 11230 29090 11282
rect 29262 11230 29314 11282
rect 29374 11230 29426 11282
rect 30942 11230 30994 11282
rect 33630 11230 33682 11282
rect 34190 11230 34242 11282
rect 38782 11230 38834 11282
rect 39118 11230 39170 11282
rect 39566 11230 39618 11282
rect 39678 11230 39730 11282
rect 40574 11230 40626 11282
rect 43262 11230 43314 11282
rect 43598 11230 43650 11282
rect 45614 11230 45666 11282
rect 47966 11230 48018 11282
rect 50318 11230 50370 11282
rect 52222 11230 52274 11282
rect 55134 11230 55186 11282
rect 55806 11230 55858 11282
rect 57486 11230 57538 11282
rect 2046 11118 2098 11170
rect 3054 11118 3106 11170
rect 3502 11118 3554 11170
rect 3950 11118 4002 11170
rect 4846 11118 4898 11170
rect 10782 11118 10834 11170
rect 11118 11118 11170 11170
rect 17614 11118 17666 11170
rect 23214 11118 23266 11170
rect 29822 11118 29874 11170
rect 30270 11118 30322 11170
rect 31278 11118 31330 11170
rect 33518 11118 33570 11170
rect 34974 11118 35026 11170
rect 40126 11118 40178 11170
rect 43374 11118 43426 11170
rect 45390 11118 45442 11170
rect 48078 11118 48130 11170
rect 48302 11118 48354 11170
rect 50206 11118 50258 11170
rect 51662 11118 51714 11170
rect 51998 11118 52050 11170
rect 54574 11118 54626 11170
rect 54686 11118 54738 11170
rect 54910 11118 54962 11170
rect 57374 11118 57426 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 50558 10950 50610 11002
rect 50662 10950 50714 11002
rect 50766 10950 50818 11002
rect 1822 10782 1874 10834
rect 3166 10782 3218 10834
rect 3502 10782 3554 10834
rect 3838 10782 3890 10834
rect 13918 10782 13970 10834
rect 14478 10782 14530 10834
rect 16382 10782 16434 10834
rect 20414 10782 20466 10834
rect 23550 10782 23602 10834
rect 28030 10782 28082 10834
rect 28254 10782 28306 10834
rect 28478 10782 28530 10834
rect 29598 10782 29650 10834
rect 34190 10782 34242 10834
rect 36654 10782 36706 10834
rect 37886 10782 37938 10834
rect 38110 10782 38162 10834
rect 39902 10782 39954 10834
rect 41806 10782 41858 10834
rect 53230 10782 53282 10834
rect 56702 10782 56754 10834
rect 2494 10670 2546 10722
rect 4510 10670 4562 10722
rect 5070 10670 5122 10722
rect 7758 10670 7810 10722
rect 9662 10670 9714 10722
rect 11118 10670 11170 10722
rect 19966 10670 20018 10722
rect 27134 10670 27186 10722
rect 30606 10670 30658 10722
rect 32510 10670 32562 10722
rect 33966 10670 34018 10722
rect 34526 10670 34578 10722
rect 35086 10670 35138 10722
rect 36766 10670 36818 10722
rect 38222 10670 38274 10722
rect 39118 10670 39170 10722
rect 41022 10670 41074 10722
rect 41582 10670 41634 10722
rect 44494 10670 44546 10722
rect 47742 10670 47794 10722
rect 48750 10670 48802 10722
rect 51102 10670 51154 10722
rect 52334 10670 52386 10722
rect 55694 10670 55746 10722
rect 2270 10558 2322 10610
rect 2830 10558 2882 10610
rect 4286 10558 4338 10610
rect 5294 10558 5346 10610
rect 5854 10558 5906 10610
rect 6414 10558 6466 10610
rect 7982 10558 8034 10610
rect 9774 10558 9826 10610
rect 9886 10558 9938 10610
rect 11230 10558 11282 10610
rect 12462 10558 12514 10610
rect 14590 10558 14642 10610
rect 17838 10558 17890 10610
rect 19182 10558 19234 10610
rect 22318 10558 22370 10610
rect 25678 10558 25730 10610
rect 26462 10558 26514 10610
rect 27470 10558 27522 10610
rect 28590 10558 28642 10610
rect 29934 10558 29986 10610
rect 31166 10558 31218 10610
rect 32062 10558 32114 10610
rect 33630 10558 33682 10610
rect 35982 10558 36034 10610
rect 38782 10558 38834 10610
rect 39342 10558 39394 10610
rect 40238 10558 40290 10610
rect 40910 10558 40962 10610
rect 41246 10558 41298 10610
rect 41470 10558 41522 10610
rect 43598 10558 43650 10610
rect 46062 10558 46114 10610
rect 47518 10558 47570 10610
rect 47966 10558 48018 10610
rect 48190 10558 48242 10610
rect 49198 10558 49250 10610
rect 51550 10558 51602 10610
rect 52222 10558 52274 10610
rect 53342 10558 53394 10610
rect 53678 10558 53730 10610
rect 53902 10558 53954 10610
rect 54574 10558 54626 10610
rect 55582 10558 55634 10610
rect 55918 10558 55970 10610
rect 56478 10558 56530 10610
rect 56814 10558 56866 10610
rect 57038 10558 57090 10610
rect 8990 10446 9042 10498
rect 11902 10446 11954 10498
rect 14030 10446 14082 10498
rect 14926 10446 14978 10498
rect 16494 10446 16546 10498
rect 17726 10446 17778 10498
rect 22766 10446 22818 10498
rect 26350 10446 26402 10498
rect 27694 10446 27746 10498
rect 29150 10446 29202 10498
rect 35870 10446 35922 10498
rect 43038 10446 43090 10498
rect 43486 10446 43538 10498
rect 45726 10446 45778 10498
rect 46398 10446 46450 10498
rect 49646 10446 49698 10498
rect 54238 10446 54290 10498
rect 6190 10334 6242 10386
rect 8206 10334 8258 10386
rect 8430 10334 8482 10386
rect 10334 10334 10386 10386
rect 13694 10334 13746 10386
rect 14478 10334 14530 10386
rect 15038 10334 15090 10386
rect 16158 10334 16210 10386
rect 36542 10334 36594 10386
rect 44382 10334 44434 10386
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 11790 9998 11842 10050
rect 12126 9998 12178 10050
rect 26462 9998 26514 10050
rect 30606 9998 30658 10050
rect 31166 9998 31218 10050
rect 55022 9998 55074 10050
rect 57486 9998 57538 10050
rect 4958 9886 5010 9938
rect 6750 9886 6802 9938
rect 9550 9886 9602 9938
rect 12350 9886 12402 9938
rect 14366 9886 14418 9938
rect 15038 9886 15090 9938
rect 23326 9886 23378 9938
rect 25566 9886 25618 9938
rect 37102 9886 37154 9938
rect 38334 9886 38386 9938
rect 42590 9886 42642 9938
rect 43038 9886 43090 9938
rect 44046 9886 44098 9938
rect 45278 9886 45330 9938
rect 50430 9886 50482 9938
rect 53342 9886 53394 9938
rect 54126 9886 54178 9938
rect 55582 9886 55634 9938
rect 1710 9774 1762 9826
rect 3278 9774 3330 9826
rect 4174 9774 4226 9826
rect 4846 9774 4898 9826
rect 6302 9774 6354 9826
rect 6974 9774 7026 9826
rect 8206 9774 8258 9826
rect 8430 9774 8482 9826
rect 9326 9774 9378 9826
rect 10334 9774 10386 9826
rect 13806 9774 13858 9826
rect 14030 9774 14082 9826
rect 15150 9774 15202 9826
rect 17614 9774 17666 9826
rect 19070 9774 19122 9826
rect 19742 9774 19794 9826
rect 20414 9774 20466 9826
rect 21422 9774 21474 9826
rect 21534 9774 21586 9826
rect 23774 9774 23826 9826
rect 25790 9774 25842 9826
rect 26014 9774 26066 9826
rect 29262 9774 29314 9826
rect 29710 9774 29762 9826
rect 32062 9774 32114 9826
rect 35646 9774 35698 9826
rect 35982 9774 36034 9826
rect 36542 9774 36594 9826
rect 37662 9774 37714 9826
rect 37886 9774 37938 9826
rect 38446 9774 38498 9826
rect 38670 9774 38722 9826
rect 39902 9774 39954 9826
rect 40798 9774 40850 9826
rect 43150 9774 43202 9826
rect 44270 9774 44322 9826
rect 47182 9774 47234 9826
rect 48526 9774 48578 9826
rect 50542 9774 50594 9826
rect 50990 9774 51042 9826
rect 51774 9774 51826 9826
rect 52110 9774 52162 9826
rect 52670 9774 52722 9826
rect 53678 9774 53730 9826
rect 54350 9774 54402 9826
rect 54574 9774 54626 9826
rect 56030 9774 56082 9826
rect 57150 9774 57202 9826
rect 2046 9662 2098 9714
rect 2718 9662 2770 9714
rect 3838 9662 3890 9714
rect 4958 9662 5010 9714
rect 6190 9662 6242 9714
rect 6750 9662 6802 9714
rect 9662 9662 9714 9714
rect 10446 9662 10498 9714
rect 11006 9662 11058 9714
rect 14814 9662 14866 9714
rect 17726 9662 17778 9714
rect 18734 9662 18786 9714
rect 23214 9662 23266 9714
rect 23550 9662 23602 9714
rect 28590 9662 28642 9714
rect 30718 9662 30770 9714
rect 31054 9662 31106 9714
rect 31726 9662 31778 9714
rect 31838 9662 31890 9714
rect 34750 9662 34802 9714
rect 34974 9662 35026 9714
rect 35310 9662 35362 9714
rect 36206 9662 36258 9714
rect 36318 9662 36370 9714
rect 38894 9662 38946 9714
rect 40126 9662 40178 9714
rect 41694 9662 41746 9714
rect 43934 9662 43986 9714
rect 45614 9662 45666 9714
rect 45726 9662 45778 9714
rect 46846 9662 46898 9714
rect 48190 9662 48242 9714
rect 49870 9662 49922 9714
rect 51886 9662 51938 9714
rect 52782 9662 52834 9714
rect 11118 9550 11170 9602
rect 17950 9550 18002 9602
rect 22766 9550 22818 9602
rect 27918 9550 27970 9602
rect 28254 9550 28306 9602
rect 30606 9550 30658 9602
rect 31166 9550 31218 9602
rect 34414 9550 34466 9602
rect 35086 9550 35138 9602
rect 35758 9550 35810 9602
rect 38334 9550 38386 9602
rect 39342 9550 39394 9602
rect 40910 9550 40962 9602
rect 41358 9550 41410 9602
rect 45950 9550 46002 9602
rect 46174 9550 46226 9602
rect 46510 9550 46562 9602
rect 46958 9550 47010 9602
rect 49758 9550 49810 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 50558 9382 50610 9434
rect 50662 9382 50714 9434
rect 50766 9382 50818 9434
rect 2718 9214 2770 9266
rect 3166 9214 3218 9266
rect 5406 9214 5458 9266
rect 6638 9214 6690 9266
rect 7310 9214 7362 9266
rect 8654 9214 8706 9266
rect 9886 9214 9938 9266
rect 1710 9102 1762 9154
rect 2046 9102 2098 9154
rect 4286 9102 4338 9154
rect 4510 9102 4562 9154
rect 5294 9102 5346 9154
rect 7758 9102 7810 9154
rect 11342 9102 11394 9154
rect 12238 9102 12290 9154
rect 13918 9102 13970 9154
rect 14590 9102 14642 9154
rect 14702 9158 14754 9210
rect 20974 9214 21026 9266
rect 22318 9214 22370 9266
rect 34750 9214 34802 9266
rect 35198 9214 35250 9266
rect 35534 9214 35586 9266
rect 36878 9214 36930 9266
rect 38446 9214 38498 9266
rect 38894 9214 38946 9266
rect 40238 9214 40290 9266
rect 40462 9214 40514 9266
rect 47518 9214 47570 9266
rect 48078 9214 48130 9266
rect 51774 9214 51826 9266
rect 52334 9214 52386 9266
rect 53454 9214 53506 9266
rect 53566 9214 53618 9266
rect 54238 9214 54290 9266
rect 55694 9214 55746 9266
rect 15486 9102 15538 9154
rect 19854 9102 19906 9154
rect 20862 9102 20914 9154
rect 21198 9102 21250 9154
rect 21982 9102 22034 9154
rect 22094 9102 22146 9154
rect 26350 9102 26402 9154
rect 26798 9102 26850 9154
rect 32286 9102 32338 9154
rect 35310 9102 35362 9154
rect 35982 9102 36034 9154
rect 36542 9102 36594 9154
rect 40126 9102 40178 9154
rect 42926 9102 42978 9154
rect 43038 9102 43090 9154
rect 47182 9102 47234 9154
rect 47294 9102 47346 9154
rect 47854 9102 47906 9154
rect 52894 9102 52946 9154
rect 55918 9102 55970 9154
rect 2382 8990 2434 9042
rect 4174 8990 4226 9042
rect 4622 8990 4674 9042
rect 5070 8990 5122 9042
rect 5630 8990 5682 9042
rect 6414 8990 6466 9042
rect 7086 8990 7138 9042
rect 8094 8990 8146 9042
rect 9662 8990 9714 9042
rect 10222 8990 10274 9042
rect 11118 8990 11170 9042
rect 13246 8990 13298 9042
rect 14926 8990 14978 9042
rect 15150 8990 15202 9042
rect 16270 8990 16322 9042
rect 17950 8990 18002 9042
rect 19294 8990 19346 9042
rect 25902 8990 25954 9042
rect 27582 8990 27634 9042
rect 28590 8990 28642 9042
rect 31390 8990 31442 9042
rect 31614 8990 31666 9042
rect 35086 8990 35138 9042
rect 36094 8990 36146 9042
rect 38222 8990 38274 9042
rect 39230 8990 39282 9042
rect 39790 8990 39842 9042
rect 43598 8990 43650 9042
rect 43822 8990 43874 9042
rect 44270 8990 44322 9042
rect 45166 8990 45218 9042
rect 47742 8990 47794 9042
rect 51662 8990 51714 9042
rect 52782 8990 52834 9042
rect 53118 8990 53170 9042
rect 54014 8990 54066 9042
rect 54126 8990 54178 9042
rect 54574 8990 54626 9042
rect 56030 8990 56082 9042
rect 56590 8990 56642 9042
rect 56702 8990 56754 9042
rect 57038 8990 57090 9042
rect 3614 8878 3666 8930
rect 7982 8878 8034 8930
rect 11006 8878 11058 8930
rect 11902 8878 11954 8930
rect 15710 8878 15762 8930
rect 20078 8878 20130 8930
rect 25566 8878 25618 8930
rect 29038 8878 29090 8930
rect 34190 8878 34242 8930
rect 42478 8878 42530 8930
rect 42590 8878 42642 8930
rect 45390 8878 45442 8930
rect 51326 8878 51378 8930
rect 34414 8766 34466 8818
rect 43038 8766 43090 8818
rect 45278 8766 45330 8818
rect 51774 8766 51826 8818
rect 53678 8766 53730 8818
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 24670 8430 24722 8482
rect 30382 8430 30434 8482
rect 2494 8318 2546 8370
rect 7982 8318 8034 8370
rect 10222 8318 10274 8370
rect 13582 8318 13634 8370
rect 14478 8318 14530 8370
rect 15038 8318 15090 8370
rect 15374 8318 15426 8370
rect 18174 8318 18226 8370
rect 25006 8318 25058 8370
rect 28142 8318 28194 8370
rect 31950 8318 32002 8370
rect 42142 8318 42194 8370
rect 49646 8318 49698 8370
rect 51214 8318 51266 8370
rect 52110 8318 52162 8370
rect 4398 8206 4450 8258
rect 4734 8206 4786 8258
rect 5742 8206 5794 8258
rect 5966 8206 6018 8258
rect 6638 8206 6690 8258
rect 7310 8206 7362 8258
rect 8318 8206 8370 8258
rect 9438 8206 9490 8258
rect 11118 8206 11170 8258
rect 13806 8206 13858 8258
rect 16830 8206 16882 8258
rect 18846 8206 18898 8258
rect 19406 8206 19458 8258
rect 20190 8206 20242 8258
rect 24670 8206 24722 8258
rect 25230 8206 25282 8258
rect 27470 8206 27522 8258
rect 28702 8206 28754 8258
rect 31838 8206 31890 8258
rect 32510 8206 32562 8258
rect 33070 8206 33122 8258
rect 34638 8206 34690 8258
rect 35310 8206 35362 8258
rect 38782 8206 38834 8258
rect 39118 8206 39170 8258
rect 39902 8206 39954 8258
rect 40350 8206 40402 8258
rect 43598 8206 43650 8258
rect 46398 8206 46450 8258
rect 50990 8206 51042 8258
rect 52894 8206 52946 8258
rect 53678 8206 53730 8258
rect 54014 8206 54066 8258
rect 54238 8206 54290 8258
rect 54462 8206 54514 8258
rect 55918 8206 55970 8258
rect 56590 8206 56642 8258
rect 57262 8206 57314 8258
rect 1710 8094 1762 8146
rect 2942 8094 2994 8146
rect 4510 8094 4562 8146
rect 7086 8094 7138 8146
rect 11454 8094 11506 8146
rect 11678 8094 11730 8146
rect 15822 8094 15874 8146
rect 19518 8094 19570 8146
rect 19854 8094 19906 8146
rect 19966 8094 20018 8146
rect 24334 8094 24386 8146
rect 27134 8094 27186 8146
rect 27246 8094 27298 8146
rect 30494 8094 30546 8146
rect 31166 8094 31218 8146
rect 31614 8094 31666 8146
rect 33294 8094 33346 8146
rect 34078 8094 34130 8146
rect 35534 8094 35586 8146
rect 35870 8094 35922 8146
rect 35982 8094 36034 8146
rect 36990 8094 37042 8146
rect 37774 8094 37826 8146
rect 38894 8094 38946 8146
rect 40798 8094 40850 8146
rect 42590 8094 42642 8146
rect 45950 8094 46002 8146
rect 47518 8094 47570 8146
rect 50206 8094 50258 8146
rect 53118 8094 53170 8146
rect 53230 8094 53282 8146
rect 54574 8094 54626 8146
rect 57486 8094 57538 8146
rect 2046 7982 2098 8034
rect 7422 7982 7474 8034
rect 7534 7982 7586 8034
rect 11902 7982 11954 8034
rect 25566 7982 25618 8034
rect 26910 7982 26962 8034
rect 28030 7982 28082 8034
rect 28254 7982 28306 8034
rect 30382 7982 30434 8034
rect 30830 7982 30882 8034
rect 36206 7982 36258 8034
rect 37102 7982 37154 8034
rect 37326 7982 37378 8034
rect 37886 7982 37938 8034
rect 38110 7982 38162 8034
rect 39454 7982 39506 8034
rect 41246 7982 41298 8034
rect 43934 7982 43986 8034
rect 47406 7982 47458 8034
rect 49870 7982 49922 8034
rect 50654 7982 50706 8034
rect 51774 7982 51826 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 50558 7814 50610 7866
rect 50662 7814 50714 7866
rect 50766 7814 50818 7866
rect 1822 7646 1874 7698
rect 8878 7646 8930 7698
rect 10110 7646 10162 7698
rect 16494 7646 16546 7698
rect 26238 7646 26290 7698
rect 27246 7646 27298 7698
rect 31390 7646 31442 7698
rect 33854 7646 33906 7698
rect 35310 7646 35362 7698
rect 5406 7534 5458 7586
rect 14702 7534 14754 7586
rect 14814 7534 14866 7586
rect 24670 7534 24722 7586
rect 26462 7534 26514 7586
rect 26910 7534 26962 7586
rect 27022 7534 27074 7586
rect 29822 7534 29874 7586
rect 30606 7534 30658 7586
rect 31726 7534 31778 7586
rect 34302 7534 34354 7586
rect 36654 7534 36706 7586
rect 36766 7534 36818 7586
rect 5630 7422 5682 7474
rect 7982 7422 8034 7474
rect 8430 7422 8482 7474
rect 9550 7422 9602 7474
rect 9774 7422 9826 7474
rect 11902 7422 11954 7474
rect 12574 7422 12626 7474
rect 13806 7422 13858 7474
rect 14478 7422 14530 7474
rect 15934 7422 15986 7474
rect 16158 7422 16210 7474
rect 22878 7422 22930 7474
rect 23214 7422 23266 7474
rect 24222 7422 24274 7474
rect 26574 7422 26626 7474
rect 27694 7422 27746 7474
rect 29038 7422 29090 7474
rect 30382 7422 30434 7474
rect 30718 7422 30770 7474
rect 31166 7422 31218 7474
rect 32062 7422 32114 7474
rect 34638 7422 34690 7474
rect 35086 7422 35138 7474
rect 35758 7422 35810 7474
rect 36318 7422 36370 7474
rect 36990 7422 37042 7474
rect 15262 7310 15314 7362
rect 15710 7310 15762 7362
rect 27582 7310 27634 7362
rect 33182 7310 33234 7362
rect 33630 7310 33682 7362
rect 33966 7310 34018 7362
rect 5966 7198 6018 7250
rect 37214 7646 37266 7698
rect 41022 7646 41074 7698
rect 49310 7646 49362 7698
rect 50654 7646 50706 7698
rect 56702 7646 56754 7698
rect 38894 7534 38946 7586
rect 40126 7534 40178 7586
rect 41582 7534 41634 7586
rect 41694 7534 41746 7586
rect 44606 7534 44658 7586
rect 47630 7534 47682 7586
rect 48750 7534 48802 7586
rect 51998 7534 52050 7586
rect 53454 7534 53506 7586
rect 55918 7534 55970 7586
rect 57262 7534 57314 7586
rect 38110 7422 38162 7474
rect 39230 7422 39282 7474
rect 39902 7422 39954 7474
rect 40798 7422 40850 7474
rect 41134 7422 41186 7474
rect 41358 7422 41410 7474
rect 44158 7422 44210 7474
rect 47182 7422 47234 7474
rect 47518 7422 47570 7474
rect 50206 7422 50258 7474
rect 50430 7422 50482 7474
rect 50878 7422 50930 7474
rect 51662 7422 51714 7474
rect 54686 7422 54738 7474
rect 56590 7422 56642 7474
rect 57150 7422 57202 7474
rect 37550 7310 37602 7362
rect 38334 7310 38386 7362
rect 43710 7310 43762 7362
rect 50766 7310 50818 7362
rect 51550 7310 51602 7362
rect 53342 7310 53394 7362
rect 8206 7198 8258 7250
rect 14030 7198 14082 7250
rect 37102 7198 37154 7250
rect 48974 7198 49026 7250
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 24334 6862 24386 6914
rect 29262 6862 29314 6914
rect 33406 6862 33458 6914
rect 37886 6862 37938 6914
rect 13582 6750 13634 6802
rect 24670 6750 24722 6802
rect 28254 6750 28306 6802
rect 35758 6750 35810 6802
rect 37438 6750 37490 6802
rect 40910 6750 40962 6802
rect 43150 6750 43202 6802
rect 48974 6750 49026 6802
rect 51102 6750 51154 6802
rect 13918 6638 13970 6690
rect 14702 6638 14754 6690
rect 15038 6638 15090 6690
rect 24446 6638 24498 6690
rect 27918 6638 27970 6690
rect 28366 6638 28418 6690
rect 29150 6638 29202 6690
rect 29374 6638 29426 6690
rect 29598 6638 29650 6690
rect 29822 6638 29874 6690
rect 32174 6638 32226 6690
rect 32510 6638 32562 6690
rect 35870 6638 35922 6690
rect 36542 6638 36594 6690
rect 36990 6638 37042 6690
rect 37214 6638 37266 6690
rect 38110 6638 38162 6690
rect 39118 6638 39170 6690
rect 39902 6638 39954 6690
rect 41022 6638 41074 6690
rect 42366 6638 42418 6690
rect 47854 6638 47906 6690
rect 48190 6638 48242 6690
rect 49086 6638 49138 6690
rect 50878 6638 50930 6690
rect 51438 6638 51490 6690
rect 53006 6638 53058 6690
rect 53902 6638 53954 6690
rect 14814 6526 14866 6578
rect 26126 6526 26178 6578
rect 26798 6526 26850 6578
rect 27470 6526 27522 6578
rect 31838 6526 31890 6578
rect 32286 6526 32338 6578
rect 32734 6526 32786 6578
rect 33294 6526 33346 6578
rect 34414 6526 34466 6578
rect 35198 6526 35250 6578
rect 35422 6526 35474 6578
rect 36206 6526 36258 6578
rect 38222 6526 38274 6578
rect 47406 6526 47458 6578
rect 49758 6526 49810 6578
rect 51326 6526 51378 6578
rect 53118 6526 53170 6578
rect 25790 6414 25842 6466
rect 26462 6414 26514 6466
rect 27134 6414 27186 6466
rect 28030 6414 28082 6466
rect 28254 6414 28306 6466
rect 30942 6414 30994 6466
rect 31502 6414 31554 6466
rect 32846 6414 32898 6466
rect 33070 6414 33122 6466
rect 33406 6414 33458 6466
rect 34078 6414 34130 6466
rect 34862 6414 34914 6466
rect 35646 6414 35698 6466
rect 36318 6414 36370 6466
rect 39118 6414 39170 6466
rect 39678 6414 39730 6466
rect 40238 6414 40290 6466
rect 40462 6414 40514 6466
rect 40574 6414 40626 6466
rect 45502 6414 45554 6466
rect 48302 6414 48354 6466
rect 50094 6414 50146 6466
rect 50206 6414 50258 6466
rect 50318 6414 50370 6466
rect 50542 6414 50594 6466
rect 54014 6414 54066 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 50558 6246 50610 6298
rect 50662 6246 50714 6298
rect 50766 6246 50818 6298
rect 25342 6078 25394 6130
rect 25566 6078 25618 6130
rect 26798 6078 26850 6130
rect 27022 6078 27074 6130
rect 27358 6078 27410 6130
rect 27582 6078 27634 6130
rect 31166 6078 31218 6130
rect 33742 6078 33794 6130
rect 35422 6078 35474 6130
rect 35870 6078 35922 6130
rect 40014 6078 40066 6130
rect 41918 6078 41970 6130
rect 47742 6078 47794 6130
rect 52558 6078 52610 6130
rect 53342 6078 53394 6130
rect 53566 6078 53618 6130
rect 26686 5966 26738 6018
rect 27246 5966 27298 6018
rect 32174 5966 32226 6018
rect 33070 5966 33122 6018
rect 37214 5966 37266 6018
rect 37550 5966 37602 6018
rect 40350 5966 40402 6018
rect 41022 5966 41074 6018
rect 45278 5966 45330 6018
rect 49198 5966 49250 6018
rect 49646 5966 49698 6018
rect 53230 5966 53282 6018
rect 25678 5854 25730 5906
rect 29934 5854 29986 5906
rect 31502 5854 31554 5906
rect 31838 5854 31890 5906
rect 33294 5854 33346 5906
rect 34078 5854 34130 5906
rect 34526 5854 34578 5906
rect 34638 5854 34690 5906
rect 34750 5854 34802 5906
rect 35198 5854 35250 5906
rect 36318 5854 36370 5906
rect 36766 5854 36818 5906
rect 37774 5854 37826 5906
rect 39790 5854 39842 5906
rect 40126 5854 40178 5906
rect 40910 5854 40962 5906
rect 41806 5854 41858 5906
rect 42366 5854 42418 5906
rect 42590 5854 42642 5906
rect 44382 5854 44434 5906
rect 44830 5854 44882 5906
rect 46286 5854 46338 5906
rect 47182 5854 47234 5906
rect 50430 5854 50482 5906
rect 51102 5854 51154 5906
rect 51438 5854 51490 5906
rect 52782 5854 52834 5906
rect 30942 5742 30994 5794
rect 37102 5742 37154 5794
rect 38222 5742 38274 5794
rect 38894 5742 38946 5794
rect 43374 5742 43426 5794
rect 43822 5742 43874 5794
rect 44942 5742 44994 5794
rect 46510 5742 46562 5794
rect 47854 5742 47906 5794
rect 49310 5742 49362 5794
rect 28030 5630 28082 5682
rect 38446 5630 38498 5682
rect 38670 5630 38722 5682
rect 39342 5630 39394 5682
rect 42926 5630 42978 5682
rect 47518 5630 47570 5682
rect 48974 5630 49026 5682
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 39678 5294 39730 5346
rect 40910 5294 40962 5346
rect 41246 5294 41298 5346
rect 44382 5294 44434 5346
rect 48078 5294 48130 5346
rect 50318 5294 50370 5346
rect 50766 5294 50818 5346
rect 28702 5182 28754 5234
rect 30606 5182 30658 5234
rect 33518 5182 33570 5234
rect 36430 5182 36482 5234
rect 38894 5182 38946 5234
rect 39342 5182 39394 5234
rect 40686 5182 40738 5234
rect 44942 5182 44994 5234
rect 47070 5182 47122 5234
rect 48414 5182 48466 5234
rect 49870 5182 49922 5234
rect 50094 5182 50146 5234
rect 29822 5070 29874 5122
rect 30942 5070 30994 5122
rect 31950 5070 32002 5122
rect 32622 5070 32674 5122
rect 32846 5070 32898 5122
rect 33182 5070 33234 5122
rect 33742 5070 33794 5122
rect 34638 5070 34690 5122
rect 34974 5070 35026 5122
rect 35870 5070 35922 5122
rect 36094 5070 36146 5122
rect 37214 5070 37266 5122
rect 37662 5070 37714 5122
rect 38670 5070 38722 5122
rect 39790 5070 39842 5122
rect 43710 5070 43762 5122
rect 44046 5070 44098 5122
rect 44718 5070 44770 5122
rect 45166 5070 45218 5122
rect 45390 5070 45442 5122
rect 45726 5070 45778 5122
rect 46958 5070 47010 5122
rect 47518 5070 47570 5122
rect 48190 5070 48242 5122
rect 48526 5070 48578 5122
rect 29374 4958 29426 5010
rect 29486 4958 29538 5010
rect 30158 4958 30210 5010
rect 31278 4958 31330 5010
rect 32174 4958 32226 5010
rect 32734 4958 32786 5010
rect 33966 4958 34018 5010
rect 35198 4958 35250 5010
rect 36318 4958 36370 5010
rect 36990 4958 37042 5010
rect 37998 4958 38050 5010
rect 43150 4958 43202 5010
rect 44270 4958 44322 5010
rect 45950 4958 46002 5010
rect 46062 4958 46114 5010
rect 46622 4958 46674 5010
rect 29150 4846 29202 4898
rect 35422 4846 35474 4898
rect 42030 4846 42082 4898
rect 42254 4846 42306 4898
rect 42366 4846 42418 4898
rect 42478 4846 42530 4898
rect 42814 4846 42866 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 50558 4678 50610 4730
rect 50662 4678 50714 4730
rect 50766 4678 50818 4730
rect 31390 4510 31442 4562
rect 31726 4510 31778 4562
rect 32062 4510 32114 4562
rect 32398 4510 32450 4562
rect 33070 4510 33122 4562
rect 33406 4510 33458 4562
rect 40910 4510 40962 4562
rect 37214 4398 37266 4450
rect 42142 4398 42194 4450
rect 45726 4398 45778 4450
rect 47966 4398 48018 4450
rect 30606 4286 30658 4338
rect 33854 4286 33906 4338
rect 36990 4286 37042 4338
rect 37886 4286 37938 4338
rect 39342 4286 39394 4338
rect 40014 4286 40066 4338
rect 42366 4286 42418 4338
rect 44046 4286 44098 4338
rect 44942 4286 44994 4338
rect 45950 4286 46002 4338
rect 47182 4286 47234 4338
rect 26910 4174 26962 4226
rect 28254 4174 28306 4226
rect 37438 4174 37490 4226
rect 37550 4174 37602 4226
rect 39118 4174 39170 4226
rect 41358 4174 41410 4226
rect 44158 4174 44210 4226
rect 44718 4174 44770 4226
rect 28702 4062 28754 4114
rect 34862 4062 34914 4114
rect 44606 4062 44658 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 35086 3726 35138 3778
rect 40350 3726 40402 3778
rect 42366 3726 42418 3778
rect 42590 3726 42642 3778
rect 43038 3726 43090 3778
rect 48190 3726 48242 3778
rect 29262 3614 29314 3666
rect 36206 3614 36258 3666
rect 39790 3614 39842 3666
rect 42142 3614 42194 3666
rect 25118 3502 25170 3554
rect 26014 3502 26066 3554
rect 31166 3502 31218 3554
rect 32510 3502 32562 3554
rect 32958 3502 33010 3554
rect 33518 3502 33570 3554
rect 34302 3502 34354 3554
rect 34862 3502 34914 3554
rect 38110 3502 38162 3554
rect 39118 3502 39170 3554
rect 40014 3502 40066 3554
rect 40910 3502 40962 3554
rect 41582 3502 41634 3554
rect 43822 3502 43874 3554
rect 45166 3502 45218 3554
rect 45614 3502 45666 3554
rect 45950 3502 46002 3554
rect 46286 3502 46338 3554
rect 47406 3502 47458 3554
rect 47630 3502 47682 3554
rect 47742 3502 47794 3554
rect 14142 3390 14194 3442
rect 14366 3390 14418 3442
rect 14702 3390 14754 3442
rect 25566 3390 25618 3442
rect 25790 3390 25842 3442
rect 26462 3390 26514 3442
rect 26798 3390 26850 3442
rect 27134 3390 27186 3442
rect 27470 3390 27522 3442
rect 28366 3390 28418 3442
rect 28702 3390 28754 3442
rect 32174 3390 32226 3442
rect 33182 3390 33234 3442
rect 33742 3390 33794 3442
rect 35534 3390 35586 3442
rect 38894 3390 38946 3442
rect 40686 3390 40738 3442
rect 41358 3390 41410 3442
rect 43598 3390 43650 3442
rect 44270 3390 44322 3442
rect 44606 3390 44658 3442
rect 44942 3390 44994 3442
rect 45726 3390 45778 3442
rect 46734 3390 46786 3442
rect 21758 3278 21810 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
rect 50558 3110 50610 3162
rect 50662 3110 50714 3162
rect 50766 3110 50818 3162
<< metal2 >>
rect 9408 49200 9520 50000
rect 10080 49200 10192 50000
rect 12096 49200 12208 50000
rect 12768 49200 12880 50000
rect 16800 49200 16912 50000
rect 17472 49200 17584 50000
rect 18144 49200 18256 50000
rect 26208 49200 26320 50000
rect 26880 49200 26992 50000
rect 28224 49200 28336 50000
rect 28896 49200 29008 50000
rect 29568 49200 29680 50000
rect 30240 49200 30352 50000
rect 34272 49200 34384 50000
rect 36960 49200 37072 50000
rect 37632 49200 37744 50000
rect 38304 49200 38416 50000
rect 38976 49200 39088 50000
rect 39648 49200 39760 50000
rect 40320 49200 40432 50000
rect 40992 49200 41104 50000
rect 41664 49200 41776 50000
rect 42336 49200 42448 50000
rect 43008 49200 43120 50000
rect 43680 49200 43792 50000
rect 44352 49200 44464 50000
rect 45024 49200 45136 50000
rect 45696 49200 45808 50000
rect 46368 49200 46480 50000
rect 8764 46450 8820 46462
rect 8764 46398 8766 46450
rect 8818 46398 8820 46450
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 8764 45890 8820 46398
rect 8764 45838 8766 45890
rect 8818 45838 8820 45890
rect 8764 45826 8820 45838
rect 9100 46450 9156 46462
rect 9100 46398 9102 46450
rect 9154 46398 9156 46450
rect 8204 45780 8260 45790
rect 8204 45686 8260 45724
rect 8428 45666 8484 45678
rect 8428 45614 8430 45666
rect 8482 45614 8484 45666
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 7980 44436 8036 44446
rect 1708 44210 1764 44222
rect 1708 44158 1710 44210
rect 1762 44158 1764 44210
rect 1708 43764 1764 44158
rect 7980 44210 8036 44380
rect 7980 44158 7982 44210
rect 8034 44158 8036 44210
rect 7980 44146 8036 44158
rect 2044 44100 2100 44110
rect 2044 44006 2100 44044
rect 2492 44098 2548 44110
rect 2492 44046 2494 44098
rect 2546 44046 2548 44098
rect 1708 43698 1764 43708
rect 2492 43764 2548 44046
rect 2492 43698 2548 43708
rect 7084 44100 7140 44110
rect 7084 43762 7140 44044
rect 7644 44100 7700 44110
rect 7644 44006 7700 44044
rect 8316 44100 8372 44110
rect 7084 43710 7086 43762
rect 7138 43710 7140 43762
rect 7084 43698 7140 43710
rect 8316 43708 8372 44044
rect 7756 43652 8372 43708
rect 7196 43540 7252 43550
rect 7196 43446 7252 43484
rect 2156 43426 2212 43438
rect 2156 43374 2158 43426
rect 2210 43374 2212 43426
rect 1820 42754 1876 42766
rect 1820 42702 1822 42754
rect 1874 42702 1876 42754
rect 1708 41972 1764 41982
rect 1596 41916 1708 41972
rect 1596 41524 1652 41916
rect 1708 41878 1764 41916
rect 1708 41748 1764 41758
rect 1820 41748 1876 42702
rect 2156 42644 2212 43374
rect 7084 43316 7140 43326
rect 7084 43222 7140 43260
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 7644 42756 7700 42766
rect 7756 42756 7812 43652
rect 7868 43538 7924 43550
rect 7868 43486 7870 43538
rect 7922 43486 7924 43538
rect 7868 43316 7924 43486
rect 8428 43540 8484 45614
rect 9100 45330 9156 46398
rect 9436 46450 9492 49200
rect 10108 46562 10164 49200
rect 10108 46510 10110 46562
rect 10162 46510 10164 46562
rect 10108 46498 10164 46510
rect 10780 46562 10836 46574
rect 10780 46510 10782 46562
rect 10834 46510 10836 46562
rect 9436 46398 9438 46450
rect 9490 46398 9492 46450
rect 9436 46386 9492 46398
rect 9660 46004 9716 46014
rect 9660 45910 9716 45948
rect 9996 45892 10052 45902
rect 10780 45892 10836 46510
rect 11900 46004 11956 46014
rect 9996 45890 10164 45892
rect 9996 45838 9998 45890
rect 10050 45838 10164 45890
rect 9996 45836 10164 45838
rect 9996 45826 10052 45836
rect 9100 45278 9102 45330
rect 9154 45278 9156 45330
rect 9100 45266 9156 45278
rect 10108 45668 10164 45836
rect 10780 45798 10836 45836
rect 11564 45892 11620 45902
rect 11564 45778 11620 45836
rect 11900 45892 11956 45948
rect 12124 45892 12180 49200
rect 12796 47012 12852 49200
rect 11900 45890 12180 45892
rect 11900 45838 11902 45890
rect 11954 45838 12180 45890
rect 11900 45836 12180 45838
rect 12348 46956 12852 47012
rect 12348 46004 12404 46956
rect 12348 45890 12404 45948
rect 14476 46004 14532 46014
rect 14476 45910 14532 45948
rect 16044 46004 16100 46014
rect 16044 45910 16100 45948
rect 16828 46004 16884 49200
rect 12348 45838 12350 45890
rect 12402 45838 12404 45890
rect 11900 45826 11956 45836
rect 12348 45826 12404 45838
rect 13132 45892 13188 45902
rect 13132 45798 13188 45836
rect 13804 45890 13860 45902
rect 13804 45838 13806 45890
rect 13858 45838 13860 45890
rect 11564 45726 11566 45778
rect 11618 45726 11620 45778
rect 9884 45220 9940 45230
rect 9884 45126 9940 45164
rect 9660 45108 9716 45118
rect 9660 45106 9828 45108
rect 9660 45054 9662 45106
rect 9714 45054 9828 45106
rect 9660 45052 9828 45054
rect 9660 45042 9716 45052
rect 8428 43474 8484 43484
rect 8652 44436 8708 44446
rect 7868 42868 7924 43260
rect 8204 43426 8260 43438
rect 8204 43374 8206 43426
rect 8258 43374 8260 43426
rect 8204 42978 8260 43374
rect 8540 43428 8596 43438
rect 8540 43334 8596 43372
rect 8204 42926 8206 42978
rect 8258 42926 8260 42978
rect 7980 42868 8036 42878
rect 7868 42866 8036 42868
rect 7868 42814 7982 42866
rect 8034 42814 8036 42866
rect 7868 42812 8036 42814
rect 7980 42802 8036 42812
rect 7644 42754 7812 42756
rect 7644 42702 7646 42754
rect 7698 42702 7812 42754
rect 7644 42700 7812 42702
rect 7644 42690 7700 42700
rect 2380 42644 2436 42654
rect 2156 42642 2436 42644
rect 2156 42590 2382 42642
rect 2434 42590 2436 42642
rect 2156 42588 2436 42590
rect 2044 42530 2100 42542
rect 2044 42478 2046 42530
rect 2098 42478 2100 42530
rect 2044 42308 2100 42478
rect 2380 42420 2436 42588
rect 7308 42644 7364 42654
rect 7308 42550 7364 42588
rect 8204 42644 8260 42926
rect 8652 42868 8708 44380
rect 9660 44436 9716 44446
rect 9772 44436 9828 45052
rect 9772 44380 9940 44436
rect 9660 44322 9716 44380
rect 9660 44270 9662 44322
rect 9714 44270 9716 44322
rect 9660 44258 9716 44270
rect 9884 44324 9940 44380
rect 9884 44322 10052 44324
rect 9884 44270 9886 44322
rect 9938 44270 10052 44322
rect 9884 44268 10052 44270
rect 9884 44258 9940 44268
rect 9772 44212 9828 44222
rect 8764 44100 8820 44110
rect 8764 44006 8820 44044
rect 9100 44098 9156 44110
rect 9100 44046 9102 44098
rect 9154 44046 9156 44098
rect 8204 42578 8260 42588
rect 8428 42812 8708 42868
rect 8876 43540 8932 43550
rect 2716 42532 2772 42542
rect 3164 42532 3220 42542
rect 2716 42438 2772 42476
rect 3052 42530 3220 42532
rect 3052 42478 3166 42530
rect 3218 42478 3220 42530
rect 3052 42476 3220 42478
rect 2380 42354 2436 42364
rect 2044 42242 2100 42252
rect 1764 41692 1876 41748
rect 2044 42082 2100 42094
rect 2044 42030 2046 42082
rect 2098 42030 2100 42082
rect 1708 41682 1764 41692
rect 2044 41636 2100 42030
rect 2716 42082 2772 42094
rect 2716 42030 2718 42082
rect 2770 42030 2772 42082
rect 2044 41570 2100 41580
rect 2380 41970 2436 41982
rect 2380 41918 2382 41970
rect 2434 41918 2436 41970
rect 2380 41860 2436 41918
rect 1596 41468 1764 41524
rect 1708 40404 1764 41468
rect 2268 41188 2324 41198
rect 2268 41094 2324 41132
rect 2380 41076 2436 41804
rect 2380 41010 2436 41020
rect 2604 41186 2660 41198
rect 2604 41134 2606 41186
rect 2658 41134 2660 41186
rect 1708 40338 1764 40348
rect 2604 40402 2660 41134
rect 2716 41076 2772 42030
rect 2940 41748 2996 41758
rect 3052 41748 3108 42476
rect 3164 42466 3220 42476
rect 7532 42532 7588 42542
rect 4396 42308 4452 42318
rect 4396 42196 4452 42252
rect 4396 42194 4900 42196
rect 4396 42142 4398 42194
rect 4450 42142 4900 42194
rect 4396 42140 4900 42142
rect 4396 42130 4452 42140
rect 3612 41972 3668 41982
rect 4508 41972 4564 41982
rect 3612 41878 3668 41916
rect 4284 41970 4564 41972
rect 4284 41918 4510 41970
rect 4562 41918 4564 41970
rect 4284 41916 4564 41918
rect 3164 41860 3220 41870
rect 3164 41766 3220 41804
rect 2996 41692 3108 41748
rect 3388 41748 3444 41758
rect 2940 41682 2996 41692
rect 3388 41188 3444 41692
rect 4284 41636 4340 41916
rect 4508 41906 4564 41916
rect 4396 41748 4452 41786
rect 4396 41682 4452 41692
rect 4284 41570 4340 41580
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 4844 41188 4900 42140
rect 7420 41972 7476 41982
rect 7532 41972 7588 42476
rect 8428 42420 8484 42812
rect 8876 42754 8932 43484
rect 8876 42702 8878 42754
rect 8930 42702 8932 42754
rect 8876 42690 8932 42702
rect 9100 42756 9156 44046
rect 9772 43764 9828 44156
rect 9884 43764 9940 43774
rect 9772 43762 9940 43764
rect 9772 43710 9886 43762
rect 9938 43710 9940 43762
rect 9772 43708 9940 43710
rect 9884 43698 9940 43708
rect 9996 43764 10052 44268
rect 10108 44322 10164 45612
rect 10220 45666 10276 45678
rect 10220 45614 10222 45666
rect 10274 45614 10276 45666
rect 10220 45332 10276 45614
rect 10556 45668 10612 45678
rect 10556 45574 10612 45612
rect 10444 45332 10500 45342
rect 10220 45276 10444 45332
rect 10444 45238 10500 45276
rect 11116 45220 11172 45230
rect 11564 45220 11620 45726
rect 12572 45780 12628 45790
rect 12572 45686 12628 45724
rect 13244 45780 13300 45790
rect 13244 45686 13300 45724
rect 13468 45778 13524 45790
rect 13468 45726 13470 45778
rect 13522 45726 13524 45778
rect 10220 45106 10276 45118
rect 10220 45054 10222 45106
rect 10274 45054 10276 45106
rect 10220 44436 10276 45054
rect 11116 45106 11172 45164
rect 11116 45054 11118 45106
rect 11170 45054 11172 45106
rect 11116 45042 11172 45054
rect 11340 45218 11620 45220
rect 11340 45166 11566 45218
rect 11618 45166 11620 45218
rect 11340 45164 11620 45166
rect 10220 44370 10276 44380
rect 10556 44436 10612 44446
rect 10556 44342 10612 44380
rect 10108 44270 10110 44322
rect 10162 44270 10164 44322
rect 10108 44100 10164 44270
rect 11340 44212 11396 45164
rect 11564 45154 11620 45164
rect 12124 45332 12180 45342
rect 12124 45106 12180 45276
rect 12236 45220 12292 45230
rect 12236 45126 12292 45164
rect 13468 45220 13524 45726
rect 13804 45332 13860 45838
rect 16492 45892 16548 45902
rect 16828 45892 16884 45948
rect 17052 45892 17108 45902
rect 16828 45890 17108 45892
rect 16828 45838 17054 45890
rect 17106 45838 17108 45890
rect 16828 45836 17108 45838
rect 16492 45798 16548 45836
rect 17052 45826 17108 45836
rect 17500 45892 17556 49200
rect 18172 46900 18228 49200
rect 18172 46844 18676 46900
rect 18620 46004 18676 46844
rect 26236 46116 26292 49200
rect 26908 47124 26964 49200
rect 26908 47068 27300 47124
rect 26236 46050 26292 46060
rect 19180 46004 19236 46014
rect 26796 46004 26852 46014
rect 18620 46002 19236 46004
rect 18620 45950 19182 46002
rect 19234 45950 19236 46002
rect 18620 45948 19236 45950
rect 17724 45892 17780 45902
rect 17556 45890 17780 45892
rect 17556 45838 17726 45890
rect 17778 45838 17780 45890
rect 17556 45836 17780 45838
rect 17500 45798 17556 45836
rect 17724 45826 17780 45836
rect 18620 45890 18676 45948
rect 19180 45938 19236 45948
rect 21196 45948 21812 46004
rect 18620 45838 18622 45890
rect 18674 45838 18676 45890
rect 18620 45826 18676 45838
rect 21084 45892 21140 45902
rect 21196 45892 21252 45948
rect 21084 45890 21252 45892
rect 21084 45838 21086 45890
rect 21138 45838 21252 45890
rect 21084 45836 21252 45838
rect 21084 45826 21140 45836
rect 13804 45266 13860 45276
rect 13916 45780 13972 45790
rect 13468 45154 13524 45164
rect 13916 45218 13972 45724
rect 15372 45778 15428 45790
rect 15372 45726 15374 45778
rect 15426 45726 15428 45778
rect 14140 45668 14196 45678
rect 14140 45666 14308 45668
rect 14140 45614 14142 45666
rect 14194 45614 14308 45666
rect 14140 45612 14308 45614
rect 14140 45602 14196 45612
rect 13916 45166 13918 45218
rect 13970 45166 13972 45218
rect 12124 45054 12126 45106
rect 12178 45054 12180 45106
rect 12124 45042 12180 45054
rect 12684 45106 12740 45118
rect 12684 45054 12686 45106
rect 12738 45054 12740 45106
rect 11564 44996 11620 45006
rect 11564 44902 11620 44940
rect 12460 44996 12516 45006
rect 11900 44882 11956 44894
rect 11900 44830 11902 44882
rect 11954 44830 11956 44882
rect 11340 44146 11396 44156
rect 11452 44322 11508 44334
rect 11452 44270 11454 44322
rect 11506 44270 11508 44322
rect 10108 44034 10164 44044
rect 9996 43698 10052 43708
rect 10220 43650 10276 43662
rect 10220 43598 10222 43650
rect 10274 43598 10276 43650
rect 10220 43540 10276 43598
rect 10668 43650 10724 43662
rect 10668 43598 10670 43650
rect 10722 43598 10724 43650
rect 10556 43540 10612 43550
rect 10220 43538 10612 43540
rect 10220 43486 10558 43538
rect 10610 43486 10612 43538
rect 10220 43484 10612 43486
rect 10332 43204 10388 43214
rect 9100 42690 9156 42700
rect 9436 42756 9492 42766
rect 10108 42756 10164 42766
rect 8316 42364 8484 42420
rect 8540 42530 8596 42542
rect 8540 42478 8542 42530
rect 8594 42478 8596 42530
rect 7308 41970 7588 41972
rect 7308 41918 7422 41970
rect 7474 41918 7588 41970
rect 7308 41916 7588 41918
rect 7644 42082 7700 42094
rect 7644 42030 7646 42082
rect 7698 42030 7700 42082
rect 5964 41748 6020 41758
rect 5292 41412 5348 41422
rect 2716 41010 2772 41020
rect 2940 41186 3444 41188
rect 2940 41134 3390 41186
rect 3442 41134 3444 41186
rect 2940 41132 3444 41134
rect 2604 40350 2606 40402
rect 2658 40350 2660 40402
rect 2044 40292 2100 40302
rect 2604 40292 2660 40350
rect 2940 40402 2996 41132
rect 3388 41122 3444 41132
rect 4508 41186 4900 41188
rect 4508 41134 4846 41186
rect 4898 41134 4900 41186
rect 4508 41132 4900 41134
rect 4060 41076 4116 41086
rect 4060 41074 4340 41076
rect 4060 41022 4062 41074
rect 4114 41022 4340 41074
rect 4060 41020 4340 41022
rect 4060 41010 4116 41020
rect 3500 40514 3556 40526
rect 3500 40462 3502 40514
rect 3554 40462 3556 40514
rect 2940 40350 2942 40402
rect 2994 40350 2996 40402
rect 2940 40338 2996 40350
rect 3276 40402 3332 40414
rect 3276 40350 3278 40402
rect 3330 40350 3332 40402
rect 2044 40290 2212 40292
rect 2044 40238 2046 40290
rect 2098 40238 2212 40290
rect 2044 40236 2212 40238
rect 2044 40226 2100 40236
rect 1708 39732 1764 39742
rect 1764 39676 1876 39732
rect 1708 39666 1764 39676
rect 1708 39394 1764 39406
rect 1708 39342 1710 39394
rect 1762 39342 1764 39394
rect 1708 39060 1764 39342
rect 1708 37492 1764 39004
rect 1820 38834 1876 39676
rect 2044 39060 2100 39070
rect 2044 38966 2100 39004
rect 1820 38782 1822 38834
rect 1874 38782 1876 38834
rect 1820 38162 1876 38782
rect 1820 38110 1822 38162
rect 1874 38110 1876 38162
rect 1820 38098 1876 38110
rect 2156 38164 2212 40236
rect 2604 40226 2660 40236
rect 3276 40292 3332 40350
rect 3276 40226 3332 40236
rect 2940 39844 2996 39854
rect 2268 39620 2324 39630
rect 2268 39526 2324 39564
rect 2940 39506 2996 39788
rect 2940 39454 2942 39506
rect 2994 39454 2996 39506
rect 2940 39442 2996 39454
rect 3052 39506 3108 39518
rect 3052 39454 3054 39506
rect 3106 39454 3108 39506
rect 2716 39396 2772 39406
rect 2604 39394 2772 39396
rect 2604 39342 2718 39394
rect 2770 39342 2772 39394
rect 2604 39340 2772 39342
rect 2156 38050 2212 38108
rect 2156 37998 2158 38050
rect 2210 37998 2212 38050
rect 2156 37986 2212 37998
rect 2268 38162 2324 38174
rect 2604 38164 2660 39340
rect 2716 39330 2772 39340
rect 3052 39284 3108 39454
rect 3500 39396 3556 40462
rect 3612 40404 3668 40414
rect 3612 40402 3780 40404
rect 3612 40350 3614 40402
rect 3666 40350 3780 40402
rect 3612 40348 3780 40350
rect 3612 40338 3668 40348
rect 3724 39620 3780 40348
rect 4060 40290 4116 40302
rect 4060 40238 4062 40290
rect 4114 40238 4116 40290
rect 4060 39844 4116 40238
rect 4060 39778 4116 39788
rect 3724 39554 3780 39564
rect 3836 39620 3892 39630
rect 3836 39618 4004 39620
rect 3836 39566 3838 39618
rect 3890 39566 4004 39618
rect 3836 39564 4004 39566
rect 3836 39554 3892 39564
rect 3500 39340 3780 39396
rect 2268 38110 2270 38162
rect 2322 38110 2324 38162
rect 2268 37716 2324 38110
rect 2492 38108 2660 38164
rect 2716 39172 2772 39182
rect 2716 39058 2772 39116
rect 2716 39006 2718 39058
rect 2770 39006 2772 39058
rect 2380 37828 2436 37838
rect 2380 37734 2436 37772
rect 2268 37650 2324 37660
rect 2268 37492 2324 37502
rect 1708 37490 2324 37492
rect 1708 37438 2270 37490
rect 2322 37438 2324 37490
rect 1708 37436 2324 37438
rect 2268 37426 2324 37436
rect 1820 37156 1876 37166
rect 1708 37154 1876 37156
rect 1708 37102 1822 37154
rect 1874 37102 1876 37154
rect 1708 37100 1876 37102
rect 1708 36370 1764 37100
rect 1820 37090 1876 37100
rect 2492 36484 2548 38108
rect 2716 37940 2772 39006
rect 3052 39058 3108 39228
rect 3052 39006 3054 39058
rect 3106 39006 3108 39058
rect 3052 38994 3108 39006
rect 3724 39060 3780 39340
rect 3724 38966 3780 39004
rect 3948 38836 4004 39564
rect 4284 39060 4340 41020
rect 4508 40626 4564 41132
rect 4844 41122 4900 41132
rect 5068 41300 5124 41310
rect 5068 41074 5124 41244
rect 5068 41022 5070 41074
rect 5122 41022 5124 41074
rect 4508 40574 4510 40626
rect 4562 40574 4564 40626
rect 4508 40562 4564 40574
rect 4956 40628 5012 40638
rect 5068 40628 5124 41022
rect 4956 40626 5124 40628
rect 4956 40574 4958 40626
rect 5010 40574 5124 40626
rect 4956 40572 5124 40574
rect 5292 40628 5348 41356
rect 5964 41188 6020 41692
rect 4956 40562 5012 40572
rect 5292 40534 5348 40572
rect 5516 41186 6020 41188
rect 5516 41134 5966 41186
rect 6018 41134 6020 41186
rect 5516 41132 6020 41134
rect 5516 40514 5572 41132
rect 5964 41122 6020 41132
rect 6412 41300 6468 41310
rect 6412 41186 6468 41244
rect 6412 41134 6414 41186
rect 6466 41134 6468 41186
rect 6412 41122 6468 41134
rect 6972 41188 7028 41198
rect 6972 41094 7028 41132
rect 7308 41186 7364 41916
rect 7420 41906 7476 41916
rect 7644 41748 7700 42030
rect 7644 41682 7700 41692
rect 8316 41188 8372 42364
rect 8540 42308 8596 42478
rect 8540 42242 8596 42252
rect 9212 42532 9268 42542
rect 8988 41972 9044 41982
rect 7308 41134 7310 41186
rect 7362 41134 7364 41186
rect 7308 41122 7364 41134
rect 7868 41186 8372 41188
rect 7868 41134 8318 41186
rect 8370 41134 8372 41186
rect 7868 41132 8372 41134
rect 7196 41076 7252 41086
rect 5516 40462 5518 40514
rect 5570 40462 5572 40514
rect 5516 40450 5572 40462
rect 5628 40962 5684 40974
rect 5628 40910 5630 40962
rect 5682 40910 5684 40962
rect 5068 40404 5124 40414
rect 4956 40402 5124 40404
rect 4956 40350 5070 40402
rect 5122 40350 5124 40402
rect 4956 40348 5124 40350
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 4396 39844 4452 39854
rect 4396 39618 4452 39788
rect 4396 39566 4398 39618
rect 4450 39566 4452 39618
rect 4396 39554 4452 39566
rect 4732 39732 4788 39742
rect 4732 39060 4788 39676
rect 4844 39508 4900 39518
rect 4844 39414 4900 39452
rect 4956 39060 5012 40348
rect 5068 40338 5124 40348
rect 5180 40290 5236 40302
rect 5180 40238 5182 40290
rect 5234 40238 5236 40290
rect 4172 39004 4676 39060
rect 4060 38836 4116 38846
rect 3948 38780 4060 38836
rect 4060 38770 4116 38780
rect 3500 38724 3556 38734
rect 4172 38668 4228 39004
rect 4620 38946 4676 39004
rect 4732 39058 4900 39060
rect 4732 39006 4734 39058
rect 4786 39006 4900 39058
rect 4732 39004 4900 39006
rect 4732 38994 4788 39004
rect 4620 38894 4622 38946
rect 4674 38894 4676 38946
rect 4620 38882 4676 38894
rect 4284 38836 4340 38846
rect 4284 38742 4340 38780
rect 3164 38612 3220 38622
rect 2828 38164 2884 38174
rect 2884 38108 3108 38164
rect 2828 38098 2884 38108
rect 2604 37884 2884 37940
rect 2604 37826 2660 37884
rect 2604 37774 2606 37826
rect 2658 37774 2660 37826
rect 2604 37762 2660 37774
rect 1708 36318 1710 36370
rect 1762 36318 1764 36370
rect 1708 35700 1764 36318
rect 2380 36428 2548 36484
rect 2716 37716 2772 37726
rect 2044 36258 2100 36270
rect 2044 36206 2046 36258
rect 2098 36206 2100 36258
rect 2044 36036 2100 36206
rect 2044 35970 2100 35980
rect 1708 35634 1764 35644
rect 2044 34356 2100 34366
rect 2044 34262 2100 34300
rect 1708 34130 1764 34142
rect 1708 34078 1710 34130
rect 1762 34078 1764 34130
rect 1708 33684 1764 34078
rect 1708 33618 1764 33628
rect 2380 33346 2436 36428
rect 2716 36370 2772 37660
rect 2828 37378 2884 37884
rect 2828 37326 2830 37378
rect 2882 37326 2884 37378
rect 2828 37314 2884 37326
rect 2940 37828 2996 37838
rect 2940 37378 2996 37772
rect 2940 37326 2942 37378
rect 2994 37326 2996 37378
rect 2940 37314 2996 37326
rect 3052 37378 3108 38108
rect 3052 37326 3054 37378
rect 3106 37326 3108 37378
rect 3052 37314 3108 37326
rect 3164 36596 3220 38556
rect 3388 38612 3556 38668
rect 3836 38612 4228 38668
rect 4844 38724 4900 39004
rect 4956 38994 5012 39004
rect 5068 40180 5124 40190
rect 5068 39618 5124 40124
rect 5180 39956 5236 40238
rect 5628 40180 5684 40910
rect 6636 40962 6692 40974
rect 6636 40910 6638 40962
rect 6690 40910 6692 40962
rect 5852 40628 5908 40638
rect 5852 40534 5908 40572
rect 5628 40114 5684 40124
rect 6188 40514 6244 40526
rect 6188 40462 6190 40514
rect 6242 40462 6244 40514
rect 6188 40068 6244 40462
rect 6188 40012 6468 40068
rect 5180 39900 6356 39956
rect 5740 39732 5796 39742
rect 5740 39638 5796 39676
rect 5068 39566 5070 39618
rect 5122 39566 5124 39618
rect 5068 38724 5124 39566
rect 5180 39620 5236 39630
rect 5516 39620 5572 39630
rect 5180 39618 5572 39620
rect 5180 39566 5182 39618
rect 5234 39566 5518 39618
rect 5570 39566 5572 39618
rect 5180 39564 5572 39566
rect 5180 39554 5236 39564
rect 5516 39554 5572 39564
rect 6300 39618 6356 39900
rect 6300 39566 6302 39618
rect 6354 39566 6356 39618
rect 6300 39554 6356 39566
rect 5852 39508 5908 39518
rect 5852 39060 5908 39452
rect 6412 39508 6468 40012
rect 6524 39732 6580 39742
rect 6524 39638 6580 39676
rect 6412 39442 6468 39452
rect 5852 39058 6020 39060
rect 5852 39006 5854 39058
rect 5906 39006 6020 39058
rect 5852 39004 6020 39006
rect 5852 38994 5908 39004
rect 3388 38050 3444 38612
rect 3388 37998 3390 38050
rect 3442 37998 3444 38050
rect 3388 37986 3444 37998
rect 3836 38050 3892 38612
rect 3836 37998 3838 38050
rect 3890 37998 3892 38050
rect 3836 37986 3892 37998
rect 3948 37938 4004 37950
rect 3948 37886 3950 37938
rect 4002 37886 4004 37938
rect 2828 36540 3220 36596
rect 3500 37042 3556 37054
rect 3500 36990 3502 37042
rect 3554 36990 3556 37042
rect 2828 36482 2884 36540
rect 2828 36430 2830 36482
rect 2882 36430 2884 36482
rect 2828 36418 2884 36430
rect 2716 36318 2718 36370
rect 2770 36318 2772 36370
rect 2492 36260 2548 36270
rect 2492 36258 2660 36260
rect 2492 36206 2494 36258
rect 2546 36206 2660 36258
rect 2492 36204 2660 36206
rect 2492 36194 2548 36204
rect 2492 35812 2548 35822
rect 2492 35718 2548 35756
rect 2604 35698 2660 36204
rect 2604 35646 2606 35698
rect 2658 35646 2660 35698
rect 2604 35634 2660 35646
rect 2716 34804 2772 36318
rect 3052 34914 3108 36540
rect 3500 36482 3556 36990
rect 3836 37042 3892 37054
rect 3836 36990 3838 37042
rect 3890 36990 3892 37042
rect 3836 36594 3892 36990
rect 3836 36542 3838 36594
rect 3890 36542 3892 36594
rect 3836 36530 3892 36542
rect 3500 36430 3502 36482
rect 3554 36430 3556 36482
rect 3500 36418 3556 36430
rect 3948 35924 4004 37886
rect 4172 37266 4228 38612
rect 4732 38612 4788 38622
rect 4732 38518 4788 38556
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 4844 38276 4900 38668
rect 4620 38220 4900 38276
rect 4956 38612 5124 38668
rect 5740 38834 5796 38846
rect 5740 38782 5742 38834
rect 5794 38782 5796 38834
rect 5740 38724 5796 38782
rect 5740 38658 5796 38668
rect 5852 38836 5908 38846
rect 4172 37214 4174 37266
rect 4226 37214 4228 37266
rect 4172 37202 4228 37214
rect 4396 37268 4452 37278
rect 4620 37268 4676 38220
rect 4732 38052 4788 38062
rect 4956 38052 5012 38612
rect 4732 38050 5012 38052
rect 4732 37998 4734 38050
rect 4786 37998 5012 38050
rect 4732 37996 5012 37998
rect 4732 37986 4788 37996
rect 5068 37940 5124 37950
rect 5068 37846 5124 37884
rect 4396 37266 4676 37268
rect 4396 37214 4398 37266
rect 4450 37214 4676 37266
rect 4396 37212 4676 37214
rect 4396 37202 4452 37212
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4396 36596 4452 36606
rect 4396 36594 4788 36596
rect 4396 36542 4398 36594
rect 4450 36542 4788 36594
rect 4396 36540 4788 36542
rect 4396 36530 4452 36540
rect 4172 36484 4228 36494
rect 3948 35858 4004 35868
rect 4060 36482 4228 36484
rect 4060 36430 4174 36482
rect 4226 36430 4228 36482
rect 4060 36428 4228 36430
rect 3164 35700 3220 35710
rect 3164 35138 3220 35644
rect 3164 35086 3166 35138
rect 3218 35086 3220 35138
rect 3164 35074 3220 35086
rect 3612 35698 3668 35710
rect 3612 35646 3614 35698
rect 3666 35646 3668 35698
rect 3052 34862 3054 34914
rect 3106 34862 3108 34914
rect 3052 34850 3108 34862
rect 2828 34804 2884 34814
rect 2716 34802 2884 34804
rect 2716 34750 2830 34802
rect 2882 34750 2884 34802
rect 2716 34748 2884 34750
rect 2828 34738 2884 34748
rect 3276 34802 3332 34814
rect 3276 34750 3278 34802
rect 3330 34750 3332 34802
rect 3276 34356 3332 34750
rect 3612 34356 3668 35646
rect 3276 34300 3668 34356
rect 2492 34018 2548 34030
rect 2492 33966 2494 34018
rect 2546 33966 2548 34018
rect 2492 33684 2548 33966
rect 2492 33618 2548 33628
rect 2380 33294 2382 33346
rect 2434 33294 2436 33346
rect 2380 32674 2436 33294
rect 2716 33346 2772 33358
rect 2716 33294 2718 33346
rect 2770 33294 2772 33346
rect 2716 33124 2772 33294
rect 2380 32622 2382 32674
rect 2434 32622 2436 32674
rect 2380 32610 2436 32622
rect 2604 33068 2716 33124
rect 2604 32562 2660 33068
rect 2716 33058 2772 33068
rect 3276 33124 3332 33134
rect 2604 32510 2606 32562
rect 2658 32510 2660 32562
rect 2604 32498 2660 32510
rect 3276 31778 3332 33068
rect 3612 32786 3668 34300
rect 4060 33570 4116 36428
rect 4172 36418 4228 36428
rect 4732 35924 4788 36540
rect 4732 35922 4900 35924
rect 4732 35870 4734 35922
rect 4786 35870 4900 35922
rect 4732 35868 4900 35870
rect 4732 35858 4788 35868
rect 4396 35700 4452 35710
rect 4396 35606 4452 35644
rect 4172 35588 4228 35598
rect 4172 35586 4340 35588
rect 4172 35534 4174 35586
rect 4226 35534 4340 35586
rect 4172 35532 4340 35534
rect 4172 35522 4228 35532
rect 4172 35364 4228 35374
rect 4172 34916 4228 35308
rect 4284 35028 4340 35532
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4844 35140 4900 35868
rect 4956 35812 5012 35850
rect 4956 35746 5012 35756
rect 4732 35084 4900 35140
rect 4956 35586 5012 35598
rect 4956 35534 4958 35586
rect 5010 35534 5012 35586
rect 4508 35028 4564 35038
rect 4284 35026 4564 35028
rect 4284 34974 4510 35026
rect 4562 34974 4564 35026
rect 4284 34972 4564 34974
rect 4172 34914 4452 34916
rect 4172 34862 4174 34914
rect 4226 34862 4452 34914
rect 4172 34860 4452 34862
rect 4172 34850 4228 34860
rect 4060 33518 4062 33570
rect 4114 33518 4116 33570
rect 4060 33506 4116 33518
rect 4172 34242 4228 34254
rect 4172 34190 4174 34242
rect 4226 34190 4228 34242
rect 3612 32734 3614 32786
rect 3666 32734 3668 32786
rect 3612 32722 3668 32734
rect 3724 33460 3780 33470
rect 3724 33346 3780 33404
rect 3724 33294 3726 33346
rect 3778 33294 3780 33346
rect 3724 32674 3780 33294
rect 3724 32622 3726 32674
rect 3778 32622 3780 32674
rect 3724 32564 3780 32622
rect 3276 31726 3278 31778
rect 3330 31726 3332 31778
rect 3276 31714 3332 31726
rect 3612 32508 3780 32564
rect 3612 31778 3668 32508
rect 4172 32116 4228 34190
rect 4396 34130 4452 34860
rect 4396 34078 4398 34130
rect 4450 34078 4452 34130
rect 4396 34066 4452 34078
rect 4508 34018 4564 34972
rect 4508 33966 4510 34018
rect 4562 33966 4564 34018
rect 4508 33954 4564 33966
rect 4732 33908 4788 35084
rect 4956 34132 5012 35534
rect 5068 34916 5124 34926
rect 5068 34822 5124 34860
rect 5068 34132 5124 34142
rect 4956 34130 5124 34132
rect 4956 34078 5070 34130
rect 5122 34078 5124 34130
rect 4956 34076 5124 34078
rect 5068 34066 5124 34076
rect 5852 34132 5908 38780
rect 5964 37492 6020 39004
rect 6412 38948 6468 38958
rect 6300 38946 6468 38948
rect 6300 38894 6414 38946
rect 6466 38894 6468 38946
rect 6300 38892 6468 38894
rect 6076 38834 6132 38846
rect 6076 38782 6078 38834
rect 6130 38782 6132 38834
rect 6076 38162 6132 38782
rect 6076 38110 6078 38162
rect 6130 38110 6132 38162
rect 6076 38098 6132 38110
rect 6076 37492 6132 37502
rect 5964 37490 6132 37492
rect 5964 37438 6078 37490
rect 6130 37438 6132 37490
rect 5964 37436 6132 37438
rect 6076 37426 6132 37436
rect 6076 35812 6132 35822
rect 6076 35718 6132 35756
rect 6188 34802 6244 34814
rect 6188 34750 6190 34802
rect 6242 34750 6244 34802
rect 6188 34356 6244 34750
rect 5852 34130 6132 34132
rect 5852 34078 5854 34130
rect 5906 34078 6132 34130
rect 5852 34076 6132 34078
rect 5852 34066 5908 34076
rect 4732 33852 4900 33908
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4172 32060 4340 32116
rect 4476 32106 4740 32116
rect 4172 31892 4228 31902
rect 4060 31890 4228 31892
rect 4060 31838 4174 31890
rect 4226 31838 4228 31890
rect 4060 31836 4228 31838
rect 3612 31726 3614 31778
rect 3666 31726 3668 31778
rect 3612 31714 3668 31726
rect 3724 31780 3780 31790
rect 3948 31780 4004 31790
rect 3724 31778 4004 31780
rect 3724 31726 3726 31778
rect 3778 31726 3950 31778
rect 4002 31726 4004 31778
rect 3724 31724 4004 31726
rect 3724 31714 3780 31724
rect 3948 31714 4004 31724
rect 2716 31556 2772 31566
rect 2716 31218 2772 31500
rect 2716 31166 2718 31218
rect 2770 31166 2772 31218
rect 2716 31154 2772 31166
rect 3164 31556 3220 31566
rect 2828 31108 2884 31118
rect 2828 31014 2884 31052
rect 2492 30994 2548 31006
rect 2492 30942 2494 30994
rect 2546 30942 2548 30994
rect 2380 30324 2436 30334
rect 2380 30098 2436 30268
rect 2492 30210 2548 30942
rect 2492 30158 2494 30210
rect 2546 30158 2548 30210
rect 2492 30146 2548 30158
rect 2380 30046 2382 30098
rect 2434 30046 2436 30098
rect 2380 30034 2436 30046
rect 3164 29538 3220 31500
rect 3724 31556 3780 31566
rect 3724 31332 3780 31500
rect 4060 31332 4116 31836
rect 4172 31826 4228 31836
rect 4284 31780 4340 32060
rect 4508 31892 4564 31902
rect 4284 31724 4452 31780
rect 3724 31276 4116 31332
rect 4172 31668 4228 31678
rect 3164 29486 3166 29538
rect 3218 29486 3220 29538
rect 3164 29474 3220 29486
rect 3276 31108 3332 31118
rect 3276 29538 3332 31052
rect 3500 30996 3556 31006
rect 3500 30212 3556 30940
rect 3724 30994 3780 31276
rect 4172 31108 4228 31612
rect 4284 31554 4340 31566
rect 4284 31502 4286 31554
rect 4338 31502 4340 31554
rect 4284 31220 4340 31502
rect 4284 31154 4340 31164
rect 3724 30942 3726 30994
rect 3778 30942 3780 30994
rect 3724 30930 3780 30942
rect 4060 30996 4116 31006
rect 4172 30996 4228 31052
rect 4060 30994 4228 30996
rect 4060 30942 4062 30994
rect 4114 30942 4228 30994
rect 4060 30940 4228 30942
rect 4284 30994 4340 31006
rect 4284 30942 4286 30994
rect 4338 30942 4340 30994
rect 4060 30930 4116 30940
rect 3836 30882 3892 30894
rect 4284 30884 4340 30942
rect 3836 30830 3838 30882
rect 3890 30830 3892 30882
rect 3836 30436 3892 30830
rect 4172 30828 4340 30884
rect 4172 30772 4228 30828
rect 4396 30772 4452 31724
rect 4508 31666 4564 31836
rect 4844 31780 4900 33852
rect 4844 31714 4900 31724
rect 5068 33684 5124 33694
rect 5068 31892 5124 33628
rect 5964 33460 6020 33498
rect 5964 33394 6020 33404
rect 5964 33234 6020 33246
rect 5964 33182 5966 33234
rect 6018 33182 6020 33234
rect 5964 33012 6020 33182
rect 5964 32946 6020 32956
rect 6076 32674 6132 34076
rect 6188 33796 6244 34300
rect 6300 34018 6356 38892
rect 6412 38882 6468 38892
rect 6524 38948 6580 38958
rect 6636 38948 6692 40910
rect 7084 40514 7140 40526
rect 7084 40462 7086 40514
rect 7138 40462 7140 40514
rect 7084 39732 7140 40462
rect 7196 40516 7252 41020
rect 7868 40740 7924 41132
rect 8316 41122 8372 41132
rect 8876 41300 8932 41310
rect 8876 41186 8932 41244
rect 8876 41134 8878 41186
rect 8930 41134 8932 41186
rect 8876 41122 8932 41134
rect 8988 41186 9044 41916
rect 8988 41134 8990 41186
rect 9042 41134 9044 41186
rect 8988 41122 9044 41134
rect 9212 41074 9268 42476
rect 9436 41186 9492 42700
rect 9772 42700 10108 42756
rect 9772 42194 9828 42700
rect 10108 42662 10164 42700
rect 9772 42142 9774 42194
rect 9826 42142 9828 42194
rect 9772 42130 9828 42142
rect 10332 42532 10388 43148
rect 10444 42644 10500 43484
rect 10556 43474 10612 43484
rect 10668 43204 10724 43598
rect 11340 43652 11396 43662
rect 11340 43538 11396 43596
rect 11340 43486 11342 43538
rect 11394 43486 11396 43538
rect 11340 43474 11396 43486
rect 11340 43316 11396 43326
rect 11452 43316 11508 44270
rect 11788 44212 11844 44222
rect 11900 44212 11956 44830
rect 12124 44436 12180 44474
rect 12124 44370 12180 44380
rect 12460 44322 12516 44940
rect 12460 44270 12462 44322
rect 12514 44270 12516 44322
rect 12460 44258 12516 44270
rect 11788 44210 11956 44212
rect 11788 44158 11790 44210
rect 11842 44158 11956 44210
rect 11788 44156 11956 44158
rect 12124 44212 12180 44222
rect 11788 44146 11844 44156
rect 12124 44118 12180 44156
rect 12684 44100 12740 45054
rect 13356 45106 13412 45118
rect 13356 45054 13358 45106
rect 13410 45054 13412 45106
rect 13356 44996 13412 45054
rect 13804 44996 13860 45006
rect 13356 44994 13860 44996
rect 13356 44942 13806 44994
rect 13858 44942 13860 44994
rect 13356 44940 13860 44942
rect 13804 44660 13860 44940
rect 13804 44594 13860 44604
rect 12124 43652 12180 43662
rect 11788 43540 11844 43550
rect 11340 43314 11508 43316
rect 11340 43262 11342 43314
rect 11394 43262 11508 43314
rect 11340 43260 11508 43262
rect 11676 43538 11844 43540
rect 11676 43486 11790 43538
rect 11842 43486 11844 43538
rect 11676 43484 11844 43486
rect 11340 43250 11396 43260
rect 10668 43138 10724 43148
rect 11452 42868 11508 42878
rect 10780 42812 11172 42868
rect 10556 42756 10612 42766
rect 10780 42756 10836 42812
rect 10556 42754 10836 42756
rect 10556 42702 10558 42754
rect 10610 42702 10836 42754
rect 10556 42700 10836 42702
rect 10556 42690 10612 42700
rect 10444 42578 10500 42588
rect 10332 42196 10388 42476
rect 10556 42196 10612 42206
rect 10332 42194 10612 42196
rect 10332 42142 10558 42194
rect 10610 42142 10612 42194
rect 10332 42140 10612 42142
rect 9548 41970 9604 41982
rect 9548 41918 9550 41970
rect 9602 41918 9604 41970
rect 9548 41300 9604 41918
rect 9996 41972 10052 41982
rect 9996 41878 10052 41916
rect 10220 41972 10276 41982
rect 10332 41972 10388 42140
rect 10556 42130 10612 42140
rect 10220 41970 10388 41972
rect 10220 41918 10222 41970
rect 10274 41918 10388 41970
rect 10220 41916 10388 41918
rect 10220 41906 10276 41916
rect 9884 41858 9940 41870
rect 9884 41806 9886 41858
rect 9938 41806 9940 41858
rect 9884 41524 9940 41806
rect 9884 41468 10388 41524
rect 10332 41410 10388 41468
rect 10332 41358 10334 41410
rect 10386 41358 10388 41410
rect 10332 41346 10388 41358
rect 9548 41234 9604 41244
rect 10668 41300 10724 41310
rect 10668 41206 10724 41244
rect 9436 41134 9438 41186
rect 9490 41134 9492 41186
rect 9436 41122 9492 41134
rect 9212 41022 9214 41074
rect 9266 41022 9268 41074
rect 9212 41010 9268 41022
rect 9772 41076 9828 41086
rect 10108 41076 10164 41086
rect 9772 41074 10164 41076
rect 9772 41022 9774 41074
rect 9826 41022 10110 41074
rect 10162 41022 10164 41074
rect 9772 41020 10164 41022
rect 9772 41010 9828 41020
rect 7980 40964 8036 40974
rect 8036 40908 8260 40964
rect 7980 40870 8036 40908
rect 7868 40684 8036 40740
rect 7196 40404 7252 40460
rect 7868 40516 7924 40526
rect 7868 40422 7924 40460
rect 7980 40514 8036 40684
rect 7980 40462 7982 40514
rect 8034 40462 8036 40514
rect 7980 40450 8036 40462
rect 7308 40404 7364 40414
rect 7196 40402 7364 40404
rect 7196 40350 7310 40402
rect 7362 40350 7364 40402
rect 7196 40348 7364 40350
rect 7308 40338 7364 40348
rect 7644 40402 7700 40414
rect 7644 40350 7646 40402
rect 7698 40350 7700 40402
rect 7644 39732 7700 40350
rect 7084 39676 7364 39732
rect 6524 38946 6692 38948
rect 6524 38894 6526 38946
rect 6578 38894 6692 38946
rect 6524 38892 6692 38894
rect 6524 38882 6580 38892
rect 6412 38610 6468 38622
rect 6412 38558 6414 38610
rect 6466 38558 6468 38610
rect 6412 37938 6468 38558
rect 6412 37886 6414 37938
rect 6466 37886 6468 37938
rect 6412 37874 6468 37886
rect 6524 37716 6580 37726
rect 6412 37378 6468 37390
rect 6412 37326 6414 37378
rect 6466 37326 6468 37378
rect 6412 36372 6468 37326
rect 6412 36306 6468 36316
rect 6412 35700 6468 35710
rect 6524 35700 6580 37660
rect 6636 37044 6692 38892
rect 6860 39508 6916 39518
rect 7084 39508 7140 39518
rect 6860 38946 6916 39452
rect 6972 39452 7084 39508
rect 6972 39058 7028 39452
rect 7084 39442 7140 39452
rect 6972 39006 6974 39058
rect 7026 39006 7028 39058
rect 6972 38994 7028 39006
rect 7308 39284 7364 39676
rect 6860 38894 6862 38946
rect 6914 38894 6916 38946
rect 6860 38882 6916 38894
rect 6748 38724 6804 38734
rect 6748 37490 6804 38668
rect 7308 38668 7364 39228
rect 6972 38612 7028 38622
rect 7308 38612 7588 38668
rect 6748 37438 6750 37490
rect 6802 37438 6804 37490
rect 6748 37426 6804 37438
rect 6860 38610 7028 38612
rect 6860 38558 6974 38610
rect 7026 38558 7028 38610
rect 6860 38556 7028 38558
rect 6636 36988 6804 37044
rect 6412 35698 6580 35700
rect 6412 35646 6414 35698
rect 6466 35646 6580 35698
rect 6412 35644 6580 35646
rect 6636 36036 6692 36046
rect 6636 35698 6692 35980
rect 6636 35646 6638 35698
rect 6690 35646 6692 35698
rect 6412 35634 6468 35644
rect 6636 35634 6692 35646
rect 6524 34692 6580 34702
rect 6524 34690 6692 34692
rect 6524 34638 6526 34690
rect 6578 34638 6692 34690
rect 6524 34636 6692 34638
rect 6524 34626 6580 34636
rect 6300 33966 6302 34018
rect 6354 33966 6356 34018
rect 6300 33908 6356 33966
rect 6300 33852 6580 33908
rect 6188 33740 6356 33796
rect 6188 33124 6244 33134
rect 6188 32786 6244 33068
rect 6188 32734 6190 32786
rect 6242 32734 6244 32786
rect 6188 32722 6244 32734
rect 6076 32622 6078 32674
rect 6130 32622 6132 32674
rect 6076 32610 6132 32622
rect 5068 31778 5124 31836
rect 5068 31726 5070 31778
rect 5122 31726 5124 31778
rect 5068 31714 5124 31726
rect 5964 32564 6020 32574
rect 4508 31614 4510 31666
rect 4562 31614 4564 31666
rect 4508 31602 4564 31614
rect 4732 31556 4788 31566
rect 4732 31554 4900 31556
rect 4732 31502 4734 31554
rect 4786 31502 4900 31554
rect 4732 31500 4900 31502
rect 4732 31490 4788 31500
rect 4620 31108 4676 31118
rect 4620 31014 4676 31052
rect 4172 30706 4228 30716
rect 4284 30716 4452 30772
rect 4284 30436 4340 30716
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4508 30436 4564 30446
rect 4284 30380 4452 30436
rect 3836 30370 3892 30380
rect 4284 30212 4340 30222
rect 3276 29486 3278 29538
rect 3330 29486 3332 29538
rect 3276 29474 3332 29486
rect 3388 30210 3556 30212
rect 3388 30158 3502 30210
rect 3554 30158 3556 30210
rect 3388 30156 3556 30158
rect 3388 29538 3444 30156
rect 3500 30146 3556 30156
rect 3836 30210 4340 30212
rect 3836 30158 4286 30210
rect 4338 30158 4340 30210
rect 3836 30156 4340 30158
rect 3388 29486 3390 29538
rect 3442 29486 3444 29538
rect 3388 29474 3444 29486
rect 3612 29986 3668 29998
rect 3612 29934 3614 29986
rect 3666 29934 3668 29986
rect 3612 29428 3668 29934
rect 3836 29650 3892 30156
rect 4284 30146 4340 30156
rect 3836 29598 3838 29650
rect 3890 29598 3892 29650
rect 3836 29586 3892 29598
rect 4396 29540 4452 30380
rect 4508 30342 4564 30380
rect 4732 30436 4788 30446
rect 4844 30436 4900 31500
rect 4956 31554 5012 31566
rect 4956 31502 4958 31554
rect 5010 31502 5012 31554
rect 4956 31444 5012 31502
rect 5964 31556 6020 32508
rect 6300 32562 6356 33740
rect 6412 33348 6468 33358
rect 6412 33254 6468 33292
rect 6412 33012 6468 33022
rect 6524 33012 6580 33852
rect 6468 32956 6580 33012
rect 6636 33012 6692 34636
rect 6748 34356 6804 36988
rect 6860 35588 6916 38556
rect 6972 38546 7028 38556
rect 7084 37716 7140 37726
rect 7084 37490 7140 37660
rect 7084 37438 7086 37490
rect 7138 37438 7140 37490
rect 7084 37426 7140 37438
rect 7420 36484 7476 36494
rect 7420 36390 7476 36428
rect 7084 36258 7140 36270
rect 7084 36206 7086 36258
rect 7138 36206 7140 36258
rect 6860 35522 6916 35532
rect 6972 36036 7028 36046
rect 6972 34916 7028 35980
rect 7084 35812 7140 36206
rect 7308 36258 7364 36270
rect 7308 36206 7310 36258
rect 7362 36206 7364 36258
rect 7308 36036 7364 36206
rect 7308 35970 7364 35980
rect 7084 35746 7140 35756
rect 7420 35924 7476 35934
rect 7308 35700 7364 35710
rect 7308 35606 7364 35644
rect 7196 35588 7252 35598
rect 7084 34916 7140 34926
rect 6972 34914 7140 34916
rect 6972 34862 7086 34914
rect 7138 34862 7140 34914
rect 6972 34860 7140 34862
rect 7084 34850 7140 34860
rect 6860 34804 6916 34842
rect 6860 34738 6916 34748
rect 7196 34692 7252 35532
rect 7420 35588 7476 35868
rect 7420 35494 7476 35532
rect 7420 34692 7476 34702
rect 6972 34636 7252 34692
rect 7308 34636 7420 34692
rect 6860 34356 6916 34366
rect 6748 34354 6916 34356
rect 6748 34302 6862 34354
rect 6914 34302 6916 34354
rect 6748 34300 6916 34302
rect 6860 33348 6916 34300
rect 6860 33282 6916 33292
rect 6972 33348 7028 34636
rect 7196 34356 7252 34366
rect 7308 34356 7364 34636
rect 7420 34626 7476 34636
rect 7196 34354 7364 34356
rect 7196 34302 7198 34354
rect 7250 34302 7364 34354
rect 7196 34300 7364 34302
rect 7196 33684 7252 34300
rect 7196 33618 7252 33628
rect 7532 33572 7588 38612
rect 7644 38050 7700 39676
rect 8204 39620 8260 40908
rect 9772 40628 9828 40638
rect 8652 39620 8708 39630
rect 8204 39564 8484 39620
rect 8316 39396 8372 39406
rect 8316 39302 8372 39340
rect 8428 39060 8484 39564
rect 8652 39526 8708 39564
rect 9660 39620 9716 39630
rect 9660 39526 9716 39564
rect 8988 39396 9044 39406
rect 8764 39284 8820 39294
rect 8764 39060 8820 39228
rect 8316 39058 8484 39060
rect 8316 39006 8430 39058
rect 8482 39006 8484 39058
rect 8316 39004 8484 39006
rect 8316 38668 8372 39004
rect 8428 38994 8484 39004
rect 8540 39058 8820 39060
rect 8540 39006 8766 39058
rect 8818 39006 8820 39058
rect 8540 39004 8820 39006
rect 7644 37998 7646 38050
rect 7698 37998 7700 38050
rect 7644 37986 7700 37998
rect 7980 38612 8372 38668
rect 8540 38668 8596 39004
rect 8764 38994 8820 39004
rect 8988 38668 9044 39340
rect 8540 38612 8820 38668
rect 8988 38612 9604 38668
rect 7980 36484 8036 38612
rect 8764 38388 8820 38612
rect 8764 38332 9044 38388
rect 8876 38162 8932 38174
rect 8876 38110 8878 38162
rect 8930 38110 8932 38162
rect 8204 38052 8260 38062
rect 8764 38052 8820 38062
rect 8204 38050 8820 38052
rect 8204 37998 8206 38050
rect 8258 37998 8766 38050
rect 8818 37998 8820 38050
rect 8204 37996 8820 37998
rect 8204 37986 8260 37996
rect 8540 37490 8596 37996
rect 8764 37986 8820 37996
rect 8540 37438 8542 37490
rect 8594 37438 8596 37490
rect 8540 37426 8596 37438
rect 8764 37380 8820 37390
rect 8876 37380 8932 38110
rect 8764 37378 8932 37380
rect 8764 37326 8766 37378
rect 8818 37326 8878 37378
rect 8930 37326 8932 37378
rect 8764 37324 8932 37326
rect 8764 37314 8820 37324
rect 8876 37286 8932 37324
rect 8652 37154 8708 37166
rect 8652 37102 8654 37154
rect 8706 37102 8708 37154
rect 8652 36708 8708 37102
rect 8652 36652 8820 36708
rect 7980 36418 8036 36428
rect 8316 36482 8372 36494
rect 8316 36430 8318 36482
rect 8370 36430 8372 36482
rect 8204 35812 8260 35822
rect 8204 35718 8260 35756
rect 8092 34356 8148 34366
rect 8316 34356 8372 36430
rect 8652 36482 8708 36494
rect 8652 36430 8654 36482
rect 8706 36430 8708 36482
rect 8652 35812 8708 36430
rect 8428 35756 8652 35812
rect 8428 35026 8484 35756
rect 8652 35746 8708 35756
rect 8764 36370 8820 36652
rect 8764 36318 8766 36370
rect 8818 36318 8820 36370
rect 8428 34974 8430 35026
rect 8482 34974 8484 35026
rect 8428 34962 8484 34974
rect 8540 35588 8596 35598
rect 8092 34354 8372 34356
rect 8092 34302 8094 34354
rect 8146 34302 8372 34354
rect 8092 34300 8372 34302
rect 8092 34290 8148 34300
rect 8540 34242 8596 35532
rect 8764 34914 8820 36318
rect 8876 36594 8932 36606
rect 8876 36542 8878 36594
rect 8930 36542 8932 36594
rect 8876 35476 8932 36542
rect 8876 35410 8932 35420
rect 8764 34862 8766 34914
rect 8818 34862 8820 34914
rect 8764 34850 8820 34862
rect 8988 34692 9044 38332
rect 9100 37380 9156 37390
rect 9100 37378 9492 37380
rect 9100 37326 9102 37378
rect 9154 37326 9492 37378
rect 9100 37324 9492 37326
rect 9100 37314 9156 37324
rect 9436 36482 9492 37324
rect 9436 36430 9438 36482
rect 9490 36430 9492 36482
rect 9436 36418 9492 36430
rect 9548 35308 9604 38612
rect 9660 38052 9716 38062
rect 9660 37958 9716 37996
rect 9772 37434 9828 40572
rect 10108 40516 10164 41020
rect 10668 40628 10724 40638
rect 10780 40628 10836 42700
rect 11116 42754 11172 42812
rect 11452 42774 11508 42812
rect 11116 42702 11118 42754
rect 11170 42702 11172 42754
rect 11116 42690 11172 42702
rect 11676 42756 11732 43484
rect 11788 43474 11844 43484
rect 11676 42690 11732 42700
rect 12124 42754 12180 43596
rect 12684 43652 12740 44044
rect 13244 44436 13300 44446
rect 13244 43762 13300 44380
rect 13804 44324 13860 44334
rect 13916 44324 13972 45166
rect 14140 45220 14196 45230
rect 14140 45126 14196 45164
rect 14252 44884 14308 45612
rect 15036 45666 15092 45678
rect 15036 45614 15038 45666
rect 15090 45614 15092 45666
rect 14364 45332 14420 45342
rect 14364 45106 14420 45276
rect 14812 45332 14868 45342
rect 14812 45238 14868 45276
rect 14364 45054 14366 45106
rect 14418 45054 14420 45106
rect 14364 45042 14420 45054
rect 14252 44818 14308 44828
rect 13804 44322 13972 44324
rect 13804 44270 13806 44322
rect 13858 44270 13972 44322
rect 13804 44268 13972 44270
rect 14924 44324 14980 44334
rect 15036 44324 15092 45614
rect 15372 45106 15428 45726
rect 20748 45778 20804 45790
rect 20748 45726 20750 45778
rect 20802 45726 20804 45778
rect 17388 45666 17444 45678
rect 17388 45614 17390 45666
rect 17442 45614 17444 45666
rect 16828 45444 16884 45454
rect 16268 45332 16324 45342
rect 15372 45054 15374 45106
rect 15426 45054 15428 45106
rect 15372 44436 15428 45054
rect 15596 45108 15652 45118
rect 15596 45014 15652 45052
rect 15708 44996 15764 45006
rect 15708 44902 15764 44940
rect 15596 44772 15652 44782
rect 15372 44370 15428 44380
rect 15484 44716 15596 44772
rect 14980 44268 15092 44324
rect 15484 44324 15540 44716
rect 15596 44706 15652 44716
rect 16268 44546 16324 45276
rect 16604 45220 16660 45230
rect 16604 45126 16660 45164
rect 16828 45106 16884 45388
rect 16828 45054 16830 45106
rect 16882 45054 16884 45106
rect 16492 44884 16548 44894
rect 16492 44790 16548 44828
rect 16268 44494 16270 44546
rect 16322 44494 16324 44546
rect 16268 44482 16324 44494
rect 16828 44548 16884 45054
rect 16828 44482 16884 44492
rect 13804 44258 13860 44268
rect 13244 43710 13246 43762
rect 13298 43710 13300 43762
rect 13244 43698 13300 43710
rect 13356 44212 13412 44222
rect 13356 43708 13412 44156
rect 13468 44100 13524 44110
rect 13468 44006 13524 44044
rect 13468 43764 13524 43774
rect 14924 43708 14980 44268
rect 15260 44210 15316 44222
rect 15260 44158 15262 44210
rect 15314 44158 15316 44210
rect 13356 43652 13524 43708
rect 14364 43652 14420 43662
rect 12684 43586 12740 43596
rect 12796 43538 12852 43550
rect 12796 43486 12798 43538
rect 12850 43486 12852 43538
rect 12796 43428 12852 43486
rect 13468 43538 13524 43652
rect 13468 43486 13470 43538
rect 13522 43486 13524 43538
rect 13468 43474 13524 43486
rect 13916 43650 14420 43652
rect 13916 43598 14366 43650
rect 14418 43598 14420 43650
rect 13916 43596 14420 43598
rect 12796 43362 12852 43372
rect 13356 43426 13412 43438
rect 13356 43374 13358 43426
rect 13410 43374 13412 43426
rect 12124 42702 12126 42754
rect 12178 42702 12180 42754
rect 12124 42690 12180 42702
rect 10892 42644 10948 42654
rect 10892 42550 10948 42588
rect 11340 42530 11396 42542
rect 11340 42478 11342 42530
rect 11394 42478 11396 42530
rect 11340 42420 11396 42478
rect 10108 40450 10164 40460
rect 10220 40572 10612 40628
rect 10220 40290 10276 40572
rect 10220 40238 10222 40290
rect 10274 40238 10276 40290
rect 10220 40226 10276 40238
rect 10332 40404 10388 40414
rect 10332 40068 10388 40348
rect 10556 40180 10612 40572
rect 10668 40626 10836 40628
rect 10668 40574 10670 40626
rect 10722 40574 10836 40626
rect 10668 40572 10836 40574
rect 10668 40562 10724 40572
rect 10556 40124 10724 40180
rect 10220 40012 10388 40068
rect 9660 37380 9716 37418
rect 9772 37382 9774 37434
rect 9826 37382 9828 37434
rect 9772 37370 9828 37382
rect 9884 39172 9940 39182
rect 9884 38836 9940 39116
rect 10108 38946 10164 38958
rect 10108 38894 10110 38946
rect 10162 38894 10164 38946
rect 10108 38836 10164 38894
rect 10220 38946 10276 40012
rect 10220 38894 10222 38946
rect 10274 38894 10276 38946
rect 10220 38882 10276 38894
rect 10556 39396 10612 39406
rect 10556 38946 10612 39340
rect 10556 38894 10558 38946
rect 10610 38894 10612 38946
rect 10556 38882 10612 38894
rect 9884 38780 10164 38836
rect 9660 37314 9716 37324
rect 9772 37156 9828 37166
rect 9660 37044 9716 37054
rect 9660 36950 9716 36988
rect 9772 36596 9828 37100
rect 8540 34190 8542 34242
rect 8594 34190 8596 34242
rect 8540 34178 8596 34190
rect 8652 34636 9044 34692
rect 9100 35252 9156 35262
rect 9100 34804 9156 35196
rect 9436 35252 9604 35308
rect 9660 36540 9828 36596
rect 9660 36370 9716 36540
rect 9660 36318 9662 36370
rect 9714 36318 9716 36370
rect 9660 35252 9716 36318
rect 9772 36370 9828 36382
rect 9772 36318 9774 36370
rect 9826 36318 9828 36370
rect 9772 36260 9828 36318
rect 9772 36194 9828 36204
rect 9212 35140 9268 35150
rect 9212 35026 9268 35084
rect 9212 34974 9214 35026
rect 9266 34974 9268 35026
rect 9212 34962 9268 34974
rect 8652 34242 8708 34636
rect 8652 34190 8654 34242
rect 8706 34190 8708 34242
rect 8652 34020 8708 34190
rect 8988 34356 9044 34366
rect 8652 33954 8708 33964
rect 8764 34130 8820 34142
rect 8764 34078 8766 34130
rect 8818 34078 8820 34130
rect 7532 33516 8148 33572
rect 7980 33348 8036 33358
rect 6972 33346 7812 33348
rect 6972 33294 6974 33346
rect 7026 33294 7812 33346
rect 6972 33292 7812 33294
rect 6972 33282 7028 33292
rect 7308 33124 7364 33134
rect 7308 33030 7364 33068
rect 7420 33122 7476 33134
rect 7420 33070 7422 33122
rect 7474 33070 7476 33122
rect 6636 32956 6916 33012
rect 6412 32946 6468 32956
rect 6860 32788 6916 32956
rect 7420 32788 7476 33070
rect 7532 33124 7588 33134
rect 7532 33030 7588 33068
rect 6748 32564 6804 32574
rect 6300 32510 6302 32562
rect 6354 32510 6356 32562
rect 6300 32498 6356 32510
rect 6636 32562 6804 32564
rect 6636 32510 6750 32562
rect 6802 32510 6804 32562
rect 6636 32508 6804 32510
rect 6636 31892 6692 32508
rect 6748 32498 6804 32508
rect 6076 31890 6692 31892
rect 6076 31838 6638 31890
rect 6690 31838 6692 31890
rect 6076 31836 6692 31838
rect 6076 31778 6132 31836
rect 6636 31826 6692 31836
rect 6076 31726 6078 31778
rect 6130 31726 6132 31778
rect 6076 31714 6132 31726
rect 6860 31780 6916 32732
rect 7308 32732 7476 32788
rect 7084 32564 7140 32574
rect 7308 32564 7364 32732
rect 7756 32674 7812 33292
rect 7980 33254 8036 33292
rect 7980 32788 8036 32798
rect 7980 32694 8036 32732
rect 7756 32622 7758 32674
rect 7810 32622 7812 32674
rect 7756 32610 7812 32622
rect 7140 32508 7364 32564
rect 7420 32562 7476 32574
rect 7420 32510 7422 32562
rect 7474 32510 7476 32562
rect 7084 32470 7140 32508
rect 6972 32450 7028 32462
rect 6972 32398 6974 32450
rect 7026 32398 7028 32450
rect 6972 32004 7028 32398
rect 7420 32116 7476 32510
rect 7868 32450 7924 32462
rect 7868 32398 7870 32450
rect 7922 32398 7924 32450
rect 7868 32116 7924 32398
rect 7420 32060 7924 32116
rect 7308 32004 7364 32014
rect 6972 31948 7140 32004
rect 6972 31780 7028 31790
rect 6860 31778 7028 31780
rect 6860 31726 6974 31778
rect 7026 31726 7028 31778
rect 6860 31724 7028 31726
rect 6972 31714 7028 31724
rect 6188 31556 6244 31566
rect 5964 31554 6244 31556
rect 5964 31502 6190 31554
rect 6242 31502 6244 31554
rect 5964 31500 6244 31502
rect 6188 31490 6244 31500
rect 6412 31556 6468 31566
rect 6412 31462 6468 31500
rect 4956 31378 5012 31388
rect 7084 31108 7140 31948
rect 7196 31892 7252 31902
rect 7196 31798 7252 31836
rect 7196 31108 7252 31118
rect 7084 31106 7252 31108
rect 7084 31054 7198 31106
rect 7250 31054 7252 31106
rect 7084 31052 7252 31054
rect 5404 30996 5460 31006
rect 5404 30902 5460 30940
rect 6300 30996 6356 31006
rect 6860 30996 6916 31006
rect 6300 30994 7140 30996
rect 6300 30942 6302 30994
rect 6354 30942 6862 30994
rect 6914 30942 7140 30994
rect 6300 30940 7140 30942
rect 6300 30930 6356 30940
rect 6860 30930 6916 30940
rect 6188 30884 6244 30894
rect 6188 30790 6244 30828
rect 6860 30772 6916 30782
rect 6300 30770 6916 30772
rect 6300 30718 6862 30770
rect 6914 30718 6916 30770
rect 6300 30716 6916 30718
rect 4732 30434 4900 30436
rect 4732 30382 4734 30434
rect 4786 30382 4900 30434
rect 4732 30380 4900 30382
rect 6076 30436 6132 30446
rect 4732 30324 4788 30380
rect 4732 30258 4788 30268
rect 6076 30322 6132 30380
rect 6076 30270 6078 30322
rect 6130 30270 6132 30322
rect 6076 30258 6132 30270
rect 6300 30210 6356 30716
rect 6860 30706 6916 30716
rect 6972 30772 7028 30782
rect 6300 30158 6302 30210
rect 6354 30158 6356 30210
rect 6300 30146 6356 30158
rect 6636 30212 6692 30222
rect 6636 30118 6692 30156
rect 4284 29538 4452 29540
rect 4284 29486 4398 29538
rect 4450 29486 4452 29538
rect 4284 29484 4452 29486
rect 4172 29428 4228 29438
rect 3612 29426 4228 29428
rect 3612 29374 4174 29426
rect 4226 29374 4228 29426
rect 3612 29372 4228 29374
rect 4172 28754 4228 29372
rect 4172 28702 4174 28754
rect 4226 28702 4228 28754
rect 4172 28690 4228 28702
rect 4284 28642 4340 29484
rect 4396 29474 4452 29484
rect 4844 30098 4900 30110
rect 4844 30046 4846 30098
rect 4898 30046 4900 30098
rect 4844 29428 4900 30046
rect 6972 30100 7028 30716
rect 7084 30434 7140 30940
rect 7196 30884 7252 31052
rect 7196 30818 7252 30828
rect 7084 30382 7086 30434
rect 7138 30382 7140 30434
rect 7084 30370 7140 30382
rect 7196 30212 7252 30222
rect 7308 30212 7364 31948
rect 8092 31892 8148 33516
rect 8652 33236 8708 33246
rect 7756 31836 8148 31892
rect 8204 33180 8652 33236
rect 8204 32004 8260 33180
rect 8652 33142 8708 33180
rect 8764 32676 8820 34078
rect 8988 33348 9044 34300
rect 8988 33254 9044 33292
rect 7644 31556 7700 31566
rect 7196 30210 7364 30212
rect 7196 30158 7198 30210
rect 7250 30158 7364 30210
rect 7196 30156 7364 30158
rect 7420 31554 7700 31556
rect 7420 31502 7646 31554
rect 7698 31502 7700 31554
rect 7420 31500 7700 31502
rect 7196 30146 7252 30156
rect 7084 30100 7140 30110
rect 6972 30098 7140 30100
rect 6972 30046 7086 30098
rect 7138 30046 7140 30098
rect 6972 30044 7140 30046
rect 7084 30034 7140 30044
rect 7420 29876 7476 31500
rect 7644 31490 7700 31500
rect 7756 30772 7812 31836
rect 7868 31668 7924 31678
rect 7868 31574 7924 31612
rect 7980 31668 8036 31678
rect 8204 31668 8260 31948
rect 7980 31666 8260 31668
rect 7980 31614 7982 31666
rect 8034 31614 8260 31666
rect 7980 31612 8260 31614
rect 8428 32620 8820 32676
rect 8428 31668 8484 32620
rect 8764 31780 8820 31790
rect 7980 31602 8036 31612
rect 8428 31602 8484 31612
rect 8652 31724 8764 31780
rect 8652 31666 8708 31724
rect 8764 31714 8820 31724
rect 8652 31614 8654 31666
rect 8706 31614 8708 31666
rect 8652 31602 8708 31614
rect 8316 31556 8372 31566
rect 8092 31554 8372 31556
rect 8092 31502 8318 31554
rect 8370 31502 8372 31554
rect 8092 31500 8372 31502
rect 7756 30706 7812 30716
rect 7980 30996 8036 31006
rect 8092 30996 8148 31500
rect 8316 31490 8372 31500
rect 8540 31556 8596 31566
rect 7980 30994 8148 30996
rect 7980 30942 7982 30994
rect 8034 30942 8148 30994
rect 7980 30940 8148 30942
rect 7756 30212 7812 30222
rect 7812 30156 7924 30212
rect 7756 30146 7812 30156
rect 7308 29820 7476 29876
rect 5068 29428 5124 29438
rect 4844 29426 5124 29428
rect 4844 29374 5070 29426
rect 5122 29374 5124 29426
rect 4844 29372 5124 29374
rect 5068 29362 5124 29372
rect 6524 29428 6580 29438
rect 4732 29316 4788 29326
rect 4732 29222 4788 29260
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4956 28868 5012 28878
rect 4956 28754 5012 28812
rect 4956 28702 4958 28754
rect 5010 28702 5012 28754
rect 4956 28690 5012 28702
rect 4284 28590 4286 28642
rect 4338 28590 4340 28642
rect 4284 28578 4340 28590
rect 6524 28530 6580 29372
rect 7308 29428 7364 29820
rect 7308 29334 7364 29372
rect 7756 29428 7812 29438
rect 7756 29334 7812 29372
rect 7420 29314 7476 29326
rect 7420 29262 7422 29314
rect 7474 29262 7476 29314
rect 7084 28756 7140 28766
rect 6524 28478 6526 28530
rect 6578 28478 6580 28530
rect 6524 28466 6580 28478
rect 6972 28644 7028 28654
rect 6860 27860 6916 27870
rect 6972 27860 7028 28588
rect 6860 27858 7028 27860
rect 6860 27806 6862 27858
rect 6914 27806 7028 27858
rect 6860 27804 7028 27806
rect 7084 27858 7140 28700
rect 7420 28082 7476 29262
rect 7868 28756 7924 30156
rect 7980 30210 8036 30940
rect 8540 30882 8596 31500
rect 9100 31444 9156 34748
rect 9436 34356 9492 35252
rect 9660 35186 9716 35196
rect 9772 35138 9828 35150
rect 9772 35086 9774 35138
rect 9826 35086 9828 35138
rect 9772 34916 9828 35086
rect 9884 35028 9940 38780
rect 9996 38612 10052 38622
rect 9996 38050 10052 38556
rect 10108 38610 10164 38622
rect 10108 38558 10110 38610
rect 10162 38558 10164 38610
rect 10108 38164 10164 38558
rect 10668 38276 10724 40124
rect 10780 39508 10836 40572
rect 11004 42364 11396 42420
rect 11452 42530 11508 42542
rect 11452 42478 11454 42530
rect 11506 42478 11508 42530
rect 11004 42084 11060 42364
rect 11452 42308 11508 42478
rect 11004 40628 11060 42028
rect 11004 40562 11060 40572
rect 11116 42252 11508 42308
rect 11676 42532 11732 42542
rect 11116 41858 11172 42252
rect 11116 41806 11118 41858
rect 11170 41806 11172 41858
rect 11116 40404 11172 41806
rect 11452 42082 11508 42094
rect 11452 42030 11454 42082
rect 11506 42030 11508 42082
rect 11452 41972 11508 42030
rect 11452 40404 11508 41916
rect 11676 41970 11732 42476
rect 11676 41918 11678 41970
rect 11730 41918 11732 41970
rect 11676 41906 11732 41918
rect 11900 42530 11956 42542
rect 11900 42478 11902 42530
rect 11954 42478 11956 42530
rect 11900 42084 11956 42478
rect 13356 42308 13412 43374
rect 13916 42754 13972 43596
rect 14364 43586 14420 43596
rect 14812 43652 14980 43708
rect 15036 43764 15092 43774
rect 15260 43764 15316 44158
rect 15484 44210 15540 44268
rect 15484 44158 15486 44210
rect 15538 44158 15540 44210
rect 15484 44146 15540 44158
rect 15596 44434 15652 44446
rect 15596 44382 15598 44434
rect 15650 44382 15652 44434
rect 15092 43708 15316 43764
rect 14140 43428 14196 43438
rect 14140 43334 14196 43372
rect 14812 42866 14868 43652
rect 15036 42978 15092 43708
rect 15596 43538 15652 44382
rect 16380 44324 16436 44334
rect 16380 44230 16436 44268
rect 17052 44324 17108 44334
rect 17388 44324 17444 45614
rect 18060 45666 18116 45678
rect 18396 45668 18452 45678
rect 18060 45614 18062 45666
rect 18114 45614 18116 45666
rect 17724 45220 17780 45230
rect 17724 45126 17780 45164
rect 17612 44660 17668 44670
rect 17500 44324 17556 44334
rect 17108 44322 17556 44324
rect 17108 44270 17502 44322
rect 17554 44270 17556 44322
rect 17108 44268 17556 44270
rect 17052 44230 17108 44268
rect 17500 44258 17556 44268
rect 17612 44212 17668 44604
rect 18060 44660 18116 45614
rect 18284 45666 18452 45668
rect 18284 45614 18398 45666
rect 18450 45614 18452 45666
rect 18284 45612 18452 45614
rect 18172 45332 18228 45342
rect 18172 45106 18228 45276
rect 18172 45054 18174 45106
rect 18226 45054 18228 45106
rect 18172 45042 18228 45054
rect 18060 44594 18116 44604
rect 17836 44212 17892 44222
rect 17612 44210 17780 44212
rect 17612 44158 17614 44210
rect 17666 44158 17780 44210
rect 17612 44156 17780 44158
rect 17612 44146 17668 44156
rect 16268 44100 16324 44110
rect 16268 44006 16324 44044
rect 16716 44098 16772 44110
rect 16716 44046 16718 44098
rect 16770 44046 16772 44098
rect 15596 43486 15598 43538
rect 15650 43486 15652 43538
rect 15596 43474 15652 43486
rect 15036 42926 15038 42978
rect 15090 42926 15092 42978
rect 15036 42914 15092 42926
rect 15260 43428 15316 43438
rect 15260 42978 15316 43372
rect 16268 43428 16324 43438
rect 16268 43334 16324 43372
rect 15260 42926 15262 42978
rect 15314 42926 15316 42978
rect 15260 42914 15316 42926
rect 14812 42814 14814 42866
rect 14866 42814 14868 42866
rect 14812 42802 14868 42814
rect 16716 42868 16772 44046
rect 17724 43540 17780 44156
rect 17836 44118 17892 44156
rect 17836 43540 17892 43550
rect 17724 43538 17892 43540
rect 17724 43486 17838 43538
rect 17890 43486 17892 43538
rect 17724 43484 17892 43486
rect 17836 43474 17892 43484
rect 17500 43426 17556 43438
rect 17500 43374 17502 43426
rect 17554 43374 17556 43426
rect 16716 42812 16884 42868
rect 13916 42702 13918 42754
rect 13970 42702 13972 42754
rect 13916 42690 13972 42702
rect 15708 42756 15764 42766
rect 16156 42756 16212 42766
rect 15708 42754 16772 42756
rect 15708 42702 15710 42754
rect 15762 42702 16158 42754
rect 16210 42702 16772 42754
rect 15708 42700 16772 42702
rect 15708 42690 15764 42700
rect 16156 42690 16212 42700
rect 13580 42642 13636 42654
rect 13580 42590 13582 42642
rect 13634 42590 13636 42642
rect 11900 40628 11956 42028
rect 12460 42252 13412 42308
rect 12460 41970 12516 42252
rect 12460 41918 12462 41970
rect 12514 41918 12516 41970
rect 12460 41906 12516 41918
rect 12684 42082 12740 42094
rect 12684 42030 12686 42082
rect 12738 42030 12740 42082
rect 12684 41524 12740 42030
rect 12908 42084 12964 42094
rect 12796 41524 12852 41534
rect 12684 41468 12796 41524
rect 12796 41458 12852 41468
rect 12908 41186 12964 42028
rect 13244 42084 13300 42094
rect 12908 41134 12910 41186
rect 12962 41134 12964 41186
rect 12908 41122 12964 41134
rect 13132 41860 13188 41870
rect 12572 41076 12628 41086
rect 12572 40982 12628 41020
rect 12796 40964 12852 40974
rect 12796 40870 12852 40908
rect 11900 40562 11956 40572
rect 12236 40514 12292 40526
rect 12236 40462 12238 40514
rect 12290 40462 12292 40514
rect 11116 40402 11284 40404
rect 11116 40350 11118 40402
rect 11170 40350 11284 40402
rect 11116 40348 11284 40350
rect 11116 40338 11172 40348
rect 11116 39844 11172 39854
rect 11116 39508 11172 39788
rect 10780 39058 10836 39452
rect 10780 39006 10782 39058
rect 10834 39006 10836 39058
rect 10780 38994 10836 39006
rect 11004 39506 11172 39508
rect 11004 39454 11118 39506
rect 11170 39454 11172 39506
rect 11004 39452 11172 39454
rect 11004 39058 11060 39452
rect 11116 39442 11172 39452
rect 11228 39620 11284 40348
rect 11452 40338 11508 40348
rect 11564 40404 11620 40414
rect 11900 40404 11956 40414
rect 12236 40404 12292 40462
rect 13020 40516 13076 40526
rect 11564 40402 11732 40404
rect 11564 40350 11566 40402
rect 11618 40350 11732 40402
rect 11564 40348 11732 40350
rect 11564 40338 11620 40348
rect 11564 39620 11620 39630
rect 11228 39618 11620 39620
rect 11228 39566 11566 39618
rect 11618 39566 11620 39618
rect 11228 39564 11620 39566
rect 11004 39006 11006 39058
rect 11058 39006 11060 39058
rect 11004 38994 11060 39006
rect 11228 38834 11284 39564
rect 11564 39554 11620 39564
rect 11228 38782 11230 38834
rect 11282 38782 11284 38834
rect 11228 38770 11284 38782
rect 10892 38724 10948 38734
rect 11676 38668 11732 40348
rect 11900 40310 11956 40348
rect 12124 40348 12236 40404
rect 12012 39508 12068 39518
rect 12012 39414 12068 39452
rect 12012 38836 12068 38846
rect 12012 38742 12068 38780
rect 10892 38630 10948 38668
rect 11452 38612 11732 38668
rect 11900 38724 11956 38734
rect 11900 38630 11956 38668
rect 10668 38220 11060 38276
rect 10108 38098 10164 38108
rect 9996 37998 9998 38050
rect 10050 37998 10052 38050
rect 9996 37940 10052 37998
rect 10332 38052 10388 38062
rect 10892 38052 10948 38062
rect 10332 38050 10948 38052
rect 10332 37998 10334 38050
rect 10386 37998 10894 38050
rect 10946 37998 10948 38050
rect 10332 37996 10948 37998
rect 10332 37986 10388 37996
rect 10892 37986 10948 37996
rect 9996 37874 10052 37884
rect 10108 37826 10164 37838
rect 10108 37774 10110 37826
rect 10162 37774 10164 37826
rect 9884 34972 10052 35028
rect 9772 34850 9828 34860
rect 9660 34804 9716 34814
rect 9660 34692 9716 34748
rect 9884 34804 9940 34814
rect 9884 34710 9940 34748
rect 9772 34692 9828 34702
rect 9660 34690 9828 34692
rect 9660 34638 9774 34690
rect 9826 34638 9828 34690
rect 9660 34636 9828 34638
rect 9772 34626 9828 34636
rect 9884 34468 9940 34478
rect 9436 34290 9492 34300
rect 9772 34356 9828 34366
rect 9772 34262 9828 34300
rect 9884 34242 9940 34412
rect 9884 34190 9886 34242
rect 9938 34190 9940 34242
rect 9884 34178 9940 34190
rect 9548 34132 9604 34142
rect 9548 34038 9604 34076
rect 9996 33348 10052 34972
rect 9772 33292 10052 33348
rect 9660 33124 9716 33134
rect 9548 33068 9660 33124
rect 9436 32788 9492 32798
rect 9548 32788 9604 33068
rect 9660 33030 9716 33068
rect 9492 32732 9604 32788
rect 9660 32788 9716 32798
rect 9772 32788 9828 33292
rect 9996 33124 10052 33134
rect 9660 32786 9828 32788
rect 9660 32734 9662 32786
rect 9714 32734 9828 32786
rect 9660 32732 9828 32734
rect 9884 33068 9996 33124
rect 9436 32722 9492 32732
rect 9660 32722 9716 32732
rect 9772 32564 9828 32574
rect 9884 32564 9940 33068
rect 9996 33030 10052 33068
rect 10108 33012 10164 37774
rect 11004 37828 11060 38220
rect 11116 38164 11172 38174
rect 11116 38070 11172 38108
rect 11116 37828 11172 37838
rect 11004 37772 11116 37828
rect 10332 37266 10388 37278
rect 10332 37214 10334 37266
rect 10386 37214 10388 37266
rect 10220 37154 10276 37166
rect 10220 37102 10222 37154
rect 10274 37102 10276 37154
rect 10220 37044 10276 37102
rect 10220 36978 10276 36988
rect 10332 36706 10388 37214
rect 10332 36654 10334 36706
rect 10386 36654 10388 36706
rect 10332 36642 10388 36654
rect 10220 36484 10276 36494
rect 10220 36390 10276 36428
rect 10332 36372 10388 36382
rect 10332 36278 10388 36316
rect 10780 36372 10836 36382
rect 10668 34916 10724 34926
rect 10668 34822 10724 34860
rect 10556 34804 10612 34814
rect 10556 34130 10612 34748
rect 10556 34078 10558 34130
rect 10610 34078 10612 34130
rect 10556 34066 10612 34078
rect 10668 34244 10724 34254
rect 10556 33348 10612 33358
rect 10668 33348 10724 34188
rect 10556 33346 10724 33348
rect 10556 33294 10558 33346
rect 10610 33294 10724 33346
rect 10556 33292 10724 33294
rect 10556 33124 10612 33292
rect 10556 33058 10612 33068
rect 10332 33012 10388 33022
rect 10108 32956 10332 33012
rect 10332 32674 10388 32956
rect 10780 32900 10836 36316
rect 10892 36260 10948 36270
rect 10892 36166 10948 36204
rect 11004 34804 11060 37772
rect 11116 37762 11172 37772
rect 11452 37156 11508 38612
rect 11564 37938 11620 37950
rect 11564 37886 11566 37938
rect 11618 37886 11620 37938
rect 11564 37268 11620 37886
rect 11676 37268 11732 37278
rect 11564 37266 11732 37268
rect 11564 37214 11678 37266
rect 11730 37214 11732 37266
rect 11564 37212 11732 37214
rect 11676 37202 11732 37212
rect 11004 34738 11060 34748
rect 11116 34914 11172 34926
rect 11116 34862 11118 34914
rect 11170 34862 11172 34914
rect 11116 34132 11172 34862
rect 11452 34468 11508 37100
rect 11564 36484 11620 36494
rect 11564 35026 11620 36428
rect 11564 34974 11566 35026
rect 11618 34974 11620 35026
rect 11564 34962 11620 34974
rect 11900 36260 11956 36270
rect 12124 36260 12180 40348
rect 12236 40338 12292 40348
rect 12684 40402 12740 40414
rect 12684 40350 12686 40402
rect 12738 40350 12740 40402
rect 12572 40180 12628 40190
rect 12236 40178 12628 40180
rect 12236 40126 12574 40178
rect 12626 40126 12628 40178
rect 12236 40124 12628 40126
rect 12236 38834 12292 40124
rect 12572 40114 12628 40124
rect 12684 39732 12740 40350
rect 12236 38782 12238 38834
rect 12290 38782 12292 38834
rect 12236 38770 12292 38782
rect 12348 39730 12740 39732
rect 12348 39678 12686 39730
rect 12738 39678 12740 39730
rect 12348 39676 12740 39678
rect 12348 38668 12404 39676
rect 12684 39666 12740 39676
rect 13020 39620 13076 40460
rect 13132 40514 13188 41804
rect 13132 40462 13134 40514
rect 13186 40462 13188 40514
rect 13132 40450 13188 40462
rect 13244 41524 13300 42028
rect 13356 41970 13412 42252
rect 13356 41918 13358 41970
rect 13410 41918 13412 41970
rect 13356 41906 13412 41918
rect 13468 42308 13524 42318
rect 13468 42082 13524 42252
rect 13580 42196 13636 42590
rect 13692 42532 13748 42542
rect 13692 42438 13748 42476
rect 16268 42530 16324 42542
rect 16268 42478 16270 42530
rect 16322 42478 16324 42530
rect 14588 42308 14644 42318
rect 13580 42130 13636 42140
rect 14028 42196 14084 42206
rect 14028 42194 14420 42196
rect 14028 42142 14030 42194
rect 14082 42142 14420 42194
rect 14028 42140 14420 42142
rect 14028 42130 14084 42140
rect 13468 42030 13470 42082
rect 13522 42030 13524 42082
rect 13468 41860 13524 42030
rect 13468 41794 13524 41804
rect 14028 41970 14084 41982
rect 14028 41918 14030 41970
rect 14082 41918 14084 41970
rect 13244 40514 13300 41468
rect 13580 41300 13636 41310
rect 13244 40462 13246 40514
rect 13298 40462 13300 40514
rect 13244 40450 13300 40462
rect 13356 41244 13580 41300
rect 13356 40514 13412 41244
rect 13580 41206 13636 41244
rect 14028 41300 14084 41918
rect 14028 41234 14084 41244
rect 13804 41076 13860 41086
rect 13804 40982 13860 41020
rect 13356 40462 13358 40514
rect 13410 40462 13412 40514
rect 13356 40450 13412 40462
rect 14252 40964 14308 40974
rect 13804 40404 13860 40414
rect 14140 40404 14196 40414
rect 13804 40402 14196 40404
rect 13804 40350 13806 40402
rect 13858 40350 14142 40402
rect 14194 40350 14196 40402
rect 13804 40348 14196 40350
rect 13804 40338 13860 40348
rect 14140 40338 14196 40348
rect 13916 39842 13972 39854
rect 13916 39790 13918 39842
rect 13970 39790 13972 39842
rect 13916 39732 13972 39790
rect 13916 39676 14196 39732
rect 13020 39060 13076 39564
rect 14028 39506 14084 39518
rect 14028 39454 14030 39506
rect 14082 39454 14084 39506
rect 13916 39396 13972 39406
rect 13804 39394 13972 39396
rect 13804 39342 13918 39394
rect 13970 39342 13972 39394
rect 13804 39340 13972 39342
rect 13244 39060 13300 39070
rect 13020 39058 13300 39060
rect 13020 39006 13246 39058
rect 13298 39006 13300 39058
rect 13020 39004 13300 39006
rect 13244 38994 13300 39004
rect 13468 39060 13524 39070
rect 13692 39060 13748 39070
rect 13468 39058 13692 39060
rect 13468 39006 13470 39058
rect 13522 39006 13692 39058
rect 13468 39004 13692 39006
rect 13468 38994 13524 39004
rect 13692 38994 13748 39004
rect 12796 38836 12852 38846
rect 12796 38742 12852 38780
rect 11956 36204 12180 36260
rect 12236 38612 12404 38668
rect 13356 38722 13412 38734
rect 13356 38670 13358 38722
rect 13410 38670 13412 38722
rect 12236 37604 12292 38612
rect 12236 36482 12292 37548
rect 13356 37492 13412 38670
rect 13804 38724 13860 39340
rect 13916 39330 13972 39340
rect 13804 38658 13860 38668
rect 13916 38836 13972 38846
rect 13916 38722 13972 38780
rect 13916 38670 13918 38722
rect 13970 38670 13972 38722
rect 13916 38658 13972 38670
rect 14028 38724 14084 39454
rect 14140 38946 14196 39676
rect 14140 38894 14142 38946
rect 14194 38894 14196 38946
rect 14140 38882 14196 38894
rect 14252 38724 14308 40908
rect 14028 38668 14308 38724
rect 14364 40290 14420 42140
rect 14588 42194 14644 42252
rect 14588 42142 14590 42194
rect 14642 42142 14644 42194
rect 14588 42130 14644 42142
rect 14476 42084 14532 42094
rect 14476 41990 14532 42028
rect 15372 42084 15428 42094
rect 15372 41990 15428 42028
rect 16268 42084 16324 42478
rect 16268 42018 16324 42028
rect 16380 42530 16436 42542
rect 16380 42478 16382 42530
rect 16434 42478 16436 42530
rect 14812 41970 14868 41982
rect 14812 41918 14814 41970
rect 14866 41918 14868 41970
rect 14812 41188 14868 41918
rect 15596 41972 15652 41982
rect 15596 41878 15652 41916
rect 16156 41970 16212 41982
rect 16156 41918 16158 41970
rect 16210 41918 16212 41970
rect 15036 41188 15092 41198
rect 14812 41186 15092 41188
rect 14812 41134 15038 41186
rect 15090 41134 15092 41186
rect 14812 41132 15092 41134
rect 15036 41122 15092 41132
rect 14588 41076 14644 41086
rect 14588 40402 14644 41020
rect 16156 40964 16212 41918
rect 16380 41300 16436 42478
rect 16492 42530 16548 42542
rect 16492 42478 16494 42530
rect 16546 42478 16548 42530
rect 16492 41972 16548 42478
rect 16492 41906 16548 41916
rect 16604 42530 16660 42542
rect 16604 42478 16606 42530
rect 16658 42478 16660 42530
rect 16604 42196 16660 42478
rect 16604 41748 16660 42140
rect 16716 41970 16772 42700
rect 16716 41918 16718 41970
rect 16770 41918 16772 41970
rect 16716 41906 16772 41918
rect 16828 41748 16884 42812
rect 16604 41692 16884 41748
rect 16380 41234 16436 41244
rect 16604 41412 16660 41422
rect 16380 41076 16436 41086
rect 16380 40982 16436 41020
rect 16156 40898 16212 40908
rect 16604 40628 16660 41356
rect 16716 40964 16772 40974
rect 16828 40964 16884 41692
rect 16940 41746 16996 41758
rect 16940 41694 16942 41746
rect 16994 41694 16996 41746
rect 16940 41188 16996 41694
rect 17388 41188 17444 41198
rect 16940 41186 17444 41188
rect 16940 41134 17390 41186
rect 17442 41134 17444 41186
rect 16940 41132 17444 41134
rect 17388 41122 17444 41132
rect 17500 41188 17556 43374
rect 18060 41300 18116 41310
rect 18060 41206 18116 41244
rect 17500 41122 17556 41132
rect 17948 41076 18004 41086
rect 17052 40964 17108 40974
rect 16828 40962 17108 40964
rect 16828 40910 17054 40962
rect 17106 40910 17108 40962
rect 16828 40908 17108 40910
rect 16716 40870 16772 40908
rect 17052 40898 17108 40908
rect 14588 40350 14590 40402
rect 14642 40350 14644 40402
rect 14588 40338 14644 40350
rect 14700 40404 14756 40414
rect 14700 40310 14756 40348
rect 14364 40238 14366 40290
rect 14418 40238 14420 40290
rect 14364 39842 14420 40238
rect 14364 39790 14366 39842
rect 14418 39790 14420 39842
rect 14364 39060 14420 39790
rect 14700 39730 14756 39742
rect 14700 39678 14702 39730
rect 14754 39678 14756 39730
rect 14588 39620 14644 39630
rect 14588 39508 14644 39564
rect 13468 37492 13524 37502
rect 13356 37436 13468 37492
rect 14028 37492 14084 38668
rect 14364 38274 14420 39004
rect 14364 38222 14366 38274
rect 14418 38222 14420 38274
rect 14364 38210 14420 38222
rect 14476 39506 14644 39508
rect 14476 39454 14590 39506
rect 14642 39454 14644 39506
rect 14476 39452 14644 39454
rect 14140 38164 14196 38174
rect 14140 38162 14308 38164
rect 14140 38110 14142 38162
rect 14194 38110 14308 38162
rect 14140 38108 14308 38110
rect 14140 38098 14196 38108
rect 14252 38052 14308 38108
rect 14476 38052 14532 39452
rect 14588 39442 14644 39452
rect 14700 39396 14756 39678
rect 14700 39330 14756 39340
rect 15372 39396 15428 39406
rect 14588 38836 14644 38846
rect 14588 38274 14644 38780
rect 15372 38834 15428 39340
rect 15372 38782 15374 38834
rect 15426 38782 15428 38834
rect 15372 38770 15428 38782
rect 16604 38834 16660 40572
rect 17388 40404 17444 40414
rect 17388 40310 17444 40348
rect 17948 40402 18004 41020
rect 17948 40350 17950 40402
rect 18002 40350 18004 40402
rect 17948 40338 18004 40350
rect 18284 40852 18340 45612
rect 18396 45602 18452 45612
rect 19628 45668 19684 45678
rect 19628 45220 19684 45612
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 20748 45332 20804 45726
rect 21308 45778 21364 45790
rect 21308 45726 21310 45778
rect 21362 45726 21364 45778
rect 21084 45668 21140 45678
rect 21084 45574 21140 45612
rect 20748 45266 20804 45276
rect 21084 45332 21140 45342
rect 21308 45332 21364 45726
rect 21084 45330 21364 45332
rect 21084 45278 21086 45330
rect 21138 45278 21364 45330
rect 21084 45276 21364 45278
rect 21756 45332 21812 45948
rect 26796 45910 26852 45948
rect 27132 45892 27188 45902
rect 21868 45332 21924 45342
rect 21756 45330 21924 45332
rect 21756 45278 21870 45330
rect 21922 45278 21924 45330
rect 21756 45276 21924 45278
rect 21084 45266 21140 45276
rect 21868 45266 21924 45276
rect 19628 45164 19796 45220
rect 18956 45108 19012 45118
rect 18956 45014 19012 45052
rect 19292 45108 19348 45118
rect 18956 44884 19012 44894
rect 18956 44322 19012 44828
rect 18956 44270 18958 44322
rect 19010 44270 19012 44322
rect 18956 44258 19012 44270
rect 19292 44210 19348 45052
rect 19628 44994 19684 45006
rect 19628 44942 19630 44994
rect 19682 44942 19684 44994
rect 19628 44324 19684 44942
rect 19628 44258 19684 44268
rect 19740 44322 19796 45164
rect 22540 45218 22596 45230
rect 22540 45166 22542 45218
rect 22594 45166 22596 45218
rect 20188 45108 20244 45118
rect 20188 45014 20244 45052
rect 20748 45108 20804 45118
rect 21756 45108 21812 45118
rect 20804 45052 20916 45108
rect 20748 45042 20804 45052
rect 19964 44994 20020 45006
rect 19964 44942 19966 44994
rect 20018 44942 20020 44994
rect 19964 44548 20020 44942
rect 20636 44996 20692 45006
rect 20636 44902 20692 44940
rect 20412 44884 20468 44894
rect 20412 44790 20468 44828
rect 19964 44482 20020 44492
rect 20524 44548 20580 44558
rect 19740 44270 19742 44322
rect 19794 44270 19796 44322
rect 19740 44258 19796 44270
rect 20412 44324 20468 44334
rect 20412 44230 20468 44268
rect 19292 44158 19294 44210
rect 19346 44158 19348 44210
rect 19292 44146 19348 44158
rect 19740 44100 19796 44110
rect 19404 44098 19796 44100
rect 19404 44046 19742 44098
rect 19794 44046 19796 44098
rect 19404 44044 19796 44046
rect 19404 42980 19460 44044
rect 19740 44034 19796 44044
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 20524 43538 20580 44492
rect 20748 44210 20804 44222
rect 20748 44158 20750 44210
rect 20802 44158 20804 44210
rect 20748 44100 20804 44158
rect 20748 44034 20804 44044
rect 20524 43486 20526 43538
rect 20578 43486 20580 43538
rect 20524 43474 20580 43486
rect 20748 43540 20804 43550
rect 20860 43540 20916 45052
rect 21644 45106 21812 45108
rect 21644 45054 21758 45106
rect 21810 45054 21812 45106
rect 21644 45052 21812 45054
rect 21308 44996 21364 45006
rect 21308 44902 21364 44940
rect 21532 44994 21588 45006
rect 21532 44942 21534 44994
rect 21586 44942 21588 44994
rect 21532 44884 21588 44942
rect 21532 44818 21588 44828
rect 21308 44548 21364 44558
rect 21308 44322 21364 44492
rect 21308 44270 21310 44322
rect 21362 44270 21364 44322
rect 21308 44258 21364 44270
rect 21644 44098 21700 45052
rect 21756 45042 21812 45052
rect 21980 45108 22036 45118
rect 22428 45108 22484 45118
rect 22036 45106 22484 45108
rect 22036 45054 22430 45106
rect 22482 45054 22484 45106
rect 22036 45052 22484 45054
rect 21980 45014 22036 45052
rect 22428 45042 22484 45052
rect 21644 44046 21646 44098
rect 21698 44046 21700 44098
rect 21644 43764 21700 44046
rect 21644 43698 21700 43708
rect 21868 44324 21924 44334
rect 20748 43538 20916 43540
rect 20748 43486 20750 43538
rect 20802 43486 20916 43538
rect 20748 43484 20916 43486
rect 20748 43474 20804 43484
rect 19180 42924 19460 42980
rect 19516 43428 19572 43438
rect 19180 42756 19236 42924
rect 18620 42754 19236 42756
rect 18620 42702 19182 42754
rect 19234 42702 19236 42754
rect 18620 42700 19236 42702
rect 18620 41858 18676 42700
rect 19180 42690 19236 42700
rect 19516 42754 19572 43372
rect 21868 43426 21924 44268
rect 22092 44322 22148 44334
rect 22092 44270 22094 44322
rect 22146 44270 22148 44322
rect 22092 44212 22148 44270
rect 22092 44146 22148 44156
rect 22204 44100 22260 44110
rect 22204 43538 22260 44044
rect 22540 43764 22596 45166
rect 22764 45108 22820 45118
rect 26796 45108 26852 45118
rect 22764 45106 22932 45108
rect 22764 45054 22766 45106
rect 22818 45054 22932 45106
rect 22764 45052 22932 45054
rect 22764 45042 22820 45052
rect 22876 44324 22932 45052
rect 23212 44324 23268 44334
rect 22876 44322 23380 44324
rect 22876 44270 23214 44322
rect 23266 44270 23380 44322
rect 22876 44268 23380 44270
rect 23212 44258 23268 44268
rect 22540 43698 22596 43708
rect 22764 44210 22820 44222
rect 22764 44158 22766 44210
rect 22818 44158 22820 44210
rect 22204 43486 22206 43538
rect 22258 43486 22260 43538
rect 22204 43474 22260 43486
rect 21868 43374 21870 43426
rect 21922 43374 21924 43426
rect 21868 43362 21924 43374
rect 22652 43426 22708 43438
rect 22652 43374 22654 43426
rect 22706 43374 22708 43426
rect 20972 43314 21028 43326
rect 20972 43262 20974 43314
rect 21026 43262 21028 43314
rect 20972 42868 21028 43262
rect 21420 43316 21476 43326
rect 21420 43222 21476 43260
rect 20972 42802 21028 42812
rect 19516 42702 19518 42754
rect 19570 42702 19572 42754
rect 19516 42308 19572 42702
rect 22652 42756 22708 43374
rect 22764 43316 22820 44158
rect 22764 43250 22820 43260
rect 22652 42700 23044 42756
rect 19516 42242 19572 42252
rect 19628 42642 19684 42654
rect 19628 42590 19630 42642
rect 19682 42590 19684 42642
rect 19628 42196 19684 42590
rect 22988 42644 23044 42700
rect 23324 42754 23380 44268
rect 23436 44212 23492 44222
rect 23436 43538 23492 44156
rect 23436 43486 23438 43538
rect 23490 43486 23492 43538
rect 23436 43474 23492 43486
rect 24332 43764 24388 43774
rect 23660 43426 23716 43438
rect 23660 43374 23662 43426
rect 23714 43374 23716 43426
rect 23324 42702 23326 42754
rect 23378 42702 23380 42754
rect 23324 42690 23380 42702
rect 23436 43316 23492 43326
rect 22988 42642 23268 42644
rect 22988 42590 22990 42642
rect 23042 42590 23268 42642
rect 22988 42588 23268 42590
rect 22988 42578 23044 42588
rect 22652 42530 22708 42542
rect 22652 42478 22654 42530
rect 22706 42478 22708 42530
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 19964 42196 20020 42206
rect 19628 42140 19796 42196
rect 19068 42084 19124 42094
rect 19068 42082 19684 42084
rect 19068 42030 19070 42082
rect 19122 42030 19684 42082
rect 19068 42028 19684 42030
rect 19068 42018 19124 42028
rect 18620 41806 18622 41858
rect 18674 41806 18676 41858
rect 18508 41188 18564 41198
rect 18620 41188 18676 41806
rect 18508 41186 18676 41188
rect 18508 41134 18510 41186
rect 18562 41134 18676 41186
rect 18508 41132 18676 41134
rect 18732 41188 18788 41198
rect 18508 41122 18564 41132
rect 17724 39732 17780 39742
rect 16604 38782 16606 38834
rect 16658 38782 16660 38834
rect 16604 38770 16660 38782
rect 16828 39508 16884 39518
rect 16828 39058 16884 39452
rect 16828 39006 16830 39058
rect 16882 39006 16884 39058
rect 16044 38724 16100 38762
rect 16044 38658 16100 38668
rect 16828 38668 16884 39006
rect 17724 38834 17780 39676
rect 18284 39618 18340 40796
rect 18396 41074 18452 41086
rect 18396 41022 18398 41074
rect 18450 41022 18452 41074
rect 18396 40628 18452 41022
rect 18396 40514 18452 40572
rect 18396 40462 18398 40514
rect 18450 40462 18452 40514
rect 18396 40450 18452 40462
rect 18284 39566 18286 39618
rect 18338 39566 18340 39618
rect 18284 39554 18340 39566
rect 18396 40290 18452 40302
rect 18396 40238 18398 40290
rect 18450 40238 18452 40290
rect 17948 39394 18004 39406
rect 17948 39342 17950 39394
rect 18002 39342 18004 39394
rect 17948 39172 18004 39342
rect 18172 39394 18228 39406
rect 18172 39342 18174 39394
rect 18226 39342 18228 39394
rect 18172 39284 18228 39342
rect 18172 39218 18228 39228
rect 17948 39106 18004 39116
rect 17724 38782 17726 38834
rect 17778 38782 17780 38834
rect 17724 38668 17780 38782
rect 17948 38946 18004 38958
rect 17948 38894 17950 38946
rect 18002 38894 18004 38946
rect 17948 38668 18004 38894
rect 18396 38722 18452 40238
rect 18732 39844 18788 41132
rect 19292 41188 19348 41198
rect 19180 41076 19236 41086
rect 18732 39778 18788 39788
rect 18844 41074 19236 41076
rect 18844 41022 19182 41074
rect 19234 41022 19236 41074
rect 18844 41020 19236 41022
rect 18844 40626 18900 41020
rect 19180 41010 19236 41020
rect 19292 41074 19348 41132
rect 19516 41188 19572 41198
rect 19516 41094 19572 41132
rect 19628 41186 19684 42028
rect 19628 41134 19630 41186
rect 19682 41134 19684 41186
rect 19628 41122 19684 41134
rect 19292 41022 19294 41074
rect 19346 41022 19348 41074
rect 19292 41010 19348 41022
rect 19740 40964 19796 42140
rect 19964 41970 20020 42140
rect 19964 41918 19966 41970
rect 20018 41918 20020 41970
rect 19964 41906 20020 41918
rect 20636 41972 20692 41982
rect 20636 41878 20692 41916
rect 22204 41972 22260 41982
rect 22204 41878 22260 41916
rect 22652 41970 22708 42478
rect 22652 41918 22654 41970
rect 22706 41918 22708 41970
rect 21196 41860 21252 41870
rect 19964 41412 20020 41422
rect 19964 41186 20020 41356
rect 19964 41134 19966 41186
rect 20018 41134 20020 41186
rect 19964 41122 20020 41134
rect 19404 40908 19796 40964
rect 19852 40964 19908 41002
rect 18844 40574 18846 40626
rect 18898 40574 18900 40626
rect 18844 39732 18900 40574
rect 19068 40852 19124 40862
rect 19068 40404 19124 40796
rect 19404 40628 19460 40908
rect 19852 40898 19908 40908
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 19068 40310 19124 40348
rect 19292 40572 19460 40628
rect 20972 40628 21028 40638
rect 19292 40068 19348 40572
rect 19516 40514 19572 40526
rect 19516 40462 19518 40514
rect 19570 40462 19572 40514
rect 19404 40404 19460 40414
rect 19516 40404 19572 40462
rect 19628 40516 19684 40526
rect 19628 40422 19684 40460
rect 19852 40516 19908 40526
rect 19852 40422 19908 40460
rect 19460 40348 19572 40404
rect 20188 40404 20244 40414
rect 19404 40338 19460 40348
rect 20188 40310 20244 40348
rect 20972 40290 21028 40572
rect 20972 40238 20974 40290
rect 21026 40238 21028 40290
rect 20972 40226 21028 40238
rect 18844 39666 18900 39676
rect 19068 40012 19348 40068
rect 19068 39618 19124 40012
rect 19180 39844 19236 39854
rect 19180 39732 19236 39788
rect 19180 39676 19348 39732
rect 19068 39566 19070 39618
rect 19122 39566 19124 39618
rect 19068 39554 19124 39566
rect 18620 39508 18676 39518
rect 18620 39414 18676 39452
rect 18956 39506 19012 39518
rect 18956 39454 18958 39506
rect 19010 39454 19012 39506
rect 18844 39396 18900 39406
rect 18844 39302 18900 39340
rect 18620 39172 18676 39182
rect 18620 38946 18676 39116
rect 18620 38894 18622 38946
rect 18674 38894 18676 38946
rect 18620 38882 18676 38894
rect 18396 38670 18398 38722
rect 18450 38670 18452 38722
rect 16828 38612 17220 38668
rect 17724 38612 17892 38668
rect 17948 38612 18228 38668
rect 14588 38222 14590 38274
rect 14642 38222 14644 38274
rect 14588 38210 14644 38222
rect 16268 38500 16324 38510
rect 14252 37996 14532 38052
rect 16268 37940 16324 38444
rect 16044 37938 16324 37940
rect 16044 37886 16270 37938
rect 16322 37886 16324 37938
rect 16044 37884 16324 37886
rect 15036 37826 15092 37838
rect 15036 37774 15038 37826
rect 15090 37774 15092 37826
rect 14476 37604 14532 37614
rect 14028 37436 14420 37492
rect 13468 37398 13524 37436
rect 12460 37380 12516 37390
rect 12460 37286 12516 37324
rect 12236 36430 12238 36482
rect 12290 36430 12292 36482
rect 11228 34356 11284 34366
rect 11228 34262 11284 34300
rect 11452 34244 11508 34412
rect 11676 34244 11732 34254
rect 11452 34242 11732 34244
rect 11452 34190 11678 34242
rect 11730 34190 11732 34242
rect 11452 34188 11732 34190
rect 11676 34178 11732 34188
rect 11788 34244 11844 34254
rect 11788 34150 11844 34188
rect 11116 34038 11172 34076
rect 11228 34020 11284 34030
rect 11284 33964 11396 34020
rect 11228 33954 11284 33964
rect 11004 33348 11060 33358
rect 11004 33346 11284 33348
rect 11004 33294 11006 33346
rect 11058 33294 11284 33346
rect 11004 33292 11284 33294
rect 11004 33282 11060 33292
rect 10332 32622 10334 32674
rect 10386 32622 10388 32674
rect 10332 32610 10388 32622
rect 10556 32844 10836 32900
rect 9772 32562 9940 32564
rect 9772 32510 9774 32562
rect 9826 32510 9940 32562
rect 9772 32508 9940 32510
rect 9772 32498 9828 32508
rect 9660 32338 9716 32350
rect 9660 32286 9662 32338
rect 9714 32286 9716 32338
rect 9660 31780 9716 32286
rect 10556 31892 10612 32844
rect 11228 32788 11284 33292
rect 11228 32722 11284 32732
rect 10668 32676 10724 32686
rect 11116 32676 11172 32686
rect 10668 32674 11172 32676
rect 10668 32622 10670 32674
rect 10722 32622 11118 32674
rect 11170 32622 11172 32674
rect 10668 32620 11172 32622
rect 10668 32610 10724 32620
rect 11004 31892 11060 32620
rect 11116 32610 11172 32620
rect 11228 32564 11284 32574
rect 11340 32564 11396 33964
rect 11900 33908 11956 36204
rect 12236 35924 12292 36430
rect 12348 37268 12404 37278
rect 12348 36482 12404 37212
rect 13244 37268 13300 37278
rect 12348 36430 12350 36482
rect 12402 36430 12404 36482
rect 12348 36418 12404 36430
rect 12460 36484 12516 36494
rect 12460 36390 12516 36428
rect 12908 36260 12964 36270
rect 12908 36166 12964 36204
rect 12236 35868 13076 35924
rect 13020 35810 13076 35868
rect 13020 35758 13022 35810
rect 13074 35758 13076 35810
rect 13020 35746 13076 35758
rect 13244 35698 13300 37212
rect 14028 37268 14084 37278
rect 14028 37174 14084 37212
rect 14252 37266 14308 37278
rect 14252 37214 14254 37266
rect 14306 37214 14308 37266
rect 14140 36484 14196 36494
rect 14028 36370 14084 36382
rect 14028 36318 14030 36370
rect 14082 36318 14084 36370
rect 13916 35924 13972 35962
rect 13916 35858 13972 35868
rect 13244 35646 13246 35698
rect 13298 35646 13300 35698
rect 13244 35634 13300 35646
rect 14028 35476 14084 36318
rect 14140 35698 14196 36428
rect 14252 36482 14308 37214
rect 14252 36430 14254 36482
rect 14306 36430 14308 36482
rect 14252 36418 14308 36430
rect 14140 35646 14142 35698
rect 14194 35646 14196 35698
rect 14140 35634 14196 35646
rect 14364 35700 14420 37436
rect 14476 37490 14532 37548
rect 14476 37438 14478 37490
rect 14530 37438 14532 37490
rect 14476 37426 14532 37438
rect 14588 37492 14644 37502
rect 14588 37378 14644 37436
rect 14588 37326 14590 37378
rect 14642 37326 14644 37378
rect 14588 37314 14644 37326
rect 15036 37044 15092 37774
rect 15820 37380 15876 37390
rect 15820 37156 15876 37324
rect 15820 37090 15876 37100
rect 15036 36978 15092 36988
rect 15148 36484 15204 36494
rect 15148 36390 15204 36428
rect 14028 34914 14084 35420
rect 14028 34862 14030 34914
rect 14082 34862 14084 34914
rect 14028 34850 14084 34862
rect 14364 34914 14420 35644
rect 14476 36260 14532 36270
rect 14476 35698 14532 36204
rect 14476 35646 14478 35698
rect 14530 35646 14532 35698
rect 14476 35634 14532 35646
rect 14700 35924 14756 35934
rect 14700 35698 14756 35868
rect 14700 35646 14702 35698
rect 14754 35646 14756 35698
rect 14364 34862 14366 34914
rect 14418 34862 14420 34914
rect 14364 34850 14420 34862
rect 14252 34692 14308 34702
rect 14252 34598 14308 34636
rect 13132 34356 13188 34366
rect 12012 34132 12068 34142
rect 12684 34132 12740 34142
rect 12012 34130 12740 34132
rect 12012 34078 12014 34130
rect 12066 34078 12686 34130
rect 12738 34078 12740 34130
rect 12012 34076 12740 34078
rect 12012 34066 12068 34076
rect 11900 33852 12068 33908
rect 11788 32788 11844 32798
rect 11844 32732 11956 32788
rect 11788 32722 11844 32732
rect 11228 32562 11396 32564
rect 11228 32510 11230 32562
rect 11282 32510 11396 32562
rect 11228 32508 11396 32510
rect 11228 32498 11284 32508
rect 10612 31836 10948 31892
rect 10556 31826 10612 31836
rect 9660 31714 9716 31724
rect 9884 31668 9940 31678
rect 9100 31378 9156 31388
rect 9548 31554 9604 31566
rect 9548 31502 9550 31554
rect 9602 31502 9604 31554
rect 9548 31444 9604 31502
rect 9548 31378 9604 31388
rect 9884 31554 9940 31612
rect 9884 31502 9886 31554
rect 9938 31502 9940 31554
rect 8652 30996 8708 31006
rect 9548 30996 9604 31006
rect 8652 30994 9604 30996
rect 8652 30942 8654 30994
rect 8706 30942 9550 30994
rect 9602 30942 9604 30994
rect 8652 30940 9604 30942
rect 8652 30930 8708 30940
rect 9548 30930 9604 30940
rect 9660 30996 9716 31006
rect 9660 30902 9716 30940
rect 8540 30830 8542 30882
rect 8594 30830 8596 30882
rect 8540 30818 8596 30830
rect 7980 30158 7982 30210
rect 8034 30158 8036 30210
rect 7980 30146 8036 30158
rect 8652 30770 8708 30782
rect 8652 30718 8654 30770
rect 8706 30718 8708 30770
rect 8652 30210 8708 30718
rect 9884 30772 9940 31502
rect 10892 31556 10948 31836
rect 11004 31826 11060 31836
rect 11116 32338 11172 32350
rect 11116 32286 11118 32338
rect 11170 32286 11172 32338
rect 11116 31778 11172 32286
rect 11340 31892 11396 31902
rect 11340 31890 11844 31892
rect 11340 31838 11342 31890
rect 11394 31838 11844 31890
rect 11340 31836 11844 31838
rect 11340 31826 11396 31836
rect 11116 31726 11118 31778
rect 11170 31726 11172 31778
rect 11116 31714 11172 31726
rect 11788 31778 11844 31836
rect 11788 31726 11790 31778
rect 11842 31726 11844 31778
rect 11788 31714 11844 31726
rect 11564 31668 11620 31678
rect 11564 31574 11620 31612
rect 10892 31218 10948 31500
rect 10892 31166 10894 31218
rect 10946 31166 10948 31218
rect 10892 31154 10948 31166
rect 11228 31332 11284 31342
rect 11228 31218 11284 31276
rect 11228 31166 11230 31218
rect 11282 31166 11284 31218
rect 11228 31154 11284 31166
rect 11676 31106 11732 31118
rect 11676 31054 11678 31106
rect 11730 31054 11732 31106
rect 11452 30996 11508 31006
rect 9884 30706 9940 30716
rect 11004 30994 11508 30996
rect 11004 30942 11454 30994
rect 11506 30942 11508 30994
rect 11004 30940 11508 30942
rect 11004 30660 11060 30940
rect 11452 30930 11508 30940
rect 11676 30772 11732 31054
rect 11788 31108 11844 31118
rect 11900 31108 11956 32732
rect 12012 31780 12068 33852
rect 12684 33460 12740 34076
rect 13132 34130 13188 34300
rect 14364 34356 14420 34366
rect 13132 34078 13134 34130
rect 13186 34078 13188 34130
rect 13132 34066 13188 34078
rect 13580 34132 13636 34142
rect 13580 34038 13636 34076
rect 13916 34130 13972 34142
rect 13916 34078 13918 34130
rect 13970 34078 13972 34130
rect 12684 33394 12740 33404
rect 13132 33460 13188 33470
rect 13132 32450 13188 33404
rect 13580 33460 13636 33470
rect 13580 33366 13636 33404
rect 13916 33460 13972 34078
rect 14364 34130 14420 34300
rect 14364 34078 14366 34130
rect 14418 34078 14420 34130
rect 14364 34066 14420 34078
rect 14700 34132 14756 35646
rect 14924 35588 14980 35598
rect 14812 35586 14980 35588
rect 14812 35534 14926 35586
rect 14978 35534 14980 35586
rect 14812 35532 14980 35534
rect 14812 35476 14868 35532
rect 14924 35522 14980 35532
rect 14812 35410 14868 35420
rect 15036 35474 15092 35486
rect 15036 35422 15038 35474
rect 15090 35422 15092 35474
rect 15036 34916 15092 35422
rect 15036 34850 15092 34860
rect 14700 34038 14756 34076
rect 15260 34132 15316 34142
rect 13916 33394 13972 33404
rect 14924 34018 14980 34030
rect 14924 33966 14926 34018
rect 14978 33966 14980 34018
rect 14028 33348 14084 33358
rect 13692 32676 13748 32686
rect 14028 32676 14084 33292
rect 13692 32674 14084 32676
rect 13692 32622 13694 32674
rect 13746 32622 14084 32674
rect 13692 32620 14084 32622
rect 14924 33348 14980 33966
rect 15036 33348 15092 33358
rect 14924 33346 15092 33348
rect 14924 33294 15038 33346
rect 15090 33294 15092 33346
rect 14924 33292 15092 33294
rect 14924 32676 14980 33292
rect 15036 33282 15092 33292
rect 13692 32610 13748 32620
rect 14924 32582 14980 32620
rect 15148 33012 15204 33022
rect 13132 32398 13134 32450
rect 13186 32398 13188 32450
rect 13132 32386 13188 32398
rect 14924 31892 14980 31902
rect 12124 31780 12180 31790
rect 12012 31724 12124 31780
rect 12124 31686 12180 31724
rect 12572 31780 12628 31790
rect 12572 31686 12628 31724
rect 14140 31668 14196 31678
rect 14140 31574 14196 31612
rect 14476 31668 14532 31678
rect 12012 31556 12068 31566
rect 12012 31462 12068 31500
rect 13916 31554 13972 31566
rect 13916 31502 13918 31554
rect 13970 31502 13972 31554
rect 11788 31106 11956 31108
rect 11788 31054 11790 31106
rect 11842 31054 11956 31106
rect 11788 31052 11956 31054
rect 12348 31106 12404 31118
rect 12348 31054 12350 31106
rect 12402 31054 12404 31106
rect 11788 31042 11844 31052
rect 12348 30996 12404 31054
rect 12460 31108 12516 31118
rect 12460 31014 12516 31052
rect 13916 31106 13972 31502
rect 13916 31054 13918 31106
rect 13970 31054 13972 31106
rect 13020 30996 13076 31006
rect 12348 30930 12404 30940
rect 12572 30994 13076 30996
rect 12572 30942 13022 30994
rect 13074 30942 13076 30994
rect 12572 30940 13076 30942
rect 11676 30706 11732 30716
rect 12348 30772 12404 30782
rect 12572 30772 12628 30940
rect 13020 30930 13076 30940
rect 13468 30996 13524 31006
rect 13132 30882 13188 30894
rect 13132 30830 13134 30882
rect 13186 30830 13188 30882
rect 12348 30770 12628 30772
rect 12348 30718 12350 30770
rect 12402 30718 12628 30770
rect 12348 30716 12628 30718
rect 12684 30772 12740 30782
rect 12348 30706 12404 30716
rect 10332 30604 11060 30660
rect 8988 30436 9044 30446
rect 8988 30342 9044 30380
rect 9884 30436 9940 30446
rect 9884 30322 9940 30380
rect 9884 30270 9886 30322
rect 9938 30270 9940 30322
rect 9884 30258 9940 30270
rect 8652 30158 8654 30210
rect 8706 30158 8708 30210
rect 8428 29426 8484 29438
rect 8428 29374 8430 29426
rect 8482 29374 8484 29426
rect 7868 28642 7924 28700
rect 7868 28590 7870 28642
rect 7922 28590 7924 28642
rect 7868 28578 7924 28590
rect 8092 29316 8148 29326
rect 7420 28030 7422 28082
rect 7474 28030 7476 28082
rect 7420 28018 7476 28030
rect 7084 27806 7086 27858
rect 7138 27806 7140 27858
rect 6860 27794 6916 27804
rect 7084 27794 7140 27806
rect 8092 27858 8148 29260
rect 8316 29204 8372 29214
rect 8316 29110 8372 29148
rect 8092 27806 8094 27858
rect 8146 27806 8148 27858
rect 8092 27794 8148 27806
rect 8428 28754 8484 29374
rect 8540 29316 8596 29326
rect 8540 29222 8596 29260
rect 8428 28702 8430 28754
rect 8482 28702 8484 28754
rect 8428 27746 8484 28702
rect 8652 28644 8708 30158
rect 9212 30212 9268 30222
rect 8764 29428 8820 29438
rect 8764 28866 8820 29372
rect 8764 28814 8766 28866
rect 8818 28814 8820 28866
rect 8764 28802 8820 28814
rect 9100 28868 9156 28878
rect 9212 28868 9268 30156
rect 10332 30210 10388 30604
rect 10332 30158 10334 30210
rect 10386 30158 10388 30210
rect 10332 30146 10388 30158
rect 10444 30436 10500 30446
rect 10444 29426 10500 30380
rect 10668 29538 10724 30604
rect 12684 30210 12740 30716
rect 12684 30158 12686 30210
rect 12738 30158 12740 30210
rect 12684 30146 12740 30158
rect 13020 30212 13076 30222
rect 13132 30212 13188 30830
rect 13020 30210 13188 30212
rect 13020 30158 13022 30210
rect 13074 30158 13188 30210
rect 13020 30156 13188 30158
rect 13468 30210 13524 30940
rect 13468 30158 13470 30210
rect 13522 30158 13524 30210
rect 13020 30146 13076 30156
rect 13468 30146 13524 30158
rect 13804 30884 13860 30894
rect 13804 30210 13860 30828
rect 13804 30158 13806 30210
rect 13858 30158 13860 30210
rect 13804 30146 13860 30158
rect 13916 30210 13972 31054
rect 13916 30158 13918 30210
rect 13970 30158 13972 30210
rect 13916 30146 13972 30158
rect 14028 31554 14084 31566
rect 14364 31556 14420 31566
rect 14028 31502 14030 31554
rect 14082 31502 14084 31554
rect 10668 29486 10670 29538
rect 10722 29486 10724 29538
rect 10668 29474 10724 29486
rect 10780 30098 10836 30110
rect 10780 30046 10782 30098
rect 10834 30046 10836 30098
rect 10444 29374 10446 29426
rect 10498 29374 10500 29426
rect 10444 29362 10500 29374
rect 9100 28866 9268 28868
rect 9100 28814 9102 28866
rect 9154 28814 9268 28866
rect 9100 28812 9268 28814
rect 10556 29204 10612 29214
rect 9100 28802 9156 28812
rect 8764 28644 8820 28654
rect 10556 28644 10612 29148
rect 10780 28756 10836 30046
rect 12796 29988 12852 29998
rect 12796 29894 12852 29932
rect 13580 29988 13636 29998
rect 13580 29894 13636 29932
rect 11452 29876 11508 29886
rect 11452 29650 11508 29820
rect 11452 29598 11454 29650
rect 11506 29598 11508 29650
rect 11452 29586 11508 29598
rect 11340 29428 11396 29438
rect 8708 28642 8820 28644
rect 8708 28590 8766 28642
rect 8818 28590 8820 28642
rect 8708 28588 8820 28590
rect 8652 28550 8708 28588
rect 8764 28578 8820 28588
rect 10332 28642 10612 28644
rect 10332 28590 10558 28642
rect 10610 28590 10612 28642
rect 10332 28588 10612 28590
rect 8988 27860 9044 27870
rect 8988 27766 9044 27804
rect 10332 27858 10388 28588
rect 10556 28578 10612 28588
rect 10668 28754 10836 28756
rect 10668 28702 10782 28754
rect 10834 28702 10836 28754
rect 10668 28700 10836 28702
rect 10332 27806 10334 27858
rect 10386 27806 10388 27858
rect 10332 27794 10388 27806
rect 10556 27860 10612 27870
rect 10668 27860 10724 28700
rect 10780 28690 10836 28700
rect 10892 29426 11396 29428
rect 10892 29374 11342 29426
rect 11394 29374 11396 29426
rect 10892 29372 11396 29374
rect 10892 28082 10948 29372
rect 11340 29362 11396 29372
rect 13132 29314 13188 29326
rect 13132 29262 13134 29314
rect 13186 29262 13188 29314
rect 11228 28644 11284 28654
rect 11228 28550 11284 28588
rect 12124 28644 12180 28654
rect 12012 28530 12068 28542
rect 12012 28478 12014 28530
rect 12066 28478 12068 28530
rect 11788 28420 11844 28430
rect 12012 28420 12068 28478
rect 12124 28530 12180 28588
rect 12572 28644 12628 28654
rect 12124 28478 12126 28530
rect 12178 28478 12180 28530
rect 12124 28466 12180 28478
rect 12348 28532 12404 28542
rect 12348 28438 12404 28476
rect 11788 28418 12012 28420
rect 11788 28366 11790 28418
rect 11842 28366 12012 28418
rect 11788 28364 12012 28366
rect 11788 28354 11844 28364
rect 12012 28354 12068 28364
rect 10892 28030 10894 28082
rect 10946 28030 10948 28082
rect 10892 28018 10948 28030
rect 12572 27970 12628 28588
rect 12796 28644 12852 28654
rect 12796 28550 12852 28588
rect 12908 28532 12964 28542
rect 13132 28532 13188 29262
rect 14028 29316 14084 31502
rect 14252 31554 14420 31556
rect 14252 31502 14366 31554
rect 14418 31502 14420 31554
rect 14252 31500 14420 31502
rect 14252 29986 14308 31500
rect 14364 31490 14420 31500
rect 14364 30884 14420 30894
rect 14364 30790 14420 30828
rect 14364 30212 14420 30222
rect 14476 30212 14532 31612
rect 14924 31666 14980 31836
rect 14924 31614 14926 31666
rect 14978 31614 14980 31666
rect 14924 31602 14980 31614
rect 15036 31668 15092 31678
rect 15036 31574 15092 31612
rect 14700 31554 14756 31566
rect 14700 31502 14702 31554
rect 14754 31502 14756 31554
rect 14700 30994 14756 31502
rect 14700 30942 14702 30994
rect 14754 30942 14756 30994
rect 14700 30930 14756 30942
rect 14364 30210 14532 30212
rect 14364 30158 14366 30210
rect 14418 30158 14532 30210
rect 14364 30156 14532 30158
rect 14364 30146 14420 30156
rect 14588 30100 14644 30110
rect 14588 30006 14644 30044
rect 14252 29934 14254 29986
rect 14306 29934 14308 29986
rect 14252 29922 14308 29934
rect 15036 29652 15092 29662
rect 15148 29652 15204 32956
rect 15260 32674 15316 34076
rect 15708 33572 15764 33582
rect 15708 33478 15764 33516
rect 15260 32622 15262 32674
rect 15314 32622 15316 32674
rect 15260 32610 15316 32622
rect 15708 32564 15764 32574
rect 15708 32470 15764 32508
rect 16044 32340 16100 37884
rect 16268 37874 16324 37884
rect 16716 38050 16772 38062
rect 16716 37998 16718 38050
rect 16770 37998 16772 38050
rect 16492 37604 16548 37614
rect 16492 37490 16548 37548
rect 16492 37438 16494 37490
rect 16546 37438 16548 37490
rect 16492 37426 16548 37438
rect 16716 37380 16772 37998
rect 16156 37266 16212 37278
rect 16156 37214 16158 37266
rect 16210 37214 16212 37266
rect 16156 37044 16212 37214
rect 16268 37268 16324 37278
rect 16268 37174 16324 37212
rect 16604 37266 16660 37278
rect 16604 37214 16606 37266
rect 16658 37214 16660 37266
rect 16380 37156 16436 37166
rect 16380 37062 16436 37100
rect 16156 36978 16212 36988
rect 16492 36370 16548 36382
rect 16492 36318 16494 36370
rect 16546 36318 16548 36370
rect 16268 35700 16324 35710
rect 16268 35606 16324 35644
rect 16492 35476 16548 36318
rect 16604 35812 16660 37214
rect 16604 35718 16660 35756
rect 16492 35410 16548 35420
rect 16716 35252 16772 37324
rect 16268 35196 16772 35252
rect 17164 38050 17220 38612
rect 17164 37998 17166 38050
rect 17218 37998 17220 38050
rect 16268 32562 16324 35196
rect 16604 34242 16660 34254
rect 16604 34190 16606 34242
rect 16658 34190 16660 34242
rect 16604 34132 16660 34190
rect 16380 34076 16660 34132
rect 16716 34130 16772 34142
rect 16716 34078 16718 34130
rect 16770 34078 16772 34130
rect 16380 33236 16436 34076
rect 16604 33906 16660 33918
rect 16604 33854 16606 33906
rect 16658 33854 16660 33906
rect 16492 33460 16548 33470
rect 16492 33366 16548 33404
rect 16604 33348 16660 33854
rect 16716 33796 16772 34078
rect 16716 33730 16772 33740
rect 16828 33348 16884 33358
rect 16604 33292 16828 33348
rect 16828 33254 16884 33292
rect 16380 32900 16436 33180
rect 16492 32900 16548 32910
rect 16380 32844 16492 32900
rect 16492 32834 16548 32844
rect 16380 32676 16436 32686
rect 16380 32582 16436 32620
rect 16268 32510 16270 32562
rect 16322 32510 16324 32562
rect 16268 32498 16324 32510
rect 16716 32564 16772 32574
rect 16716 32450 16772 32508
rect 16716 32398 16718 32450
rect 16770 32398 16772 32450
rect 16716 32386 16772 32398
rect 16044 32284 16436 32340
rect 16268 31892 16324 31902
rect 15596 31780 15652 31790
rect 15484 31668 15540 31678
rect 15484 31574 15540 31612
rect 15596 31108 15652 31724
rect 15932 31220 15988 31230
rect 15932 31126 15988 31164
rect 15596 31014 15652 31052
rect 16268 31108 16324 31836
rect 16380 31780 16436 32284
rect 16716 31780 16772 31790
rect 16380 31778 16772 31780
rect 16380 31726 16718 31778
rect 16770 31726 16772 31778
rect 16380 31724 16772 31726
rect 16716 31714 16772 31724
rect 17164 31780 17220 37998
rect 17388 37828 17444 37838
rect 17388 37734 17444 37772
rect 17500 37826 17556 37838
rect 17500 37774 17502 37826
rect 17554 37774 17556 37826
rect 17500 37716 17556 37774
rect 17500 37650 17556 37660
rect 17500 37266 17556 37278
rect 17500 37214 17502 37266
rect 17554 37214 17556 37266
rect 17388 37044 17444 37054
rect 17388 35698 17444 36988
rect 17500 35922 17556 37214
rect 17500 35870 17502 35922
rect 17554 35870 17556 35922
rect 17500 35858 17556 35870
rect 17612 37268 17668 37278
rect 17612 35810 17668 37212
rect 17612 35758 17614 35810
rect 17666 35758 17668 35810
rect 17612 35746 17668 35758
rect 17836 36484 17892 38612
rect 18060 37604 18116 37614
rect 17948 37156 18004 37166
rect 17948 37062 18004 37100
rect 17948 36484 18004 36494
rect 17836 36482 18004 36484
rect 17836 36430 17950 36482
rect 18002 36430 18004 36482
rect 17836 36428 18004 36430
rect 17388 35646 17390 35698
rect 17442 35646 17444 35698
rect 17388 35634 17444 35646
rect 17836 35252 17892 36428
rect 17948 36418 18004 36428
rect 18060 36370 18116 37548
rect 18060 36318 18062 36370
rect 18114 36318 18116 36370
rect 17948 35812 18004 35822
rect 17948 35698 18004 35756
rect 17948 35646 17950 35698
rect 18002 35646 18004 35698
rect 17948 35634 18004 35646
rect 18060 35700 18116 36318
rect 18060 35634 18116 35644
rect 18172 37268 18228 38612
rect 17836 35186 17892 35196
rect 17948 35476 18004 35486
rect 17836 35026 17892 35038
rect 17836 34974 17838 35026
rect 17890 34974 17892 35026
rect 17388 34916 17444 34926
rect 17388 34822 17444 34860
rect 17500 34018 17556 34030
rect 17500 33966 17502 34018
rect 17554 33966 17556 34018
rect 17388 33570 17444 33582
rect 17388 33518 17390 33570
rect 17442 33518 17444 33570
rect 17276 33348 17332 33358
rect 17276 33254 17332 33292
rect 17388 32674 17444 33518
rect 17500 33572 17556 33966
rect 17500 33506 17556 33516
rect 17836 34020 17892 34974
rect 17948 34914 18004 35420
rect 17948 34862 17950 34914
rect 18002 34862 18004 34914
rect 17948 34850 18004 34862
rect 17948 34130 18004 34142
rect 17948 34078 17950 34130
rect 18002 34078 18004 34130
rect 17948 34020 18004 34078
rect 17836 33964 17948 34020
rect 17836 33458 17892 33964
rect 17948 33954 18004 33964
rect 17836 33406 17838 33458
rect 17890 33406 17892 33458
rect 17836 33394 17892 33406
rect 17948 33572 18004 33582
rect 17948 33346 18004 33516
rect 17948 33294 17950 33346
rect 18002 33294 18004 33346
rect 17948 33282 18004 33294
rect 17836 33236 17892 33246
rect 17388 32622 17390 32674
rect 17442 32622 17444 32674
rect 17388 31890 17444 32622
rect 17388 31838 17390 31890
rect 17442 31838 17444 31890
rect 17388 31826 17444 31838
rect 17724 33124 17780 33134
rect 17724 32562 17780 33068
rect 17724 32510 17726 32562
rect 17778 32510 17780 32562
rect 17164 31714 17220 31724
rect 17724 31778 17780 32510
rect 17836 32564 17892 33180
rect 17836 32470 17892 32508
rect 18060 32450 18116 32462
rect 18060 32398 18062 32450
rect 18114 32398 18116 32450
rect 18060 32340 18116 32398
rect 18172 32340 18228 37212
rect 18396 37268 18452 38670
rect 18508 38724 18564 38734
rect 18508 38162 18564 38668
rect 18508 38110 18510 38162
rect 18562 38110 18564 38162
rect 18508 38098 18564 38110
rect 18732 38050 18788 38062
rect 18732 37998 18734 38050
rect 18786 37998 18788 38050
rect 18732 37268 18788 37998
rect 18396 37266 18788 37268
rect 18396 37214 18398 37266
rect 18450 37214 18788 37266
rect 18396 37212 18788 37214
rect 18956 37268 19012 39454
rect 19180 39284 19236 39294
rect 19180 38276 19236 39228
rect 19292 38500 19348 39676
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 19852 38834 19908 38846
rect 19852 38782 19854 38834
rect 19906 38782 19908 38834
rect 19852 38724 19908 38782
rect 20524 38836 20580 38846
rect 20860 38836 20916 38846
rect 20524 38834 20916 38836
rect 20524 38782 20526 38834
rect 20578 38782 20862 38834
rect 20914 38782 20916 38834
rect 20524 38780 20916 38782
rect 20524 38770 20580 38780
rect 19852 38658 19908 38668
rect 20412 38724 20468 38734
rect 19292 38434 19348 38444
rect 20076 38500 20132 38510
rect 19180 38220 19348 38276
rect 19068 37268 19124 37278
rect 18956 37212 19068 37268
rect 18396 37202 18452 37212
rect 19068 37174 19124 37212
rect 19292 37266 19348 38220
rect 19404 37940 19460 37950
rect 19404 37938 19572 37940
rect 19404 37886 19406 37938
rect 19458 37886 19572 37938
rect 19404 37884 19572 37886
rect 19404 37874 19460 37884
rect 19292 37214 19294 37266
rect 19346 37214 19348 37266
rect 19292 37202 19348 37214
rect 19516 37266 19572 37884
rect 20076 37828 20132 38444
rect 20076 37772 20244 37828
rect 19628 37716 19684 37726
rect 19628 37380 19684 37660
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 20076 37492 20132 37502
rect 20188 37492 20244 37772
rect 20076 37490 20244 37492
rect 20076 37438 20078 37490
rect 20130 37438 20244 37490
rect 20076 37436 20244 37438
rect 20076 37426 20132 37436
rect 19964 37380 20020 37390
rect 19628 37378 20020 37380
rect 19628 37326 19966 37378
rect 20018 37326 20020 37378
rect 19628 37324 20020 37326
rect 19964 37314 20020 37324
rect 19516 37214 19518 37266
rect 19570 37214 19572 37266
rect 19516 37202 19572 37214
rect 20300 37268 20356 37278
rect 20300 37174 20356 37212
rect 19180 37154 19236 37166
rect 19180 37102 19182 37154
rect 19234 37102 19236 37154
rect 18396 37042 18452 37054
rect 18396 36990 18398 37042
rect 18450 36990 18452 37042
rect 18396 36596 18452 36990
rect 19180 36708 19236 37102
rect 19180 36642 19236 36652
rect 18620 36596 18676 36606
rect 18396 36540 18620 36596
rect 18284 36372 18340 36382
rect 18284 36278 18340 36316
rect 18396 36036 18452 36540
rect 18620 36502 18676 36540
rect 19516 36596 19572 36606
rect 18956 36372 19012 36382
rect 18956 36278 19012 36316
rect 18284 35980 18452 36036
rect 18284 34802 18340 35980
rect 18508 35812 18564 35822
rect 18284 34750 18286 34802
rect 18338 34750 18340 34802
rect 18284 34738 18340 34750
rect 18396 34804 18452 34814
rect 18396 34242 18452 34748
rect 18396 34190 18398 34242
rect 18450 34190 18452 34242
rect 18396 34178 18452 34190
rect 18508 33796 18564 35756
rect 18620 35700 18676 35710
rect 18620 35606 18676 35644
rect 19516 35698 19572 36540
rect 20188 36482 20244 36494
rect 20188 36430 20190 36482
rect 20242 36430 20244 36482
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 20188 35924 20244 36430
rect 19516 35646 19518 35698
rect 19570 35646 19572 35698
rect 19516 35634 19572 35646
rect 20076 35868 20244 35924
rect 19292 35586 19348 35598
rect 19292 35534 19294 35586
rect 19346 35534 19348 35586
rect 19292 35476 19348 35534
rect 19292 35410 19348 35420
rect 20076 35476 20132 35868
rect 20188 35700 20244 35710
rect 20188 35606 20244 35644
rect 20076 35410 20132 35420
rect 18844 35252 18900 35262
rect 18844 34914 18900 35196
rect 18844 34862 18846 34914
rect 18898 34862 18900 34914
rect 18844 34850 18900 34862
rect 19404 34972 19796 35028
rect 18956 34692 19012 34702
rect 18956 34598 19012 34636
rect 19180 34692 19236 34702
rect 19404 34692 19460 34972
rect 19740 34914 19796 34972
rect 19740 34862 19742 34914
rect 19794 34862 19796 34914
rect 19740 34850 19796 34862
rect 19516 34804 19572 34814
rect 19516 34710 19572 34748
rect 20076 34804 20132 34814
rect 20076 34710 20132 34748
rect 19180 34690 19460 34692
rect 19180 34638 19182 34690
rect 19234 34638 19460 34690
rect 19180 34636 19460 34638
rect 19628 34690 19684 34702
rect 19628 34638 19630 34690
rect 19682 34638 19684 34690
rect 19180 34242 19236 34636
rect 19180 34190 19182 34242
rect 19234 34190 19236 34242
rect 19180 34178 19236 34190
rect 18844 34020 18900 34030
rect 18844 33926 18900 33964
rect 18508 33730 18564 33740
rect 18844 33796 18900 33806
rect 18844 33346 18900 33740
rect 18844 33294 18846 33346
rect 18898 33294 18900 33346
rect 18844 33282 18900 33294
rect 19180 33346 19236 33358
rect 19180 33294 19182 33346
rect 19234 33294 19236 33346
rect 19068 33124 19124 33134
rect 19068 33030 19124 33068
rect 18620 32900 18676 32910
rect 18396 32788 18452 32798
rect 18396 32694 18452 32732
rect 18284 32676 18340 32686
rect 18284 32582 18340 32620
rect 18060 32284 18340 32340
rect 17724 31726 17726 31778
rect 17778 31726 17780 31778
rect 17724 31714 17780 31726
rect 18172 31780 18228 31790
rect 18284 31780 18340 32284
rect 18508 31780 18564 31790
rect 18284 31778 18564 31780
rect 18284 31726 18510 31778
rect 18562 31726 18564 31778
rect 18284 31724 18564 31726
rect 18172 31686 18228 31724
rect 18508 31714 18564 31724
rect 18620 31666 18676 32844
rect 19180 32676 19236 33294
rect 19404 33348 19460 33358
rect 19404 33254 19460 33292
rect 19628 33124 19684 34638
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 20300 34132 20356 34142
rect 20300 34038 20356 34076
rect 20412 33124 20468 38668
rect 20860 38164 20916 38780
rect 20860 38098 20916 38108
rect 20748 36596 20804 36606
rect 20748 36502 20804 36540
rect 20636 36372 20692 36382
rect 20636 35922 20692 36316
rect 20636 35870 20638 35922
rect 20690 35870 20692 35922
rect 20636 35858 20692 35870
rect 20524 35700 20580 35710
rect 20524 35606 20580 35644
rect 20860 35698 20916 35710
rect 20860 35646 20862 35698
rect 20914 35646 20916 35698
rect 19628 33068 20244 33124
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 19180 32610 19236 32620
rect 20076 32674 20132 32686
rect 20076 32622 20078 32674
rect 20130 32622 20132 32674
rect 19964 32564 20020 32574
rect 19964 32470 20020 32508
rect 20076 32116 20132 32622
rect 19516 32060 20132 32116
rect 19516 31892 19572 32060
rect 18844 31836 19572 31892
rect 18844 31778 18900 31836
rect 18844 31726 18846 31778
rect 18898 31726 18900 31778
rect 18844 31714 18900 31726
rect 18620 31614 18622 31666
rect 18674 31614 18676 31666
rect 18620 31602 18676 31614
rect 19292 31668 19348 31678
rect 16268 30994 16324 31052
rect 16268 30942 16270 30994
rect 16322 30942 16324 30994
rect 16268 30930 16324 30942
rect 16492 31554 16548 31566
rect 16492 31502 16494 31554
rect 16546 31502 16548 31554
rect 16492 30996 16548 31502
rect 16828 31332 16884 31342
rect 16884 31276 16996 31332
rect 16828 31266 16884 31276
rect 15260 30882 15316 30894
rect 15260 30830 15262 30882
rect 15314 30830 15316 30882
rect 15260 30212 15316 30830
rect 16492 30772 16548 30940
rect 16268 30770 16548 30772
rect 16268 30718 16494 30770
rect 16546 30718 16548 30770
rect 16268 30716 16548 30718
rect 15260 30146 15316 30156
rect 16044 30324 16100 30334
rect 14588 29650 15204 29652
rect 14588 29598 15038 29650
rect 15090 29598 15204 29650
rect 14588 29596 15204 29598
rect 14588 29594 14644 29596
rect 14476 29538 14532 29550
rect 14476 29486 14478 29538
rect 14530 29486 14532 29538
rect 14588 29542 14590 29594
rect 14642 29542 14644 29594
rect 15036 29586 15092 29596
rect 14588 29530 14644 29542
rect 14476 29428 14532 29486
rect 14476 29372 14644 29428
rect 14028 29250 14084 29260
rect 14140 29204 14196 29214
rect 14140 28754 14196 29148
rect 14140 28702 14142 28754
rect 14194 28702 14196 28754
rect 14140 28690 14196 28702
rect 14476 29202 14532 29214
rect 14476 29150 14478 29202
rect 14530 29150 14532 29202
rect 13916 28642 13972 28654
rect 13916 28590 13918 28642
rect 13970 28590 13972 28642
rect 12908 28530 13188 28532
rect 12908 28478 12910 28530
rect 12962 28478 13188 28530
rect 12908 28476 13188 28478
rect 13580 28532 13636 28542
rect 12908 28420 12964 28476
rect 13580 28438 13636 28476
rect 12572 27918 12574 27970
rect 12626 27918 12628 27970
rect 12572 27906 12628 27918
rect 12796 28364 12908 28420
rect 10556 27858 10724 27860
rect 10556 27806 10558 27858
rect 10610 27806 10724 27858
rect 10556 27804 10724 27806
rect 12796 27858 12852 28364
rect 12908 28354 12964 28364
rect 13804 28420 13860 28430
rect 12796 27806 12798 27858
rect 12850 27806 12852 27858
rect 10556 27794 10612 27804
rect 12796 27794 12852 27806
rect 8428 27694 8430 27746
rect 8482 27694 8484 27746
rect 8428 27682 8484 27694
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 1932 27188 1988 27198
rect 13804 27188 13860 28364
rect 13916 27972 13972 28590
rect 14364 28644 14420 28654
rect 14364 28550 14420 28588
rect 13916 27970 14308 27972
rect 13916 27918 13918 27970
rect 13970 27918 14308 27970
rect 13916 27916 14308 27918
rect 13916 27906 13972 27916
rect 14140 27746 14196 27758
rect 14140 27694 14142 27746
rect 14194 27694 14196 27746
rect 14140 27300 14196 27694
rect 14140 27234 14196 27244
rect 13916 27188 13972 27198
rect 13804 27186 13972 27188
rect 13804 27134 13918 27186
rect 13970 27134 13972 27186
rect 13804 27132 13972 27134
rect 1932 27094 1988 27132
rect 13916 27122 13972 27132
rect 14252 27186 14308 27916
rect 14252 27134 14254 27186
rect 14306 27134 14308 27186
rect 14252 27122 14308 27134
rect 4284 27074 4340 27086
rect 4284 27022 4286 27074
rect 4338 27022 4340 27074
rect 4284 26516 4340 27022
rect 12012 26962 12068 26974
rect 12012 26910 12014 26962
rect 12066 26910 12068 26962
rect 12012 26908 12068 26910
rect 11676 26852 12068 26908
rect 12348 26964 12404 27002
rect 12348 26898 12404 26908
rect 14476 26962 14532 29150
rect 14588 28644 14644 29372
rect 15148 28868 15204 29596
rect 15596 29652 15652 29662
rect 15932 29652 15988 29662
rect 15596 29650 15932 29652
rect 15596 29598 15598 29650
rect 15650 29598 15932 29650
rect 15596 29596 15932 29598
rect 15596 29586 15652 29596
rect 15932 29558 15988 29596
rect 16044 29538 16100 30268
rect 16268 29988 16324 30716
rect 16492 30706 16548 30716
rect 16604 31220 16660 31230
rect 16604 30436 16660 31164
rect 16268 29922 16324 29932
rect 16492 30380 16660 30436
rect 16828 30770 16884 30782
rect 16828 30718 16830 30770
rect 16882 30718 16884 30770
rect 16492 29652 16548 30380
rect 16604 30212 16660 30222
rect 16604 30118 16660 30156
rect 16828 29988 16884 30718
rect 16716 29932 16884 29988
rect 16940 30436 16996 31276
rect 16940 30210 16996 30380
rect 16940 30158 16942 30210
rect 16994 30158 16996 30210
rect 16604 29652 16660 29662
rect 16492 29650 16660 29652
rect 16492 29598 16606 29650
rect 16658 29598 16660 29650
rect 16492 29596 16660 29598
rect 16604 29586 16660 29596
rect 16044 29486 16046 29538
rect 16098 29486 16100 29538
rect 16044 29474 16100 29486
rect 16380 29540 16436 29550
rect 15708 29428 15764 29438
rect 15708 29334 15764 29372
rect 16380 29426 16436 29484
rect 16716 29540 16772 29932
rect 16828 29652 16884 29662
rect 16940 29652 16996 30158
rect 17164 31220 17220 31230
rect 17164 30210 17220 31164
rect 17612 31220 17668 31230
rect 17612 31126 17668 31164
rect 17388 31108 17444 31118
rect 17388 31014 17444 31052
rect 17836 30996 17892 31006
rect 17836 30902 17892 30940
rect 17948 30994 18004 31006
rect 17948 30942 17950 30994
rect 18002 30942 18004 30994
rect 17724 30882 17780 30894
rect 17724 30830 17726 30882
rect 17778 30830 17780 30882
rect 17612 30324 17668 30334
rect 17612 30230 17668 30268
rect 17164 30158 17166 30210
rect 17218 30158 17220 30210
rect 17052 29986 17108 29998
rect 17052 29934 17054 29986
rect 17106 29934 17108 29986
rect 17052 29764 17108 29934
rect 17164 29988 17220 30158
rect 17388 30212 17444 30222
rect 17724 30212 17780 30830
rect 17948 30436 18004 30942
rect 19292 30996 19348 31612
rect 19292 30930 19348 30940
rect 19516 31666 19572 31836
rect 19628 31892 19684 31902
rect 19628 31890 20020 31892
rect 19628 31838 19630 31890
rect 19682 31838 20020 31890
rect 19628 31836 20020 31838
rect 19628 31826 19684 31836
rect 19964 31778 20020 31836
rect 19964 31726 19966 31778
rect 20018 31726 20020 31778
rect 19964 31714 20020 31726
rect 20188 31778 20244 33068
rect 20412 33058 20468 33068
rect 20524 35364 20580 35374
rect 20188 31726 20190 31778
rect 20242 31726 20244 31778
rect 19516 31614 19518 31666
rect 19570 31614 19572 31666
rect 19516 30882 19572 31614
rect 20076 31556 20132 31594
rect 20076 31490 20132 31500
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 20076 31108 20132 31118
rect 20188 31108 20244 31726
rect 20300 32562 20356 32574
rect 20300 32510 20302 32562
rect 20354 32510 20356 32562
rect 20300 31668 20356 32510
rect 20412 31668 20468 31678
rect 20300 31666 20468 31668
rect 20300 31614 20414 31666
rect 20466 31614 20468 31666
rect 20300 31612 20468 31614
rect 20412 31602 20468 31612
rect 20076 31106 20244 31108
rect 20076 31054 20078 31106
rect 20130 31054 20244 31106
rect 20076 31052 20244 31054
rect 20076 31042 20132 31052
rect 19516 30830 19518 30882
rect 19570 30830 19572 30882
rect 19516 30818 19572 30830
rect 17724 30156 17892 30212
rect 17388 30118 17444 30156
rect 17724 29988 17780 29998
rect 17164 29986 17780 29988
rect 17164 29934 17726 29986
rect 17778 29934 17780 29986
rect 17164 29932 17780 29934
rect 17724 29922 17780 29932
rect 17052 29708 17668 29764
rect 16828 29650 16996 29652
rect 16828 29598 16830 29650
rect 16882 29598 16996 29650
rect 16828 29596 16996 29598
rect 17612 29650 17668 29708
rect 17612 29598 17614 29650
rect 17666 29598 17668 29650
rect 16828 29586 16884 29596
rect 17612 29586 17668 29598
rect 16716 29474 16772 29484
rect 16380 29374 16382 29426
rect 16434 29374 16436 29426
rect 15260 28868 15316 28878
rect 15148 28866 15764 28868
rect 15148 28814 15262 28866
rect 15314 28814 15764 28866
rect 15148 28812 15764 28814
rect 15260 28802 15316 28812
rect 14924 28644 14980 28654
rect 14588 28642 14980 28644
rect 14588 28590 14926 28642
rect 14978 28590 14980 28642
rect 14588 28588 14980 28590
rect 14924 27860 14980 28588
rect 14924 27766 14980 27804
rect 15148 28418 15204 28430
rect 15148 28366 15150 28418
rect 15202 28366 15204 28418
rect 14700 27524 14756 27534
rect 14700 27074 14756 27468
rect 14700 27022 14702 27074
rect 14754 27022 14756 27074
rect 14700 27010 14756 27022
rect 15148 27074 15204 28366
rect 15148 27022 15150 27074
rect 15202 27022 15204 27074
rect 15148 27010 15204 27022
rect 15260 28308 15316 28318
rect 14476 26910 14478 26962
rect 14530 26910 14532 26962
rect 14476 26898 14532 26910
rect 12236 26852 12292 26862
rect 4284 26450 4340 26460
rect 8652 26516 8708 26526
rect 4284 26290 4340 26302
rect 4284 26238 4286 26290
rect 4338 26238 4340 26290
rect 1932 26180 1988 26190
rect 1932 26086 1988 26124
rect 4284 26180 4340 26238
rect 4284 26114 4340 26124
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 1932 25620 1988 25630
rect 1932 25526 1988 25564
rect 8652 25618 8708 26460
rect 11676 26402 11732 26852
rect 12236 26758 12292 26796
rect 13580 26852 13636 26862
rect 11676 26350 11678 26402
rect 11730 26350 11732 26402
rect 11676 26338 11732 26350
rect 12908 26404 12964 26414
rect 11564 26292 11620 26302
rect 8652 25566 8654 25618
rect 8706 25566 8708 25618
rect 4284 25508 4340 25518
rect 4284 25414 4340 25452
rect 8652 25284 8708 25566
rect 9548 26178 9604 26190
rect 9548 26126 9550 26178
rect 9602 26126 9604 26178
rect 9548 25508 9604 26126
rect 9548 25442 9604 25452
rect 11564 25506 11620 26236
rect 12460 26292 12516 26302
rect 12460 26198 12516 26236
rect 12908 26180 12964 26348
rect 12908 26086 12964 26124
rect 12124 25732 12180 25742
rect 12124 25730 12740 25732
rect 12124 25678 12126 25730
rect 12178 25678 12740 25730
rect 12124 25676 12740 25678
rect 12124 25666 12180 25676
rect 11564 25454 11566 25506
rect 11618 25454 11620 25506
rect 11564 25442 11620 25454
rect 10780 25396 10836 25406
rect 10780 25302 10836 25340
rect 12236 25394 12292 25406
rect 12236 25342 12238 25394
rect 12290 25342 12292 25394
rect 8652 25218 8708 25228
rect 12124 25284 12180 25294
rect 12236 25284 12292 25342
rect 12460 25396 12516 25406
rect 12460 25302 12516 25340
rect 12684 25394 12740 25676
rect 13580 25730 13636 26796
rect 15036 26180 15092 26190
rect 14924 26178 15092 26180
rect 14924 26126 15038 26178
rect 15090 26126 15092 26178
rect 14924 26124 15092 26126
rect 14252 25844 14308 25854
rect 13580 25678 13582 25730
rect 13634 25678 13636 25730
rect 13580 25666 13636 25678
rect 14140 25732 14196 25742
rect 13468 25620 13524 25630
rect 14140 25620 14196 25676
rect 12796 25508 12852 25518
rect 12796 25414 12852 25452
rect 12684 25342 12686 25394
rect 12738 25342 12740 25394
rect 12684 25330 12740 25342
rect 13468 25396 13524 25564
rect 13692 25618 14196 25620
rect 13692 25566 14142 25618
rect 14194 25566 14196 25618
rect 13692 25564 14196 25566
rect 13692 25506 13748 25564
rect 14140 25554 14196 25564
rect 13692 25454 13694 25506
rect 13746 25454 13748 25506
rect 13580 25396 13636 25406
rect 13468 25394 13636 25396
rect 13468 25342 13582 25394
rect 13634 25342 13636 25394
rect 13468 25340 13636 25342
rect 13580 25330 13636 25340
rect 12348 25284 12404 25294
rect 12236 25228 12348 25284
rect 12124 25190 12180 25228
rect 12348 25218 12404 25228
rect 13132 25284 13188 25294
rect 1932 24948 1988 24958
rect 1932 24610 1988 24892
rect 4284 24948 4340 24958
rect 4284 24722 4340 24892
rect 4732 24948 4788 24958
rect 4732 24854 4788 24892
rect 13132 24946 13188 25228
rect 13692 25284 13748 25454
rect 13692 25218 13748 25228
rect 13132 24894 13134 24946
rect 13186 24894 13188 24946
rect 13132 24882 13188 24894
rect 14252 24948 14308 25788
rect 14924 25506 14980 26124
rect 15036 26114 15092 26124
rect 15260 26068 15316 28252
rect 15596 28196 15652 28812
rect 15708 28754 15764 28812
rect 15708 28702 15710 28754
rect 15762 28702 15764 28754
rect 15708 28690 15764 28702
rect 16380 28756 16436 29374
rect 17388 29428 17444 29438
rect 17388 29334 17444 29372
rect 16380 28662 16436 28700
rect 16716 29314 16772 29326
rect 16716 29262 16718 29314
rect 16770 29262 16772 29314
rect 16716 28532 16772 29262
rect 16716 28466 16772 28476
rect 17052 29316 17108 29326
rect 16940 28420 16996 28430
rect 16940 28326 16996 28364
rect 15596 28140 16324 28196
rect 15596 27858 15652 28140
rect 16268 28082 16324 28140
rect 16268 28030 16270 28082
rect 16322 28030 16324 28082
rect 16268 28018 16324 28030
rect 15820 27972 15876 27982
rect 15820 27878 15876 27916
rect 15596 27806 15598 27858
rect 15650 27806 15652 27858
rect 15596 27794 15652 27806
rect 16268 27300 16324 27310
rect 16268 27206 16324 27244
rect 15260 26002 15316 26012
rect 15484 27188 15540 27198
rect 14924 25454 14926 25506
rect 14978 25454 14980 25506
rect 14924 25442 14980 25454
rect 15260 25508 15316 25518
rect 15484 25508 15540 27132
rect 16604 27186 16660 27198
rect 16604 27134 16606 27186
rect 16658 27134 16660 27186
rect 16492 26962 16548 26974
rect 16492 26910 16494 26962
rect 16546 26910 16548 26962
rect 16268 26404 16324 26414
rect 16268 26310 16324 26348
rect 16492 26404 16548 26910
rect 16492 26338 16548 26348
rect 15708 26292 15764 26302
rect 15708 26198 15764 26236
rect 16044 26290 16100 26302
rect 16044 26238 16046 26290
rect 16098 26238 16100 26290
rect 15260 25506 15540 25508
rect 15260 25454 15262 25506
rect 15314 25454 15540 25506
rect 15260 25452 15540 25454
rect 15260 25442 15316 25452
rect 15148 25284 15204 25294
rect 16044 25284 16100 26238
rect 15148 25282 16100 25284
rect 15148 25230 15150 25282
rect 15202 25230 16100 25282
rect 15148 25228 16100 25230
rect 16380 26290 16436 26302
rect 16380 26238 16382 26290
rect 16434 26238 16436 26290
rect 16380 25284 16436 26238
rect 16604 25508 16660 27134
rect 17052 27074 17108 29260
rect 17500 29316 17556 29326
rect 17500 29222 17556 29260
rect 17836 29092 17892 30156
rect 17948 30098 18004 30380
rect 20188 30436 20244 30446
rect 20188 30322 20244 30380
rect 20188 30270 20190 30322
rect 20242 30270 20244 30322
rect 20188 30258 20244 30270
rect 19740 30212 19796 30222
rect 19628 30156 19740 30212
rect 17948 30046 17950 30098
rect 18002 30046 18004 30098
rect 17948 30034 18004 30046
rect 19292 30098 19348 30110
rect 19292 30046 19294 30098
rect 19346 30046 19348 30098
rect 18732 29652 18788 29662
rect 17500 29036 17892 29092
rect 18060 29426 18116 29438
rect 18060 29374 18062 29426
rect 18114 29374 18116 29426
rect 17500 28530 17556 29036
rect 18060 28980 18116 29374
rect 18396 29428 18452 29438
rect 18396 29334 18452 29372
rect 18620 29426 18676 29438
rect 18620 29374 18622 29426
rect 18674 29374 18676 29426
rect 18060 28914 18116 28924
rect 18508 29314 18564 29326
rect 18508 29262 18510 29314
rect 18562 29262 18564 29314
rect 18172 28866 18228 28878
rect 18508 28868 18564 29262
rect 18620 29204 18676 29374
rect 18620 29138 18676 29148
rect 18172 28814 18174 28866
rect 18226 28814 18228 28866
rect 18172 28756 18228 28814
rect 17724 28700 18228 28756
rect 18284 28812 18564 28868
rect 17724 28642 17780 28700
rect 17724 28590 17726 28642
rect 17778 28590 17780 28642
rect 17724 28578 17780 28590
rect 17500 28478 17502 28530
rect 17554 28478 17556 28530
rect 17500 28466 17556 28478
rect 18060 28532 18116 28542
rect 18060 28438 18116 28476
rect 17052 27022 17054 27074
rect 17106 27022 17108 27074
rect 17052 27010 17108 27022
rect 17276 28420 17332 28430
rect 17276 28084 17332 28364
rect 17612 28420 17668 28430
rect 18172 28420 18228 28430
rect 17612 28418 17780 28420
rect 17612 28366 17614 28418
rect 17666 28366 17780 28418
rect 17612 28364 17780 28366
rect 17612 28354 17668 28364
rect 17500 28084 17556 28094
rect 17276 28028 17500 28084
rect 17164 26908 17220 26918
rect 17276 26908 17332 28028
rect 17500 27990 17556 28028
rect 17164 26906 17332 26908
rect 17164 26854 17166 26906
rect 17218 26854 17332 26906
rect 17388 26964 17444 26974
rect 17612 26964 17668 26974
rect 17388 26962 17668 26964
rect 17388 26910 17390 26962
rect 17442 26910 17614 26962
rect 17666 26910 17668 26962
rect 17388 26908 17668 26910
rect 17388 26898 17444 26908
rect 17612 26898 17668 26908
rect 17164 26852 17332 26854
rect 17164 26842 17220 26852
rect 17164 26628 17220 26638
rect 16828 26404 16884 26414
rect 16828 26310 16884 26348
rect 16604 25442 16660 25452
rect 16716 25732 16772 25742
rect 16604 25284 16660 25294
rect 16716 25284 16772 25676
rect 17164 25394 17220 26572
rect 17724 26402 17780 28364
rect 18172 28326 18228 28364
rect 18284 28196 18340 28812
rect 18732 28754 18788 29596
rect 18956 29426 19012 29438
rect 18956 29374 18958 29426
rect 19010 29374 19012 29426
rect 18956 29204 19012 29374
rect 19292 29428 19348 30046
rect 19628 29876 19684 30156
rect 19740 30118 19796 30156
rect 19628 29810 19684 29820
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 19964 29540 20020 29550
rect 19292 29334 19348 29372
rect 19516 29426 19572 29438
rect 19964 29428 20020 29484
rect 19516 29374 19518 29426
rect 19570 29374 19572 29426
rect 19404 29314 19460 29326
rect 19404 29262 19406 29314
rect 19458 29262 19460 29314
rect 19404 29204 19460 29262
rect 18956 29148 19460 29204
rect 19516 29204 19572 29374
rect 19516 29138 19572 29148
rect 19628 29426 20020 29428
rect 19628 29374 19966 29426
rect 20018 29374 20020 29426
rect 19628 29372 20020 29374
rect 19628 28868 19684 29372
rect 19964 29362 20020 29372
rect 20524 29092 20580 35308
rect 20860 34244 20916 35646
rect 20860 34178 20916 34188
rect 20972 34018 21028 34030
rect 20972 33966 20974 34018
rect 21026 33966 21028 34018
rect 20972 33348 21028 33966
rect 20972 33282 21028 33292
rect 20972 30996 21028 31006
rect 20972 30902 21028 30940
rect 21196 29764 21252 41804
rect 21980 41860 22036 41870
rect 21980 41766 22036 41804
rect 22652 41860 22708 41918
rect 22652 41794 22708 41804
rect 22876 42530 22932 42542
rect 22876 42478 22878 42530
rect 22930 42478 22932 42530
rect 21420 41186 21476 41198
rect 21420 41134 21422 41186
rect 21474 41134 21476 41186
rect 21420 41076 21476 41134
rect 21420 41010 21476 41020
rect 21644 41186 21700 41198
rect 21644 41134 21646 41186
rect 21698 41134 21700 41186
rect 21644 40628 21700 41134
rect 22876 41188 22932 42478
rect 23212 41298 23268 42588
rect 23436 42642 23492 43260
rect 23660 42754 23716 43374
rect 23996 43316 24052 43326
rect 23996 43314 24276 43316
rect 23996 43262 23998 43314
rect 24050 43262 24276 43314
rect 23996 43260 24276 43262
rect 23996 43250 24052 43260
rect 23660 42702 23662 42754
rect 23714 42702 23716 42754
rect 23660 42690 23716 42702
rect 23436 42590 23438 42642
rect 23490 42590 23492 42642
rect 23436 42578 23492 42590
rect 23324 41972 23380 41982
rect 23324 41878 23380 41916
rect 23660 41972 23716 41982
rect 23660 41878 23716 41916
rect 23212 41246 23214 41298
rect 23266 41246 23268 41298
rect 23212 41234 23268 41246
rect 23436 41858 23492 41870
rect 23436 41806 23438 41858
rect 23490 41806 23492 41858
rect 23100 41188 23156 41198
rect 22876 41132 23100 41188
rect 23100 41094 23156 41132
rect 22316 41076 22372 41086
rect 22316 40982 22372 41020
rect 21644 40562 21700 40572
rect 22428 40964 22484 40974
rect 21532 40516 21588 40526
rect 21532 40422 21588 40460
rect 22428 40402 22484 40908
rect 22764 40626 22820 40638
rect 22764 40574 22766 40626
rect 22818 40574 22820 40626
rect 22428 40350 22430 40402
rect 22482 40350 22484 40402
rect 22428 40338 22484 40350
rect 22652 40404 22708 40414
rect 22540 39730 22596 39742
rect 22540 39678 22542 39730
rect 22594 39678 22596 39730
rect 21980 39620 22036 39630
rect 21868 39508 21924 39518
rect 21868 38834 21924 39452
rect 21980 39506 22036 39564
rect 21980 39454 21982 39506
rect 22034 39454 22036 39506
rect 21980 38946 22036 39454
rect 22540 39508 22596 39678
rect 22540 39442 22596 39452
rect 21980 38894 21982 38946
rect 22034 38894 22036 38946
rect 21980 38882 22036 38894
rect 22204 39394 22260 39406
rect 22204 39342 22206 39394
rect 22258 39342 22260 39394
rect 21868 38782 21870 38834
rect 21922 38782 21924 38834
rect 21868 38770 21924 38782
rect 21532 38722 21588 38734
rect 21532 38670 21534 38722
rect 21586 38670 21588 38722
rect 21308 36708 21364 36718
rect 21308 36594 21364 36652
rect 21308 36542 21310 36594
rect 21362 36542 21364 36594
rect 21308 36530 21364 36542
rect 21532 36484 21588 38670
rect 21868 38162 21924 38174
rect 21868 38110 21870 38162
rect 21922 38110 21924 38162
rect 21532 36390 21588 36428
rect 21756 36596 21812 36606
rect 21756 36482 21812 36540
rect 21756 36430 21758 36482
rect 21810 36430 21812 36482
rect 21756 35698 21812 36430
rect 21756 35646 21758 35698
rect 21810 35646 21812 35698
rect 21756 35634 21812 35646
rect 21868 35364 21924 38110
rect 21980 38164 22036 38174
rect 21980 38070 22036 38108
rect 22204 38050 22260 39342
rect 22316 39396 22372 39406
rect 22316 38834 22372 39340
rect 22316 38782 22318 38834
rect 22370 38782 22372 38834
rect 22316 38770 22372 38782
rect 22540 38836 22596 38846
rect 22652 38836 22708 40348
rect 22540 38834 22708 38836
rect 22540 38782 22542 38834
rect 22594 38782 22708 38834
rect 22540 38780 22708 38782
rect 22764 39618 22820 40574
rect 23324 40402 23380 40414
rect 23324 40350 23326 40402
rect 23378 40350 23380 40402
rect 22764 39566 22766 39618
rect 22818 39566 22820 39618
rect 22764 38834 22820 39566
rect 23100 39618 23156 39630
rect 23100 39566 23102 39618
rect 23154 39566 23156 39618
rect 23100 39396 23156 39566
rect 23324 39620 23380 40350
rect 23436 40404 23492 41806
rect 23660 41076 23716 41086
rect 23548 40516 23604 40526
rect 23548 40422 23604 40460
rect 23660 40514 23716 41020
rect 23660 40462 23662 40514
rect 23714 40462 23716 40514
rect 23660 40450 23716 40462
rect 23996 41074 24052 41086
rect 23996 41022 23998 41074
rect 24050 41022 24052 41074
rect 23436 39730 23492 40348
rect 23436 39678 23438 39730
rect 23490 39678 23492 39730
rect 23436 39666 23492 39678
rect 23324 39554 23380 39564
rect 23100 39330 23156 39340
rect 23660 39508 23716 39518
rect 23660 38946 23716 39452
rect 23660 38894 23662 38946
rect 23714 38894 23716 38946
rect 23660 38882 23716 38894
rect 22764 38782 22766 38834
rect 22818 38782 22820 38834
rect 22540 38770 22596 38780
rect 22764 38770 22820 38782
rect 23212 38836 23268 38846
rect 23436 38836 23492 38846
rect 23212 38834 23492 38836
rect 23212 38782 23214 38834
rect 23266 38782 23438 38834
rect 23490 38782 23492 38834
rect 23212 38780 23492 38782
rect 23212 38770 23268 38780
rect 23436 38770 23492 38780
rect 23548 38724 23604 38762
rect 23996 38668 24052 41022
rect 23548 38658 23604 38668
rect 22204 37998 22206 38050
rect 22258 37998 22260 38050
rect 22204 37986 22260 37998
rect 23660 38612 24052 38668
rect 23212 37492 23268 37502
rect 22092 36708 22148 36718
rect 21980 36484 22036 36494
rect 21980 35586 22036 36428
rect 22092 35698 22148 36652
rect 23212 36594 23268 37436
rect 23548 37492 23604 37502
rect 23324 37268 23380 37278
rect 23380 37212 23492 37268
rect 23324 37174 23380 37212
rect 23436 36706 23492 37212
rect 23548 37266 23604 37436
rect 23548 37214 23550 37266
rect 23602 37214 23604 37266
rect 23548 37202 23604 37214
rect 23436 36654 23438 36706
rect 23490 36654 23492 36706
rect 23436 36642 23492 36654
rect 23212 36542 23214 36594
rect 23266 36542 23268 36594
rect 23212 36530 23268 36542
rect 22204 36484 22260 36494
rect 22652 36484 22708 36494
rect 22204 36482 22708 36484
rect 22204 36430 22206 36482
rect 22258 36430 22654 36482
rect 22706 36430 22708 36482
rect 22204 36428 22708 36430
rect 22204 36418 22260 36428
rect 22652 36418 22708 36428
rect 22316 36260 22372 36270
rect 22092 35646 22094 35698
rect 22146 35646 22148 35698
rect 22092 35634 22148 35646
rect 22204 36258 22372 36260
rect 22204 36206 22318 36258
rect 22370 36206 22372 36258
rect 22204 36204 22372 36206
rect 21980 35534 21982 35586
rect 22034 35534 22036 35586
rect 21980 35522 22036 35534
rect 21868 35298 21924 35308
rect 22204 34916 22260 36204
rect 22316 36194 22372 36204
rect 22540 36258 22596 36270
rect 22540 36206 22542 36258
rect 22594 36206 22596 36258
rect 22540 35810 22596 36206
rect 23660 36036 23716 38612
rect 23884 38050 23940 38062
rect 23884 37998 23886 38050
rect 23938 37998 23940 38050
rect 23884 37828 23940 37998
rect 24108 38052 24164 38062
rect 24108 37958 24164 37996
rect 23884 37762 23940 37772
rect 23996 37044 24052 37054
rect 23996 36950 24052 36988
rect 23772 36372 23828 36382
rect 23996 36372 24052 36382
rect 23772 36370 24052 36372
rect 23772 36318 23774 36370
rect 23826 36318 23998 36370
rect 24050 36318 24052 36370
rect 23772 36316 24052 36318
rect 23772 36306 23828 36316
rect 23996 36306 24052 36316
rect 23436 35980 23716 36036
rect 24220 36036 24276 43260
rect 24332 38948 24388 43708
rect 24332 38274 24388 38892
rect 25452 38948 25508 38958
rect 25452 38854 25508 38892
rect 24332 38222 24334 38274
rect 24386 38222 24388 38274
rect 24332 38210 24388 38222
rect 25228 38722 25284 38734
rect 25228 38670 25230 38722
rect 25282 38670 25284 38722
rect 25004 38052 25060 38062
rect 25004 37958 25060 37996
rect 24444 37938 24500 37950
rect 24444 37886 24446 37938
rect 24498 37886 24500 37938
rect 24444 37268 24500 37886
rect 25228 37828 25284 38670
rect 25564 38610 25620 38622
rect 25564 38558 25566 38610
rect 25618 38558 25620 38610
rect 25564 38162 25620 38558
rect 25564 38110 25566 38162
rect 25618 38110 25620 38162
rect 25564 38098 25620 38110
rect 25228 37762 25284 37772
rect 25900 37938 25956 37950
rect 25900 37886 25902 37938
rect 25954 37886 25956 37938
rect 25900 37378 25956 37886
rect 25900 37326 25902 37378
rect 25954 37326 25956 37378
rect 24444 37202 24500 37212
rect 25228 37268 25284 37278
rect 25228 37174 25284 37212
rect 25788 37266 25844 37278
rect 25788 37214 25790 37266
rect 25842 37214 25844 37266
rect 24556 37044 24612 37054
rect 24556 36706 24612 36988
rect 24556 36654 24558 36706
rect 24610 36654 24612 36706
rect 24556 36642 24612 36654
rect 25340 37044 25396 37054
rect 25340 36594 25396 36988
rect 25788 37044 25844 37214
rect 25788 36978 25844 36988
rect 25340 36542 25342 36594
rect 25394 36542 25396 36594
rect 25340 36530 25396 36542
rect 24332 36482 24388 36494
rect 24332 36430 24334 36482
rect 24386 36430 24388 36482
rect 24332 36370 24388 36430
rect 24780 36484 24836 36494
rect 25788 36484 25844 36494
rect 25900 36484 25956 37326
rect 24780 36482 24948 36484
rect 24780 36430 24782 36482
rect 24834 36430 24948 36482
rect 24780 36428 24948 36430
rect 24780 36418 24836 36428
rect 24332 36318 24334 36370
rect 24386 36318 24388 36370
rect 24332 36306 24388 36318
rect 24444 36260 24500 36270
rect 24444 36258 24724 36260
rect 24444 36206 24446 36258
rect 24498 36206 24724 36258
rect 24444 36204 24724 36206
rect 24444 36194 24500 36204
rect 24220 35980 24612 36036
rect 23436 35924 23492 35980
rect 22540 35758 22542 35810
rect 22594 35758 22596 35810
rect 21868 34860 22260 34916
rect 22316 35028 22372 35038
rect 22316 34916 22372 34972
rect 22428 34916 22484 34926
rect 22316 34914 22484 34916
rect 22316 34862 22430 34914
rect 22482 34862 22484 34914
rect 22316 34860 22484 34862
rect 21644 34804 21700 34814
rect 21644 34354 21700 34748
rect 21644 34302 21646 34354
rect 21698 34302 21700 34354
rect 21644 34290 21700 34302
rect 21532 34244 21588 34254
rect 21532 34150 21588 34188
rect 21420 34130 21476 34142
rect 21420 34078 21422 34130
rect 21474 34078 21476 34130
rect 21420 33348 21476 34078
rect 21420 33282 21476 33292
rect 21420 31108 21476 31118
rect 21420 30436 21476 31052
rect 21868 31108 21924 34860
rect 22092 34692 22148 34702
rect 22316 34692 22372 34860
rect 22428 34850 22484 34860
rect 22092 34690 22372 34692
rect 22092 34638 22094 34690
rect 22146 34638 22372 34690
rect 22092 34636 22372 34638
rect 22092 34626 22148 34636
rect 21980 34412 22484 34468
rect 21980 34130 22036 34412
rect 22316 34244 22372 34254
rect 22316 34150 22372 34188
rect 22428 34244 22484 34412
rect 22540 34244 22596 35758
rect 23324 35922 23492 35924
rect 23324 35870 23438 35922
rect 23490 35870 23492 35922
rect 23324 35868 23492 35870
rect 22764 35026 22820 35038
rect 22764 34974 22766 35026
rect 22818 34974 22820 35026
rect 22764 34916 22820 34974
rect 22764 34850 22820 34860
rect 22988 35028 23044 35038
rect 22652 34804 22708 34814
rect 22652 34710 22708 34748
rect 22988 34356 23044 34972
rect 23324 34804 23380 35868
rect 23436 35858 23492 35868
rect 24556 35922 24612 35980
rect 24556 35870 24558 35922
rect 24610 35870 24612 35922
rect 23548 35698 23604 35710
rect 23548 35646 23550 35698
rect 23602 35646 23604 35698
rect 23548 35588 23604 35646
rect 24444 35698 24500 35710
rect 24444 35646 24446 35698
rect 24498 35646 24500 35698
rect 23996 35588 24052 35598
rect 23548 35586 24052 35588
rect 23548 35534 23998 35586
rect 24050 35534 24052 35586
rect 23548 35532 24052 35534
rect 23436 35474 23492 35486
rect 23436 35422 23438 35474
rect 23490 35422 23492 35474
rect 23436 34914 23492 35422
rect 23548 35028 23604 35532
rect 23996 35522 24052 35532
rect 24444 35140 24500 35646
rect 24444 35074 24500 35084
rect 23548 34962 23604 34972
rect 23436 34862 23438 34914
rect 23490 34862 23492 34914
rect 23436 34850 23492 34862
rect 23772 34916 23828 34926
rect 23772 34822 23828 34860
rect 24332 34914 24388 34926
rect 24332 34862 24334 34914
rect 24386 34862 24388 34914
rect 23324 34692 23380 34748
rect 23884 34802 23940 34814
rect 23884 34750 23886 34802
rect 23938 34750 23940 34802
rect 23324 34636 23716 34692
rect 22988 34354 23492 34356
rect 22988 34302 22990 34354
rect 23042 34302 23492 34354
rect 22988 34300 23492 34302
rect 22988 34290 23044 34300
rect 22428 34242 22596 34244
rect 22428 34190 22430 34242
rect 22482 34190 22596 34242
rect 22428 34188 22596 34190
rect 22428 34178 22484 34188
rect 21980 34078 21982 34130
rect 22034 34078 22036 34130
rect 21980 34066 22036 34078
rect 23436 34130 23492 34300
rect 23436 34078 23438 34130
rect 23490 34078 23492 34130
rect 23436 34066 23492 34078
rect 23660 34130 23716 34636
rect 23660 34078 23662 34130
rect 23714 34078 23716 34130
rect 23660 34066 23716 34078
rect 22316 33906 22372 33918
rect 22316 33854 22318 33906
rect 22370 33854 22372 33906
rect 22316 33346 22372 33854
rect 22316 33294 22318 33346
rect 22370 33294 22372 33346
rect 22316 32562 22372 33294
rect 22316 32510 22318 32562
rect 22370 32510 22372 32562
rect 22316 32498 22372 32510
rect 22540 33348 22596 33358
rect 22540 32562 22596 33292
rect 22764 33236 22820 33246
rect 22764 33234 23156 33236
rect 22764 33182 22766 33234
rect 22818 33182 23156 33234
rect 22764 33180 23156 33182
rect 22764 33170 22820 33180
rect 22540 32510 22542 32562
rect 22594 32510 22596 32562
rect 22540 32498 22596 32510
rect 22764 32450 22820 32462
rect 22764 32398 22766 32450
rect 22818 32398 22820 32450
rect 21980 31108 22036 31118
rect 21924 31106 22036 31108
rect 21924 31054 21982 31106
rect 22034 31054 22036 31106
rect 21924 31052 22036 31054
rect 21868 31014 21924 31052
rect 21980 31042 22036 31052
rect 22092 31106 22148 31118
rect 22092 31054 22094 31106
rect 22146 31054 22148 31106
rect 22092 30996 22148 31054
rect 22652 30996 22708 31006
rect 22092 30940 22484 30996
rect 21644 30884 21700 30894
rect 21644 30790 21700 30828
rect 22092 30772 22148 30782
rect 22092 30770 22260 30772
rect 22092 30718 22094 30770
rect 22146 30718 22260 30770
rect 22092 30716 22260 30718
rect 22092 30706 22148 30716
rect 21420 30342 21476 30380
rect 21756 30322 21812 30334
rect 21756 30270 21758 30322
rect 21810 30270 21812 30322
rect 21532 30212 21588 30222
rect 21756 30212 21812 30270
rect 22092 30212 22148 30222
rect 21756 30210 22148 30212
rect 21756 30158 22094 30210
rect 22146 30158 22148 30210
rect 21756 30156 22148 30158
rect 21532 29988 21588 30156
rect 21644 29988 21700 29998
rect 21532 29986 21700 29988
rect 21532 29934 21646 29986
rect 21698 29934 21700 29986
rect 21532 29932 21700 29934
rect 21644 29922 21700 29932
rect 21196 29708 21812 29764
rect 21420 29426 21476 29438
rect 21420 29374 21422 29426
rect 21474 29374 21476 29426
rect 18732 28702 18734 28754
rect 18786 28702 18788 28754
rect 18732 28644 18788 28702
rect 18732 28578 18788 28588
rect 19404 28812 19684 28868
rect 20076 29036 20580 29092
rect 20636 29316 20692 29326
rect 21084 29316 21140 29326
rect 21420 29316 21476 29374
rect 20636 29314 21420 29316
rect 20636 29262 20638 29314
rect 20690 29262 21086 29314
rect 21138 29262 21420 29314
rect 20636 29260 21420 29262
rect 18172 28140 18340 28196
rect 18060 27972 18116 27982
rect 18060 27878 18116 27916
rect 17948 27860 18004 27870
rect 17948 27766 18004 27804
rect 17948 27188 18004 27198
rect 17948 27094 18004 27132
rect 18172 27074 18228 28140
rect 18956 27972 19012 27982
rect 18956 27878 19012 27916
rect 18508 27860 18564 27870
rect 18732 27860 18788 27870
rect 18508 27858 18788 27860
rect 18508 27806 18510 27858
rect 18562 27806 18734 27858
rect 18786 27806 18788 27858
rect 18508 27804 18788 27806
rect 18508 27794 18564 27804
rect 18172 27022 18174 27074
rect 18226 27022 18228 27074
rect 18172 27010 18228 27022
rect 18284 27746 18340 27758
rect 18284 27694 18286 27746
rect 18338 27694 18340 27746
rect 17724 26350 17726 26402
rect 17778 26350 17780 26402
rect 17724 26338 17780 26350
rect 17836 26292 17892 26302
rect 17388 25620 17444 25630
rect 17388 25526 17444 25564
rect 17836 25620 17892 26236
rect 18284 26290 18340 27694
rect 18732 27748 18788 27804
rect 18844 27860 18900 27870
rect 18844 27766 18900 27804
rect 19404 27858 19460 28812
rect 20076 28532 20132 29036
rect 20188 28868 20244 28878
rect 20636 28868 20692 29260
rect 21084 29250 21140 29260
rect 21420 29222 21476 29260
rect 21532 29092 21588 29708
rect 21756 29538 21812 29708
rect 21756 29486 21758 29538
rect 21810 29486 21812 29538
rect 20244 28812 20692 28868
rect 20188 28754 20244 28812
rect 20188 28702 20190 28754
rect 20242 28702 20244 28754
rect 20188 28690 20244 28702
rect 20412 28644 20468 28654
rect 20412 28550 20468 28588
rect 20076 28466 20132 28476
rect 20636 28530 20692 28812
rect 20748 29036 21588 29092
rect 21644 29314 21700 29326
rect 21644 29262 21646 29314
rect 21698 29262 21700 29314
rect 20748 28642 20804 29036
rect 20748 28590 20750 28642
rect 20802 28590 20804 28642
rect 20748 28578 20804 28590
rect 20636 28478 20638 28530
rect 20690 28478 20692 28530
rect 20636 28466 20692 28478
rect 21420 28418 21476 28430
rect 21420 28366 21422 28418
rect 21474 28366 21476 28418
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 20748 28084 20804 28094
rect 21420 28084 21476 28366
rect 20748 28082 21476 28084
rect 20748 28030 20750 28082
rect 20802 28030 21422 28082
rect 21474 28030 21476 28082
rect 20748 28028 21476 28030
rect 20748 28018 20804 28028
rect 21420 28018 21476 28028
rect 21644 28420 21700 29262
rect 21756 28866 21812 29486
rect 22092 29428 22148 30156
rect 22204 30100 22260 30716
rect 22204 29650 22260 30044
rect 22204 29598 22206 29650
rect 22258 29598 22260 29650
rect 22204 29586 22260 29598
rect 22316 30210 22372 30222
rect 22316 30158 22318 30210
rect 22370 30158 22372 30210
rect 22316 29428 22372 30158
rect 22428 30212 22484 30940
rect 22428 30146 22484 30156
rect 22540 30940 22652 30996
rect 22764 30996 22820 32398
rect 22988 32116 23044 32126
rect 22876 30996 22932 31006
rect 22764 30994 22932 30996
rect 22764 30942 22878 30994
rect 22930 30942 22932 30994
rect 22764 30940 22932 30942
rect 22540 29650 22596 30940
rect 22652 30930 22708 30940
rect 22876 30930 22932 30940
rect 22540 29598 22542 29650
rect 22594 29598 22596 29650
rect 22540 29586 22596 29598
rect 22428 29428 22484 29438
rect 22316 29426 22484 29428
rect 22316 29374 22430 29426
rect 22482 29374 22484 29426
rect 22316 29372 22484 29374
rect 22092 29362 22148 29372
rect 21756 28814 21758 28866
rect 21810 28814 21812 28866
rect 21756 28802 21812 28814
rect 21980 29316 22036 29326
rect 21980 28754 22036 29260
rect 22428 29204 22484 29372
rect 22652 29428 22708 29438
rect 22652 29334 22708 29372
rect 22428 29138 22484 29148
rect 22988 28980 23044 32060
rect 23100 30210 23156 33180
rect 23212 32788 23268 32798
rect 23212 32674 23268 32732
rect 23884 32676 23940 34750
rect 24332 34804 24388 34862
rect 24556 34916 24612 35870
rect 24556 34850 24612 34860
rect 24332 34738 24388 34748
rect 24332 34132 24388 34142
rect 24332 34038 24388 34076
rect 23212 32622 23214 32674
rect 23266 32622 23268 32674
rect 23212 32610 23268 32622
rect 23660 32620 23940 32676
rect 24668 32676 24724 36204
rect 24780 35700 24836 35710
rect 24780 35606 24836 35644
rect 24892 35028 24948 36428
rect 25788 36482 25956 36484
rect 25788 36430 25790 36482
rect 25842 36430 25956 36482
rect 25788 36428 25956 36430
rect 26012 37154 26068 37166
rect 26012 37102 26014 37154
rect 26066 37102 26068 37154
rect 25788 36418 25844 36428
rect 25340 35700 25396 35710
rect 25340 35606 25396 35644
rect 26012 35588 26068 37102
rect 26236 36372 26292 36382
rect 26236 36278 26292 36316
rect 25900 35586 26068 35588
rect 25900 35534 26014 35586
rect 26066 35534 26068 35586
rect 25900 35532 26068 35534
rect 25564 35474 25620 35486
rect 25564 35422 25566 35474
rect 25618 35422 25620 35474
rect 25116 35140 25172 35150
rect 25172 35084 25284 35140
rect 25116 35074 25172 35084
rect 24892 34962 24948 34972
rect 25228 35026 25284 35084
rect 25228 34974 25230 35026
rect 25282 34974 25284 35026
rect 25228 34962 25284 34974
rect 25340 34916 25396 34926
rect 25340 34822 25396 34860
rect 25564 34804 25620 35422
rect 25452 34356 25508 34366
rect 25564 34356 25620 34748
rect 25900 34468 25956 35532
rect 26012 35522 26068 35532
rect 26124 35698 26180 35710
rect 26124 35646 26126 35698
rect 26178 35646 26180 35698
rect 26012 34916 26068 34926
rect 26124 34916 26180 35646
rect 26012 34914 26124 34916
rect 26012 34862 26014 34914
rect 26066 34862 26124 34914
rect 26012 34860 26124 34862
rect 26012 34850 26068 34860
rect 25900 34402 25956 34412
rect 25452 34354 25620 34356
rect 25452 34302 25454 34354
rect 25506 34302 25620 34354
rect 25452 34300 25620 34302
rect 25452 34290 25508 34300
rect 24892 34132 24948 34142
rect 24892 33346 24948 34076
rect 25228 34132 25284 34142
rect 25228 34038 25284 34076
rect 25340 34018 25396 34030
rect 25340 33966 25342 34018
rect 25394 33966 25396 34018
rect 25340 33572 25396 33966
rect 25340 33516 25508 33572
rect 24892 33294 24894 33346
rect 24946 33294 24948 33346
rect 24892 33282 24948 33294
rect 25452 33346 25508 33516
rect 25452 33294 25454 33346
rect 25506 33294 25508 33346
rect 25452 33282 25508 33294
rect 25340 33234 25396 33246
rect 25340 33182 25342 33234
rect 25394 33182 25396 33234
rect 25116 33122 25172 33134
rect 25116 33070 25118 33122
rect 25170 33070 25172 33122
rect 24668 32620 24836 32676
rect 23324 32452 23380 32462
rect 23324 32358 23380 32396
rect 23100 30158 23102 30210
rect 23154 30158 23156 30210
rect 23100 30146 23156 30158
rect 23212 31218 23268 31230
rect 23212 31166 23214 31218
rect 23266 31166 23268 31218
rect 23212 30212 23268 31166
rect 23548 31108 23604 31118
rect 23548 31014 23604 31052
rect 23324 30996 23380 31006
rect 23324 30902 23380 30940
rect 23548 30324 23604 30334
rect 23548 30230 23604 30268
rect 23212 30146 23268 30156
rect 23324 30210 23380 30222
rect 23324 30158 23326 30210
rect 23378 30158 23380 30210
rect 23324 30100 23380 30158
rect 23324 30034 23380 30044
rect 21980 28702 21982 28754
rect 22034 28702 22036 28754
rect 21980 28690 22036 28702
rect 22204 28924 23044 28980
rect 19404 27806 19406 27858
rect 19458 27806 19460 27858
rect 19404 27794 19460 27806
rect 21644 27970 21700 28364
rect 21644 27918 21646 27970
rect 21698 27918 21700 27970
rect 18732 27682 18788 27692
rect 20636 27748 20692 27758
rect 20636 27654 20692 27692
rect 21532 27748 21588 27758
rect 21532 27654 21588 27692
rect 20972 27636 21028 27646
rect 20972 27634 21476 27636
rect 20972 27582 20974 27634
rect 21026 27582 21476 27634
rect 20972 27580 21476 27582
rect 20972 27570 21028 27580
rect 18620 27074 18676 27086
rect 18620 27022 18622 27074
rect 18674 27022 18676 27074
rect 18620 26292 18676 27022
rect 19180 27076 19236 27086
rect 18284 26238 18286 26290
rect 18338 26238 18340 26290
rect 18284 26226 18340 26238
rect 18396 26290 18676 26292
rect 18396 26238 18622 26290
rect 18674 26238 18676 26290
rect 18396 26236 18676 26238
rect 17276 25508 17332 25518
rect 17276 25414 17332 25452
rect 17164 25342 17166 25394
rect 17218 25342 17220 25394
rect 17164 25330 17220 25342
rect 16380 25282 16772 25284
rect 16380 25230 16606 25282
rect 16658 25230 16772 25282
rect 16380 25228 16772 25230
rect 15148 25218 15204 25228
rect 16604 25218 16660 25228
rect 14252 24882 14308 24892
rect 11900 24724 11956 24734
rect 4284 24670 4286 24722
rect 4338 24670 4340 24722
rect 4284 24658 4340 24670
rect 11788 24722 11956 24724
rect 11788 24670 11902 24722
rect 11954 24670 11956 24722
rect 11788 24668 11956 24670
rect 1932 24558 1934 24610
rect 1986 24558 1988 24610
rect 1932 24546 1988 24558
rect 5292 24610 5348 24622
rect 5292 24558 5294 24610
rect 5346 24558 5348 24610
rect 5292 24388 5348 24558
rect 4476 24332 4740 24342
rect 1932 24276 1988 24286
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 1932 24162 1988 24220
rect 1932 24110 1934 24162
rect 1986 24110 1988 24162
rect 1932 24098 1988 24110
rect 4284 24052 4340 24062
rect 4284 23938 4340 23996
rect 4284 23886 4286 23938
rect 4338 23886 4340 23938
rect 4284 23874 4340 23886
rect 4956 24050 5012 24062
rect 4956 23998 4958 24050
rect 5010 23998 5012 24050
rect 3052 23828 3108 23838
rect 1932 23604 1988 23614
rect 1932 23042 1988 23548
rect 1932 22990 1934 23042
rect 1986 22990 1988 23042
rect 1932 22978 1988 22990
rect 3052 22594 3108 23772
rect 4620 23828 4676 23838
rect 4620 23734 4676 23772
rect 4284 23716 4340 23726
rect 4172 23660 4284 23716
rect 3052 22542 3054 22594
rect 3106 22542 3108 22594
rect 2268 22372 2324 22382
rect 2268 22278 2324 22316
rect 2828 22372 2884 22382
rect 2828 22278 2884 22316
rect 2492 22260 2548 22270
rect 2492 22166 2548 22204
rect 2268 21700 2324 21710
rect 2268 21606 2324 21644
rect 3052 21700 3108 22542
rect 3388 23044 3444 23054
rect 3388 22594 3444 22988
rect 3388 22542 3390 22594
rect 3442 22542 3444 22594
rect 3388 22530 3444 22542
rect 4060 22372 4116 22382
rect 3948 22370 4116 22372
rect 3948 22318 4062 22370
rect 4114 22318 4116 22370
rect 3948 22316 4116 22318
rect 3052 21634 3108 21644
rect 3164 21812 3220 21822
rect 2716 21588 2772 21598
rect 2492 21532 2716 21588
rect 2492 19458 2548 21532
rect 2716 21494 2772 21532
rect 3164 21586 3220 21756
rect 3948 21810 4004 22316
rect 4060 22306 4116 22316
rect 3948 21758 3950 21810
rect 4002 21758 4004 21810
rect 3948 21746 4004 21758
rect 4172 22260 4228 23660
rect 4284 23650 4340 23660
rect 4844 23716 4900 23726
rect 4844 23622 4900 23660
rect 4284 23156 4340 23166
rect 4284 23062 4340 23100
rect 4732 23044 4788 23054
rect 4732 22950 4788 22988
rect 4844 22932 4900 22942
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4732 22596 4788 22606
rect 4508 22484 4564 22494
rect 4508 22390 4564 22428
rect 3612 21700 3668 21710
rect 3164 21534 3166 21586
rect 3218 21534 3220 21586
rect 2940 21476 2996 21486
rect 2492 19406 2494 19458
rect 2546 19406 2548 19458
rect 2492 19394 2548 19406
rect 2716 20018 2772 20030
rect 2716 19966 2718 20018
rect 2770 19966 2772 20018
rect 1708 19122 1764 19134
rect 1708 19070 1710 19122
rect 1762 19070 1764 19122
rect 1708 18900 1764 19070
rect 2044 19012 2100 19022
rect 2044 18918 2100 18956
rect 1764 18844 1876 18900
rect 1708 18834 1764 18844
rect 1820 18674 1876 18844
rect 2716 18788 2772 19966
rect 2828 19906 2884 19918
rect 2828 19854 2830 19906
rect 2882 19854 2884 19906
rect 2828 19234 2884 19854
rect 2828 19182 2830 19234
rect 2882 19182 2884 19234
rect 2828 19124 2884 19182
rect 2828 19058 2884 19068
rect 2940 18788 2996 21420
rect 3164 21140 3220 21534
rect 3052 21084 3220 21140
rect 3276 21588 3332 21598
rect 3052 20244 3108 21084
rect 3164 20916 3220 20926
rect 3276 20916 3332 21532
rect 3612 21586 3668 21644
rect 4060 21700 4116 21710
rect 4172 21700 4228 22204
rect 4732 21810 4788 22540
rect 4844 22482 4900 22876
rect 4844 22430 4846 22482
rect 4898 22430 4900 22482
rect 4844 22418 4900 22430
rect 4956 22370 5012 23998
rect 5068 23716 5124 23726
rect 5068 23714 5236 23716
rect 5068 23662 5070 23714
rect 5122 23662 5236 23714
rect 5068 23660 5236 23662
rect 5068 23650 5124 23660
rect 5180 23154 5236 23660
rect 5180 23102 5182 23154
rect 5234 23102 5236 23154
rect 4956 22318 4958 22370
rect 5010 22318 5012 22370
rect 4956 22306 5012 22318
rect 5068 22484 5124 22494
rect 5068 22036 5124 22428
rect 4732 21758 4734 21810
rect 4786 21758 4788 21810
rect 4732 21746 4788 21758
rect 4956 21980 5124 22036
rect 4060 21698 4228 21700
rect 4060 21646 4062 21698
rect 4114 21646 4228 21698
rect 4060 21644 4228 21646
rect 4060 21634 4116 21644
rect 3612 21534 3614 21586
rect 3666 21534 3668 21586
rect 3612 21522 3668 21534
rect 4284 21586 4340 21598
rect 4284 21534 4286 21586
rect 4338 21534 4340 21586
rect 4284 21364 4340 21534
rect 4620 21588 4676 21598
rect 4620 21494 4676 21532
rect 4844 21588 4900 21598
rect 4844 21494 4900 21532
rect 4284 21298 4340 21308
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 3388 21028 3444 21038
rect 3388 21026 4004 21028
rect 3388 20974 3390 21026
rect 3442 20974 4004 21026
rect 3388 20972 4004 20974
rect 3388 20962 3444 20972
rect 3164 20914 3332 20916
rect 3164 20862 3166 20914
rect 3218 20862 3332 20914
rect 3164 20860 3332 20862
rect 3164 20850 3220 20860
rect 3612 20802 3668 20814
rect 3612 20750 3614 20802
rect 3666 20750 3668 20802
rect 3052 20178 3108 20188
rect 3500 20244 3556 20254
rect 2716 18722 2772 18732
rect 2828 18732 2996 18788
rect 3052 19234 3108 19246
rect 3052 19182 3054 19234
rect 3106 19182 3108 19234
rect 3052 18788 3108 19182
rect 1820 18622 1822 18674
rect 1874 18622 1876 18674
rect 1820 18610 1876 18622
rect 2044 18564 2100 18574
rect 1708 18226 1764 18238
rect 1708 18174 1710 18226
rect 1762 18174 1764 18226
rect 1708 17556 1764 18174
rect 1708 17106 1764 17500
rect 1708 17054 1710 17106
rect 1762 17054 1764 17106
rect 1708 17042 1764 17054
rect 2044 17106 2100 18508
rect 2716 18452 2772 18462
rect 2380 18450 2772 18452
rect 2380 18398 2718 18450
rect 2770 18398 2772 18450
rect 2380 18396 2772 18398
rect 2268 18338 2324 18350
rect 2268 18286 2270 18338
rect 2322 18286 2324 18338
rect 2268 18226 2324 18286
rect 2268 18174 2270 18226
rect 2322 18174 2324 18226
rect 2268 18162 2324 18174
rect 2268 17668 2324 17678
rect 2380 17668 2436 18396
rect 2716 18386 2772 18396
rect 2268 17666 2436 17668
rect 2268 17614 2270 17666
rect 2322 17614 2436 17666
rect 2268 17612 2436 17614
rect 2604 17666 2660 17678
rect 2604 17614 2606 17666
rect 2658 17614 2660 17666
rect 2268 17602 2324 17612
rect 2044 17054 2046 17106
rect 2098 17054 2100 17106
rect 2044 17042 2100 17054
rect 2604 16772 2660 17614
rect 2604 16706 2660 16716
rect 1708 16212 1764 16222
rect 1708 16098 1764 16156
rect 2828 16210 2884 18732
rect 3052 18722 3108 18732
rect 3388 19124 3444 19134
rect 2940 18564 2996 18574
rect 2940 18470 2996 18508
rect 3052 18450 3108 18462
rect 3052 18398 3054 18450
rect 3106 18398 3108 18450
rect 3052 17108 3108 18398
rect 3388 17892 3444 19068
rect 3500 17892 3556 20188
rect 3612 19346 3668 20750
rect 3948 20020 4004 20972
rect 4956 21026 5012 21980
rect 5068 21812 5124 21822
rect 5068 21718 5124 21756
rect 5180 21364 5236 23102
rect 5292 23156 5348 24332
rect 10332 24610 10388 24622
rect 10332 24558 10334 24610
rect 10386 24558 10388 24610
rect 10332 24276 10388 24558
rect 9996 24220 10388 24276
rect 10556 24498 10612 24510
rect 10556 24446 10558 24498
rect 10610 24446 10612 24498
rect 6412 23940 6468 23950
rect 5852 23938 6468 23940
rect 5852 23886 6414 23938
rect 6466 23886 6468 23938
rect 5852 23884 6468 23886
rect 5292 23090 5348 23100
rect 5628 23826 5684 23838
rect 5628 23774 5630 23826
rect 5682 23774 5684 23826
rect 5628 22596 5684 23774
rect 5628 22530 5684 22540
rect 5740 23716 5796 23726
rect 5852 23716 5908 23884
rect 6412 23874 6468 23884
rect 6972 23940 7028 23950
rect 6636 23826 6692 23838
rect 6636 23774 6638 23826
rect 6690 23774 6692 23826
rect 5740 23714 5908 23716
rect 5740 23662 5742 23714
rect 5794 23662 5908 23714
rect 5740 23660 5908 23662
rect 5964 23714 6020 23726
rect 5964 23662 5966 23714
rect 6018 23662 6020 23714
rect 5180 21298 5236 21308
rect 4956 20974 4958 21026
rect 5010 20974 5012 21026
rect 4956 20962 5012 20974
rect 4060 20804 4116 20814
rect 4396 20804 4452 20814
rect 4060 20802 4452 20804
rect 4060 20750 4062 20802
rect 4114 20750 4398 20802
rect 4450 20750 4452 20802
rect 4060 20748 4452 20750
rect 4060 20738 4116 20748
rect 4396 20738 4452 20748
rect 4620 20804 4676 20814
rect 4620 20802 4900 20804
rect 4620 20750 4622 20802
rect 4674 20750 4900 20802
rect 4620 20748 4900 20750
rect 4620 20738 4676 20748
rect 4620 20580 4676 20590
rect 3948 20018 4228 20020
rect 3948 19966 3950 20018
rect 4002 19966 4228 20018
rect 3948 19964 4228 19966
rect 3948 19954 4004 19964
rect 3612 19294 3614 19346
rect 3666 19294 3668 19346
rect 3612 19282 3668 19294
rect 3724 19234 3780 19246
rect 3724 19182 3726 19234
rect 3778 19182 3780 19234
rect 3724 18788 3780 19182
rect 4172 19234 4228 19964
rect 4620 19796 4676 20524
rect 4844 20132 4900 20748
rect 5740 20580 5796 23660
rect 5964 22482 6020 23662
rect 6636 23716 6692 23774
rect 6748 23828 6804 23838
rect 6748 23826 6916 23828
rect 6748 23774 6750 23826
rect 6802 23774 6916 23826
rect 6748 23772 6916 23774
rect 6748 23762 6804 23772
rect 6636 23604 6692 23660
rect 6636 23548 6804 23604
rect 5964 22430 5966 22482
rect 6018 22430 6020 22482
rect 5964 22418 6020 22430
rect 6188 23154 6244 23166
rect 6188 23102 6190 23154
rect 6242 23102 6244 23154
rect 6188 22484 6244 23102
rect 6188 22418 6244 22428
rect 6524 22260 6580 22270
rect 6524 22166 6580 22204
rect 6636 22036 6692 22046
rect 5740 20514 5796 20524
rect 6188 21364 6244 21374
rect 5516 20244 5572 20254
rect 5404 20188 5516 20244
rect 5180 20132 5236 20142
rect 4844 20130 5236 20132
rect 4844 20078 5182 20130
rect 5234 20078 5236 20130
rect 4844 20076 5236 20078
rect 5180 20066 5236 20076
rect 5404 20130 5460 20188
rect 5516 20178 5572 20188
rect 5404 20078 5406 20130
rect 5458 20078 5460 20130
rect 5404 20066 5460 20078
rect 4732 20020 4788 20030
rect 4732 19926 4788 19964
rect 5516 20020 5572 20030
rect 5516 19926 5572 19964
rect 4620 19740 4900 19796
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4172 19182 4174 19234
rect 4226 19182 4228 19234
rect 4172 19170 4228 19182
rect 4508 19236 4564 19246
rect 4508 19142 4564 19180
rect 4396 19124 4452 19134
rect 4396 19030 4452 19068
rect 3724 18722 3780 18732
rect 4844 18674 4900 19740
rect 6188 19460 6244 21308
rect 6636 21028 6692 21980
rect 6748 21588 6804 23548
rect 6860 22484 6916 23772
rect 6972 23266 7028 23884
rect 7868 23938 7924 23950
rect 7868 23886 7870 23938
rect 7922 23886 7924 23938
rect 6972 23214 6974 23266
rect 7026 23214 7028 23266
rect 6972 23202 7028 23214
rect 7196 23714 7252 23726
rect 7196 23662 7198 23714
rect 7250 23662 7252 23714
rect 7196 22596 7252 23662
rect 7868 23266 7924 23886
rect 7868 23214 7870 23266
rect 7922 23214 7924 23266
rect 7868 22932 7924 23214
rect 8316 23938 8372 23950
rect 8316 23886 8318 23938
rect 8370 23886 8372 23938
rect 8316 23156 8372 23886
rect 9996 23938 10052 24220
rect 9996 23886 9998 23938
rect 10050 23886 10052 23938
rect 8540 23828 8596 23838
rect 8540 23734 8596 23772
rect 9996 23604 10052 23886
rect 10108 24052 10164 24062
rect 10556 24052 10612 24446
rect 10108 24050 10612 24052
rect 10108 23998 10110 24050
rect 10162 23998 10612 24050
rect 10108 23996 10612 23998
rect 10892 24498 10948 24510
rect 10892 24446 10894 24498
rect 10946 24446 10948 24498
rect 10892 24052 10948 24446
rect 10892 23996 11284 24052
rect 10108 23940 10164 23996
rect 10108 23874 10164 23884
rect 10668 23828 10724 23838
rect 11004 23828 11060 23838
rect 10668 23826 11060 23828
rect 10668 23774 10670 23826
rect 10722 23774 11006 23826
rect 11058 23774 11060 23826
rect 10668 23772 11060 23774
rect 10668 23762 10724 23772
rect 11004 23762 11060 23772
rect 11116 23716 11172 23726
rect 11116 23622 11172 23660
rect 9996 23548 10164 23604
rect 7868 22866 7924 22876
rect 8092 23154 8372 23156
rect 8092 23102 8318 23154
rect 8370 23102 8372 23154
rect 8092 23100 8372 23102
rect 7196 22530 7252 22540
rect 6860 22428 7140 22484
rect 7084 22372 7140 22428
rect 8092 22482 8148 23100
rect 8316 23090 8372 23100
rect 8988 23154 9044 23166
rect 8988 23102 8990 23154
rect 9042 23102 9044 23154
rect 8540 23042 8596 23054
rect 8540 22990 8542 23042
rect 8594 22990 8596 23042
rect 8092 22430 8094 22482
rect 8146 22430 8148 22482
rect 8092 22418 8148 22430
rect 8428 22596 8484 22606
rect 7420 22372 7476 22382
rect 7084 22370 8036 22372
rect 7084 22318 7422 22370
rect 7474 22318 8036 22370
rect 7084 22316 8036 22318
rect 7420 22306 7476 22316
rect 7196 21698 7252 21710
rect 7196 21646 7198 21698
rect 7250 21646 7252 21698
rect 7084 21588 7140 21598
rect 6748 21586 7140 21588
rect 6748 21534 7086 21586
rect 7138 21534 7140 21586
rect 6748 21532 7140 21534
rect 7084 21522 7140 21532
rect 6636 20972 6804 21028
rect 6748 20914 6804 20972
rect 6748 20862 6750 20914
rect 6802 20862 6804 20914
rect 6748 20850 6804 20862
rect 6300 20804 6356 20814
rect 6300 20802 6468 20804
rect 6300 20750 6302 20802
rect 6354 20750 6468 20802
rect 6300 20748 6468 20750
rect 6300 20738 6356 20748
rect 6412 20244 6468 20748
rect 6412 19906 6468 20188
rect 6636 20802 6692 20814
rect 6636 20750 6638 20802
rect 6690 20750 6692 20802
rect 6412 19854 6414 19906
rect 6466 19854 6468 19906
rect 6412 19842 6468 19854
rect 6524 20130 6580 20142
rect 6524 20078 6526 20130
rect 6578 20078 6580 20130
rect 6524 19908 6580 20078
rect 6636 20020 6692 20750
rect 7084 20580 7140 20590
rect 7196 20580 7252 21646
rect 7980 21586 8036 22316
rect 8428 22370 8484 22540
rect 8428 22318 8430 22370
rect 8482 22318 8484 22370
rect 8428 22306 8484 22318
rect 8316 22260 8372 22270
rect 7980 21534 7982 21586
rect 8034 21534 8036 21586
rect 7980 20802 8036 21534
rect 8092 21810 8148 21822
rect 8092 21758 8094 21810
rect 8146 21758 8148 21810
rect 8092 21476 8148 21758
rect 8092 21410 8148 21420
rect 7980 20750 7982 20802
rect 8034 20750 8036 20802
rect 7980 20738 8036 20750
rect 7140 20524 7252 20580
rect 7084 20514 7140 20524
rect 8204 20468 8260 20478
rect 8204 20130 8260 20412
rect 8204 20078 8206 20130
rect 8258 20078 8260 20130
rect 8204 20066 8260 20078
rect 6636 19954 6692 19964
rect 7756 20018 7812 20030
rect 7756 19966 7758 20018
rect 7810 19966 7812 20018
rect 6524 19842 6580 19852
rect 7420 19906 7476 19918
rect 7420 19854 7422 19906
rect 7474 19854 7476 19906
rect 6748 19796 6804 19806
rect 7420 19796 7476 19854
rect 6748 19794 7476 19796
rect 6748 19742 6750 19794
rect 6802 19742 7476 19794
rect 6748 19740 7476 19742
rect 7756 19908 7812 19966
rect 6748 19730 6804 19740
rect 6636 19460 6692 19470
rect 6188 19458 6692 19460
rect 6188 19406 6638 19458
rect 6690 19406 6692 19458
rect 6188 19404 6692 19406
rect 6636 19394 6692 19404
rect 5068 19236 5124 19246
rect 5068 19012 5124 19180
rect 6972 19234 7028 19246
rect 6972 19182 6974 19234
rect 7026 19182 7028 19234
rect 5628 19124 5684 19134
rect 5628 19030 5684 19068
rect 5964 19012 6020 19022
rect 5068 19010 5348 19012
rect 5068 18958 5070 19010
rect 5122 18958 5348 19010
rect 5068 18956 5348 18958
rect 5068 18946 5124 18956
rect 4844 18622 4846 18674
rect 4898 18622 4900 18674
rect 4844 18610 4900 18622
rect 4956 18900 5012 18910
rect 4172 18562 4228 18574
rect 4172 18510 4174 18562
rect 4226 18510 4228 18562
rect 4060 18452 4116 18462
rect 3836 18450 4116 18452
rect 3836 18398 4062 18450
rect 4114 18398 4116 18450
rect 3836 18396 4116 18398
rect 3724 17892 3780 17902
rect 3500 17890 3780 17892
rect 3500 17838 3726 17890
rect 3778 17838 3780 17890
rect 3500 17836 3780 17838
rect 3388 17826 3444 17836
rect 3724 17826 3780 17836
rect 3052 17042 3108 17052
rect 3388 17666 3444 17678
rect 3388 17614 3390 17666
rect 3442 17614 3444 17666
rect 2940 16882 2996 16894
rect 2940 16830 2942 16882
rect 2994 16830 2996 16882
rect 2940 16772 2996 16830
rect 2940 16706 2996 16716
rect 3388 16882 3444 17614
rect 3388 16830 3390 16882
rect 3442 16830 3444 16882
rect 3388 16772 3444 16830
rect 3388 16706 3444 16716
rect 3500 17668 3556 17678
rect 2828 16158 2830 16210
rect 2882 16158 2884 16210
rect 2828 16146 2884 16158
rect 1708 16046 1710 16098
rect 1762 16046 1764 16098
rect 1708 14644 1764 16046
rect 3388 16100 3444 16110
rect 2044 15988 2100 15998
rect 2044 15894 2100 15932
rect 2940 15986 2996 15998
rect 2940 15934 2942 15986
rect 2994 15934 2996 15986
rect 2156 15876 2212 15886
rect 2156 15314 2212 15820
rect 2716 15876 2772 15886
rect 2716 15782 2772 15820
rect 2156 15262 2158 15314
rect 2210 15262 2212 15314
rect 2156 15250 2212 15262
rect 2604 15316 2660 15326
rect 1820 14868 1876 14878
rect 1876 14812 1988 14868
rect 1820 14802 1876 14812
rect 1820 14644 1876 14654
rect 1708 14642 1876 14644
rect 1708 14590 1822 14642
rect 1874 14590 1876 14642
rect 1708 14588 1876 14590
rect 1820 14578 1876 14588
rect 1820 13748 1876 13758
rect 1932 13748 1988 14812
rect 2604 14530 2660 15260
rect 2940 14754 2996 15934
rect 3388 15540 3444 16044
rect 3388 15474 3444 15484
rect 2940 14702 2942 14754
rect 2994 14702 2996 14754
rect 2940 14690 2996 14702
rect 3388 15314 3444 15326
rect 3388 15262 3390 15314
rect 3442 15262 3444 15314
rect 3052 14644 3108 14654
rect 3388 14644 3444 15262
rect 3500 15090 3556 17612
rect 3836 17556 3892 18396
rect 4060 18386 4116 18396
rect 4172 17892 4228 18510
rect 4956 18562 5012 18844
rect 4956 18510 4958 18562
rect 5010 18510 5012 18562
rect 4172 17826 4228 17836
rect 4284 18452 4340 18462
rect 4284 17668 4340 18396
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 4396 17892 4452 17902
rect 4452 17836 4564 17892
rect 4396 17826 4452 17836
rect 4396 17668 4452 17678
rect 3612 17500 3892 17556
rect 4060 17666 4452 17668
rect 4060 17614 4398 17666
rect 4450 17614 4452 17666
rect 4060 17612 4452 17614
rect 3612 16994 3668 17500
rect 3612 16942 3614 16994
rect 3666 16942 3668 16994
rect 3612 16930 3668 16942
rect 3948 17108 4004 17118
rect 3612 15874 3668 15886
rect 3612 15822 3614 15874
rect 3666 15822 3668 15874
rect 3612 15764 3668 15822
rect 3836 15876 3892 15886
rect 3836 15782 3892 15820
rect 3612 15698 3668 15708
rect 3948 15148 4004 17052
rect 4060 15986 4116 17612
rect 4396 17602 4452 17612
rect 4508 16882 4564 17836
rect 4732 17556 4788 17566
rect 4956 17556 5012 18510
rect 5180 18788 5236 18798
rect 5292 18788 5348 18956
rect 5964 18918 6020 18956
rect 5292 18732 5796 18788
rect 5180 18116 5236 18732
rect 5180 18060 5348 18116
rect 4732 17554 5012 17556
rect 4732 17502 4734 17554
rect 4786 17502 5012 17554
rect 4732 17500 5012 17502
rect 4732 17490 4788 17500
rect 5180 17108 5236 17118
rect 4508 16830 4510 16882
rect 4562 16830 4564 16882
rect 4508 16818 4564 16830
rect 4844 17106 5236 17108
rect 4844 17054 5182 17106
rect 5234 17054 5236 17106
rect 4844 17052 5236 17054
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 4620 16100 4676 16110
rect 4620 16006 4676 16044
rect 4060 15934 4062 15986
rect 4114 15934 4116 15986
rect 4060 15922 4116 15934
rect 4172 15986 4228 15998
rect 4172 15934 4174 15986
rect 4226 15934 4228 15986
rect 3500 15038 3502 15090
rect 3554 15038 3556 15090
rect 3500 15026 3556 15038
rect 3836 15092 4004 15148
rect 3052 14642 3556 14644
rect 3052 14590 3054 14642
rect 3106 14590 3556 14642
rect 3052 14588 3556 14590
rect 3052 14578 3108 14588
rect 2604 14478 2606 14530
rect 2658 14478 2660 14530
rect 2604 14466 2660 14478
rect 3500 14530 3556 14588
rect 3500 14478 3502 14530
rect 3554 14478 3556 14530
rect 3500 14466 3556 14478
rect 3836 14530 3892 15092
rect 3836 14478 3838 14530
rect 3890 14478 3892 14530
rect 2044 14308 2100 14318
rect 2044 13970 2100 14252
rect 3724 14308 3780 14318
rect 3724 14214 3780 14252
rect 2044 13918 2046 13970
rect 2098 13918 2100 13970
rect 2044 13906 2100 13918
rect 2380 14196 2436 14206
rect 2380 13858 2436 14140
rect 3164 14196 3220 14206
rect 2716 14084 2772 14094
rect 2716 13970 2772 14028
rect 2716 13918 2718 13970
rect 2770 13918 2772 13970
rect 2716 13906 2772 13918
rect 3164 13970 3220 14140
rect 3724 13972 3780 13982
rect 3836 13972 3892 14478
rect 4172 14084 4228 15934
rect 4844 15538 4900 17052
rect 5180 17042 5236 17052
rect 4956 16884 5012 16894
rect 4956 16790 5012 16828
rect 5068 16884 5124 16894
rect 5292 16884 5348 18060
rect 5068 16882 5348 16884
rect 5068 16830 5070 16882
rect 5122 16830 5348 16882
rect 5068 16828 5348 16830
rect 5068 16818 5124 16828
rect 4844 15486 4846 15538
rect 4898 15486 4900 15538
rect 4844 15474 4900 15486
rect 4956 15540 5012 15550
rect 4956 15446 5012 15484
rect 4508 15316 4564 15326
rect 4284 15314 4564 15316
rect 4284 15262 4510 15314
rect 4562 15262 4564 15314
rect 4284 15260 4564 15262
rect 4284 15092 4340 15260
rect 4508 15250 4564 15260
rect 4732 15314 4788 15326
rect 4732 15262 4734 15314
rect 4786 15262 4788 15314
rect 4732 15148 4788 15262
rect 5180 15314 5236 15326
rect 5180 15262 5182 15314
rect 5234 15262 5236 15314
rect 4732 15092 4900 15148
rect 4284 14308 4340 15036
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 4844 14532 4900 15092
rect 4956 14532 5012 14542
rect 4844 14476 4956 14532
rect 4284 14242 4340 14252
rect 4620 14418 4676 14430
rect 4620 14366 4622 14418
rect 4674 14366 4676 14418
rect 4620 14084 4676 14366
rect 4956 14418 5012 14476
rect 4956 14366 4958 14418
rect 5010 14366 5012 14418
rect 4956 14354 5012 14366
rect 4172 14028 4676 14084
rect 3164 13918 3166 13970
rect 3218 13918 3220 13970
rect 3164 13906 3220 13918
rect 3388 13970 3892 13972
rect 3388 13918 3726 13970
rect 3778 13918 3892 13970
rect 3388 13916 3892 13918
rect 2380 13806 2382 13858
rect 2434 13806 2436 13858
rect 2380 13794 2436 13806
rect 1820 13746 1932 13748
rect 1820 13694 1822 13746
rect 1874 13694 1932 13746
rect 1820 13692 1932 13694
rect 1820 13682 1876 13692
rect 1932 13654 1988 13692
rect 1708 13524 1764 13534
rect 1708 12964 1764 13468
rect 2044 13524 2100 13534
rect 1708 12962 1876 12964
rect 1708 12910 1710 12962
rect 1762 12910 1876 12962
rect 1708 12908 1876 12910
rect 1708 12898 1764 12908
rect 1708 12740 1764 12750
rect 1708 12402 1764 12684
rect 1708 12350 1710 12402
rect 1762 12350 1764 12402
rect 1708 12180 1764 12350
rect 1708 12114 1764 12124
rect 1708 11282 1764 11294
rect 1708 11230 1710 11282
rect 1762 11230 1764 11282
rect 1708 10836 1764 11230
rect 1708 10388 1764 10780
rect 1820 10834 1876 12908
rect 2044 12850 2100 13468
rect 2044 12798 2046 12850
rect 2098 12798 2100 12850
rect 2044 12786 2100 12798
rect 2380 12852 2436 12862
rect 3388 12852 3444 13916
rect 3724 13906 3780 13916
rect 3724 13748 3780 13758
rect 3948 13748 4004 13758
rect 4396 13748 4452 13758
rect 3780 13692 3892 13748
rect 3724 13682 3780 13692
rect 3836 13300 3892 13692
rect 3948 13746 4452 13748
rect 3948 13694 3950 13746
rect 4002 13694 4398 13746
rect 4450 13694 4452 13746
rect 3948 13692 4452 13694
rect 3948 13524 4004 13692
rect 4396 13682 4452 13692
rect 4620 13524 4676 14028
rect 4732 13972 4788 13982
rect 4732 13878 4788 13916
rect 5180 13972 5236 15262
rect 5180 13906 5236 13916
rect 3948 13458 4004 13468
rect 4284 13468 4676 13524
rect 3836 13244 4116 13300
rect 3500 13188 3556 13198
rect 3500 13186 3780 13188
rect 3500 13134 3502 13186
rect 3554 13134 3780 13186
rect 3500 13132 3780 13134
rect 3500 13122 3556 13132
rect 3500 12852 3556 12862
rect 3388 12850 3556 12852
rect 3388 12798 3502 12850
rect 3554 12798 3556 12850
rect 3388 12796 3556 12798
rect 2380 12758 2436 12796
rect 3500 12786 3556 12796
rect 3612 12850 3668 12862
rect 3612 12798 3614 12850
rect 3666 12798 3668 12850
rect 2716 12738 2772 12750
rect 2716 12686 2718 12738
rect 2770 12686 2772 12738
rect 2716 12628 2772 12686
rect 3388 12628 3444 12638
rect 2716 12572 3388 12628
rect 2044 12292 2100 12302
rect 2044 12198 2100 12236
rect 2716 12290 2772 12302
rect 2716 12238 2718 12290
rect 2770 12238 2772 12290
rect 2380 12178 2436 12190
rect 2380 12126 2382 12178
rect 2434 12126 2436 12178
rect 2380 12068 2436 12126
rect 2380 11508 2436 12012
rect 2380 11442 2436 11452
rect 1820 10782 1822 10834
rect 1874 10782 1876 10834
rect 1820 10770 1876 10782
rect 2044 11170 2100 11182
rect 2044 11118 2046 11170
rect 2098 11118 2100 11170
rect 2044 10836 2100 11118
rect 2716 11172 2772 12238
rect 3388 11508 3444 12572
rect 3500 12178 3556 12190
rect 3500 12126 3502 12178
rect 3554 12126 3556 12178
rect 3500 11732 3556 12126
rect 3612 11956 3668 12798
rect 3724 12068 3780 13132
rect 4060 13074 4116 13244
rect 4060 13022 4062 13074
rect 4114 13022 4116 13074
rect 4060 13010 4116 13022
rect 4284 12628 4340 13468
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 4508 12852 4564 12862
rect 4508 12758 4564 12796
rect 4956 12740 5012 12750
rect 4956 12646 5012 12684
rect 4284 12562 4340 12572
rect 4620 12404 4676 12414
rect 4620 12310 4676 12348
rect 3836 12068 3892 12078
rect 3724 12066 3892 12068
rect 3724 12014 3838 12066
rect 3890 12014 3892 12066
rect 3724 12012 3892 12014
rect 3612 11890 3668 11900
rect 3500 11676 3780 11732
rect 3612 11508 3668 11518
rect 3388 11452 3556 11508
rect 2716 11106 2772 11116
rect 2828 11394 2884 11406
rect 2828 11342 2830 11394
rect 2882 11342 2884 11394
rect 2044 10770 2100 10780
rect 2828 10836 2884 11342
rect 3388 11284 3444 11294
rect 3164 11228 3388 11284
rect 2828 10770 2884 10780
rect 3052 11170 3108 11182
rect 3052 11118 3054 11170
rect 3106 11118 3108 11170
rect 2492 10724 2548 10734
rect 2492 10630 2548 10668
rect 2268 10610 2324 10622
rect 2268 10558 2270 10610
rect 2322 10558 2324 10610
rect 2268 10500 2324 10558
rect 2828 10610 2884 10622
rect 2828 10558 2830 10610
rect 2882 10558 2884 10610
rect 2828 10500 2884 10558
rect 2044 10444 2884 10500
rect 1820 10388 1876 10398
rect 1708 10332 1820 10388
rect 1820 10322 1876 10332
rect 1708 10164 1764 10174
rect 1708 9826 1764 10108
rect 1708 9774 1710 9826
rect 1762 9774 1764 9826
rect 1708 9762 1764 9774
rect 2044 9714 2100 10444
rect 2044 9662 2046 9714
rect 2098 9662 2100 9714
rect 2044 9650 2100 9662
rect 2492 10164 2548 10174
rect 1708 9492 1764 9502
rect 1708 9154 1764 9436
rect 1708 9102 1710 9154
rect 1762 9102 1764 9154
rect 1708 8428 1764 9102
rect 2044 9156 2100 9166
rect 2044 9062 2100 9100
rect 2380 9042 2436 9054
rect 2380 8990 2382 9042
rect 2434 8990 2436 9042
rect 2380 8820 2436 8990
rect 2380 8754 2436 8764
rect 1708 8372 1876 8428
rect 1708 8148 1764 8158
rect 1708 8054 1764 8092
rect 1820 7698 1876 8372
rect 2492 8370 2548 10108
rect 3052 10164 3108 11118
rect 3164 10834 3220 11228
rect 3388 11190 3444 11228
rect 3500 11170 3556 11452
rect 3500 11118 3502 11170
rect 3554 11118 3556 11170
rect 3500 11060 3556 11118
rect 3164 10782 3166 10834
rect 3218 10782 3220 10834
rect 3164 10770 3220 10782
rect 3388 11004 3556 11060
rect 3052 10098 3108 10108
rect 3164 10388 3220 10398
rect 2716 9716 2772 9726
rect 2716 9266 2772 9660
rect 2716 9214 2718 9266
rect 2770 9214 2772 9266
rect 2716 9202 2772 9214
rect 3164 9266 3220 10332
rect 3276 9826 3332 9838
rect 3276 9774 3278 9826
rect 3330 9774 3332 9826
rect 3276 9380 3332 9774
rect 3276 9314 3332 9324
rect 3164 9214 3166 9266
rect 3218 9214 3220 9266
rect 3164 9202 3220 9214
rect 3388 9268 3444 11004
rect 3500 10836 3556 10846
rect 3612 10836 3668 11452
rect 3724 11396 3780 11676
rect 3836 11508 3892 12012
rect 5180 12068 5236 12078
rect 5180 11974 5236 12012
rect 4844 11844 4900 11854
rect 5404 11844 5460 18732
rect 5628 18564 5684 18574
rect 5628 18470 5684 18508
rect 5740 18564 5796 18732
rect 6188 18564 6244 18574
rect 5740 18562 6244 18564
rect 5740 18510 5742 18562
rect 5794 18510 6190 18562
rect 6242 18510 6244 18562
rect 5740 18508 6244 18510
rect 5740 18498 5796 18508
rect 6188 18498 6244 18508
rect 6748 18562 6804 18574
rect 6748 18510 6750 18562
rect 6802 18510 6804 18562
rect 6524 18452 6580 18462
rect 6300 18450 6580 18452
rect 6300 18398 6526 18450
rect 6578 18398 6580 18450
rect 6300 18396 6580 18398
rect 5628 18226 5684 18238
rect 5628 18174 5630 18226
rect 5682 18174 5684 18226
rect 5628 17668 5684 18174
rect 6300 17892 6356 18396
rect 6524 18386 6580 18396
rect 6188 17836 6356 17892
rect 6636 18116 6692 18126
rect 5516 16882 5572 16894
rect 5516 16830 5518 16882
rect 5570 16830 5572 16882
rect 5516 15538 5572 16830
rect 5628 16884 5684 17612
rect 5852 17778 5908 17790
rect 5852 17726 5854 17778
rect 5906 17726 5908 17778
rect 5852 17106 5908 17726
rect 6188 17554 6244 17836
rect 6188 17502 6190 17554
rect 6242 17502 6244 17554
rect 6188 17490 6244 17502
rect 5852 17054 5854 17106
rect 5906 17054 5908 17106
rect 5852 17042 5908 17054
rect 5628 16818 5684 16828
rect 6076 16994 6132 17006
rect 6076 16942 6078 16994
rect 6130 16942 6132 16994
rect 6076 16324 6132 16942
rect 6188 16884 6244 16894
rect 6188 16882 6468 16884
rect 6188 16830 6190 16882
rect 6242 16830 6468 16882
rect 6188 16828 6468 16830
rect 6188 16818 6244 16828
rect 5740 16268 6076 16324
rect 5516 15486 5518 15538
rect 5570 15486 5572 15538
rect 5516 15474 5572 15486
rect 5628 15988 5684 15998
rect 5628 15540 5684 15932
rect 5516 15316 5572 15326
rect 5628 15316 5684 15484
rect 5740 15538 5796 16268
rect 6076 16258 6132 16268
rect 6188 16100 6244 16110
rect 5740 15486 5742 15538
rect 5794 15486 5796 15538
rect 5740 15474 5796 15486
rect 5964 16098 6244 16100
rect 5964 16046 6190 16098
rect 6242 16046 6244 16098
rect 5964 16044 6244 16046
rect 5964 15538 6020 16044
rect 6188 16034 6244 16044
rect 6300 15988 6356 15998
rect 6300 15894 6356 15932
rect 5964 15486 5966 15538
rect 6018 15486 6020 15538
rect 5516 15314 5684 15316
rect 5516 15262 5518 15314
rect 5570 15262 5684 15314
rect 5516 15260 5684 15262
rect 5516 15250 5572 15260
rect 5964 13972 6020 15486
rect 6188 15428 6244 15438
rect 6412 15428 6468 16828
rect 6524 16324 6580 16334
rect 6524 15538 6580 16268
rect 6524 15486 6526 15538
rect 6578 15486 6580 15538
rect 6524 15474 6580 15486
rect 6188 15426 6468 15428
rect 6188 15374 6190 15426
rect 6242 15374 6468 15426
rect 6188 15372 6468 15374
rect 6188 15362 6244 15372
rect 6300 14532 6356 15372
rect 6636 15148 6692 18060
rect 6748 17220 6804 18510
rect 6860 18450 6916 18462
rect 6860 18398 6862 18450
rect 6914 18398 6916 18450
rect 6860 17892 6916 18398
rect 6972 18116 7028 19182
rect 7196 19234 7252 19246
rect 7196 19182 7198 19234
rect 7250 19182 7252 19234
rect 7196 19124 7252 19182
rect 7196 19058 7252 19068
rect 7308 18674 7364 19740
rect 7308 18622 7310 18674
rect 7362 18622 7364 18674
rect 7308 18610 7364 18622
rect 7532 19012 7588 19022
rect 7532 18564 7588 18956
rect 7756 18788 7812 19852
rect 8316 19458 8372 22204
rect 8540 21700 8596 22990
rect 8988 22594 9044 23102
rect 8988 22542 8990 22594
rect 9042 22542 9044 22594
rect 8988 22530 9044 22542
rect 9884 22482 9940 22494
rect 9884 22430 9886 22482
rect 9938 22430 9940 22482
rect 8540 21634 8596 21644
rect 8652 22370 8708 22382
rect 8652 22318 8654 22370
rect 8706 22318 8708 22370
rect 8652 21476 8708 22318
rect 8876 22370 8932 22382
rect 8876 22318 8878 22370
rect 8930 22318 8932 22370
rect 8876 22260 8932 22318
rect 8876 22194 8932 22204
rect 9548 22258 9604 22270
rect 9548 22206 9550 22258
rect 9602 22206 9604 22258
rect 8652 21410 8708 21420
rect 9548 21028 9604 22206
rect 9772 22148 9828 22158
rect 8764 20972 9604 21028
rect 9660 22146 9828 22148
rect 9660 22094 9774 22146
rect 9826 22094 9828 22146
rect 9660 22092 9828 22094
rect 8764 20914 8820 20972
rect 9660 20916 9716 22092
rect 9772 22082 9828 22092
rect 8764 20862 8766 20914
rect 8818 20862 8820 20914
rect 8316 19406 8318 19458
rect 8370 19406 8372 19458
rect 8316 19394 8372 19406
rect 8652 19458 8708 19470
rect 8652 19406 8654 19458
rect 8706 19406 8708 19458
rect 8428 19124 8484 19134
rect 8652 19124 8708 19406
rect 8428 19122 8708 19124
rect 8428 19070 8430 19122
rect 8482 19070 8708 19122
rect 8428 19068 8708 19070
rect 7868 19012 7924 19022
rect 7868 18918 7924 18956
rect 8316 19010 8372 19022
rect 8316 18958 8318 19010
rect 8370 18958 8372 19010
rect 7756 18732 7924 18788
rect 7532 18470 7588 18508
rect 7644 18452 7700 18462
rect 7644 18450 7812 18452
rect 7644 18398 7646 18450
rect 7698 18398 7812 18450
rect 7644 18396 7812 18398
rect 7644 18386 7700 18396
rect 6972 18050 7028 18060
rect 6860 17826 6916 17836
rect 7308 17668 7364 17678
rect 7308 17574 7364 17612
rect 6972 17220 7028 17230
rect 6748 17164 6972 17220
rect 6972 17106 7028 17164
rect 6972 17054 6974 17106
rect 7026 17054 7028 17106
rect 6972 17042 7028 17054
rect 7308 16884 7364 16894
rect 7308 16882 7476 16884
rect 7308 16830 7310 16882
rect 7362 16830 7476 16882
rect 7308 16828 7476 16830
rect 7308 16818 7364 16828
rect 6748 16772 6804 16782
rect 6748 16210 6804 16716
rect 6748 16158 6750 16210
rect 6802 16158 6804 16210
rect 6748 16146 6804 16158
rect 7308 16100 7364 16110
rect 7196 16044 7308 16100
rect 6300 14438 6356 14476
rect 6412 15092 6692 15148
rect 6748 15314 6804 15326
rect 6748 15262 6750 15314
rect 6802 15262 6804 15314
rect 6748 15092 6804 15262
rect 6412 14420 6468 15092
rect 6804 15036 7140 15092
rect 6748 15026 6804 15036
rect 6636 14420 6692 14430
rect 6412 14418 6692 14420
rect 6412 14366 6638 14418
rect 6690 14366 6692 14418
rect 6412 14364 6692 14366
rect 7084 14420 7140 15036
rect 7196 14754 7252 16044
rect 7308 16006 7364 16044
rect 7420 15988 7476 16828
rect 7308 15540 7364 15550
rect 7420 15540 7476 15932
rect 7308 15538 7476 15540
rect 7308 15486 7310 15538
rect 7362 15486 7476 15538
rect 7308 15484 7476 15486
rect 7532 15764 7588 15774
rect 7308 15474 7364 15484
rect 7532 15314 7588 15708
rect 7532 15262 7534 15314
rect 7586 15262 7588 15314
rect 7532 15250 7588 15262
rect 7756 15148 7812 18396
rect 7868 17778 7924 18732
rect 8316 18564 8372 18958
rect 8316 18498 8372 18508
rect 8092 18338 8148 18350
rect 8092 18286 8094 18338
rect 8146 18286 8148 18338
rect 8092 18116 8148 18286
rect 8092 18050 8148 18060
rect 7868 17726 7870 17778
rect 7922 17726 7924 17778
rect 7868 17714 7924 17726
rect 7980 17892 8036 17902
rect 7980 17668 8036 17836
rect 8316 17668 8372 17678
rect 7980 17666 8372 17668
rect 7980 17614 8318 17666
rect 8370 17614 8372 17666
rect 7980 17612 8372 17614
rect 7980 16882 8036 17612
rect 8316 17602 8372 17612
rect 8428 17444 8484 19068
rect 8652 17444 8708 17454
rect 8428 17442 8708 17444
rect 8428 17390 8654 17442
rect 8706 17390 8708 17442
rect 8428 17388 8708 17390
rect 8316 16996 8372 17006
rect 8316 16902 8372 16940
rect 7980 16830 7982 16882
rect 8034 16830 8036 16882
rect 7980 16818 8036 16830
rect 7868 16770 7924 16782
rect 7868 16718 7870 16770
rect 7922 16718 7924 16770
rect 7868 16660 7924 16718
rect 7924 16604 8036 16660
rect 7868 16594 7924 16604
rect 7980 16322 8036 16604
rect 7980 16270 7982 16322
rect 8034 16270 8036 16322
rect 7980 16258 8036 16270
rect 7868 16098 7924 16110
rect 7868 16046 7870 16098
rect 7922 16046 7924 16098
rect 7868 15876 7924 16046
rect 7868 15810 7924 15820
rect 8092 15986 8148 15998
rect 8092 15934 8094 15986
rect 8146 15934 8148 15986
rect 8092 15764 8148 15934
rect 8092 15538 8148 15708
rect 8092 15486 8094 15538
rect 8146 15486 8148 15538
rect 8092 15474 8148 15486
rect 8652 15428 8708 17388
rect 8764 16884 8820 20862
rect 8876 20860 9716 20916
rect 8876 20802 8932 20860
rect 8876 20750 8878 20802
rect 8930 20750 8932 20802
rect 8876 20738 8932 20750
rect 9436 19908 9492 19918
rect 8988 19458 9044 19470
rect 8988 19406 8990 19458
rect 9042 19406 9044 19458
rect 8988 19346 9044 19406
rect 8988 19294 8990 19346
rect 9042 19294 9044 19346
rect 8988 19282 9044 19294
rect 9100 16884 9156 16894
rect 8764 16818 8820 16828
rect 8876 16828 9100 16884
rect 8876 15538 8932 16828
rect 9100 16790 9156 16828
rect 9212 16100 9268 16110
rect 9212 16006 9268 16044
rect 8876 15486 8878 15538
rect 8930 15486 8932 15538
rect 8876 15474 8932 15486
rect 8652 15362 8708 15372
rect 7868 15316 7924 15326
rect 7868 15222 7924 15260
rect 8204 15316 8260 15326
rect 8540 15316 8596 15326
rect 8204 15314 8596 15316
rect 8204 15262 8206 15314
rect 8258 15262 8542 15314
rect 8594 15262 8596 15314
rect 8204 15260 8596 15262
rect 7196 14702 7198 14754
rect 7250 14702 7252 14754
rect 7196 14690 7252 14702
rect 7644 15092 7812 15148
rect 7196 14420 7252 14430
rect 7084 14418 7252 14420
rect 7084 14366 7198 14418
rect 7250 14366 7252 14418
rect 7084 14364 7252 14366
rect 6636 14354 6692 14364
rect 7196 14354 7252 14364
rect 7308 14418 7364 14430
rect 7308 14366 7310 14418
rect 7362 14366 7364 14418
rect 7308 14084 7364 14366
rect 7644 14308 7700 15092
rect 7644 14242 7700 14252
rect 7308 14018 7364 14028
rect 8204 14084 8260 15260
rect 8540 15250 8596 15260
rect 9436 15148 9492 19852
rect 9660 19234 9716 20860
rect 9884 21586 9940 22430
rect 10108 22148 10164 23548
rect 10780 23154 10836 23166
rect 10780 23102 10782 23154
rect 10834 23102 10836 23154
rect 10220 22148 10276 22158
rect 10108 22092 10220 22148
rect 10220 22082 10276 22092
rect 10220 21812 10276 21822
rect 10220 21810 10724 21812
rect 10220 21758 10222 21810
rect 10274 21758 10724 21810
rect 10220 21756 10724 21758
rect 10220 21746 10276 21756
rect 9884 21534 9886 21586
rect 9938 21534 9940 21586
rect 9884 20802 9940 21534
rect 10332 21586 10388 21598
rect 10332 21534 10334 21586
rect 10386 21534 10388 21586
rect 9884 20750 9886 20802
rect 9938 20750 9940 20802
rect 9884 20738 9940 20750
rect 10108 21476 10164 21486
rect 10108 21362 10164 21420
rect 10108 21310 10110 21362
rect 10162 21310 10164 21362
rect 10108 20802 10164 21310
rect 10108 20750 10110 20802
rect 10162 20750 10164 20802
rect 10108 20738 10164 20750
rect 10220 20690 10276 20702
rect 10220 20638 10222 20690
rect 10274 20638 10276 20690
rect 10220 20580 10276 20638
rect 10220 20514 10276 20524
rect 9660 19182 9662 19234
rect 9714 19182 9716 19234
rect 9660 19170 9716 19182
rect 9996 19122 10052 19134
rect 9996 19070 9998 19122
rect 10050 19070 10052 19122
rect 9884 19010 9940 19022
rect 9884 18958 9886 19010
rect 9938 18958 9940 19010
rect 9884 18788 9940 18958
rect 9996 18900 10052 19070
rect 9996 18834 10052 18844
rect 9884 18722 9940 18732
rect 10332 18676 10388 21534
rect 10668 20802 10724 21756
rect 10780 21588 10836 23102
rect 11228 23156 11284 23996
rect 11228 23090 11284 23100
rect 11788 23716 11844 24668
rect 11900 24658 11956 24668
rect 14588 24722 14644 24734
rect 14588 24670 14590 24722
rect 14642 24670 14644 24722
rect 12124 24612 12180 24622
rect 11788 23154 11844 23660
rect 11788 23102 11790 23154
rect 11842 23102 11844 23154
rect 11788 23090 11844 23102
rect 12012 24610 12180 24612
rect 12012 24558 12126 24610
rect 12178 24558 12180 24610
rect 12012 24556 12180 24558
rect 12012 23266 12068 24556
rect 12124 24546 12180 24556
rect 12572 24612 12628 24622
rect 12572 24518 12628 24556
rect 14364 24610 14420 24622
rect 14364 24558 14366 24610
rect 14418 24558 14420 24610
rect 14028 23940 14084 23950
rect 14028 23846 14084 23884
rect 14252 23828 14308 23838
rect 14252 23734 14308 23772
rect 14364 23828 14420 24558
rect 14588 23828 14644 24670
rect 15260 24724 15316 24734
rect 15708 24724 15764 24734
rect 15260 24722 15764 24724
rect 15260 24670 15262 24722
rect 15314 24670 15710 24722
rect 15762 24670 15764 24722
rect 15260 24668 15764 24670
rect 15260 24658 15316 24668
rect 15708 24658 15764 24668
rect 15596 24498 15652 24510
rect 15596 24446 15598 24498
rect 15650 24446 15652 24498
rect 15260 24052 15316 24062
rect 15596 24052 15652 24446
rect 15260 24050 15652 24052
rect 15260 23998 15262 24050
rect 15314 23998 15652 24050
rect 15260 23996 15652 23998
rect 16716 24050 16772 24062
rect 16716 23998 16718 24050
rect 16770 23998 16772 24050
rect 14364 23826 14532 23828
rect 14364 23774 14366 23826
rect 14418 23774 14532 23826
rect 14364 23772 14532 23774
rect 14364 23762 14420 23772
rect 13804 23380 13860 23390
rect 13804 23286 13860 23324
rect 12012 23214 12014 23266
rect 12066 23214 12068 23266
rect 11004 23042 11060 23054
rect 11004 22990 11006 23042
rect 11058 22990 11060 23042
rect 11004 22258 11060 22990
rect 11116 22932 11172 22942
rect 11116 22838 11172 22876
rect 12012 22594 12068 23214
rect 13468 23156 13524 23166
rect 14252 23156 14308 23166
rect 13468 23062 13524 23100
rect 14140 23154 14308 23156
rect 14140 23102 14254 23154
rect 14306 23102 14308 23154
rect 14140 23100 14308 23102
rect 12012 22542 12014 22594
rect 12066 22542 12068 22594
rect 12012 22530 12068 22542
rect 12124 22932 12180 22942
rect 12124 22484 12180 22876
rect 12124 22390 12180 22428
rect 13580 22484 13636 22494
rect 13580 22390 13636 22428
rect 11340 22372 11396 22382
rect 11564 22372 11620 22382
rect 11340 22370 11620 22372
rect 11340 22318 11342 22370
rect 11394 22318 11566 22370
rect 11618 22318 11620 22370
rect 11340 22316 11620 22318
rect 11340 22306 11396 22316
rect 11564 22306 11620 22316
rect 12572 22372 12628 22382
rect 12572 22278 12628 22316
rect 14028 22372 14084 22382
rect 14028 22278 14084 22316
rect 11004 22206 11006 22258
rect 11058 22206 11060 22258
rect 11004 22036 11060 22206
rect 11004 21970 11060 21980
rect 11116 22146 11172 22158
rect 11116 22094 11118 22146
rect 11170 22094 11172 22146
rect 11116 21588 11172 22094
rect 12124 22148 12180 22158
rect 10780 21532 11172 21588
rect 11228 21698 11284 21710
rect 11228 21646 11230 21698
rect 11282 21646 11284 21698
rect 10668 20750 10670 20802
rect 10722 20750 10724 20802
rect 10668 20738 10724 20750
rect 10332 18610 10388 18620
rect 10668 19234 10724 19246
rect 10668 19182 10670 19234
rect 10722 19182 10724 19234
rect 9996 18564 10052 18574
rect 9996 18470 10052 18508
rect 10108 18564 10164 18574
rect 10108 18562 10276 18564
rect 10108 18510 10110 18562
rect 10162 18510 10276 18562
rect 10108 18508 10276 18510
rect 10108 18498 10164 18508
rect 10220 18340 10276 18508
rect 10556 18452 10612 18462
rect 10668 18452 10724 19182
rect 10892 19236 10948 21532
rect 11004 21362 11060 21374
rect 11004 21310 11006 21362
rect 11058 21310 11060 21362
rect 11004 20580 11060 21310
rect 11004 20514 11060 20524
rect 11116 20802 11172 20814
rect 11116 20750 11118 20802
rect 11170 20750 11172 20802
rect 11116 20130 11172 20750
rect 11116 20078 11118 20130
rect 11170 20078 11172 20130
rect 11116 19460 11172 20078
rect 11228 20020 11284 21646
rect 11340 21364 11396 21374
rect 11340 21362 11620 21364
rect 11340 21310 11342 21362
rect 11394 21310 11620 21362
rect 11340 21308 11620 21310
rect 11340 21298 11396 21308
rect 11564 20802 11620 21308
rect 11564 20750 11566 20802
rect 11618 20750 11620 20802
rect 11564 20738 11620 20750
rect 11564 20580 11620 20590
rect 11340 20020 11396 20030
rect 11228 20018 11396 20020
rect 11228 19966 11342 20018
rect 11394 19966 11396 20018
rect 11228 19964 11396 19966
rect 11116 19394 11172 19404
rect 11340 19236 11396 19964
rect 10892 19180 11284 19236
rect 11116 18676 11172 18686
rect 10556 18450 10948 18452
rect 10556 18398 10558 18450
rect 10610 18398 10948 18450
rect 10556 18396 10948 18398
rect 10556 18386 10612 18396
rect 10276 18284 10500 18340
rect 10220 18274 10276 18284
rect 10108 18226 10164 18238
rect 10108 18174 10110 18226
rect 10162 18174 10164 18226
rect 9772 17724 10052 17780
rect 9772 16996 9828 17724
rect 9772 16902 9828 16940
rect 9884 17556 9940 17566
rect 9884 16996 9940 17500
rect 9996 17554 10052 17724
rect 10108 17668 10164 18174
rect 10108 17602 10164 17612
rect 10332 17666 10388 17678
rect 10332 17614 10334 17666
rect 10386 17614 10388 17666
rect 9996 17502 9998 17554
rect 10050 17502 10052 17554
rect 9996 17444 10052 17502
rect 10332 17556 10388 17614
rect 10332 17490 10388 17500
rect 9996 17378 10052 17388
rect 10220 17442 10276 17454
rect 10220 17390 10222 17442
rect 10274 17390 10276 17442
rect 10220 17332 10276 17390
rect 10220 17266 10276 17276
rect 10444 17220 10500 18284
rect 10780 18226 10836 18238
rect 10780 18174 10782 18226
rect 10834 18174 10836 18226
rect 10780 17778 10836 18174
rect 10780 17726 10782 17778
rect 10834 17726 10836 17778
rect 10780 17714 10836 17726
rect 10892 17668 10948 18396
rect 11116 18450 11172 18620
rect 11116 18398 11118 18450
rect 11170 18398 11172 18450
rect 11116 18386 11172 18398
rect 11116 17668 11172 17678
rect 10892 17666 11172 17668
rect 10892 17614 11118 17666
rect 11170 17614 11172 17666
rect 10892 17612 11172 17614
rect 11116 17602 11172 17612
rect 10668 17444 10724 17454
rect 10668 17350 10724 17388
rect 10892 17444 10948 17454
rect 11228 17444 11284 19180
rect 11340 19142 11396 19180
rect 11564 19908 11620 20524
rect 12012 20018 12068 20030
rect 12012 19966 12014 20018
rect 12066 19966 12068 20018
rect 12012 19908 12068 19966
rect 11564 19852 12068 19908
rect 11564 19234 11620 19852
rect 12124 19796 12180 22092
rect 12348 21700 12404 21710
rect 12348 21588 12404 21644
rect 13580 21700 13636 21710
rect 13580 21606 13636 21644
rect 12236 21586 12404 21588
rect 12236 21534 12350 21586
rect 12402 21534 12404 21586
rect 12236 21532 12404 21534
rect 12236 20914 12292 21532
rect 12348 21522 12404 21532
rect 12460 21474 12516 21486
rect 12460 21422 12462 21474
rect 12514 21422 12516 21474
rect 12348 21028 12404 21038
rect 12348 20934 12404 20972
rect 12236 20862 12238 20914
rect 12290 20862 12292 20914
rect 12236 20850 12292 20862
rect 12460 20802 12516 21422
rect 14140 21252 14196 23100
rect 14252 23090 14308 23100
rect 14476 23044 14532 23772
rect 14588 23762 14644 23772
rect 15148 23938 15204 23950
rect 15148 23886 15150 23938
rect 15202 23886 15204 23938
rect 15148 23380 15204 23886
rect 15148 23314 15204 23324
rect 15260 23154 15316 23996
rect 15260 23102 15262 23154
rect 15314 23102 15316 23154
rect 15260 23090 15316 23102
rect 15484 23380 15540 23390
rect 15484 23154 15540 23324
rect 16156 23268 16212 23278
rect 16156 23174 16212 23212
rect 15484 23102 15486 23154
rect 15538 23102 15540 23154
rect 15484 23090 15540 23102
rect 16716 23156 16772 23998
rect 16828 23940 16884 23950
rect 16828 23846 16884 23884
rect 17836 23938 17892 25564
rect 18284 25508 18340 25518
rect 18396 25508 18452 26236
rect 18620 26226 18676 26236
rect 18732 26964 18788 26974
rect 18732 26178 18788 26908
rect 18732 26126 18734 26178
rect 18786 26126 18788 26178
rect 18732 26114 18788 26126
rect 19180 25956 19236 27020
rect 18284 25506 18396 25508
rect 18284 25454 18286 25506
rect 18338 25454 18396 25506
rect 18284 25452 18396 25454
rect 18284 25442 18340 25452
rect 18396 25414 18452 25452
rect 18620 25900 19236 25956
rect 19292 27074 19348 27086
rect 19292 27022 19294 27074
rect 19346 27022 19348 27074
rect 18620 25506 18676 25900
rect 19292 25732 19348 27022
rect 19852 27076 19908 27086
rect 20188 27076 20244 27086
rect 19908 27074 20244 27076
rect 19908 27022 20190 27074
rect 20242 27022 20244 27074
rect 19908 27020 20244 27022
rect 19852 26982 19908 27020
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 20188 26404 20244 27020
rect 20748 27076 20804 27086
rect 20748 26982 20804 27020
rect 21420 26964 21476 27580
rect 21644 27524 21700 27918
rect 21532 27468 21700 27524
rect 21868 27860 21924 27870
rect 21532 27186 21588 27468
rect 21532 27134 21534 27186
rect 21586 27134 21588 27186
rect 21532 27122 21588 27134
rect 21868 27074 21924 27804
rect 21868 27022 21870 27074
rect 21922 27022 21924 27074
rect 21868 27010 21924 27022
rect 21644 26964 21700 26974
rect 21420 26962 21700 26964
rect 21420 26910 21646 26962
rect 21698 26910 21700 26962
rect 21420 26908 21700 26910
rect 21644 26898 21700 26908
rect 19964 26348 20244 26404
rect 19740 26292 19796 26302
rect 19740 26290 19908 26292
rect 19740 26238 19742 26290
rect 19794 26238 19908 26290
rect 19740 26236 19908 26238
rect 19740 26226 19796 26236
rect 18956 25676 19348 25732
rect 18620 25454 18622 25506
rect 18674 25454 18676 25506
rect 18620 25442 18676 25454
rect 18732 25506 18788 25518
rect 18732 25454 18734 25506
rect 18786 25454 18788 25506
rect 18732 24948 18788 25454
rect 18956 25508 19012 25676
rect 19628 25618 19684 25630
rect 19628 25566 19630 25618
rect 19682 25566 19684 25618
rect 18956 25452 19236 25508
rect 19068 25172 19124 25182
rect 18732 24882 18788 24892
rect 18956 25116 19068 25172
rect 18844 24836 18900 24846
rect 18844 24742 18900 24780
rect 18956 24834 19012 25116
rect 19068 25106 19124 25116
rect 18956 24782 18958 24834
rect 19010 24782 19012 24834
rect 18956 24770 19012 24782
rect 18620 24722 18676 24734
rect 18620 24670 18622 24722
rect 18674 24670 18676 24722
rect 18508 24052 18564 24062
rect 18620 24052 18676 24670
rect 19180 24500 19236 25452
rect 19292 25396 19348 25406
rect 19628 25396 19684 25566
rect 19740 25508 19796 25518
rect 19740 25414 19796 25452
rect 19292 24722 19348 25340
rect 19516 25340 19684 25396
rect 19516 25172 19572 25340
rect 19852 25284 19908 26236
rect 19964 26290 20020 26348
rect 19964 26238 19966 26290
rect 20018 26238 20020 26290
rect 19964 26226 20020 26238
rect 20076 25508 20132 25518
rect 20076 25394 20132 25452
rect 20076 25342 20078 25394
rect 20130 25342 20132 25394
rect 20076 25330 20132 25342
rect 20188 25394 20244 26348
rect 20300 26178 20356 26190
rect 20300 26126 20302 26178
rect 20354 26126 20356 26178
rect 20300 25844 20356 26126
rect 20300 25778 20356 25788
rect 21868 25620 21924 25630
rect 21868 25526 21924 25564
rect 22204 25508 22260 28924
rect 22764 28756 22820 28766
rect 22540 28532 22596 28542
rect 22316 28420 22372 28430
rect 22316 28326 22372 28364
rect 22428 28418 22484 28430
rect 22428 28366 22430 28418
rect 22482 28366 22484 28418
rect 22316 27748 22372 27758
rect 22316 27654 22372 27692
rect 22428 27524 22484 28366
rect 22540 27860 22596 28476
rect 22540 27766 22596 27804
rect 22428 27458 22484 27468
rect 22764 26740 22820 28700
rect 22876 28644 22932 28654
rect 22876 28550 22932 28588
rect 23660 28532 23716 32620
rect 24220 32562 24276 32574
rect 24220 32510 24222 32562
rect 24274 32510 24276 32562
rect 23772 32452 23828 32462
rect 23828 32396 24164 32452
rect 23772 32358 23828 32396
rect 24108 31778 24164 32396
rect 24108 31726 24110 31778
rect 24162 31726 24164 31778
rect 24108 31714 24164 31726
rect 24220 31556 24276 32510
rect 24668 32450 24724 32462
rect 24668 32398 24670 32450
rect 24722 32398 24724 32450
rect 24444 31668 24500 31678
rect 24444 31574 24500 31612
rect 24220 31462 24276 31500
rect 24668 31556 24724 32398
rect 24668 31490 24724 31500
rect 24556 31106 24612 31118
rect 24556 31054 24558 31106
rect 24610 31054 24612 31106
rect 24332 30884 24388 30894
rect 24332 30790 24388 30828
rect 24332 30324 24388 30334
rect 24556 30324 24612 31054
rect 24668 30884 24724 30894
rect 24668 30790 24724 30828
rect 24668 30436 24724 30446
rect 24780 30436 24836 32620
rect 25116 32002 25172 33070
rect 25340 33124 25396 33182
rect 25564 33124 25620 34300
rect 26124 34242 26180 34860
rect 26124 34190 26126 34242
rect 26178 34190 26180 34242
rect 26124 34178 26180 34190
rect 26348 34914 26404 34926
rect 26348 34862 26350 34914
rect 26402 34862 26404 34914
rect 26348 34468 26404 34862
rect 26684 34916 26740 34926
rect 26684 34822 26740 34860
rect 25900 34132 25956 34142
rect 25900 34038 25956 34076
rect 26348 34130 26404 34412
rect 26348 34078 26350 34130
rect 26402 34078 26404 34130
rect 26348 34066 26404 34078
rect 26572 34690 26628 34702
rect 26572 34638 26574 34690
rect 26626 34638 26628 34690
rect 25340 33068 25620 33124
rect 25116 31950 25118 32002
rect 25170 31950 25172 32002
rect 25116 31938 25172 31950
rect 26124 32674 26180 32686
rect 26124 32622 26126 32674
rect 26178 32622 26180 32674
rect 26124 31892 26180 32622
rect 25676 31890 26180 31892
rect 25676 31838 26126 31890
rect 26178 31838 26180 31890
rect 25676 31836 26180 31838
rect 24668 30434 24836 30436
rect 24668 30382 24670 30434
rect 24722 30382 24836 30434
rect 24668 30380 24836 30382
rect 24892 31778 24948 31790
rect 24892 31726 24894 31778
rect 24946 31726 24948 31778
rect 24668 30370 24724 30380
rect 24388 30268 24612 30324
rect 24108 30212 24164 30222
rect 24108 30118 24164 30156
rect 24332 30210 24388 30268
rect 24332 30158 24334 30210
rect 24386 30158 24388 30210
rect 24332 30146 24388 30158
rect 24892 30210 24948 31726
rect 25340 31778 25396 31790
rect 25340 31726 25342 31778
rect 25394 31726 25396 31778
rect 25340 31668 25396 31726
rect 25676 31778 25732 31836
rect 26124 31826 26180 31836
rect 26236 32562 26292 32574
rect 26236 32510 26238 32562
rect 26290 32510 26292 32562
rect 25676 31726 25678 31778
rect 25730 31726 25732 31778
rect 25676 31714 25732 31726
rect 25340 31602 25396 31612
rect 26012 31666 26068 31678
rect 26012 31614 26014 31666
rect 26066 31614 26068 31666
rect 25452 31554 25508 31566
rect 25452 31502 25454 31554
rect 25506 31502 25508 31554
rect 24892 30158 24894 30210
rect 24946 30158 24948 30210
rect 24892 30100 24948 30158
rect 25228 30772 25284 30782
rect 25228 30210 25284 30716
rect 25228 30158 25230 30210
rect 25282 30158 25284 30210
rect 25228 30146 25284 30158
rect 25340 30212 25396 30222
rect 24892 30034 24948 30044
rect 25340 30098 25396 30156
rect 25340 30046 25342 30098
rect 25394 30046 25396 30098
rect 25340 30034 25396 30046
rect 24220 29986 24276 29998
rect 24220 29934 24222 29986
rect 24274 29934 24276 29986
rect 24220 28868 24276 29934
rect 23660 28466 23716 28476
rect 23884 28812 24276 28868
rect 22988 27636 23044 27646
rect 22988 27542 23044 27580
rect 22988 27132 23268 27188
rect 22764 26674 22820 26684
rect 22876 26964 22932 26974
rect 22988 26964 23044 27132
rect 22876 26962 23044 26964
rect 22876 26910 22878 26962
rect 22930 26910 23044 26962
rect 22876 26908 23044 26910
rect 23100 26964 23156 27002
rect 22428 26180 22484 26190
rect 22428 26086 22484 26124
rect 22876 25844 22932 26908
rect 23100 26898 23156 26908
rect 23212 26962 23268 27132
rect 23212 26910 23214 26962
rect 23266 26910 23268 26962
rect 23212 26898 23268 26910
rect 23324 27076 23380 27086
rect 22876 25778 22932 25788
rect 23100 26292 23156 26302
rect 23324 26292 23380 27020
rect 23772 26964 23828 27002
rect 23772 26898 23828 26908
rect 23884 26908 23940 28812
rect 23996 28644 24052 28654
rect 23996 28642 24276 28644
rect 23996 28590 23998 28642
rect 24050 28590 24276 28642
rect 23996 28588 24276 28590
rect 23996 28578 24052 28588
rect 24220 27076 24276 28588
rect 24668 28530 24724 28542
rect 24668 28478 24670 28530
rect 24722 28478 24724 28530
rect 24668 28084 24724 28478
rect 24668 28018 24724 28028
rect 25340 28084 25396 28094
rect 25340 27990 25396 28028
rect 25452 28082 25508 31502
rect 25900 31556 25956 31566
rect 26012 31556 26068 31614
rect 25956 31500 26068 31556
rect 25900 30994 25956 31500
rect 26236 31218 26292 32510
rect 26572 32564 26628 34638
rect 26684 33906 26740 33918
rect 26684 33854 26686 33906
rect 26738 33854 26740 33906
rect 26684 33236 26740 33854
rect 26684 33170 26740 33180
rect 26684 32564 26740 32574
rect 26572 32562 26740 32564
rect 26572 32510 26686 32562
rect 26738 32510 26740 32562
rect 26572 32508 26740 32510
rect 26684 32498 26740 32508
rect 26348 32452 26404 32462
rect 26348 32450 26516 32452
rect 26348 32398 26350 32450
rect 26402 32398 26516 32450
rect 26348 32396 26516 32398
rect 26348 32386 26404 32396
rect 26236 31166 26238 31218
rect 26290 31166 26292 31218
rect 26236 31154 26292 31166
rect 26348 31666 26404 31678
rect 26348 31614 26350 31666
rect 26402 31614 26404 31666
rect 25900 30942 25902 30994
rect 25954 30942 25956 30994
rect 25900 30930 25956 30942
rect 25676 30884 25732 30894
rect 25676 30790 25732 30828
rect 26236 30884 26292 30894
rect 26348 30884 26404 31614
rect 26292 30828 26404 30884
rect 26236 30818 26292 30828
rect 26460 30660 26516 32396
rect 26572 31780 26628 31790
rect 26572 31686 26628 31724
rect 26572 30884 26628 30894
rect 26572 30790 26628 30828
rect 26684 30882 26740 30894
rect 26684 30830 26686 30882
rect 26738 30830 26740 30882
rect 26236 30604 26516 30660
rect 26124 30210 26180 30222
rect 26124 30158 26126 30210
rect 26178 30158 26180 30210
rect 25564 29988 25620 29998
rect 25564 29986 25956 29988
rect 25564 29934 25566 29986
rect 25618 29934 25956 29986
rect 25564 29932 25956 29934
rect 25564 29922 25620 29932
rect 25900 29876 25956 29932
rect 26124 29876 26180 30158
rect 25900 29820 26180 29876
rect 25452 28030 25454 28082
rect 25506 28030 25508 28082
rect 25452 28018 25508 28030
rect 25676 28644 25732 28654
rect 25676 28082 25732 28588
rect 25676 28030 25678 28082
rect 25730 28030 25732 28082
rect 25676 28018 25732 28030
rect 25228 27860 25284 27870
rect 24220 26982 24276 27020
rect 24556 27858 25284 27860
rect 24556 27806 25230 27858
rect 25282 27806 25284 27858
rect 24556 27804 25284 27806
rect 24332 26964 24388 26974
rect 23436 26850 23492 26862
rect 23884 26852 24052 26908
rect 23436 26798 23438 26850
rect 23490 26798 23492 26850
rect 23436 26628 23492 26798
rect 23436 26562 23492 26572
rect 23772 26516 23828 26526
rect 23996 26516 24052 26852
rect 23772 26514 24052 26516
rect 23772 26462 23774 26514
rect 23826 26462 24052 26514
rect 23772 26460 24052 26462
rect 24108 26628 24164 26638
rect 23772 26450 23828 26460
rect 23548 26292 23604 26302
rect 23100 26290 23380 26292
rect 23100 26238 23102 26290
rect 23154 26238 23380 26290
rect 23100 26236 23380 26238
rect 23436 26290 23604 26292
rect 23436 26238 23550 26290
rect 23602 26238 23604 26290
rect 23436 26236 23604 26238
rect 23100 25620 23156 26236
rect 23100 25554 23156 25564
rect 23212 25956 23268 25966
rect 22204 25442 22260 25452
rect 20188 25342 20190 25394
rect 20242 25342 20244 25394
rect 20188 25330 20244 25342
rect 22652 25396 22708 25406
rect 19516 25106 19572 25116
rect 19628 25228 19908 25284
rect 20412 25282 20468 25294
rect 20412 25230 20414 25282
rect 20466 25230 20468 25282
rect 19292 24670 19294 24722
rect 19346 24670 19348 24722
rect 19292 24658 19348 24670
rect 19516 24948 19572 24958
rect 19180 24444 19348 24500
rect 18508 24050 18676 24052
rect 18508 23998 18510 24050
rect 18562 23998 18676 24050
rect 18508 23996 18676 23998
rect 18508 23986 18564 23996
rect 17836 23886 17838 23938
rect 17890 23886 17892 23938
rect 17836 23874 17892 23886
rect 19068 23940 19124 23950
rect 18060 23266 18116 23278
rect 18060 23214 18062 23266
rect 18114 23214 18116 23266
rect 17948 23156 18004 23166
rect 16716 23090 16772 23100
rect 17836 23154 18004 23156
rect 17836 23102 17950 23154
rect 18002 23102 18004 23154
rect 17836 23100 18004 23102
rect 14364 22988 14532 23044
rect 16492 23044 16548 23054
rect 14252 22930 14308 22942
rect 14252 22878 14254 22930
rect 14306 22878 14308 22930
rect 14252 22372 14308 22878
rect 14252 22306 14308 22316
rect 14364 21252 14420 22988
rect 14588 22930 14644 22942
rect 14588 22878 14590 22930
rect 14642 22878 14644 22930
rect 14476 22372 14532 22382
rect 14476 22278 14532 22316
rect 14588 21698 14644 22878
rect 14924 22484 14980 22494
rect 14924 22258 14980 22428
rect 14924 22206 14926 22258
rect 14978 22206 14980 22258
rect 14588 21646 14590 21698
rect 14642 21646 14644 21698
rect 14588 21634 14644 21646
rect 14700 21812 14756 21822
rect 14700 21586 14756 21756
rect 14700 21534 14702 21586
rect 14754 21534 14756 21586
rect 14700 21522 14756 21534
rect 14924 21362 14980 22206
rect 15260 22482 15316 22494
rect 15260 22430 15262 22482
rect 15314 22430 15316 22482
rect 15148 22146 15204 22158
rect 15148 22094 15150 22146
rect 15202 22094 15204 22146
rect 15148 21812 15204 22094
rect 15260 22036 15316 22430
rect 15708 22484 15764 22494
rect 15708 22390 15764 22428
rect 15932 22370 15988 22382
rect 15932 22318 15934 22370
rect 15986 22318 15988 22370
rect 15260 21980 15764 22036
rect 14924 21310 14926 21362
rect 14978 21310 14980 21362
rect 14924 21252 14980 21310
rect 15036 21756 15148 21812
rect 15036 21364 15092 21756
rect 15148 21746 15204 21756
rect 15148 21588 15204 21598
rect 15596 21588 15652 21598
rect 15148 21586 15652 21588
rect 15148 21534 15150 21586
rect 15202 21534 15598 21586
rect 15650 21534 15652 21586
rect 15148 21532 15652 21534
rect 15708 21588 15764 21980
rect 15932 21812 15988 22318
rect 15932 21746 15988 21756
rect 16492 21698 16548 22988
rect 16604 22484 16660 22494
rect 16604 22390 16660 22428
rect 17500 22260 17556 22270
rect 17388 22204 17500 22260
rect 17388 22146 17444 22204
rect 17500 22194 17556 22204
rect 17724 22258 17780 22270
rect 17724 22206 17726 22258
rect 17778 22206 17780 22258
rect 17388 22094 17390 22146
rect 17442 22094 17444 22146
rect 17388 22082 17444 22094
rect 17612 22148 17668 22158
rect 17612 22054 17668 22092
rect 17724 21924 17780 22206
rect 17724 21858 17780 21868
rect 16492 21646 16494 21698
rect 16546 21646 16548 21698
rect 16492 21634 16548 21646
rect 15820 21588 15876 21598
rect 15708 21586 15876 21588
rect 15708 21534 15822 21586
rect 15874 21534 15876 21586
rect 15708 21532 15876 21534
rect 15148 21522 15204 21532
rect 15036 21308 15204 21364
rect 14364 21196 14532 21252
rect 14924 21196 15092 21252
rect 14140 21186 14196 21196
rect 13804 20916 13860 20926
rect 14364 20916 14420 20926
rect 13804 20914 14420 20916
rect 13804 20862 13806 20914
rect 13858 20862 14366 20914
rect 14418 20862 14420 20914
rect 13804 20860 14420 20862
rect 13804 20850 13860 20860
rect 14364 20850 14420 20860
rect 12460 20750 12462 20802
rect 12514 20750 12516 20802
rect 12460 20242 12516 20750
rect 13580 20802 13636 20814
rect 13580 20750 13582 20802
rect 13634 20750 13636 20802
rect 13580 20244 13636 20750
rect 13916 20692 13972 20702
rect 14476 20692 14532 21196
rect 13916 20598 13972 20636
rect 14364 20636 14532 20692
rect 14588 20802 14644 20814
rect 14812 20804 14868 20814
rect 14588 20750 14590 20802
rect 14642 20750 14644 20802
rect 12460 20190 12462 20242
rect 12514 20190 12516 20242
rect 12460 20178 12516 20190
rect 13356 20188 13636 20244
rect 13244 19908 13300 19918
rect 13356 19908 13412 20188
rect 13300 19852 13412 19908
rect 14252 20132 14308 20142
rect 13244 19814 13300 19852
rect 11564 19182 11566 19234
rect 11618 19182 11620 19234
rect 11564 19170 11620 19182
rect 12012 19740 12180 19796
rect 11676 19124 11732 19134
rect 11676 19030 11732 19068
rect 11452 18900 11508 18910
rect 11452 18450 11508 18844
rect 11452 18398 11454 18450
rect 11506 18398 11508 18450
rect 11452 18228 11508 18398
rect 11452 18162 11508 18172
rect 11788 18562 11844 18574
rect 11788 18510 11790 18562
rect 11842 18510 11844 18562
rect 11788 18452 11844 18510
rect 11452 17556 11508 17566
rect 11676 17556 11732 17566
rect 11452 17554 11732 17556
rect 11452 17502 11454 17554
rect 11506 17502 11678 17554
rect 11730 17502 11732 17554
rect 11452 17500 11732 17502
rect 11452 17490 11508 17500
rect 11676 17490 11732 17500
rect 10892 17350 10948 17388
rect 11116 17388 11284 17444
rect 11340 17442 11396 17454
rect 11340 17390 11342 17442
rect 11394 17390 11396 17442
rect 10332 17164 10500 17220
rect 10108 16996 10164 17006
rect 9884 16994 10164 16996
rect 9884 16942 10110 16994
rect 10162 16942 10164 16994
rect 9884 16940 10164 16942
rect 9548 16882 9604 16894
rect 9548 16830 9550 16882
rect 9602 16830 9604 16882
rect 9548 16322 9604 16830
rect 9548 16270 9550 16322
rect 9602 16270 9604 16322
rect 9548 16258 9604 16270
rect 9884 16322 9940 16940
rect 10108 16930 10164 16940
rect 9996 16772 10052 16782
rect 9996 16678 10052 16716
rect 9884 16270 9886 16322
rect 9938 16270 9940 16322
rect 9884 16258 9940 16270
rect 9548 16098 9604 16110
rect 9548 16046 9550 16098
rect 9602 16046 9604 16098
rect 9548 15876 9604 16046
rect 10220 16098 10276 16110
rect 10220 16046 10222 16098
rect 10274 16046 10276 16098
rect 9548 15810 9604 15820
rect 9884 15876 9940 15886
rect 9660 15764 9716 15774
rect 9660 15314 9716 15708
rect 9884 15538 9940 15820
rect 10220 15876 10276 16046
rect 10220 15810 10276 15820
rect 9884 15486 9886 15538
rect 9938 15486 9940 15538
rect 9884 15474 9940 15486
rect 9660 15262 9662 15314
rect 9714 15262 9716 15314
rect 9660 15250 9716 15262
rect 9436 15092 9716 15148
rect 8204 14018 8260 14028
rect 8316 14308 8372 14318
rect 5964 13906 6020 13916
rect 6972 13972 7028 13982
rect 6972 13878 7028 13916
rect 6524 13858 6580 13870
rect 6524 13806 6526 13858
rect 6578 13806 6580 13858
rect 6300 13748 6356 13758
rect 6524 13748 6580 13806
rect 6860 13748 6916 13758
rect 6300 13746 6468 13748
rect 6300 13694 6302 13746
rect 6354 13694 6468 13746
rect 6300 13692 6468 13694
rect 6524 13746 6916 13748
rect 6524 13694 6862 13746
rect 6914 13694 6916 13746
rect 6524 13692 6916 13694
rect 6300 13682 6356 13692
rect 5964 12852 6020 12862
rect 5740 12850 6020 12852
rect 5740 12798 5966 12850
rect 6018 12798 6020 12850
rect 5740 12796 6020 12798
rect 5516 12292 5572 12302
rect 5572 12236 5684 12292
rect 5516 12198 5572 12236
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4844 11620 4900 11788
rect 4732 11564 4900 11620
rect 5180 11788 5460 11844
rect 4620 11508 4676 11518
rect 3836 11506 4676 11508
rect 3836 11454 4622 11506
rect 4674 11454 4676 11506
rect 3836 11452 4676 11454
rect 4620 11442 4676 11452
rect 3724 11394 4228 11396
rect 3724 11342 3726 11394
rect 3778 11342 4228 11394
rect 3724 11340 4228 11342
rect 3724 11330 3780 11340
rect 3948 11172 4004 11182
rect 3836 10836 3892 10846
rect 3612 10834 3892 10836
rect 3612 10782 3838 10834
rect 3890 10782 3892 10834
rect 3612 10780 3892 10782
rect 3500 10742 3556 10780
rect 3836 10770 3892 10780
rect 3948 10612 4004 11116
rect 4172 11060 4228 11340
rect 4284 11284 4340 11294
rect 4732 11284 4788 11564
rect 4956 11508 5012 11518
rect 4956 11414 5012 11452
rect 4284 11282 4788 11284
rect 4284 11230 4286 11282
rect 4338 11230 4788 11282
rect 4284 11228 4788 11230
rect 4284 11218 4340 11228
rect 4844 11170 4900 11182
rect 4844 11118 4846 11170
rect 4898 11118 4900 11170
rect 4844 11060 4900 11118
rect 4172 11004 4900 11060
rect 4508 10722 4564 10734
rect 5068 10724 5124 10734
rect 4508 10670 4510 10722
rect 4562 10670 4564 10722
rect 4060 10612 4116 10622
rect 3948 10556 4060 10612
rect 4060 10546 4116 10556
rect 4284 10610 4340 10622
rect 4284 10558 4286 10610
rect 4338 10558 4340 10610
rect 3836 10052 3892 10062
rect 3836 9714 3892 9996
rect 3836 9662 3838 9714
rect 3890 9662 3892 9714
rect 3500 9268 3556 9278
rect 3388 9212 3500 9268
rect 3500 9202 3556 9212
rect 3836 9044 3892 9662
rect 3836 8978 3892 8988
rect 4172 9826 4228 9838
rect 4172 9774 4174 9826
rect 4226 9774 4228 9826
rect 4172 9716 4228 9774
rect 4172 9042 4228 9660
rect 4284 9156 4340 10558
rect 4508 10500 4564 10670
rect 4508 10434 4564 10444
rect 4844 10668 5068 10724
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4844 9828 4900 10668
rect 5068 10630 5124 10668
rect 5068 10500 5124 10510
rect 4956 9940 5012 9950
rect 4956 9846 5012 9884
rect 4732 9826 4900 9828
rect 4732 9774 4846 9826
rect 4898 9774 4900 9826
rect 4732 9772 4900 9774
rect 4732 9492 4788 9772
rect 4284 9062 4340 9100
rect 4508 9436 4788 9492
rect 4508 9154 4564 9436
rect 4508 9102 4510 9154
rect 4562 9102 4564 9154
rect 4508 9090 4564 9102
rect 4172 8990 4174 9042
rect 4226 8990 4228 9042
rect 3612 8930 3668 8942
rect 3612 8878 3614 8930
rect 3666 8878 3668 8930
rect 3612 8820 3668 8878
rect 3612 8754 3668 8764
rect 4172 8428 4228 8990
rect 4620 9044 4676 9054
rect 4620 8950 4676 8988
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 4844 8428 4900 9772
rect 4956 9716 5012 9726
rect 5068 9716 5124 10444
rect 4956 9714 5124 9716
rect 4956 9662 4958 9714
rect 5010 9662 5124 9714
rect 4956 9660 5124 9662
rect 4956 9604 5012 9660
rect 4956 9538 5012 9548
rect 5180 9380 5236 11788
rect 5628 11396 5684 12236
rect 5740 12068 5796 12796
rect 5964 12786 6020 12796
rect 6300 12738 6356 12750
rect 6300 12686 6302 12738
rect 6354 12686 6356 12738
rect 6300 12516 6356 12686
rect 6412 12516 6468 13692
rect 6860 13300 6916 13692
rect 6972 13524 7028 13534
rect 6972 13430 7028 13468
rect 6860 13244 7140 13300
rect 6636 12962 6692 12974
rect 6636 12910 6638 12962
rect 6690 12910 6692 12962
rect 6412 12460 6580 12516
rect 6300 12450 6356 12460
rect 5852 12290 5908 12302
rect 5852 12238 5854 12290
rect 5906 12238 5908 12290
rect 5852 12180 5908 12238
rect 6412 12292 6468 12302
rect 6300 12180 6356 12190
rect 5852 12124 6300 12180
rect 6300 12086 6356 12124
rect 6412 12178 6468 12236
rect 6412 12126 6414 12178
rect 6466 12126 6468 12178
rect 5740 11620 5796 12012
rect 6300 11844 6356 11854
rect 6412 11844 6468 12126
rect 6356 11788 6468 11844
rect 6524 12290 6580 12460
rect 6524 12238 6526 12290
rect 6578 12238 6580 12290
rect 6300 11778 6356 11788
rect 5740 11554 5796 11564
rect 6300 11618 6356 11630
rect 6300 11566 6302 11618
rect 6354 11566 6356 11618
rect 5292 11394 5684 11396
rect 5292 11342 5630 11394
rect 5682 11342 5684 11394
rect 5292 11340 5684 11342
rect 5292 10610 5348 11340
rect 5628 11330 5684 11340
rect 5740 11284 5796 11294
rect 5740 11190 5796 11228
rect 5292 10558 5294 10610
rect 5346 10558 5348 10610
rect 5292 10546 5348 10558
rect 5852 10612 5908 10622
rect 5852 10518 5908 10556
rect 6188 10386 6244 10398
rect 6188 10334 6190 10386
rect 6242 10334 6244 10386
rect 5180 9314 5236 9324
rect 5292 10164 5348 10174
rect 5292 9156 5348 10108
rect 6188 9714 6244 10334
rect 6300 9826 6356 11566
rect 6412 11396 6468 11406
rect 6412 11302 6468 11340
rect 6524 11284 6580 12238
rect 6636 12180 6692 12910
rect 6860 12852 6916 12862
rect 7084 12852 7140 13244
rect 7868 13076 7924 13086
rect 6860 12850 7028 12852
rect 6860 12798 6862 12850
rect 6914 12798 7028 12850
rect 6860 12796 7028 12798
rect 6860 12786 6916 12796
rect 6636 12114 6692 12124
rect 6748 12178 6804 12190
rect 6748 12126 6750 12178
rect 6802 12126 6804 12178
rect 6748 12068 6804 12126
rect 6804 12012 6916 12068
rect 6748 12002 6804 12012
rect 6860 11394 6916 12012
rect 6860 11342 6862 11394
rect 6914 11342 6916 11394
rect 6860 11330 6916 11342
rect 6972 11396 7028 12796
rect 7084 12758 7140 12796
rect 7420 12962 7476 12974
rect 7420 12910 7422 12962
rect 7474 12910 7476 12962
rect 7420 12516 7476 12910
rect 7420 12450 7476 12460
rect 7532 12964 7588 12974
rect 7196 12180 7252 12190
rect 7532 12180 7588 12908
rect 7644 12740 7700 12750
rect 7868 12740 7924 13020
rect 7644 12738 7924 12740
rect 7644 12686 7646 12738
rect 7698 12686 7924 12738
rect 7644 12684 7924 12686
rect 7644 12674 7700 12684
rect 7196 12178 7812 12180
rect 7196 12126 7198 12178
rect 7250 12126 7534 12178
rect 7586 12126 7812 12178
rect 7196 12124 7812 12126
rect 7196 12114 7252 12124
rect 7532 12114 7588 12124
rect 7644 11844 7700 11854
rect 7308 11788 7644 11844
rect 7028 11340 7140 11396
rect 6972 11330 7028 11340
rect 6524 11218 6580 11228
rect 6412 10610 6468 10622
rect 6412 10558 6414 10610
rect 6466 10558 6468 10610
rect 6412 10164 6468 10558
rect 6412 10098 6468 10108
rect 6748 9940 6804 9950
rect 6300 9774 6302 9826
rect 6354 9774 6356 9826
rect 6300 9762 6356 9774
rect 6412 9938 6804 9940
rect 6412 9886 6750 9938
rect 6802 9886 6804 9938
rect 6412 9884 6804 9886
rect 6188 9662 6190 9714
rect 6242 9662 6244 9714
rect 6188 9650 6244 9662
rect 5404 9268 5460 9278
rect 5404 9174 5460 9212
rect 5292 9062 5348 9100
rect 5068 9044 5124 9054
rect 5068 8950 5124 8988
rect 5628 9042 5684 9054
rect 5628 8990 5630 9042
rect 5682 8990 5684 9042
rect 4172 8372 4564 8428
rect 2492 8318 2494 8370
rect 2546 8318 2548 8370
rect 2492 8306 2548 8318
rect 4396 8258 4452 8270
rect 4396 8206 4398 8258
rect 4450 8206 4452 8258
rect 2940 8148 2996 8158
rect 2940 8054 2996 8092
rect 1820 7646 1822 7698
rect 1874 7646 1876 7698
rect 1820 7634 1876 7646
rect 2044 8034 2100 8046
rect 2044 7982 2046 8034
rect 2098 7982 2100 8034
rect 2044 7476 2100 7982
rect 4396 7924 4452 8206
rect 4508 8146 4564 8372
rect 4508 8094 4510 8146
rect 4562 8094 4564 8146
rect 4508 8082 4564 8094
rect 4620 8372 4900 8428
rect 5628 8428 5684 8990
rect 6412 9044 6468 9884
rect 6748 9874 6804 9884
rect 6972 9940 7028 9950
rect 6972 9826 7028 9884
rect 6972 9774 6974 9826
rect 7026 9774 7028 9826
rect 6972 9762 7028 9774
rect 6748 9716 6804 9726
rect 6748 9622 6804 9660
rect 7084 9604 7140 11340
rect 6636 9268 6692 9278
rect 6636 9174 6692 9212
rect 6412 8950 6468 8988
rect 7084 9042 7140 9548
rect 7308 9268 7364 11788
rect 7644 11778 7700 11788
rect 7756 10722 7812 12124
rect 7756 10670 7758 10722
rect 7810 10670 7812 10722
rect 7756 10658 7812 10670
rect 7868 10612 7924 12684
rect 8204 12292 8260 12302
rect 7980 12068 8036 12078
rect 7980 11974 8036 12012
rect 8204 12068 8260 12236
rect 8204 12002 8260 12012
rect 8316 12290 8372 14252
rect 9212 13412 9268 13422
rect 8540 13300 8596 13310
rect 8540 12516 8596 13244
rect 8652 12964 8708 12974
rect 8652 12870 8708 12908
rect 8876 12964 8932 12974
rect 9100 12964 9156 12974
rect 8876 12628 8932 12908
rect 8876 12562 8932 12572
rect 8988 12962 9156 12964
rect 8988 12910 9102 12962
rect 9154 12910 9156 12962
rect 8988 12908 9156 12910
rect 8540 12402 8596 12460
rect 8540 12350 8542 12402
rect 8594 12350 8596 12402
rect 8540 12338 8596 12350
rect 8652 12404 8708 12414
rect 8988 12404 9044 12908
rect 9100 12898 9156 12908
rect 8652 12402 9044 12404
rect 8652 12350 8654 12402
rect 8706 12350 9044 12402
rect 8652 12348 9044 12350
rect 9212 12852 9268 13356
rect 8652 12338 8708 12348
rect 8316 12238 8318 12290
rect 8370 12238 8372 12290
rect 8316 11844 8372 12238
rect 8764 12180 8820 12190
rect 8764 12086 8820 12124
rect 8988 12180 9044 12190
rect 9212 12180 9268 12796
rect 9548 12852 9604 12862
rect 9548 12758 9604 12796
rect 8988 12178 9268 12180
rect 8988 12126 8990 12178
rect 9042 12126 9268 12178
rect 8988 12124 9268 12126
rect 9548 12628 9604 12638
rect 9548 12178 9604 12572
rect 9548 12126 9550 12178
rect 9602 12126 9604 12178
rect 8988 12114 9044 12124
rect 8316 11778 8372 11788
rect 9212 11956 9268 11966
rect 9212 11506 9268 11900
rect 9212 11454 9214 11506
rect 9266 11454 9268 11506
rect 7980 10612 8036 10622
rect 7868 10610 8036 10612
rect 7868 10558 7982 10610
rect 8034 10558 8036 10610
rect 7868 10556 8036 10558
rect 7980 10546 8036 10556
rect 8988 10500 9044 10510
rect 8988 10406 9044 10444
rect 8204 10388 8260 10398
rect 8092 10386 8260 10388
rect 8092 10334 8206 10386
rect 8258 10334 8260 10386
rect 8092 10332 8260 10334
rect 7756 9716 7812 9726
rect 7308 9266 7476 9268
rect 7308 9214 7310 9266
rect 7362 9214 7476 9266
rect 7308 9212 7476 9214
rect 7308 9202 7364 9212
rect 7084 8990 7086 9042
rect 7138 8990 7140 9042
rect 7084 8978 7140 8990
rect 7196 9044 7252 9054
rect 7196 8428 7252 8988
rect 5628 8372 5796 8428
rect 7196 8372 7364 8428
rect 4620 7924 4676 8372
rect 4732 8260 4788 8270
rect 4732 8166 4788 8204
rect 5404 8260 5460 8270
rect 4396 7868 4676 7924
rect 5404 7586 5460 8204
rect 5404 7534 5406 7586
rect 5458 7534 5460 7586
rect 5404 7522 5460 7534
rect 5740 8258 5796 8372
rect 5740 8206 5742 8258
rect 5794 8206 5796 8258
rect 2044 7410 2100 7420
rect 5628 7476 5684 7486
rect 5740 7476 5796 8206
rect 5964 8260 6020 8270
rect 5964 8166 6020 8204
rect 6636 8260 6692 8270
rect 6636 8166 6692 8204
rect 7084 8260 7140 8270
rect 7084 8146 7140 8204
rect 7308 8258 7364 8372
rect 7420 8372 7476 9212
rect 7756 9154 7812 9660
rect 7756 9102 7758 9154
rect 7810 9102 7812 9154
rect 7756 8428 7812 9102
rect 8092 9604 8148 10332
rect 8204 10322 8260 10332
rect 8428 10386 8484 10398
rect 8428 10334 8430 10386
rect 8482 10334 8484 10386
rect 8428 10052 8484 10334
rect 8204 9996 8484 10052
rect 8204 9940 8260 9996
rect 8204 9826 8260 9884
rect 8428 9828 8484 9838
rect 9212 9828 9268 11454
rect 9548 9938 9604 12126
rect 9660 12402 9716 15092
rect 10108 14530 10164 14542
rect 10108 14478 10110 14530
rect 10162 14478 10164 14530
rect 9996 13412 10052 13422
rect 10108 13412 10164 14478
rect 10052 13356 10164 13412
rect 9996 13346 10052 13356
rect 10332 13300 10388 17164
rect 10444 16324 10500 16334
rect 10444 16210 10500 16268
rect 10444 16158 10446 16210
rect 10498 16158 10500 16210
rect 10444 16146 10500 16158
rect 10556 14530 10612 14542
rect 10556 14478 10558 14530
rect 10610 14478 10612 14530
rect 10556 14196 10612 14478
rect 10892 14308 10948 14318
rect 10892 14214 10948 14252
rect 10556 14130 10612 14140
rect 10108 13244 10388 13300
rect 10668 13634 10724 13646
rect 10668 13582 10670 13634
rect 10722 13582 10724 13634
rect 10108 12850 10164 13244
rect 10444 12964 10500 12974
rect 10108 12798 10110 12850
rect 10162 12798 10164 12850
rect 9660 12350 9662 12402
rect 9714 12350 9716 12402
rect 9660 11956 9716 12350
rect 9772 12738 9828 12750
rect 9772 12686 9774 12738
rect 9826 12686 9828 12738
rect 9772 12180 9828 12686
rect 9884 12292 9940 12302
rect 9884 12198 9940 12236
rect 9772 12114 9828 12124
rect 9660 11890 9716 11900
rect 9996 11394 10052 11406
rect 9996 11342 9998 11394
rect 10050 11342 10052 11394
rect 9772 11282 9828 11294
rect 9772 11230 9774 11282
rect 9826 11230 9828 11282
rect 9660 10724 9716 10734
rect 9660 10630 9716 10668
rect 9548 9886 9550 9938
rect 9602 9886 9604 9938
rect 9548 9874 9604 9886
rect 9772 10610 9828 11230
rect 9772 10558 9774 10610
rect 9826 10558 9828 10610
rect 9324 9828 9380 9838
rect 8204 9774 8206 9826
rect 8258 9774 8260 9826
rect 8204 9762 8260 9774
rect 8316 9826 8484 9828
rect 8316 9774 8430 9826
rect 8482 9774 8484 9826
rect 8316 9772 8484 9774
rect 8316 9604 8372 9772
rect 8428 9762 8484 9772
rect 8652 9826 9380 9828
rect 8652 9774 9326 9826
rect 9378 9774 9380 9826
rect 8652 9772 9380 9774
rect 8092 9548 8372 9604
rect 8092 9268 8148 9548
rect 8092 9042 8148 9212
rect 8652 9266 8708 9772
rect 9324 9762 9380 9772
rect 9660 9716 9716 9726
rect 9772 9716 9828 10558
rect 9884 10610 9940 10622
rect 9884 10558 9886 10610
rect 9938 10558 9940 10610
rect 9884 10500 9940 10558
rect 9996 10500 10052 11342
rect 10108 11284 10164 12798
rect 10332 12962 10500 12964
rect 10332 12910 10446 12962
rect 10498 12910 10500 12962
rect 10332 12908 10500 12910
rect 10332 12292 10388 12908
rect 10444 12898 10500 12908
rect 10556 12852 10612 12862
rect 10444 12404 10500 12414
rect 10556 12404 10612 12796
rect 10444 12402 10612 12404
rect 10444 12350 10446 12402
rect 10498 12350 10612 12402
rect 10444 12348 10612 12350
rect 10668 12402 10724 13582
rect 10892 13524 10948 13534
rect 11116 13524 11172 17388
rect 11340 17332 11396 17390
rect 11788 17444 11844 18396
rect 11900 18228 11956 18238
rect 11900 17554 11956 18172
rect 12012 17780 12068 19740
rect 12124 19460 12180 19470
rect 12124 19366 12180 19404
rect 12572 19236 12628 19246
rect 12572 19142 12628 19180
rect 12236 19122 12292 19134
rect 12236 19070 12238 19122
rect 12290 19070 12292 19122
rect 12124 19012 12180 19022
rect 12124 18918 12180 18956
rect 12236 18788 12292 19070
rect 12236 17892 12292 18732
rect 12684 19122 12740 19134
rect 12684 19070 12686 19122
rect 12738 19070 12740 19122
rect 12684 18676 12740 19070
rect 12684 18610 12740 18620
rect 13468 18900 13524 18910
rect 13468 18674 13524 18844
rect 13468 18622 13470 18674
rect 13522 18622 13524 18674
rect 13356 18564 13412 18574
rect 12348 18340 12404 18350
rect 12348 18338 12516 18340
rect 12348 18286 12350 18338
rect 12402 18286 12516 18338
rect 12348 18284 12516 18286
rect 12348 18274 12404 18284
rect 12460 18116 12516 18284
rect 12236 17836 12404 17892
rect 12012 17724 12292 17780
rect 11900 17502 11902 17554
rect 11954 17502 11956 17554
rect 11900 17490 11956 17502
rect 12012 17554 12068 17566
rect 12012 17502 12014 17554
rect 12066 17502 12068 17554
rect 11788 17378 11844 17388
rect 11340 17266 11396 17276
rect 12012 17220 12068 17502
rect 12012 17164 12180 17220
rect 11900 17108 11956 17118
rect 11788 16098 11844 16110
rect 11788 16046 11790 16098
rect 11842 16046 11844 16098
rect 11788 15876 11844 16046
rect 11788 15810 11844 15820
rect 11228 15092 11284 15102
rect 11228 14418 11284 15036
rect 11228 14366 11230 14418
rect 11282 14366 11284 14418
rect 11228 14354 11284 14366
rect 10892 13522 11172 13524
rect 10892 13470 10894 13522
rect 10946 13470 11172 13522
rect 10892 13468 11172 13470
rect 11340 13746 11396 13758
rect 11340 13694 11342 13746
rect 11394 13694 11396 13746
rect 10892 13458 10948 13468
rect 11340 12964 11396 13694
rect 11788 12964 11844 12974
rect 11340 12962 11844 12964
rect 11340 12910 11342 12962
rect 11394 12910 11790 12962
rect 11842 12910 11844 12962
rect 11340 12908 11844 12910
rect 11340 12898 11396 12908
rect 11788 12898 11844 12908
rect 11452 12740 11508 12750
rect 10668 12350 10670 12402
rect 10722 12350 10724 12402
rect 10444 12338 10500 12348
rect 10668 12338 10724 12350
rect 11228 12738 11732 12740
rect 11228 12686 11454 12738
rect 11506 12686 11732 12738
rect 11228 12684 11732 12686
rect 10332 12198 10388 12236
rect 10108 11218 10164 11228
rect 10668 12180 10724 12190
rect 9940 10444 10164 10500
rect 9884 10406 9940 10444
rect 10108 9828 10164 10444
rect 10332 10386 10388 10398
rect 10332 10334 10334 10386
rect 10386 10334 10388 10386
rect 10332 10052 10388 10334
rect 10332 9986 10388 9996
rect 10332 9828 10388 9838
rect 10108 9826 10388 9828
rect 10108 9774 10334 9826
rect 10386 9774 10388 9826
rect 10108 9772 10388 9774
rect 10332 9762 10388 9772
rect 9660 9714 9772 9716
rect 9660 9662 9662 9714
rect 9714 9662 9772 9714
rect 9660 9660 9772 9662
rect 9660 9650 9716 9660
rect 9772 9622 9828 9660
rect 10444 9716 10500 9726
rect 10444 9622 10500 9660
rect 10668 9380 10724 12124
rect 10892 11394 10948 11406
rect 10892 11342 10894 11394
rect 10946 11342 10948 11394
rect 10780 11172 10836 11182
rect 10892 11172 10948 11342
rect 11116 11172 11172 11182
rect 10892 11170 11172 11172
rect 10892 11118 11118 11170
rect 11170 11118 11172 11170
rect 10892 11116 11172 11118
rect 10780 11078 10836 11116
rect 11004 10724 11060 11116
rect 11116 11106 11172 11116
rect 11004 9714 11060 10668
rect 11004 9662 11006 9714
rect 11058 9662 11060 9714
rect 11004 9650 11060 9662
rect 11116 10722 11172 10734
rect 11116 10670 11118 10722
rect 11170 10670 11172 10722
rect 11116 9602 11172 10670
rect 11228 10610 11284 12684
rect 11452 12674 11508 12684
rect 11676 12178 11732 12684
rect 11676 12126 11678 12178
rect 11730 12126 11732 12178
rect 11676 12114 11732 12126
rect 11564 12066 11620 12078
rect 11564 12014 11566 12066
rect 11618 12014 11620 12066
rect 11452 11844 11508 11854
rect 11340 11284 11396 11294
rect 11340 11190 11396 11228
rect 11452 11282 11508 11788
rect 11452 11230 11454 11282
rect 11506 11230 11508 11282
rect 11228 10558 11230 10610
rect 11282 10558 11284 10610
rect 11228 10546 11284 10558
rect 11116 9550 11118 9602
rect 11170 9550 11172 9602
rect 11116 9538 11172 9550
rect 10668 9324 11284 9380
rect 8652 9214 8654 9266
rect 8706 9214 8708 9266
rect 8652 9202 8708 9214
rect 9884 9268 9940 9278
rect 9884 9174 9940 9212
rect 8092 8990 8094 9042
rect 8146 8990 8148 9042
rect 7420 8306 7476 8316
rect 7532 8372 7812 8428
rect 7980 8930 8036 8942
rect 7980 8878 7982 8930
rect 8034 8878 8036 8930
rect 7308 8206 7310 8258
rect 7362 8206 7364 8258
rect 7308 8194 7364 8206
rect 7084 8094 7086 8146
rect 7138 8094 7140 8146
rect 7084 8082 7140 8094
rect 7420 8036 7476 8046
rect 7420 7942 7476 7980
rect 7532 8034 7588 8372
rect 7980 8370 8036 8878
rect 7980 8318 7982 8370
rect 8034 8318 8036 8370
rect 7980 8306 8036 8318
rect 7532 7982 7534 8034
rect 7586 7982 7588 8034
rect 5628 7474 5796 7476
rect 5628 7422 5630 7474
rect 5682 7422 5796 7474
rect 5628 7420 5796 7422
rect 5628 7410 5684 7420
rect 5964 7252 6020 7262
rect 7532 7252 7588 7982
rect 7980 7476 8036 7486
rect 8092 7476 8148 8990
rect 9660 9042 9716 9054
rect 10220 9044 10276 9054
rect 9660 8990 9662 9042
rect 9714 8990 9716 9042
rect 9660 8428 9716 8990
rect 10108 9042 10276 9044
rect 10108 8990 10222 9042
rect 10274 8990 10276 9042
rect 10108 8988 10276 8990
rect 9548 8372 9604 8382
rect 9660 8372 9828 8428
rect 8316 8258 8372 8270
rect 8316 8206 8318 8258
rect 8370 8206 8372 8258
rect 8316 8148 8372 8206
rect 8316 8082 8372 8092
rect 8428 8260 8484 8270
rect 7980 7474 8148 7476
rect 7980 7422 7982 7474
rect 8034 7422 8148 7474
rect 7980 7420 8148 7422
rect 8428 7474 8484 8204
rect 9436 8260 9492 8270
rect 9436 8166 9492 8204
rect 8876 7700 8932 7710
rect 8876 7606 8932 7644
rect 8428 7422 8430 7474
rect 8482 7422 8484 7474
rect 7980 7410 8036 7420
rect 8428 7410 8484 7422
rect 9548 7474 9604 8316
rect 9548 7422 9550 7474
rect 9602 7422 9604 7474
rect 9548 7410 9604 7422
rect 9772 7476 9828 8372
rect 10108 8148 10164 8988
rect 10220 8978 10276 8988
rect 11116 9042 11172 9054
rect 11116 8990 11118 9042
rect 11170 8990 11172 9042
rect 11004 8930 11060 8942
rect 11004 8878 11006 8930
rect 11058 8878 11060 8930
rect 10220 8372 10276 8382
rect 10220 8278 10276 8316
rect 10108 7698 10164 8092
rect 10108 7646 10110 7698
rect 10162 7646 10164 7698
rect 10108 7634 10164 7646
rect 9772 7382 9828 7420
rect 11004 7476 11060 8878
rect 11116 8258 11172 8990
rect 11116 8206 11118 8258
rect 11170 8206 11172 8258
rect 11116 7700 11172 8206
rect 11228 7924 11284 9324
rect 11452 9268 11508 11230
rect 11564 10836 11620 12014
rect 11900 11506 11956 17052
rect 12012 16994 12068 17006
rect 12012 16942 12014 16994
rect 12066 16942 12068 16994
rect 12012 16436 12068 16942
rect 12012 16370 12068 16380
rect 12012 15988 12068 15998
rect 12124 15988 12180 17164
rect 12236 17108 12292 17724
rect 12236 17042 12292 17052
rect 12012 15986 12124 15988
rect 12012 15934 12014 15986
rect 12066 15934 12124 15986
rect 12012 15932 12124 15934
rect 12012 15922 12068 15932
rect 12124 15894 12180 15932
rect 12236 16884 12292 16894
rect 12124 15314 12180 15326
rect 12124 15262 12126 15314
rect 12178 15262 12180 15314
rect 12124 14530 12180 15262
rect 12124 14478 12126 14530
rect 12178 14478 12180 14530
rect 12124 13300 12180 14478
rect 12236 14644 12292 16828
rect 12348 16436 12404 17836
rect 12460 17556 12516 18060
rect 13356 17892 13412 18508
rect 13468 18452 13524 18622
rect 14252 18674 14308 20076
rect 14252 18622 14254 18674
rect 14306 18622 14308 18674
rect 14252 18610 14308 18622
rect 13468 18386 13524 18396
rect 13916 18450 13972 18462
rect 13916 18398 13918 18450
rect 13970 18398 13972 18450
rect 13916 18340 13972 18398
rect 14364 18340 14420 20636
rect 14588 20468 14644 20750
rect 14588 20402 14644 20412
rect 14700 20748 14812 20804
rect 13916 18274 13972 18284
rect 14252 18284 14420 18340
rect 14476 20244 14532 20254
rect 14476 20130 14532 20188
rect 14588 20244 14644 20254
rect 14700 20244 14756 20748
rect 14812 20738 14868 20748
rect 14588 20242 14756 20244
rect 14588 20190 14590 20242
rect 14642 20190 14756 20242
rect 14588 20188 14756 20190
rect 14588 20178 14644 20188
rect 14476 20078 14478 20130
rect 14530 20078 14532 20130
rect 13468 18228 13524 18238
rect 13468 18134 13524 18172
rect 12908 17836 13412 17892
rect 12684 17556 12740 17566
rect 12460 17554 12740 17556
rect 12460 17502 12686 17554
rect 12738 17502 12740 17554
rect 12460 17500 12740 17502
rect 12684 16996 12740 17500
rect 12796 17442 12852 17454
rect 12796 17390 12798 17442
rect 12850 17390 12852 17442
rect 12796 17220 12852 17390
rect 12796 17154 12852 17164
rect 12684 16940 12852 16996
rect 12348 16370 12404 16380
rect 12796 16212 12852 16940
rect 12796 16146 12852 16156
rect 12684 16100 12740 16110
rect 12460 16044 12684 16100
rect 12460 15538 12516 16044
rect 12684 16006 12740 16044
rect 12796 15876 12852 15886
rect 12796 15782 12852 15820
rect 12908 15652 12964 17836
rect 13580 17778 13636 17790
rect 13580 17726 13582 17778
rect 13634 17726 13636 17778
rect 13020 17668 13076 17678
rect 13580 17668 13636 17726
rect 13020 17666 13636 17668
rect 13020 17614 13022 17666
rect 13074 17614 13636 17666
rect 13020 17612 13636 17614
rect 13692 17668 13748 17678
rect 13020 17602 13076 17612
rect 13692 17574 13748 17612
rect 13356 17444 13412 17454
rect 12460 15486 12462 15538
rect 12514 15486 12516 15538
rect 12460 15474 12516 15486
rect 12684 15596 12964 15652
rect 13020 15874 13076 15886
rect 13020 15822 13022 15874
rect 13074 15822 13076 15874
rect 12684 15092 12740 15596
rect 12684 15026 12740 15036
rect 12796 15316 12852 15326
rect 13020 15316 13076 15822
rect 13132 15316 13188 15326
rect 13020 15314 13188 15316
rect 13020 15262 13134 15314
rect 13186 15262 13188 15314
rect 13020 15260 13188 15262
rect 12796 14754 12852 15260
rect 13132 15250 13188 15260
rect 12796 14702 12798 14754
rect 12850 14702 12852 14754
rect 12796 14690 12852 14702
rect 12236 14588 12740 14644
rect 12236 14418 12292 14588
rect 12684 14532 12740 14588
rect 12684 14476 12852 14532
rect 12236 14366 12238 14418
rect 12290 14366 12292 14418
rect 12796 14418 12852 14476
rect 12236 14354 12292 14366
rect 12684 14362 12740 14374
rect 12460 14308 12516 14318
rect 12684 14310 12686 14362
rect 12738 14310 12740 14362
rect 12796 14366 12798 14418
rect 12850 14366 12852 14418
rect 12796 14354 12852 14366
rect 12460 14306 12628 14308
rect 12460 14254 12462 14306
rect 12514 14254 12628 14306
rect 12460 14252 12628 14254
rect 12460 14242 12516 14252
rect 12572 13748 12628 14252
rect 12684 14196 12740 14310
rect 12684 14130 12740 14140
rect 13356 14196 13412 17388
rect 14028 16884 14084 16894
rect 13804 16100 13860 16110
rect 13692 16098 13860 16100
rect 13692 16046 13806 16098
rect 13858 16046 13860 16098
rect 13692 16044 13860 16046
rect 13692 15316 13748 16044
rect 13804 16034 13860 16044
rect 13692 15222 13748 15260
rect 13356 14130 13412 14140
rect 12684 13748 12740 13758
rect 12572 13692 12684 13748
rect 12684 13654 12740 13692
rect 12908 13746 12964 13758
rect 12908 13694 12910 13746
rect 12962 13694 12964 13746
rect 12908 13524 12964 13694
rect 12908 13458 12964 13468
rect 13580 13634 13636 13646
rect 13580 13582 13582 13634
rect 13634 13582 13636 13634
rect 12124 13234 12180 13244
rect 12124 12850 12180 12862
rect 12124 12798 12126 12850
rect 12178 12798 12180 12850
rect 12012 12738 12068 12750
rect 12012 12686 12014 12738
rect 12066 12686 12068 12738
rect 12012 12404 12068 12686
rect 12012 12068 12068 12348
rect 12012 12002 12068 12012
rect 12124 12740 12180 12798
rect 12124 11844 12180 12684
rect 12124 11778 12180 11788
rect 12348 12066 12404 12078
rect 12348 12014 12350 12066
rect 12402 12014 12404 12066
rect 12348 11620 12404 12014
rect 13580 11620 13636 13582
rect 13916 13634 13972 13646
rect 13916 13582 13918 13634
rect 13970 13582 13972 13634
rect 13916 13524 13972 13582
rect 13916 13458 13972 13468
rect 14028 12628 14084 16828
rect 14252 15148 14308 18284
rect 14476 17556 14532 20078
rect 14700 20020 14756 20030
rect 14700 19926 14756 19964
rect 14924 20018 14980 20030
rect 14924 19966 14926 20018
rect 14978 19966 14980 20018
rect 14476 17500 14644 17556
rect 14364 16882 14420 16894
rect 14364 16830 14366 16882
rect 14418 16830 14420 16882
rect 14364 16324 14420 16830
rect 14364 16258 14420 16268
rect 14476 16772 14532 16782
rect 14476 15988 14532 16716
rect 14588 16100 14644 17500
rect 14924 17444 14980 19966
rect 15036 19684 15092 21196
rect 15148 19796 15204 21308
rect 15260 20914 15316 21532
rect 15596 21522 15652 21532
rect 15820 21522 15876 21532
rect 17612 21586 17668 21598
rect 17612 21534 17614 21586
rect 17666 21534 17668 21586
rect 17612 21252 17668 21534
rect 17164 21196 17668 21252
rect 17724 21474 17780 21486
rect 17724 21422 17726 21474
rect 17778 21422 17780 21474
rect 16156 21028 16212 21038
rect 16156 20934 16212 20972
rect 15260 20862 15262 20914
rect 15314 20862 15316 20914
rect 15260 20850 15316 20862
rect 15596 20804 15652 20814
rect 15596 20710 15652 20748
rect 15820 20802 15876 20814
rect 15820 20750 15822 20802
rect 15874 20750 15876 20802
rect 15820 20468 15876 20750
rect 15820 20402 15876 20412
rect 16044 20802 16100 20814
rect 16044 20750 16046 20802
rect 16098 20750 16100 20802
rect 15260 20132 15316 20142
rect 15260 20038 15316 20076
rect 15372 20132 15428 20142
rect 15372 20130 15540 20132
rect 15372 20078 15374 20130
rect 15426 20078 15540 20130
rect 15372 20076 15540 20078
rect 15372 20066 15428 20076
rect 15484 19908 15540 20076
rect 15372 19796 15428 19806
rect 15148 19794 15428 19796
rect 15148 19742 15374 19794
rect 15426 19742 15428 19794
rect 15148 19740 15428 19742
rect 15372 19730 15428 19740
rect 15036 19628 15316 19684
rect 15260 19012 15316 19628
rect 15484 19460 15540 19852
rect 15932 19908 15988 19918
rect 16044 19908 16100 20750
rect 17164 20802 17220 21196
rect 17500 21028 17556 21038
rect 17724 21028 17780 21422
rect 17500 21026 17780 21028
rect 17500 20974 17502 21026
rect 17554 20974 17780 21026
rect 17500 20972 17780 20974
rect 17500 20962 17556 20972
rect 17164 20750 17166 20802
rect 17218 20750 17220 20802
rect 17164 20738 17220 20750
rect 17388 20804 17444 20814
rect 17388 20710 17444 20748
rect 16828 20690 16884 20702
rect 16828 20638 16830 20690
rect 16882 20638 16884 20690
rect 15932 19906 16100 19908
rect 15932 19854 15934 19906
rect 15986 19854 16100 19906
rect 15932 19852 16100 19854
rect 16268 20132 16324 20142
rect 15932 19796 15988 19852
rect 15932 19730 15988 19740
rect 15484 19404 15876 19460
rect 15260 18956 15652 19012
rect 15148 18452 15204 18462
rect 15148 18358 15204 18396
rect 15596 18450 15652 18956
rect 15596 18398 15598 18450
rect 15650 18398 15652 18450
rect 15596 18386 15652 18398
rect 15820 18676 15876 19404
rect 16268 19122 16324 20076
rect 16268 19070 16270 19122
rect 16322 19070 16324 19122
rect 16268 19058 16324 19070
rect 15260 18338 15316 18350
rect 15260 18286 15262 18338
rect 15314 18286 15316 18338
rect 15036 18228 15092 18238
rect 15036 17666 15092 18172
rect 15260 17890 15316 18286
rect 15260 17838 15262 17890
rect 15314 17838 15316 17890
rect 15260 17826 15316 17838
rect 15036 17614 15038 17666
rect 15090 17614 15092 17666
rect 15036 17602 15092 17614
rect 14924 17378 14980 17388
rect 14700 17108 14756 17118
rect 14700 17014 14756 17052
rect 15036 16994 15092 17006
rect 15036 16942 15038 16994
rect 15090 16942 15092 16994
rect 14924 16884 14980 16894
rect 15036 16884 15092 16942
rect 14980 16828 15092 16884
rect 15372 16994 15428 17006
rect 15372 16942 15374 16994
rect 15426 16942 15428 16994
rect 14924 16818 14980 16828
rect 15148 16324 15204 16334
rect 15372 16324 15428 16942
rect 15708 16324 15764 16334
rect 15372 16322 15764 16324
rect 15372 16270 15710 16322
rect 15762 16270 15764 16322
rect 15372 16268 15764 16270
rect 14812 16212 14868 16222
rect 14812 16118 14868 16156
rect 14588 16006 14644 16044
rect 14476 15894 14532 15932
rect 15148 15316 15204 16268
rect 15708 16258 15764 16268
rect 15820 16100 15876 18620
rect 15932 19010 15988 19022
rect 15932 18958 15934 19010
rect 15986 18958 15988 19010
rect 15932 18340 15988 18958
rect 16716 18562 16772 18574
rect 16716 18510 16718 18562
rect 16770 18510 16772 18562
rect 15932 17220 15988 18284
rect 16268 18452 16324 18462
rect 16268 17890 16324 18396
rect 16268 17838 16270 17890
rect 16322 17838 16324 17890
rect 16268 17826 16324 17838
rect 16604 18450 16660 18462
rect 16604 18398 16606 18450
rect 16658 18398 16660 18450
rect 15932 17154 15988 17164
rect 16268 17668 16324 17678
rect 16268 17442 16324 17612
rect 16268 17390 16270 17442
rect 16322 17390 16324 17442
rect 16268 17108 16324 17390
rect 16268 17042 16324 17052
rect 16380 17556 16436 17566
rect 16604 17556 16660 18398
rect 16716 18340 16772 18510
rect 16828 18564 16884 20638
rect 16940 20578 16996 20590
rect 17500 20580 17556 20590
rect 17836 20580 17892 23100
rect 17948 23090 18004 23100
rect 16940 20526 16942 20578
rect 16994 20526 16996 20578
rect 16940 20132 16996 20526
rect 16940 20066 16996 20076
rect 17388 20578 17892 20580
rect 17388 20526 17502 20578
rect 17554 20526 17892 20578
rect 17388 20524 17892 20526
rect 17948 22148 18004 22158
rect 17948 20804 18004 22092
rect 17276 20020 17332 20030
rect 17388 20020 17444 20524
rect 17500 20514 17556 20524
rect 17500 20130 17556 20142
rect 17500 20078 17502 20130
rect 17554 20078 17556 20130
rect 17500 20020 17556 20078
rect 17332 19964 17556 20020
rect 17612 20020 17668 20030
rect 17276 19954 17332 19964
rect 17500 19794 17556 19806
rect 17500 19742 17502 19794
rect 17554 19742 17556 19794
rect 16940 19234 16996 19246
rect 16940 19182 16942 19234
rect 16994 19182 16996 19234
rect 16940 18674 16996 19182
rect 17500 19234 17556 19742
rect 17500 19182 17502 19234
rect 17554 19182 17556 19234
rect 17500 19170 17556 19182
rect 17612 18900 17668 19964
rect 17612 18834 17668 18844
rect 16940 18622 16942 18674
rect 16994 18622 16996 18674
rect 16940 18610 16996 18622
rect 16828 18498 16884 18508
rect 17500 18564 17556 18574
rect 17836 18564 17892 18574
rect 17556 18562 17892 18564
rect 17556 18510 17838 18562
rect 17890 18510 17892 18562
rect 17556 18508 17892 18510
rect 16716 18274 16772 18284
rect 16380 17554 16660 17556
rect 16380 17502 16382 17554
rect 16434 17502 16660 17554
rect 16380 17500 16660 17502
rect 16044 16770 16100 16782
rect 16044 16718 16046 16770
rect 16098 16718 16100 16770
rect 16044 16324 16100 16718
rect 16268 16660 16324 16670
rect 16268 16566 16324 16604
rect 16044 16258 16100 16268
rect 16268 16324 16324 16334
rect 16380 16324 16436 17500
rect 16492 16658 16548 16670
rect 16492 16606 16494 16658
rect 16546 16606 16548 16658
rect 16492 16548 16548 16606
rect 16716 16660 16772 16670
rect 16940 16660 16996 16670
rect 16772 16604 16884 16660
rect 16716 16594 16772 16604
rect 16492 16482 16548 16492
rect 16268 16322 16436 16324
rect 16268 16270 16270 16322
rect 16322 16270 16436 16322
rect 16268 16268 16436 16270
rect 16268 16258 16324 16268
rect 15820 16044 16100 16100
rect 15148 15222 15204 15260
rect 15260 15986 15316 15998
rect 15260 15934 15262 15986
rect 15314 15934 15316 15986
rect 14700 15202 14756 15214
rect 14700 15150 14702 15202
rect 14754 15150 14756 15202
rect 14252 15092 14420 15148
rect 14140 13748 14196 13758
rect 14140 13654 14196 13692
rect 14364 13300 14420 15092
rect 14700 14532 14756 15150
rect 15260 14532 15316 15934
rect 14700 14438 14756 14476
rect 15036 14476 15316 14532
rect 15372 15874 15428 15886
rect 15372 15822 15374 15874
rect 15426 15822 15428 15874
rect 14476 14420 14532 14430
rect 14476 13524 14532 14364
rect 14476 13430 14532 13468
rect 14588 14418 14644 14430
rect 14588 14366 14590 14418
rect 14642 14366 14644 14418
rect 14364 13244 14532 13300
rect 12348 11564 12740 11620
rect 11900 11454 11902 11506
rect 11954 11454 11956 11506
rect 11900 11442 11956 11454
rect 12572 11396 12628 11406
rect 12684 11396 12740 11564
rect 13580 11554 13636 11564
rect 13692 12572 14084 12628
rect 12796 11396 12852 11406
rect 12684 11394 12852 11396
rect 12684 11342 12798 11394
rect 12850 11342 12852 11394
rect 12684 11340 12852 11342
rect 12572 11302 12628 11340
rect 12460 11172 12516 11182
rect 11564 10780 11844 10836
rect 11788 10050 11844 10780
rect 12460 10612 12516 11116
rect 12796 10948 12852 11340
rect 13692 11172 13748 12572
rect 13804 12404 13860 12414
rect 13804 12310 13860 12348
rect 13916 12180 13972 12190
rect 14364 12180 14420 12190
rect 13916 12086 13972 12124
rect 14140 12178 14420 12180
rect 14140 12126 14366 12178
rect 14418 12126 14420 12178
rect 14140 12124 14420 12126
rect 13804 11956 13860 11966
rect 14140 11956 14196 12124
rect 14364 12114 14420 12124
rect 13804 11954 14196 11956
rect 13804 11902 13806 11954
rect 13858 11902 14196 11954
rect 13804 11900 14196 11902
rect 14252 11954 14308 11966
rect 14252 11902 14254 11954
rect 14306 11902 14308 11954
rect 13804 11890 13860 11900
rect 14252 11620 14308 11902
rect 12796 10882 12852 10892
rect 13580 11116 13748 11172
rect 13916 11564 14308 11620
rect 14476 11618 14532 13244
rect 14588 12964 14644 14366
rect 14588 12898 14644 12908
rect 14812 13746 14868 13758
rect 14812 13694 14814 13746
rect 14866 13694 14868 13746
rect 14700 12740 14756 12750
rect 14700 12646 14756 12684
rect 14812 12404 14868 13694
rect 15036 13748 15092 14476
rect 15372 14420 15428 15822
rect 15596 15876 15652 15886
rect 15596 15874 15764 15876
rect 15596 15822 15598 15874
rect 15650 15822 15764 15874
rect 15596 15820 15764 15822
rect 15596 15810 15652 15820
rect 15596 15428 15652 15438
rect 15596 15334 15652 15372
rect 15484 15314 15540 15326
rect 15484 15262 15486 15314
rect 15538 15262 15540 15314
rect 15484 15148 15540 15262
rect 15484 15092 15652 15148
rect 15372 14354 15428 14364
rect 15484 14644 15540 14654
rect 15148 14306 15204 14318
rect 15148 14254 15150 14306
rect 15202 14254 15204 14306
rect 15148 14196 15204 14254
rect 15372 14196 15428 14206
rect 15148 14140 15372 14196
rect 15372 14130 15428 14140
rect 15148 13972 15204 13982
rect 15484 13972 15540 14588
rect 15148 13970 15540 13972
rect 15148 13918 15150 13970
rect 15202 13918 15540 13970
rect 15148 13916 15540 13918
rect 15148 13906 15204 13916
rect 15596 13860 15652 15092
rect 15708 14642 15764 15820
rect 15932 15874 15988 15886
rect 15932 15822 15934 15874
rect 15986 15822 15988 15874
rect 15932 15428 15988 15822
rect 15932 15362 15988 15372
rect 15708 14590 15710 14642
rect 15762 14590 15764 14642
rect 15708 14578 15764 14590
rect 15820 15314 15876 15326
rect 15820 15262 15822 15314
rect 15874 15262 15876 15314
rect 15820 14420 15876 15262
rect 16044 14644 16100 16044
rect 16156 15540 16212 15550
rect 16156 15446 16212 15484
rect 16044 14578 16100 14588
rect 16156 14420 16212 14430
rect 15820 14418 16212 14420
rect 15820 14366 16158 14418
rect 16210 14366 16212 14418
rect 15820 14364 16212 14366
rect 15484 13804 15596 13860
rect 15036 13692 15204 13748
rect 15148 12404 15204 13692
rect 15260 13076 15316 13086
rect 15484 13076 15540 13804
rect 15596 13766 15652 13804
rect 15708 14196 15764 14206
rect 15708 13746 15764 14140
rect 15708 13694 15710 13746
rect 15762 13694 15764 13746
rect 15708 13682 15764 13694
rect 16156 13746 16212 14364
rect 16156 13694 16158 13746
rect 16210 13694 16212 13746
rect 16156 13682 16212 13694
rect 16380 13636 16436 16268
rect 16716 16212 16772 16222
rect 16716 16098 16772 16156
rect 16716 16046 16718 16098
rect 16770 16046 16772 16098
rect 16716 15764 16772 16046
rect 16492 15708 16772 15764
rect 16828 16210 16884 16604
rect 16940 16566 16996 16604
rect 16828 16158 16830 16210
rect 16882 16158 16884 16210
rect 16492 15314 16548 15708
rect 16716 15316 16772 15326
rect 16828 15316 16884 16158
rect 16492 15262 16494 15314
rect 16546 15262 16548 15314
rect 16492 15250 16548 15262
rect 16604 15314 16884 15316
rect 16604 15262 16718 15314
rect 16770 15262 16884 15314
rect 16604 15260 16884 15262
rect 16604 13746 16660 15260
rect 16716 15250 16772 15260
rect 17388 14532 17444 14542
rect 16604 13694 16606 13746
rect 16658 13694 16660 13746
rect 16604 13636 16660 13694
rect 16940 13748 16996 13758
rect 16940 13654 16996 13692
rect 16604 13580 16884 13636
rect 16380 13570 16436 13580
rect 15260 13074 15540 13076
rect 15260 13022 15262 13074
rect 15314 13022 15540 13074
rect 15260 13020 15540 13022
rect 15708 13524 15764 13534
rect 15260 13010 15316 13020
rect 15596 12964 15652 12974
rect 15596 12850 15652 12908
rect 15708 12962 15764 13468
rect 16828 13074 16884 13580
rect 16828 13022 16830 13074
rect 16882 13022 16884 13074
rect 16828 13010 16884 13022
rect 15708 12910 15710 12962
rect 15762 12910 15764 12962
rect 15708 12898 15764 12910
rect 17388 12962 17444 14476
rect 17388 12910 17390 12962
rect 17442 12910 17444 12962
rect 17388 12898 17444 12910
rect 15596 12798 15598 12850
rect 15650 12798 15652 12850
rect 15596 12516 15652 12798
rect 15596 12460 15876 12516
rect 15372 12404 15428 12414
rect 15148 12348 15372 12404
rect 14812 12338 14868 12348
rect 15372 12310 15428 12348
rect 14476 11566 14478 11618
rect 14530 11566 14532 11618
rect 13916 11396 13972 11564
rect 14476 11554 14532 11566
rect 14588 12180 14644 12190
rect 14364 11506 14420 11518
rect 14364 11454 14366 11506
rect 14418 11454 14420 11506
rect 12348 10610 12516 10612
rect 12348 10558 12462 10610
rect 12514 10558 12516 10610
rect 12348 10556 12516 10558
rect 11788 9998 11790 10050
rect 11842 9998 11844 10050
rect 11788 9986 11844 9998
rect 11900 10498 11956 10510
rect 11900 10446 11902 10498
rect 11954 10446 11956 10498
rect 11452 9202 11508 9212
rect 11340 9154 11396 9166
rect 11340 9102 11342 9154
rect 11394 9102 11396 9154
rect 11340 8148 11396 9102
rect 11900 8930 11956 10446
rect 12236 10388 12292 10398
rect 12124 10052 12180 10062
rect 12124 9958 12180 9996
rect 12236 9154 12292 10332
rect 12348 9938 12404 10556
rect 12460 10546 12516 10556
rect 12348 9886 12350 9938
rect 12402 9886 12404 9938
rect 12348 9874 12404 9886
rect 13580 9380 13636 11116
rect 13692 10948 13748 10958
rect 13692 10388 13748 10892
rect 13916 10834 13972 11340
rect 13916 10782 13918 10834
rect 13970 10782 13972 10834
rect 13692 10386 13860 10388
rect 13692 10334 13694 10386
rect 13746 10334 13860 10386
rect 13692 10332 13860 10334
rect 13692 10322 13748 10332
rect 13804 9826 13860 10332
rect 13804 9774 13806 9826
rect 13858 9774 13860 9826
rect 13804 9762 13860 9774
rect 13916 9828 13972 10782
rect 14028 11394 14084 11406
rect 14028 11342 14030 11394
rect 14082 11342 14084 11394
rect 14028 10498 14084 11342
rect 14028 10446 14030 10498
rect 14082 10446 14084 10498
rect 14028 10434 14084 10446
rect 14364 9940 14420 11454
rect 14476 11172 14532 11182
rect 14476 10834 14532 11116
rect 14476 10782 14478 10834
rect 14530 10782 14532 10834
rect 14476 10770 14532 10782
rect 14588 10610 14644 12124
rect 15820 12066 15876 12460
rect 16268 12404 16324 12414
rect 16324 12348 16436 12404
rect 16268 12338 16324 12348
rect 16380 12290 16436 12348
rect 16380 12238 16382 12290
rect 16434 12238 16436 12290
rect 16380 12226 16436 12238
rect 15820 12014 15822 12066
rect 15874 12014 15876 12066
rect 15820 11956 15876 12014
rect 15820 11890 15876 11900
rect 16268 12178 16324 12190
rect 16268 12126 16270 12178
rect 16322 12126 16324 12178
rect 15932 11508 15988 11518
rect 15932 11414 15988 11452
rect 15484 11396 15540 11406
rect 15484 11302 15540 11340
rect 15708 11394 15764 11406
rect 15708 11342 15710 11394
rect 15762 11342 15764 11394
rect 14588 10558 14590 10610
rect 14642 10558 14644 10610
rect 14476 10388 14532 10398
rect 14476 10294 14532 10332
rect 14588 10052 14644 10558
rect 14924 10498 14980 10510
rect 14924 10446 14926 10498
rect 14978 10446 14980 10498
rect 14924 10388 14980 10446
rect 14924 10322 14980 10332
rect 15036 10386 15092 10398
rect 15036 10334 15038 10386
rect 15090 10334 15092 10386
rect 14140 9938 14420 9940
rect 14140 9886 14366 9938
rect 14418 9886 14420 9938
rect 14140 9884 14420 9886
rect 14028 9828 14084 9838
rect 13916 9826 14084 9828
rect 13916 9774 14030 9826
rect 14082 9774 14084 9826
rect 13916 9772 14084 9774
rect 14028 9762 14084 9772
rect 13580 9314 13636 9324
rect 12236 9102 12238 9154
rect 12290 9102 12292 9154
rect 12236 9090 12292 9102
rect 13916 9156 13972 9166
rect 14140 9156 14196 9884
rect 14364 9874 14420 9884
rect 14476 9996 14588 10052
rect 14476 9716 14532 9996
rect 14588 9986 14644 9996
rect 15036 9938 15092 10334
rect 15708 10388 15764 11342
rect 16156 10388 16212 10398
rect 16268 10388 16324 12126
rect 16492 12178 16548 12190
rect 16492 12126 16494 12178
rect 16546 12126 16548 12178
rect 16380 11620 16436 11630
rect 16380 11526 16436 11564
rect 16492 11396 16548 12126
rect 16940 12178 16996 12190
rect 16940 12126 16942 12178
rect 16994 12126 16996 12178
rect 16380 10836 16436 10846
rect 16492 10836 16548 11340
rect 16828 11956 16884 11966
rect 16828 11282 16884 11900
rect 16828 11230 16830 11282
rect 16882 11230 16884 11282
rect 16828 11218 16884 11230
rect 16940 11508 16996 12126
rect 17500 11788 17556 18508
rect 17836 18498 17892 18508
rect 17948 18562 18004 20748
rect 18060 20132 18116 23214
rect 18284 23154 18340 23166
rect 18284 23102 18286 23154
rect 18338 23102 18340 23154
rect 18172 22370 18228 22382
rect 18172 22318 18174 22370
rect 18226 22318 18228 22370
rect 18172 22260 18228 22318
rect 18284 22372 18340 23102
rect 18508 23044 18564 23054
rect 18508 22950 18564 22988
rect 18620 22932 18676 22942
rect 18620 22838 18676 22876
rect 19068 22482 19124 23884
rect 19068 22430 19070 22482
rect 19122 22430 19124 22482
rect 19068 22418 19124 22430
rect 19180 23154 19236 23166
rect 19180 23102 19182 23154
rect 19234 23102 19236 23154
rect 18396 22372 18452 22382
rect 18284 22370 18452 22372
rect 18284 22318 18398 22370
rect 18450 22318 18452 22370
rect 18284 22316 18452 22318
rect 18396 22306 18452 22316
rect 18172 22194 18228 22204
rect 18732 21924 18788 21934
rect 18508 20804 18564 20814
rect 18508 20802 18676 20804
rect 18508 20750 18510 20802
rect 18562 20750 18676 20802
rect 18508 20748 18676 20750
rect 18508 20738 18564 20748
rect 18060 20066 18116 20076
rect 18172 19234 18228 19246
rect 18172 19182 18174 19234
rect 18226 19182 18228 19234
rect 18172 18674 18228 19182
rect 18172 18622 18174 18674
rect 18226 18622 18228 18674
rect 18172 18610 18228 18622
rect 18508 19012 18564 19022
rect 17948 18510 17950 18562
rect 18002 18510 18004 18562
rect 17948 17668 18004 18510
rect 18508 18562 18564 18956
rect 18620 18676 18676 20748
rect 18732 20580 18788 21868
rect 19180 21812 19236 23102
rect 19292 22932 19348 24444
rect 19292 22838 19348 22876
rect 19180 21756 19348 21812
rect 19180 21586 19236 21598
rect 19180 21534 19182 21586
rect 19234 21534 19236 21586
rect 19180 21026 19236 21534
rect 19180 20974 19182 21026
rect 19234 20974 19236 21026
rect 19180 20962 19236 20974
rect 18732 20486 18788 20524
rect 19068 20690 19124 20702
rect 19068 20638 19070 20690
rect 19122 20638 19124 20690
rect 19068 20020 19124 20638
rect 19180 20580 19236 20590
rect 19180 20486 19236 20524
rect 19068 19954 19124 19964
rect 19292 19346 19348 21756
rect 19516 21698 19572 24892
rect 19628 23940 19684 25228
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 20300 24836 20356 24846
rect 20300 24742 20356 24780
rect 19852 24724 19908 24734
rect 19852 24630 19908 24668
rect 19740 23940 19796 23950
rect 19628 23884 19740 23940
rect 19740 23874 19796 23884
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 20412 23268 20468 25230
rect 20524 24834 20580 24846
rect 20524 24782 20526 24834
rect 20578 24782 20580 24834
rect 20524 24052 20580 24782
rect 20636 24836 20692 24846
rect 20636 24742 20692 24780
rect 21084 24836 21140 24846
rect 21084 24742 21140 24780
rect 22652 24834 22708 25340
rect 23212 24948 23268 25900
rect 22876 24946 23268 24948
rect 22876 24894 23214 24946
rect 23266 24894 23268 24946
rect 22876 24892 23268 24894
rect 22652 24782 22654 24834
rect 22706 24782 22708 24834
rect 22652 24770 22708 24782
rect 22764 24834 22820 24846
rect 22764 24782 22766 24834
rect 22818 24782 22820 24834
rect 21532 24724 21588 24734
rect 21308 24388 21364 24398
rect 20636 24052 20692 24062
rect 20524 23996 20636 24052
rect 20636 23958 20692 23996
rect 21308 24050 21364 24332
rect 21308 23998 21310 24050
rect 21362 23998 21364 24050
rect 21308 23828 21364 23998
rect 21308 23762 21364 23772
rect 21532 23604 21588 24668
rect 22764 24164 22820 24782
rect 22764 24098 22820 24108
rect 21532 23538 21588 23548
rect 22204 23324 22820 23380
rect 20412 23202 20468 23212
rect 21644 23266 21700 23278
rect 21644 23214 21646 23266
rect 21698 23214 21700 23266
rect 21532 23156 21588 23166
rect 21420 23154 21588 23156
rect 21420 23102 21534 23154
rect 21586 23102 21588 23154
rect 21420 23100 21588 23102
rect 21420 22372 21476 23100
rect 21532 23090 21588 23100
rect 21308 22370 21476 22372
rect 21308 22318 21422 22370
rect 21474 22318 21476 22370
rect 21308 22316 21476 22318
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 19516 21646 19518 21698
rect 19570 21646 19572 21698
rect 19516 21634 19572 21646
rect 20748 21700 20804 21710
rect 20748 21606 20804 21644
rect 21308 21586 21364 22316
rect 21420 22306 21476 22316
rect 21644 22370 21700 23214
rect 22204 23042 22260 23324
rect 22204 22990 22206 23042
rect 22258 22990 22260 23042
rect 21644 22318 21646 22370
rect 21698 22318 21700 22370
rect 21644 21700 21700 22318
rect 21644 21634 21700 21644
rect 22092 22594 22148 22606
rect 22092 22542 22094 22594
rect 22146 22542 22148 22594
rect 21308 21534 21310 21586
rect 21362 21534 21364 21586
rect 21308 21140 21364 21534
rect 21308 21084 21700 21140
rect 21420 20916 21476 20926
rect 19740 20692 19796 20702
rect 19292 19294 19294 19346
rect 19346 19294 19348 19346
rect 19292 19282 19348 19294
rect 19628 20636 19740 20692
rect 18732 19236 18788 19246
rect 18732 19122 18788 19180
rect 19404 19236 19460 19274
rect 19404 19170 19460 19180
rect 19180 19124 19236 19134
rect 18732 19070 18734 19122
rect 18786 19070 18788 19122
rect 18732 19058 18788 19070
rect 18844 19068 19180 19124
rect 18620 18582 18676 18620
rect 18844 18674 18900 19068
rect 19180 19058 19236 19068
rect 19404 19012 19460 19022
rect 18844 18622 18846 18674
rect 18898 18622 18900 18674
rect 18844 18610 18900 18622
rect 19180 18676 19236 18686
rect 19180 18582 19236 18620
rect 19404 18674 19460 18956
rect 19404 18622 19406 18674
rect 19458 18622 19460 18674
rect 19404 18610 19460 18622
rect 19628 18676 19684 20636
rect 19740 20626 19796 20636
rect 21196 20692 21252 20702
rect 21420 20692 21476 20860
rect 21196 20598 21252 20636
rect 21308 20690 21476 20692
rect 21308 20638 21422 20690
rect 21474 20638 21476 20690
rect 21308 20636 21476 20638
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 20412 20130 20468 20142
rect 20412 20078 20414 20130
rect 20466 20078 20468 20130
rect 20188 20018 20244 20030
rect 20188 19966 20190 20018
rect 20242 19966 20244 20018
rect 19740 19234 19796 19246
rect 19740 19182 19742 19234
rect 19794 19182 19796 19234
rect 19740 19124 19796 19182
rect 19740 19058 19796 19068
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19964 18676 20020 18686
rect 20188 18676 20244 19966
rect 19628 18620 19908 18676
rect 18508 18510 18510 18562
rect 18562 18510 18564 18562
rect 18508 18498 18564 18510
rect 19516 18564 19572 18574
rect 19516 18562 19684 18564
rect 19516 18510 19518 18562
rect 19570 18510 19684 18562
rect 19516 18508 19684 18510
rect 19516 18498 19572 18508
rect 18620 17668 18676 17678
rect 17948 17602 18004 17612
rect 18060 17666 18676 17668
rect 18060 17614 18622 17666
rect 18674 17614 18676 17666
rect 18060 17612 18676 17614
rect 17836 17444 17892 17454
rect 17612 16996 17668 17006
rect 17612 16322 17668 16940
rect 17724 16994 17780 17006
rect 17724 16942 17726 16994
rect 17778 16942 17780 16994
rect 17724 16884 17780 16942
rect 17836 16994 17892 17388
rect 17836 16942 17838 16994
rect 17890 16942 17892 16994
rect 17836 16930 17892 16942
rect 18060 17108 18116 17612
rect 18620 17602 18676 17612
rect 18844 17666 18900 17678
rect 18844 17614 18846 17666
rect 18898 17614 18900 17666
rect 18284 17444 18340 17454
rect 18284 17442 18564 17444
rect 18284 17390 18286 17442
rect 18338 17390 18564 17442
rect 18284 17388 18564 17390
rect 18284 17378 18340 17388
rect 17724 16818 17780 16828
rect 17612 16270 17614 16322
rect 17666 16270 17668 16322
rect 17612 15426 17668 16270
rect 17612 15374 17614 15426
rect 17666 15374 17668 15426
rect 17612 15362 17668 15374
rect 17724 16658 17780 16670
rect 17724 16606 17726 16658
rect 17778 16606 17780 16658
rect 17724 16548 17780 16606
rect 17724 16098 17780 16492
rect 17724 16046 17726 16098
rect 17778 16046 17780 16098
rect 17724 15204 17780 16046
rect 17836 16660 17892 16670
rect 17836 15314 17892 16604
rect 17836 15262 17838 15314
rect 17890 15262 17892 15314
rect 17836 15250 17892 15262
rect 17724 15138 17780 15148
rect 18060 13860 18116 17052
rect 18508 16994 18564 17388
rect 18508 16942 18510 16994
rect 18562 16942 18564 16994
rect 18284 16882 18340 16894
rect 18284 16830 18286 16882
rect 18338 16830 18340 16882
rect 18172 16770 18228 16782
rect 18172 16718 18174 16770
rect 18226 16718 18228 16770
rect 18172 16098 18228 16718
rect 18284 16660 18340 16830
rect 18284 16594 18340 16604
rect 18172 16046 18174 16098
rect 18226 16046 18228 16098
rect 18172 16034 18228 16046
rect 18396 16100 18452 16110
rect 18396 15538 18452 16044
rect 18396 15486 18398 15538
rect 18450 15486 18452 15538
rect 18396 15474 18452 15486
rect 18060 13746 18116 13804
rect 18060 13694 18062 13746
rect 18114 13694 18116 13746
rect 18060 13682 18116 13694
rect 18284 15316 18340 15326
rect 18284 13636 18340 15260
rect 18508 15316 18564 16942
rect 18844 16436 18900 17614
rect 19516 17666 19572 17678
rect 19516 17614 19518 17666
rect 19570 17614 19572 17666
rect 19068 16996 19124 17006
rect 19068 16902 19124 16940
rect 19516 16884 19572 17614
rect 19628 17556 19684 18508
rect 19852 18562 19908 18620
rect 19964 18674 20244 18676
rect 19964 18622 19966 18674
rect 20018 18622 20244 18674
rect 19964 18620 20244 18622
rect 20412 19236 20468 20078
rect 20524 20018 20580 20030
rect 20524 19966 20526 20018
rect 20578 19966 20580 20018
rect 20524 19348 20580 19966
rect 21308 20018 21364 20636
rect 21420 20626 21476 20636
rect 21532 20690 21588 20702
rect 21532 20638 21534 20690
rect 21586 20638 21588 20690
rect 21308 19966 21310 20018
rect 21362 19966 21364 20018
rect 21308 19954 21364 19966
rect 21532 19908 21588 20638
rect 21644 20468 21700 21084
rect 22092 20804 22148 22542
rect 22092 20738 22148 20748
rect 22204 20690 22260 22990
rect 22428 23156 22484 23166
rect 22428 21698 22484 23100
rect 22764 23154 22820 23324
rect 22764 23102 22766 23154
rect 22818 23102 22820 23154
rect 22764 23090 22820 23102
rect 22540 23044 22596 23054
rect 22540 21810 22596 22988
rect 22652 23042 22708 23054
rect 22652 22990 22654 23042
rect 22706 22990 22708 23042
rect 22652 22596 22708 22990
rect 22764 22596 22820 22606
rect 22652 22540 22764 22596
rect 22764 22530 22820 22540
rect 22876 22484 22932 24892
rect 23212 24882 23268 24892
rect 23324 24948 23380 24958
rect 23436 24948 23492 26236
rect 23548 26226 23604 26236
rect 24108 26290 24164 26572
rect 24108 26238 24110 26290
rect 24162 26238 24164 26290
rect 24108 26226 24164 26238
rect 23660 26180 23716 26190
rect 23660 26086 23716 26124
rect 23324 24946 23492 24948
rect 23324 24894 23326 24946
rect 23378 24894 23492 24946
rect 23324 24892 23492 24894
rect 23548 25172 23604 25182
rect 23324 24882 23380 24892
rect 22988 24724 23044 24734
rect 23436 24724 23492 24734
rect 23548 24724 23604 25116
rect 22988 24722 23156 24724
rect 22988 24670 22990 24722
rect 23042 24670 23156 24722
rect 22988 24668 23156 24670
rect 22988 24658 23044 24668
rect 23100 24164 23156 24668
rect 23436 24722 23604 24724
rect 23436 24670 23438 24722
rect 23490 24670 23604 24722
rect 23436 24668 23604 24670
rect 23772 24948 23828 24958
rect 23772 24722 23828 24892
rect 24220 24948 24276 24958
rect 24220 24854 24276 24892
rect 23772 24670 23774 24722
rect 23826 24670 23828 24722
rect 23436 24658 23492 24668
rect 23772 24658 23828 24670
rect 24332 24836 24388 26908
rect 24444 25172 24500 25182
rect 24444 24946 24500 25116
rect 24444 24894 24446 24946
rect 24498 24894 24500 24946
rect 24444 24882 24500 24894
rect 24556 24946 24612 27804
rect 25228 27794 25284 27804
rect 25004 26962 25060 26974
rect 25004 26910 25006 26962
rect 25058 26910 25060 26962
rect 25004 25732 25060 26910
rect 26236 26908 26292 30604
rect 26684 30436 26740 30830
rect 26348 30380 26740 30436
rect 26348 30098 26404 30380
rect 26796 30324 26852 45052
rect 27132 43708 27188 45836
rect 27244 44996 27300 47068
rect 27580 47010 27636 47022
rect 27580 46958 27582 47010
rect 27634 46958 27636 47010
rect 27580 46004 27636 46958
rect 28252 47010 28308 49200
rect 28252 46958 28254 47010
rect 28306 46958 28308 47010
rect 28252 46946 28308 46958
rect 27580 45890 27636 45948
rect 27580 45838 27582 45890
rect 27634 45838 27636 45890
rect 27580 45826 27636 45838
rect 28364 45892 28420 45902
rect 28364 45798 28420 45836
rect 27804 45666 27860 45678
rect 27804 45614 27806 45666
rect 27858 45614 27860 45666
rect 27356 44996 27412 45006
rect 27244 44994 27412 44996
rect 27244 44942 27358 44994
rect 27410 44942 27412 44994
rect 27244 44940 27412 44942
rect 27356 44930 27412 44940
rect 27132 43652 27300 43708
rect 27020 36372 27076 36382
rect 26908 35028 26964 35038
rect 26908 34914 26964 34972
rect 26908 34862 26910 34914
rect 26962 34862 26964 34914
rect 26908 34850 26964 34862
rect 26908 32676 26964 32686
rect 26908 32582 26964 32620
rect 26908 31108 26964 31118
rect 26908 30994 26964 31052
rect 26908 30942 26910 30994
rect 26962 30942 26964 30994
rect 26908 30930 26964 30942
rect 26348 30046 26350 30098
rect 26402 30046 26404 30098
rect 26348 30034 26404 30046
rect 26684 30268 26852 30324
rect 26684 28308 26740 30268
rect 27020 30210 27076 36316
rect 27020 30158 27022 30210
rect 27074 30158 27076 30210
rect 27020 30146 27076 30158
rect 27132 31556 27188 31566
rect 26908 30098 26964 30110
rect 26908 30046 26910 30098
rect 26962 30046 26964 30098
rect 26796 29538 26852 29550
rect 26796 29486 26798 29538
rect 26850 29486 26852 29538
rect 26796 29204 26852 29486
rect 26796 29138 26852 29148
rect 26908 29092 26964 30046
rect 27132 29650 27188 31500
rect 27132 29598 27134 29650
rect 27186 29598 27188 29650
rect 27132 29586 27188 29598
rect 26908 29026 26964 29036
rect 27244 28868 27300 43652
rect 27804 38668 27860 45614
rect 28700 44436 28756 44446
rect 28924 44436 28980 49200
rect 29596 46228 29652 49200
rect 30268 46674 30324 49200
rect 30268 46622 30270 46674
rect 30322 46622 30324 46674
rect 30268 46610 30324 46622
rect 31052 46674 31108 46686
rect 31052 46622 31054 46674
rect 31106 46622 31108 46674
rect 29596 46172 30100 46228
rect 29372 46116 29428 46126
rect 29372 46022 29428 46060
rect 30044 45330 30100 46172
rect 30044 45278 30046 45330
rect 30098 45278 30100 45330
rect 29260 45108 29316 45118
rect 29260 45014 29316 45052
rect 28700 44434 29428 44436
rect 28700 44382 28702 44434
rect 28754 44382 29428 44434
rect 28700 44380 29428 44382
rect 28700 44370 28756 44380
rect 29372 44322 29428 44380
rect 30044 44434 30100 45278
rect 31052 45330 31108 46622
rect 31500 46674 31556 46686
rect 31500 46622 31502 46674
rect 31554 46622 31556 46674
rect 31500 45890 31556 46622
rect 31500 45838 31502 45890
rect 31554 45838 31556 45890
rect 31500 45826 31556 45838
rect 31052 45278 31054 45330
rect 31106 45278 31108 45330
rect 31052 45266 31108 45278
rect 31276 45666 31332 45678
rect 31276 45614 31278 45666
rect 31330 45614 31332 45666
rect 30380 45220 30436 45230
rect 30044 44382 30046 44434
rect 30098 44382 30100 44434
rect 30044 44370 30100 44382
rect 30268 45218 30436 45220
rect 30268 45166 30382 45218
rect 30434 45166 30436 45218
rect 30268 45164 30436 45166
rect 29372 44270 29374 44322
rect 29426 44270 29428 44322
rect 29372 44258 29428 44270
rect 29148 44098 29204 44110
rect 29148 44046 29150 44098
rect 29202 44046 29204 44098
rect 29148 43708 29204 44046
rect 28924 43652 29204 43708
rect 28700 42420 28756 42430
rect 28364 40852 28420 40862
rect 27356 38612 27860 38668
rect 28028 40292 28084 40302
rect 28028 38668 28084 40236
rect 28364 40068 28420 40796
rect 28476 40628 28532 40638
rect 28700 40628 28756 42364
rect 28476 40626 28756 40628
rect 28476 40574 28478 40626
rect 28530 40574 28756 40626
rect 28476 40572 28756 40574
rect 28476 40562 28532 40572
rect 28700 40514 28756 40572
rect 28700 40462 28702 40514
rect 28754 40462 28756 40514
rect 28700 40180 28756 40462
rect 28812 40514 28868 40526
rect 28812 40462 28814 40514
rect 28866 40462 28868 40514
rect 28812 40292 28868 40462
rect 28812 40226 28868 40236
rect 28700 40114 28756 40124
rect 28364 40012 28532 40068
rect 28364 39506 28420 39518
rect 28364 39454 28366 39506
rect 28418 39454 28420 39506
rect 28140 39396 28196 39406
rect 28364 39396 28420 39454
rect 28476 39506 28532 40012
rect 28700 39620 28756 39630
rect 28700 39526 28756 39564
rect 28476 39454 28478 39506
rect 28530 39454 28532 39506
rect 28476 39442 28532 39454
rect 28140 39394 28420 39396
rect 28140 39342 28142 39394
rect 28194 39342 28420 39394
rect 28140 39340 28420 39342
rect 28140 39330 28196 39340
rect 28364 39060 28420 39340
rect 28700 39060 28756 39070
rect 28364 39004 28700 39060
rect 28700 38966 28756 39004
rect 28812 38948 28868 38958
rect 28028 38612 28308 38668
rect 27356 31220 27412 38612
rect 28252 38050 28308 38612
rect 28252 37998 28254 38050
rect 28306 37998 28308 38050
rect 28252 37986 28308 37998
rect 28588 37828 28644 37838
rect 28588 37734 28644 37772
rect 28476 37380 28532 37390
rect 28364 37324 28476 37380
rect 28252 36596 28308 36606
rect 28252 35922 28308 36540
rect 28252 35870 28254 35922
rect 28306 35870 28308 35922
rect 28252 35858 28308 35870
rect 27916 35252 27972 35262
rect 27804 35028 27860 35038
rect 27692 34244 27748 34254
rect 27692 34150 27748 34188
rect 27356 31154 27412 31164
rect 27468 34132 27524 34142
rect 27468 31668 27524 34076
rect 27804 33908 27860 34972
rect 27916 34354 27972 35196
rect 28364 35252 28420 37324
rect 28476 37286 28532 37324
rect 28812 37378 28868 38892
rect 28812 37326 28814 37378
rect 28866 37326 28868 37378
rect 28812 37314 28868 37326
rect 28924 36036 28980 43652
rect 30044 42642 30100 42654
rect 30044 42590 30046 42642
rect 30098 42590 30100 42642
rect 30044 42420 30100 42590
rect 30044 42354 30100 42364
rect 30156 42644 30212 42654
rect 30044 42196 30100 42206
rect 30156 42196 30212 42588
rect 30044 42194 30212 42196
rect 30044 42142 30046 42194
rect 30098 42142 30212 42194
rect 30044 42140 30212 42142
rect 30268 42196 30324 45164
rect 30380 45154 30436 45164
rect 30380 44996 30436 45006
rect 30380 44434 30436 44940
rect 30380 44382 30382 44434
rect 30434 44382 30436 44434
rect 30380 44370 30436 44382
rect 30492 42644 30548 42654
rect 30380 42532 30436 42542
rect 30380 42438 30436 42476
rect 30268 42140 30436 42196
rect 30044 42130 30100 42140
rect 29708 42082 29764 42094
rect 29708 42030 29710 42082
rect 29762 42030 29764 42082
rect 29708 41188 29764 42030
rect 30268 41970 30324 41982
rect 30268 41918 30270 41970
rect 30322 41918 30324 41970
rect 29708 40852 29764 41132
rect 29708 40786 29764 40796
rect 29820 41412 29876 41422
rect 29820 41074 29876 41356
rect 29820 41022 29822 41074
rect 29874 41022 29876 41074
rect 29036 40402 29092 40414
rect 29036 40350 29038 40402
rect 29090 40350 29092 40402
rect 29036 39620 29092 40350
rect 29820 40402 29876 41022
rect 29820 40350 29822 40402
rect 29874 40350 29876 40402
rect 29820 40338 29876 40350
rect 30044 41188 30100 41198
rect 30268 41188 30324 41918
rect 30044 41186 30324 41188
rect 30044 41134 30046 41186
rect 30098 41134 30324 41186
rect 30044 41132 30324 41134
rect 30044 40404 30100 41132
rect 30380 40628 30436 42140
rect 30492 42194 30548 42588
rect 31276 42644 31332 45614
rect 34300 44996 34356 49200
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 35084 46004 35140 46014
rect 35084 45910 35140 45948
rect 36988 46004 37044 49200
rect 37660 47012 37716 49200
rect 37660 46956 38164 47012
rect 36540 45892 36596 45902
rect 36988 45892 37044 45948
rect 37212 45892 37268 45902
rect 36988 45890 37268 45892
rect 36988 45838 37214 45890
rect 37266 45838 37268 45890
rect 36988 45836 37268 45838
rect 36540 45798 36596 45836
rect 37212 45826 37268 45836
rect 38108 45892 38164 46956
rect 38332 46452 38388 49200
rect 38332 46396 38724 46452
rect 38108 45798 38164 45836
rect 38668 45890 38724 46396
rect 38668 45838 38670 45890
rect 38722 45838 38724 45890
rect 35532 45780 35588 45790
rect 35532 45686 35588 45724
rect 36876 45666 36932 45678
rect 36876 45614 36878 45666
rect 36930 45614 36932 45666
rect 36316 45108 36372 45118
rect 34748 44996 34804 45006
rect 34300 44994 34804 44996
rect 34300 44942 34750 44994
rect 34802 44942 34804 44994
rect 34300 44940 34804 44942
rect 34748 44930 34804 44940
rect 36204 44996 36260 45006
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 32508 44434 32564 44446
rect 32508 44382 32510 44434
rect 32562 44382 32564 44434
rect 32172 44210 32228 44222
rect 32172 44158 32174 44210
rect 32226 44158 32228 44210
rect 32172 43092 32228 44158
rect 32172 43026 32228 43036
rect 31948 42756 32004 42766
rect 32508 42756 32564 44382
rect 33516 44322 33572 44334
rect 33516 44270 33518 44322
rect 33570 44270 33572 44322
rect 33516 43428 33572 44270
rect 34076 44322 34132 44334
rect 34076 44270 34078 44322
rect 34130 44270 34132 44322
rect 33628 44210 33684 44222
rect 33628 44158 33630 44210
rect 33682 44158 33684 44210
rect 33628 43708 33684 44158
rect 34076 43988 34132 44270
rect 36204 44322 36260 44940
rect 36316 44546 36372 45052
rect 36316 44494 36318 44546
rect 36370 44494 36372 44546
rect 36316 44482 36372 44494
rect 36652 45108 36708 45118
rect 36876 45108 36932 45614
rect 36652 45106 36932 45108
rect 36652 45054 36654 45106
rect 36706 45054 36932 45106
rect 36652 45052 36932 45054
rect 37212 45668 37268 45678
rect 36204 44270 36206 44322
rect 36258 44270 36260 44322
rect 36204 44258 36260 44270
rect 36316 44212 36372 44222
rect 36316 44118 36372 44156
rect 34076 43932 34692 43988
rect 34636 43708 34692 43932
rect 36652 43708 36708 45052
rect 37212 44434 37268 45612
rect 37548 45666 37604 45678
rect 37884 45668 37940 45678
rect 37548 45614 37550 45666
rect 37602 45614 37604 45666
rect 37212 44382 37214 44434
rect 37266 44382 37268 44434
rect 37212 44370 37268 44382
rect 37436 44994 37492 45006
rect 37436 44942 37438 44994
rect 37490 44942 37492 44994
rect 33628 43652 33796 43708
rect 34412 43652 34468 43662
rect 34636 43652 35028 43708
rect 33516 43362 33572 43372
rect 33628 42980 33684 42990
rect 33516 42924 33628 42980
rect 33516 42866 33572 42924
rect 33628 42914 33684 42924
rect 33516 42814 33518 42866
rect 33570 42814 33572 42866
rect 33516 42802 33572 42814
rect 31948 42754 32564 42756
rect 31948 42702 31950 42754
rect 32002 42702 32564 42754
rect 31948 42700 32564 42702
rect 33628 42754 33684 42766
rect 33628 42702 33630 42754
rect 33682 42702 33684 42754
rect 31276 42578 31332 42588
rect 31724 42644 31780 42654
rect 31724 42550 31780 42588
rect 30716 42530 30772 42542
rect 30716 42478 30718 42530
rect 30770 42478 30772 42530
rect 30716 42420 30772 42478
rect 31948 42532 32004 42700
rect 33292 42644 33348 42654
rect 31948 42466 32004 42476
rect 33180 42588 33292 42644
rect 30716 42354 30772 42364
rect 30492 42142 30494 42194
rect 30546 42142 30548 42194
rect 30492 42130 30548 42142
rect 30604 41970 30660 41982
rect 30604 41918 30606 41970
rect 30658 41918 30660 41970
rect 30604 41860 30660 41918
rect 32508 41972 32564 41982
rect 31052 41860 31108 41870
rect 30604 41858 31108 41860
rect 30604 41806 31054 41858
rect 31106 41806 31108 41858
rect 30604 41804 31108 41806
rect 31052 41300 31108 41804
rect 31052 41234 31108 41244
rect 32508 41412 32564 41916
rect 33180 41970 33236 42588
rect 33292 42578 33348 42588
rect 33404 42532 33460 42542
rect 33404 41972 33460 42476
rect 33628 42420 33684 42702
rect 33628 42354 33684 42364
rect 33180 41918 33182 41970
rect 33234 41918 33236 41970
rect 33180 41906 33236 41918
rect 33292 41970 33460 41972
rect 33292 41918 33406 41970
rect 33458 41918 33460 41970
rect 33292 41916 33460 41918
rect 33292 41636 33348 41916
rect 33404 41906 33460 41916
rect 32172 41188 32228 41198
rect 31164 41074 31220 41086
rect 31164 41022 31166 41074
rect 31218 41022 31220 41074
rect 31164 40740 31220 41022
rect 31164 40674 31220 40684
rect 31276 40962 31332 40974
rect 31276 40910 31278 40962
rect 31330 40910 31332 40962
rect 30268 40572 30436 40628
rect 30156 40404 30212 40414
rect 30044 40402 30212 40404
rect 30044 40350 30158 40402
rect 30210 40350 30212 40402
rect 30044 40348 30212 40350
rect 30156 40338 30212 40348
rect 29484 39730 29540 39742
rect 29484 39678 29486 39730
rect 29538 39678 29540 39730
rect 29372 39620 29428 39630
rect 29036 39618 29428 39620
rect 29036 39566 29374 39618
rect 29426 39566 29428 39618
rect 29036 39564 29428 39566
rect 29372 39554 29428 39564
rect 29484 39620 29540 39678
rect 29484 39554 29540 39564
rect 29932 39172 29988 39182
rect 29372 39060 29428 39070
rect 29036 38946 29092 38958
rect 29036 38894 29038 38946
rect 29090 38894 29092 38946
rect 29036 38668 29092 38894
rect 29372 38946 29428 39004
rect 29372 38894 29374 38946
rect 29426 38894 29428 38946
rect 29372 38882 29428 38894
rect 29820 38948 29876 38958
rect 29820 38854 29876 38892
rect 29932 38946 29988 39116
rect 29932 38894 29934 38946
rect 29986 38894 29988 38946
rect 29932 38882 29988 38894
rect 29036 38612 29204 38668
rect 29148 36036 29204 38612
rect 29820 38610 29876 38622
rect 29820 38558 29822 38610
rect 29874 38558 29876 38610
rect 29596 38162 29652 38174
rect 29596 38110 29598 38162
rect 29650 38110 29652 38162
rect 29372 37492 29428 37502
rect 29260 37380 29316 37390
rect 29260 37286 29316 37324
rect 29372 37378 29428 37436
rect 29596 37490 29652 38110
rect 29820 38050 29876 38558
rect 29820 37998 29822 38050
rect 29874 37998 29876 38050
rect 29820 37986 29876 37998
rect 30156 38162 30212 38174
rect 30156 38110 30158 38162
rect 30210 38110 30212 38162
rect 29708 37828 29764 37838
rect 29764 37772 29876 37828
rect 29708 37762 29764 37772
rect 29596 37438 29598 37490
rect 29650 37438 29652 37490
rect 29596 37426 29652 37438
rect 29820 37490 29876 37772
rect 29820 37438 29822 37490
rect 29874 37438 29876 37490
rect 29372 37326 29374 37378
rect 29426 37326 29428 37378
rect 29372 37314 29428 37326
rect 29260 37042 29316 37054
rect 29260 36990 29262 37042
rect 29314 36990 29316 37042
rect 29260 36484 29316 36990
rect 29484 36596 29540 36606
rect 29484 36502 29540 36540
rect 29372 36484 29428 36494
rect 29260 36482 29428 36484
rect 29260 36430 29374 36482
rect 29426 36430 29428 36482
rect 29260 36428 29428 36430
rect 29372 36418 29428 36428
rect 29820 36036 29876 37438
rect 29932 37492 29988 37502
rect 29932 37378 29988 37436
rect 29932 37326 29934 37378
rect 29986 37326 29988 37378
rect 29932 37314 29988 37326
rect 30044 36708 30100 36718
rect 28924 35980 29092 36036
rect 29148 35980 29428 36036
rect 28476 35924 28532 35934
rect 28476 35922 28756 35924
rect 28476 35870 28478 35922
rect 28530 35870 28756 35922
rect 28476 35868 28756 35870
rect 28476 35858 28532 35868
rect 28700 35812 28756 35868
rect 28924 35812 28980 35822
rect 28700 35810 28980 35812
rect 28700 35758 28926 35810
rect 28978 35758 28980 35810
rect 28700 35756 28980 35758
rect 28588 35700 28644 35710
rect 28588 35606 28644 35644
rect 28364 35186 28420 35196
rect 27916 34302 27918 34354
rect 27970 34302 27972 34354
rect 27916 34290 27972 34302
rect 28476 34692 28532 34702
rect 27804 33852 27972 33908
rect 27804 33570 27860 33582
rect 27804 33518 27806 33570
rect 27858 33518 27860 33570
rect 27580 33236 27636 33246
rect 27580 32562 27636 33180
rect 27580 32510 27582 32562
rect 27634 32510 27636 32562
rect 27580 32498 27636 32510
rect 27692 33234 27748 33246
rect 27692 33182 27694 33234
rect 27746 33182 27748 33234
rect 27692 32004 27748 33182
rect 27804 32004 27860 33518
rect 27916 33234 27972 33852
rect 28028 33906 28084 33918
rect 28028 33854 28030 33906
rect 28082 33854 28084 33906
rect 28028 33348 28084 33854
rect 28140 33906 28196 33918
rect 28140 33854 28142 33906
rect 28194 33854 28196 33906
rect 28140 33572 28196 33854
rect 28252 33572 28308 33582
rect 28140 33570 28308 33572
rect 28140 33518 28254 33570
rect 28306 33518 28308 33570
rect 28140 33516 28308 33518
rect 28252 33506 28308 33516
rect 28476 33570 28532 34636
rect 28924 34580 28980 35756
rect 28812 34356 28868 34366
rect 28812 34242 28868 34300
rect 28812 34190 28814 34242
rect 28866 34190 28868 34242
rect 28812 34178 28868 34190
rect 28924 34244 28980 34524
rect 28924 34150 28980 34188
rect 28588 34132 28644 34142
rect 28588 34038 28644 34076
rect 28476 33518 28478 33570
rect 28530 33518 28532 33570
rect 28476 33506 28532 33518
rect 28028 33292 28308 33348
rect 27916 33182 27918 33234
rect 27970 33182 27972 33234
rect 27916 32228 27972 33182
rect 28252 32676 28308 33292
rect 28364 32676 28420 32686
rect 28252 32674 28420 32676
rect 28252 32622 28366 32674
rect 28418 32622 28420 32674
rect 28252 32620 28420 32622
rect 28364 32610 28420 32620
rect 28588 32562 28644 32574
rect 28588 32510 28590 32562
rect 28642 32510 28644 32562
rect 27916 32172 28420 32228
rect 28140 32004 28196 32014
rect 27804 31948 28084 32004
rect 27692 31938 27748 31948
rect 27804 31778 27860 31790
rect 27804 31726 27806 31778
rect 27858 31726 27860 31778
rect 27804 31668 27860 31726
rect 27468 31612 27860 31668
rect 26796 28812 27300 28868
rect 26796 28754 26852 28812
rect 26796 28702 26798 28754
rect 26850 28702 26852 28754
rect 26796 28690 26852 28702
rect 27020 28644 27076 28654
rect 27020 28550 27076 28588
rect 27244 28532 27300 28812
rect 27244 28438 27300 28476
rect 27356 28530 27412 28542
rect 27356 28478 27358 28530
rect 27410 28478 27412 28530
rect 26684 28252 27300 28308
rect 27132 27188 27188 28252
rect 27244 28082 27300 28252
rect 27244 28030 27246 28082
rect 27298 28030 27300 28082
rect 27244 28018 27300 28030
rect 27356 28084 27412 28478
rect 27356 28018 27412 28028
rect 27468 27860 27524 31612
rect 27916 31220 27972 31230
rect 27916 31126 27972 31164
rect 27804 30210 27860 30222
rect 27804 30158 27806 30210
rect 27858 30158 27860 30210
rect 27132 27094 27188 27132
rect 27244 27804 27524 27860
rect 27580 29428 27636 29438
rect 26012 26852 26292 26908
rect 26460 26964 26516 26974
rect 25004 25666 25060 25676
rect 25676 26066 25732 26078
rect 25676 26014 25678 26066
rect 25730 26014 25732 26066
rect 25676 25396 25732 26014
rect 25676 25330 25732 25340
rect 25900 25732 25956 25742
rect 24556 24894 24558 24946
rect 24610 24894 24612 24946
rect 24556 24882 24612 24894
rect 25564 24948 25620 24958
rect 24332 24388 24388 24780
rect 24668 24722 24724 24734
rect 24668 24670 24670 24722
rect 24722 24670 24724 24722
rect 24668 24612 24724 24670
rect 25452 24724 25508 24734
rect 25340 24612 25396 24622
rect 24724 24556 25172 24612
rect 24668 24546 24724 24556
rect 24780 24388 24836 24398
rect 24332 24332 24780 24388
rect 24444 24164 24500 24174
rect 23100 24108 23492 24164
rect 23436 24050 23492 24108
rect 23436 23998 23438 24050
rect 23490 23998 23492 24050
rect 23436 23986 23492 23998
rect 24108 23938 24164 23950
rect 24108 23886 24110 23938
rect 24162 23886 24164 23938
rect 22876 22418 22932 22428
rect 22988 23154 23044 23166
rect 22988 23102 22990 23154
rect 23042 23102 23044 23154
rect 22540 21758 22542 21810
rect 22594 21758 22596 21810
rect 22540 21746 22596 21758
rect 22428 21646 22430 21698
rect 22482 21646 22484 21698
rect 22428 20802 22484 21646
rect 22428 20750 22430 20802
rect 22482 20750 22484 20802
rect 22428 20738 22484 20750
rect 22988 20804 23044 23102
rect 23660 23044 23716 23054
rect 24108 23044 24164 23886
rect 24444 23938 24500 24108
rect 24444 23886 24446 23938
rect 24498 23886 24500 23938
rect 24444 23874 24500 23886
rect 24780 23938 24836 24332
rect 24780 23886 24782 23938
rect 24834 23886 24836 23938
rect 24780 23874 24836 23886
rect 25004 24164 25060 24174
rect 24332 23828 24388 23838
rect 24220 23492 24276 23502
rect 24220 23378 24276 23436
rect 24220 23326 24222 23378
rect 24274 23326 24276 23378
rect 24220 23314 24276 23326
rect 23660 23042 24164 23044
rect 23660 22990 23662 23042
rect 23714 22990 24164 23042
rect 23660 22988 24164 22990
rect 22988 20738 23044 20748
rect 23100 22370 23156 22382
rect 23100 22318 23102 22370
rect 23154 22318 23156 22370
rect 23100 21698 23156 22318
rect 23100 21646 23102 21698
rect 23154 21646 23156 21698
rect 22204 20638 22206 20690
rect 22258 20638 22260 20690
rect 22204 20626 22260 20638
rect 22540 20692 22596 20702
rect 21644 20412 22372 20468
rect 21420 19906 21588 19908
rect 21420 19854 21534 19906
rect 21586 19854 21588 19906
rect 21420 19852 21588 19854
rect 21420 19796 21476 19852
rect 21532 19842 21588 19852
rect 20524 19282 20580 19292
rect 21308 19740 21476 19796
rect 21308 19346 21364 19740
rect 21308 19294 21310 19346
rect 21362 19294 21364 19346
rect 21308 19282 21364 19294
rect 21420 19348 21476 19358
rect 20412 18676 20468 19180
rect 21420 19234 21476 19292
rect 21420 19182 21422 19234
rect 21474 19182 21476 19234
rect 21420 19170 21476 19182
rect 21756 19236 21812 19246
rect 21756 19142 21812 19180
rect 19964 18610 20020 18620
rect 20412 18610 20468 18620
rect 19852 18510 19854 18562
rect 19906 18510 19908 18562
rect 19852 18498 19908 18510
rect 20300 18564 20356 18574
rect 20188 18452 20244 18462
rect 20300 18452 20356 18508
rect 20188 18450 20356 18452
rect 20188 18398 20190 18450
rect 20242 18398 20356 18450
rect 20188 18396 20356 18398
rect 20748 18450 20804 18462
rect 20748 18398 20750 18450
rect 20802 18398 20804 18450
rect 20188 18386 20244 18396
rect 19628 17490 19684 17500
rect 20636 17556 20692 17566
rect 20636 17462 20692 17500
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19516 16818 19572 16828
rect 18844 15876 18900 16380
rect 20636 16324 20692 16334
rect 20636 16230 20692 16268
rect 19180 16100 19236 16110
rect 19180 16006 19236 16044
rect 20524 16098 20580 16110
rect 20524 16046 20526 16098
rect 20578 16046 20580 16098
rect 18844 15810 18900 15820
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 20524 15540 20580 16046
rect 20524 15474 20580 15484
rect 20636 15652 20692 15662
rect 20748 15652 20804 18398
rect 21308 18450 21364 18462
rect 21308 18398 21310 18450
rect 21362 18398 21364 18450
rect 21308 17444 21364 18398
rect 22092 18450 22148 18462
rect 22092 18398 22094 18450
rect 22146 18398 22148 18450
rect 21308 17378 21364 17388
rect 21868 17666 21924 17678
rect 21868 17614 21870 17666
rect 21922 17614 21924 17666
rect 20972 17108 21028 17118
rect 20972 16994 21028 17052
rect 20972 16942 20974 16994
rect 21026 16942 21028 16994
rect 20972 16930 21028 16942
rect 21868 16100 21924 17614
rect 21980 17556 22036 17566
rect 22092 17556 22148 18398
rect 22036 17554 22148 17556
rect 22036 17502 22094 17554
rect 22146 17502 22148 17554
rect 22036 17500 22148 17502
rect 21980 16882 22036 17500
rect 22092 17490 22148 17500
rect 21980 16830 21982 16882
rect 22034 16830 22036 16882
rect 21980 16818 22036 16830
rect 21868 16034 21924 16044
rect 20692 15596 20804 15652
rect 21532 15876 21588 15886
rect 19180 15316 19236 15326
rect 18508 15314 19236 15316
rect 18508 15262 18510 15314
rect 18562 15262 19182 15314
rect 19234 15262 19236 15314
rect 18508 15260 19236 15262
rect 18508 15250 18564 15260
rect 19180 15250 19236 15260
rect 20636 15314 20692 15596
rect 20636 15262 20638 15314
rect 20690 15262 20692 15314
rect 20636 15250 20692 15262
rect 21196 15428 21252 15438
rect 19292 15204 19348 15242
rect 19292 15138 19348 15148
rect 21196 15148 21252 15372
rect 21308 15316 21364 15326
rect 21308 15222 21364 15260
rect 21532 15148 21588 15820
rect 22204 15316 22260 15354
rect 22204 15250 22260 15260
rect 22316 15148 22372 20412
rect 22540 20130 22596 20636
rect 23100 20692 23156 21646
rect 23436 22370 23492 22382
rect 23436 22318 23438 22370
rect 23490 22318 23492 22370
rect 23100 20626 23156 20636
rect 23212 21474 23268 21486
rect 23212 21422 23214 21474
rect 23266 21422 23268 21474
rect 22540 20078 22542 20130
rect 22594 20078 22596 20130
rect 22540 20066 22596 20078
rect 23212 20132 23268 21422
rect 23324 21364 23380 21374
rect 23436 21364 23492 22318
rect 23660 21700 23716 22988
rect 24108 22596 24164 22606
rect 23884 22372 23940 22382
rect 23884 21810 23940 22316
rect 24108 22370 24164 22540
rect 24108 22318 24110 22370
rect 24162 22318 24164 22370
rect 24108 22306 24164 22318
rect 23884 21758 23886 21810
rect 23938 21758 23940 21810
rect 23884 21746 23940 21758
rect 24332 21810 24388 23772
rect 24668 23828 24724 23838
rect 24668 23734 24724 23772
rect 24780 23604 24836 23614
rect 24780 23378 24836 23548
rect 24780 23326 24782 23378
rect 24834 23326 24836 23378
rect 24780 23314 24836 23326
rect 24444 23268 24500 23278
rect 24444 23174 24500 23212
rect 24556 23266 24612 23278
rect 24556 23214 24558 23266
rect 24610 23214 24612 23266
rect 24332 21758 24334 21810
rect 24386 21758 24388 21810
rect 24332 21746 24388 21758
rect 23660 21634 23716 21644
rect 24556 21476 24612 23214
rect 24892 22484 24948 22494
rect 25004 22484 25060 24108
rect 25116 23938 25172 24556
rect 25340 24518 25396 24556
rect 25116 23886 25118 23938
rect 25170 23886 25172 23938
rect 25116 23874 25172 23886
rect 25340 24052 25396 24062
rect 25340 23714 25396 23996
rect 25452 23938 25508 24668
rect 25452 23886 25454 23938
rect 25506 23886 25508 23938
rect 25452 23874 25508 23886
rect 25340 23662 25342 23714
rect 25394 23662 25396 23714
rect 25340 23650 25396 23662
rect 25228 23492 25284 23502
rect 25228 23378 25284 23436
rect 25564 23380 25620 24892
rect 25900 24946 25956 25676
rect 25900 24894 25902 24946
rect 25954 24894 25956 24946
rect 25900 24882 25956 24894
rect 26012 24946 26068 26852
rect 26012 24894 26014 24946
rect 26066 24894 26068 24946
rect 26012 24882 26068 24894
rect 26124 26290 26180 26302
rect 26124 26238 26126 26290
rect 26178 26238 26180 26290
rect 25788 24722 25844 24734
rect 25788 24670 25790 24722
rect 25842 24670 25844 24722
rect 25676 23828 25732 23838
rect 25676 23734 25732 23772
rect 25228 23326 25230 23378
rect 25282 23326 25284 23378
rect 25228 23314 25284 23326
rect 25340 23378 25620 23380
rect 25340 23326 25566 23378
rect 25618 23326 25620 23378
rect 25340 23324 25620 23326
rect 24892 22482 25060 22484
rect 24892 22430 24894 22482
rect 24946 22430 25060 22482
rect 24892 22428 25060 22430
rect 24892 22418 24948 22428
rect 25340 22258 25396 23324
rect 25564 23314 25620 23324
rect 25676 22484 25732 22494
rect 25788 22484 25844 24670
rect 26124 23826 26180 26238
rect 26348 26290 26404 26302
rect 26348 26238 26350 26290
rect 26402 26238 26404 26290
rect 26348 25396 26404 26238
rect 26124 23774 26126 23826
rect 26178 23774 26180 23826
rect 26124 23044 26180 23774
rect 26124 22978 26180 22988
rect 26236 25340 26348 25396
rect 25676 22482 25844 22484
rect 25676 22430 25678 22482
rect 25730 22430 25844 22482
rect 25676 22428 25844 22430
rect 25676 22418 25732 22428
rect 25900 22372 25956 22382
rect 25340 22206 25342 22258
rect 25394 22206 25396 22258
rect 25340 22194 25396 22206
rect 25788 22316 25900 22372
rect 25788 22258 25844 22316
rect 25900 22306 25956 22316
rect 25788 22206 25790 22258
rect 25842 22206 25844 22258
rect 25788 22194 25844 22206
rect 25564 22148 25620 22158
rect 25564 22146 25732 22148
rect 25564 22094 25566 22146
rect 25618 22094 25732 22146
rect 25564 22092 25732 22094
rect 25564 22082 25620 22092
rect 25676 22036 25732 22092
rect 26236 22036 26292 25340
rect 26348 25330 26404 25340
rect 26348 24836 26404 24846
rect 26348 23938 26404 24780
rect 26460 24722 26516 26908
rect 26684 26290 26740 26302
rect 26684 26238 26686 26290
rect 26738 26238 26740 26290
rect 26572 25506 26628 25518
rect 26572 25454 26574 25506
rect 26626 25454 26628 25506
rect 26572 25282 26628 25454
rect 26572 25230 26574 25282
rect 26626 25230 26628 25282
rect 26572 25218 26628 25230
rect 26684 24948 26740 26238
rect 26684 24882 26740 24892
rect 26796 25284 26852 25294
rect 27020 25284 27076 25294
rect 26796 25282 27076 25284
rect 26796 25230 26798 25282
rect 26850 25230 27022 25282
rect 27074 25230 27076 25282
rect 26796 25228 27076 25230
rect 26460 24670 26462 24722
rect 26514 24670 26516 24722
rect 26460 24658 26516 24670
rect 26348 23886 26350 23938
rect 26402 23886 26404 23938
rect 26348 23874 26404 23886
rect 26796 23492 26852 25228
rect 27020 25218 27076 25228
rect 27244 24948 27300 27804
rect 27580 27748 27636 29372
rect 27804 29204 27860 30158
rect 28028 29988 28084 31948
rect 27804 28756 27860 29148
rect 27804 28690 27860 28700
rect 27916 29932 28084 29988
rect 27804 28532 27860 28542
rect 27804 28438 27860 28476
rect 27468 27692 27636 27748
rect 27804 28084 27860 28094
rect 27356 26964 27412 27002
rect 27356 26898 27412 26908
rect 27244 24882 27300 24892
rect 27356 25172 27412 25182
rect 26796 23426 26852 23436
rect 26908 24834 26964 24846
rect 26908 24782 26910 24834
rect 26962 24782 26964 24834
rect 26796 23156 26852 23166
rect 26796 23062 26852 23100
rect 25676 21980 26292 22036
rect 26460 22484 26516 22494
rect 26460 22258 26516 22428
rect 26460 22206 26462 22258
rect 26514 22206 26516 22258
rect 25564 21924 25620 21934
rect 25340 21700 25396 21710
rect 25340 21586 25396 21644
rect 25340 21534 25342 21586
rect 25394 21534 25396 21586
rect 25340 21522 25396 21534
rect 24668 21476 24724 21486
rect 24556 21474 24724 21476
rect 24556 21422 24670 21474
rect 24722 21422 24724 21474
rect 24556 21420 24724 21422
rect 23324 21362 23492 21364
rect 23324 21310 23326 21362
rect 23378 21310 23492 21362
rect 23324 21308 23492 21310
rect 23324 20188 23380 21308
rect 24668 21252 24724 21420
rect 24668 21186 24724 21196
rect 23996 20804 24052 20814
rect 23996 20710 24052 20748
rect 24108 20690 24164 20702
rect 24108 20638 24110 20690
rect 24162 20638 24164 20690
rect 23884 20244 23940 20264
rect 23324 20132 23940 20188
rect 23212 20066 23268 20076
rect 22764 20018 22820 20030
rect 22764 19966 22766 20018
rect 22818 19966 22820 20018
rect 22764 19458 22820 19966
rect 23660 20018 23716 20030
rect 23660 19966 23662 20018
rect 23714 19966 23716 20018
rect 22764 19406 22766 19458
rect 22818 19406 22820 19458
rect 22764 19394 22820 19406
rect 23212 19906 23268 19918
rect 23212 19854 23214 19906
rect 23266 19854 23268 19906
rect 23212 19348 23268 19854
rect 23212 19282 23268 19292
rect 23436 19346 23492 19358
rect 23436 19294 23438 19346
rect 23490 19294 23492 19346
rect 22876 19122 22932 19134
rect 22876 19070 22878 19122
rect 22930 19070 22932 19122
rect 22764 19010 22820 19022
rect 22764 18958 22766 19010
rect 22818 18958 22820 19010
rect 22764 18564 22820 18958
rect 22764 18498 22820 18508
rect 22540 18338 22596 18350
rect 22540 18286 22542 18338
rect 22594 18286 22596 18338
rect 22540 17668 22596 18286
rect 22876 17892 22932 19070
rect 22876 17826 22932 17836
rect 23436 17892 23492 19294
rect 23548 19122 23604 19134
rect 23548 19070 23550 19122
rect 23602 19070 23604 19122
rect 23548 18564 23604 19070
rect 23660 18674 23716 19966
rect 23660 18622 23662 18674
rect 23714 18622 23716 18674
rect 23660 18610 23716 18622
rect 23548 18452 23604 18508
rect 23772 18562 23828 18574
rect 23772 18510 23774 18562
rect 23826 18510 23828 18562
rect 23772 18452 23828 18510
rect 23548 18396 23828 18452
rect 23548 18226 23604 18238
rect 23548 18174 23550 18226
rect 23602 18174 23604 18226
rect 23548 17892 23604 18174
rect 23492 17836 23604 17892
rect 23436 17826 23492 17836
rect 23212 17668 23268 17678
rect 22540 17602 22596 17612
rect 23100 17612 23212 17668
rect 23100 16882 23156 17612
rect 23212 17574 23268 17612
rect 23212 16996 23268 17006
rect 23212 16902 23268 16940
rect 23100 16830 23102 16882
rect 23154 16830 23156 16882
rect 23100 16818 23156 16830
rect 23772 16770 23828 16782
rect 23772 16718 23774 16770
rect 23826 16718 23828 16770
rect 23772 16324 23828 16718
rect 23772 16258 23828 16268
rect 22428 16100 22484 16110
rect 22484 16044 22708 16100
rect 22428 16006 22484 16044
rect 22540 15874 22596 15886
rect 22540 15822 22542 15874
rect 22594 15822 22596 15874
rect 22540 15764 22596 15822
rect 22540 15698 22596 15708
rect 21196 15092 21588 15148
rect 18396 14644 18452 14654
rect 18396 14550 18452 14588
rect 19068 14644 19124 14654
rect 19068 13860 19124 14588
rect 19068 13794 19124 13804
rect 19292 14530 19348 14542
rect 19292 14478 19294 14530
rect 19346 14478 19348 14530
rect 18732 13748 18788 13758
rect 18732 13654 18788 13692
rect 18284 13634 18452 13636
rect 18284 13582 18286 13634
rect 18338 13582 18452 13634
rect 18284 13580 18452 13582
rect 18284 13570 18340 13580
rect 17724 13524 17780 13534
rect 17724 13522 18004 13524
rect 17724 13470 17726 13522
rect 17778 13470 18004 13522
rect 17724 13468 18004 13470
rect 17724 13458 17780 13468
rect 17948 12516 18004 13468
rect 17836 12460 18340 12516
rect 17388 11732 17556 11788
rect 17724 12178 17780 12190
rect 17724 12126 17726 12178
rect 17778 12126 17780 12178
rect 16380 10834 16548 10836
rect 16380 10782 16382 10834
rect 16434 10782 16548 10834
rect 16380 10780 16548 10782
rect 16380 10770 16436 10780
rect 16940 10612 16996 11452
rect 17164 11620 17220 11630
rect 17164 11394 17220 11564
rect 17164 11342 17166 11394
rect 17218 11342 17220 11394
rect 17164 11330 17220 11342
rect 16940 10546 16996 10556
rect 16492 10500 16548 10510
rect 16492 10406 16548 10444
rect 15708 10386 16324 10388
rect 15708 10334 16158 10386
rect 16210 10334 16324 10386
rect 15708 10332 16324 10334
rect 15036 9886 15038 9938
rect 15090 9886 15092 9938
rect 15036 9874 15092 9886
rect 15148 9826 15204 9838
rect 15148 9774 15150 9826
rect 15202 9774 15204 9826
rect 13916 9154 14196 9156
rect 13916 9102 13918 9154
rect 13970 9102 14196 9154
rect 13916 9100 14196 9102
rect 14364 9660 14532 9716
rect 14812 9716 14868 9726
rect 13916 9090 13972 9100
rect 11900 8878 11902 8930
rect 11954 8878 11956 8930
rect 11900 8428 11956 8878
rect 13244 9042 13300 9054
rect 13244 8990 13246 9042
rect 13298 8990 13300 9042
rect 11900 8372 12628 8428
rect 12572 8260 12628 8372
rect 13244 8372 13300 8990
rect 13244 8306 13300 8316
rect 13580 8372 13636 8382
rect 13580 8278 13636 8316
rect 12572 8194 12628 8204
rect 13804 8260 13860 8270
rect 11452 8148 11508 8158
rect 11340 8146 11508 8148
rect 11340 8094 11454 8146
rect 11506 8094 11508 8146
rect 11340 8092 11508 8094
rect 11228 7858 11284 7868
rect 11116 7634 11172 7644
rect 11452 7588 11508 8092
rect 11676 8148 11732 8158
rect 11676 8054 11732 8092
rect 11452 7522 11508 7532
rect 11900 8034 11956 8046
rect 11900 7982 11902 8034
rect 11954 7982 11956 8034
rect 11004 7410 11060 7420
rect 11900 7474 11956 7982
rect 13580 7588 13636 7598
rect 11900 7422 11902 7474
rect 11954 7422 11956 7474
rect 11900 7410 11956 7422
rect 12572 7476 12628 7486
rect 12572 7382 12628 7420
rect 8204 7252 8260 7262
rect 7532 7250 8260 7252
rect 7532 7198 8206 7250
rect 8258 7198 8260 7250
rect 7532 7196 8260 7198
rect 5964 7158 6020 7196
rect 8204 7186 8260 7196
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 13580 6802 13636 7532
rect 13804 7474 13860 8204
rect 13804 7422 13806 7474
rect 13858 7422 13860 7474
rect 13804 7410 13860 7422
rect 13916 8036 13972 8046
rect 13580 6750 13582 6802
rect 13634 6750 13636 6802
rect 13580 6738 13636 6750
rect 13916 6804 13972 7980
rect 14028 7252 14084 7262
rect 14028 7158 14084 7196
rect 13916 6690 13972 6748
rect 13916 6638 13918 6690
rect 13970 6638 13972 6690
rect 13916 6626 13972 6638
rect 14364 5908 14420 9660
rect 14812 9622 14868 9660
rect 15148 9380 15204 9774
rect 14476 9324 15204 9380
rect 14476 8370 14532 9324
rect 14700 9210 14756 9222
rect 14588 9156 14644 9166
rect 14700 9158 14702 9210
rect 14754 9158 14756 9210
rect 14700 9156 14756 9158
rect 14812 9212 15092 9268
rect 14812 9156 14868 9212
rect 14700 9100 14812 9156
rect 14588 9062 14644 9100
rect 14812 9090 14868 9100
rect 14476 8318 14478 8370
rect 14530 8318 14532 8370
rect 14476 8306 14532 8318
rect 14924 9042 14980 9054
rect 14924 8990 14926 9042
rect 14978 8990 14980 9042
rect 14924 8148 14980 8990
rect 15036 8370 15092 9212
rect 15484 9154 15540 9166
rect 15484 9102 15486 9154
rect 15538 9102 15540 9154
rect 15036 8318 15038 8370
rect 15090 8318 15092 8370
rect 15036 8306 15092 8318
rect 15148 9042 15204 9054
rect 15148 8990 15150 9042
rect 15202 8990 15204 9042
rect 14924 8082 14980 8092
rect 14812 7924 14868 7934
rect 14588 7700 14644 7710
rect 14476 7474 14532 7486
rect 14476 7422 14478 7474
rect 14530 7422 14532 7474
rect 14476 7364 14532 7422
rect 14588 7364 14644 7644
rect 14700 7588 14756 7598
rect 14700 7494 14756 7532
rect 14812 7586 14868 7868
rect 14812 7534 14814 7586
rect 14866 7534 14868 7586
rect 14812 7522 14868 7534
rect 15148 7588 15204 8990
rect 15148 7522 15204 7532
rect 15372 8370 15428 8382
rect 15372 8318 15374 8370
rect 15426 8318 15428 8370
rect 15260 7364 15316 7402
rect 14532 7308 14868 7364
rect 14476 7298 14532 7308
rect 14700 6804 14756 6814
rect 14700 6690 14756 6748
rect 14700 6638 14702 6690
rect 14754 6638 14756 6690
rect 14700 6626 14756 6638
rect 14812 6578 14868 7308
rect 15260 7298 15316 7308
rect 15372 6916 15428 8318
rect 15484 7700 15540 9102
rect 15708 8932 15764 8942
rect 16156 8932 16212 10332
rect 17388 10052 17444 11732
rect 17724 11620 17780 12126
rect 17724 11554 17780 11564
rect 17612 11396 17668 11406
rect 17612 11170 17668 11340
rect 17724 11396 17780 11406
rect 17836 11396 17892 12460
rect 17948 12290 18004 12302
rect 17948 12238 17950 12290
rect 18002 12238 18004 12290
rect 17948 11956 18004 12238
rect 18284 12290 18340 12460
rect 18396 12404 18452 13580
rect 18732 13524 18788 13534
rect 18732 13074 18788 13468
rect 19292 13524 19348 14478
rect 19964 14420 20020 14430
rect 20300 14420 20356 14430
rect 19964 14418 20356 14420
rect 19964 14366 19966 14418
rect 20018 14366 20302 14418
rect 20354 14366 20356 14418
rect 19964 14364 20356 14366
rect 19964 14354 20020 14364
rect 20300 14354 20356 14364
rect 21420 14418 21476 14430
rect 21420 14366 21422 14418
rect 21474 14366 21476 14418
rect 19292 13458 19348 13468
rect 19628 14308 19684 14318
rect 18732 13022 18734 13074
rect 18786 13022 18788 13074
rect 18396 12338 18452 12348
rect 18508 12402 18564 12414
rect 18508 12350 18510 12402
rect 18562 12350 18564 12402
rect 18284 12238 18286 12290
rect 18338 12238 18340 12290
rect 18284 12226 18340 12238
rect 17948 11890 18004 11900
rect 17724 11394 17892 11396
rect 17724 11342 17726 11394
rect 17778 11342 17892 11394
rect 17724 11340 17892 11342
rect 17724 11330 17780 11340
rect 17612 11118 17614 11170
rect 17666 11118 17668 11170
rect 17612 11106 17668 11118
rect 17836 10610 17892 11340
rect 17836 10558 17838 10610
rect 17890 10558 17892 10610
rect 17836 10546 17892 10558
rect 18284 11844 18340 11854
rect 17724 10500 17780 10510
rect 17724 10406 17780 10444
rect 17388 9996 17780 10052
rect 17612 9828 17668 9838
rect 17612 9734 17668 9772
rect 17724 9714 17780 9996
rect 18284 9828 18340 11788
rect 18508 11394 18564 12350
rect 18732 11618 18788 13022
rect 19068 12850 19124 12862
rect 19068 12798 19070 12850
rect 19122 12798 19124 12850
rect 19068 12740 19124 12798
rect 19628 12740 19684 14252
rect 20412 14308 20468 14318
rect 20412 14214 20468 14252
rect 20636 14308 20692 14318
rect 20636 14214 20692 14252
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 20860 13972 20916 13982
rect 19740 13860 19796 13870
rect 19740 13746 19796 13804
rect 20412 13860 20468 13870
rect 19740 13694 19742 13746
rect 19794 13694 19796 13746
rect 19740 13682 19796 13694
rect 20076 13746 20132 13758
rect 20076 13694 20078 13746
rect 20130 13694 20132 13746
rect 20076 13524 20132 13694
rect 20076 13458 20132 13468
rect 20412 12850 20468 13804
rect 20748 13636 20804 13646
rect 20748 13412 20804 13580
rect 20860 13634 20916 13916
rect 20860 13582 20862 13634
rect 20914 13582 20916 13634
rect 20860 13570 20916 13582
rect 20748 13356 20916 13412
rect 20748 12964 20804 12974
rect 20748 12870 20804 12908
rect 20412 12798 20414 12850
rect 20466 12798 20468 12850
rect 20412 12786 20468 12798
rect 19068 12684 19684 12740
rect 19628 12404 19684 12684
rect 20748 12740 20804 12750
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19740 12404 19796 12414
rect 19628 12402 19796 12404
rect 19628 12350 19742 12402
rect 19794 12350 19796 12402
rect 19628 12348 19796 12350
rect 19740 12338 19796 12348
rect 19964 12404 20020 12414
rect 19516 12292 19572 12302
rect 19516 12198 19572 12236
rect 19964 12290 20020 12348
rect 19964 12238 19966 12290
rect 20018 12238 20020 12290
rect 19180 12178 19236 12190
rect 19180 12126 19182 12178
rect 19234 12126 19236 12178
rect 19180 11844 19236 12126
rect 19964 12068 20020 12238
rect 20076 12292 20132 12302
rect 20076 12198 20132 12236
rect 20748 12292 20804 12684
rect 20860 12402 20916 13356
rect 21420 13076 21476 14366
rect 21532 14308 21588 15092
rect 22092 15092 22372 15148
rect 22428 15540 22484 15550
rect 22428 15314 22484 15484
rect 22428 15262 22430 15314
rect 22482 15262 22484 15314
rect 21756 14420 21812 14430
rect 21756 14326 21812 14364
rect 21532 14306 21700 14308
rect 21532 14254 21534 14306
rect 21586 14254 21700 14306
rect 21532 14252 21700 14254
rect 21532 14242 21588 14252
rect 21644 13970 21700 14252
rect 21644 13918 21646 13970
rect 21698 13918 21700 13970
rect 21644 13906 21700 13918
rect 21420 13020 21812 13076
rect 21420 12740 21476 13020
rect 21756 12962 21812 13020
rect 21756 12910 21758 12962
rect 21810 12910 21812 12962
rect 21756 12898 21812 12910
rect 21420 12674 21476 12684
rect 20860 12350 20862 12402
rect 20914 12350 20916 12402
rect 20860 12338 20916 12350
rect 20748 12198 20804 12236
rect 21084 12178 21140 12190
rect 21084 12126 21086 12178
rect 21138 12126 21140 12178
rect 19964 12012 20468 12068
rect 19180 11778 19236 11788
rect 18732 11566 18734 11618
rect 18786 11566 18788 11618
rect 18732 11554 18788 11566
rect 20300 11620 20356 11630
rect 20188 11508 20244 11518
rect 18508 11342 18510 11394
rect 18562 11342 18564 11394
rect 18508 11330 18564 11342
rect 19180 11396 19236 11406
rect 19180 11302 19236 11340
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19964 10724 20020 10734
rect 20188 10724 20244 11452
rect 19964 10722 20244 10724
rect 19964 10670 19966 10722
rect 20018 10670 20244 10722
rect 19964 10668 20244 10670
rect 20300 11394 20356 11564
rect 20300 11342 20302 11394
rect 20354 11342 20356 11394
rect 19964 10658 20020 10668
rect 19180 10612 19236 10622
rect 20300 10612 20356 11342
rect 20412 10834 20468 12012
rect 21084 11284 21140 12126
rect 21868 12178 21924 12190
rect 21868 12126 21870 12178
rect 21922 12126 21924 12178
rect 21420 12066 21476 12078
rect 21420 12014 21422 12066
rect 21474 12014 21476 12066
rect 21420 11508 21476 12014
rect 21420 11442 21476 11452
rect 21532 11620 21588 11630
rect 21868 11620 21924 12126
rect 21588 11564 21924 11620
rect 21532 11506 21588 11564
rect 21532 11454 21534 11506
rect 21586 11454 21588 11506
rect 21532 11442 21588 11454
rect 21644 11284 21700 11294
rect 21084 11282 21700 11284
rect 21084 11230 21646 11282
rect 21698 11230 21700 11282
rect 21084 11228 21700 11230
rect 21644 11218 21700 11228
rect 22092 11172 22148 15092
rect 22204 14644 22260 14654
rect 22428 14644 22484 15262
rect 22652 15428 22708 16044
rect 22764 15988 22820 15998
rect 22764 15894 22820 15932
rect 23100 15876 23156 15886
rect 23100 15782 23156 15820
rect 23660 15876 23716 15886
rect 22652 15148 22708 15372
rect 23660 15426 23716 15820
rect 23884 15764 23940 20132
rect 24108 19796 24164 20638
rect 25452 20692 25508 20702
rect 25452 20598 25508 20636
rect 24556 20132 24612 20142
rect 24556 20038 24612 20076
rect 24108 19702 24164 19740
rect 25452 19348 25508 19358
rect 25564 19348 25620 21868
rect 26460 21924 26516 22206
rect 26460 21858 26516 21868
rect 26796 22370 26852 22382
rect 26796 22318 26798 22370
rect 26850 22318 26852 22370
rect 25676 21812 25732 21822
rect 25676 20580 25732 21756
rect 26012 21476 26068 21486
rect 26012 21474 26180 21476
rect 26012 21422 26014 21474
rect 26066 21422 26180 21474
rect 26012 21420 26180 21422
rect 26012 21410 26068 21420
rect 25676 20130 25732 20524
rect 26012 20802 26068 20814
rect 26012 20750 26014 20802
rect 26066 20750 26068 20802
rect 25900 20356 25956 20366
rect 25900 20242 25956 20300
rect 25900 20190 25902 20242
rect 25954 20190 25956 20242
rect 25900 20178 25956 20190
rect 26012 20244 26068 20750
rect 26124 20580 26180 21420
rect 26796 21252 26852 22318
rect 26796 21186 26852 21196
rect 26908 20804 26964 24782
rect 27132 24722 27188 24734
rect 27132 24670 27134 24722
rect 27186 24670 27188 24722
rect 27020 23828 27076 23838
rect 27020 23734 27076 23772
rect 27132 22596 27188 24670
rect 27356 24724 27412 25116
rect 27468 24836 27524 27692
rect 27580 27188 27636 27198
rect 27580 26962 27636 27132
rect 27580 26910 27582 26962
rect 27634 26910 27636 26962
rect 27580 26898 27636 26910
rect 27692 26908 27748 26918
rect 27804 26908 27860 28028
rect 27692 26906 27860 26908
rect 27692 26854 27694 26906
rect 27746 26854 27860 26906
rect 27692 26852 27860 26854
rect 27692 26842 27748 26852
rect 27692 26628 27748 26638
rect 27692 26290 27748 26572
rect 27916 26402 27972 29932
rect 28140 29876 28196 31948
rect 28252 31778 28308 31790
rect 28252 31726 28254 31778
rect 28306 31726 28308 31778
rect 28252 31556 28308 31726
rect 28364 31668 28420 32172
rect 28588 32004 28644 32510
rect 28700 32450 28756 32462
rect 28700 32398 28702 32450
rect 28754 32398 28756 32450
rect 28700 32116 28756 32398
rect 28700 32050 28756 32060
rect 28588 31938 28644 31948
rect 28364 31602 28420 31612
rect 28252 31490 28308 31500
rect 28364 31220 28420 31230
rect 28252 30996 28308 31006
rect 28252 30902 28308 30940
rect 28364 30436 28420 31164
rect 28924 31220 28980 31258
rect 28924 31154 28980 31164
rect 28476 31106 28532 31118
rect 28476 31054 28478 31106
rect 28530 31054 28532 31106
rect 28476 30884 28532 31054
rect 28924 30996 28980 31006
rect 29036 30996 29092 35980
rect 29260 35698 29316 35710
rect 29260 35646 29262 35698
rect 29314 35646 29316 35698
rect 29260 35476 29316 35646
rect 29260 35410 29316 35420
rect 29148 35252 29204 35262
rect 29148 34914 29204 35196
rect 29148 34862 29150 34914
rect 29202 34862 29204 34914
rect 29148 34130 29204 34862
rect 29148 34078 29150 34130
rect 29202 34078 29204 34130
rect 29148 34066 29204 34078
rect 29372 35252 29428 35980
rect 29484 35980 29876 36036
rect 29932 36652 30044 36708
rect 29484 35476 29540 35980
rect 29820 35812 29876 35850
rect 29820 35746 29876 35756
rect 29708 35698 29764 35710
rect 29708 35646 29710 35698
rect 29762 35646 29764 35698
rect 29708 35588 29764 35646
rect 29708 35532 29876 35588
rect 29484 35420 29764 35476
rect 29372 34914 29428 35196
rect 29372 34862 29374 34914
rect 29426 34862 29428 34914
rect 29372 34244 29428 34862
rect 29708 34914 29764 35420
rect 29820 35252 29876 35532
rect 29820 35186 29876 35196
rect 29708 34862 29710 34914
rect 29762 34862 29764 34914
rect 29484 34692 29540 34702
rect 29484 34598 29540 34636
rect 29596 34690 29652 34702
rect 29596 34638 29598 34690
rect 29650 34638 29652 34690
rect 29596 34580 29652 34638
rect 29596 34514 29652 34524
rect 29596 34356 29652 34366
rect 29708 34356 29764 34862
rect 29652 34300 29764 34356
rect 29596 34262 29652 34300
rect 29484 34244 29540 34254
rect 29372 34242 29540 34244
rect 29372 34190 29486 34242
rect 29538 34190 29540 34242
rect 29372 34188 29540 34190
rect 29372 34132 29428 34188
rect 29484 34178 29540 34188
rect 29372 34066 29428 34076
rect 29820 34132 29876 34142
rect 29820 34038 29876 34076
rect 29372 33122 29428 33134
rect 29372 33070 29374 33122
rect 29426 33070 29428 33122
rect 29372 32676 29428 33070
rect 29428 32620 29540 32676
rect 29372 32610 29428 32620
rect 29372 31778 29428 31790
rect 29372 31726 29374 31778
rect 29426 31726 29428 31778
rect 29148 31668 29204 31678
rect 29148 31574 29204 31612
rect 29372 30996 29428 31726
rect 28980 30940 29092 30996
rect 29148 30940 29428 30996
rect 28924 30902 28980 30940
rect 28476 30818 28532 30828
rect 29036 30770 29092 30782
rect 29036 30718 29038 30770
rect 29090 30718 29092 30770
rect 28364 30212 28420 30380
rect 28588 30436 28644 30446
rect 29036 30436 29092 30718
rect 28588 30434 29092 30436
rect 28588 30382 28590 30434
rect 28642 30382 29092 30434
rect 28588 30380 29092 30382
rect 28588 30370 28644 30380
rect 29036 30324 29092 30380
rect 29036 30258 29092 30268
rect 28364 30156 28532 30212
rect 28476 30098 28532 30156
rect 28476 30046 28478 30098
rect 28530 30046 28532 30098
rect 28028 29820 28196 29876
rect 28252 29986 28308 29998
rect 28252 29934 28254 29986
rect 28306 29934 28308 29986
rect 28028 29428 28084 29820
rect 28140 29652 28196 29662
rect 28140 29558 28196 29596
rect 28028 29372 28196 29428
rect 27916 26350 27918 26402
rect 27970 26350 27972 26402
rect 27916 26338 27972 26350
rect 28028 28868 28084 28878
rect 28028 27186 28084 28812
rect 28140 27972 28196 29372
rect 28140 27906 28196 27916
rect 28028 27134 28030 27186
rect 28082 27134 28084 27186
rect 27692 26238 27694 26290
rect 27746 26238 27748 26290
rect 27692 26226 27748 26238
rect 27916 25620 27972 25658
rect 27468 24770 27524 24780
rect 27580 25564 27916 25620
rect 27356 24630 27412 24668
rect 27244 24500 27300 24510
rect 27244 24406 27300 24444
rect 27580 24052 27636 25564
rect 27916 25554 27972 25564
rect 28028 25284 28084 27134
rect 28252 26516 28308 29934
rect 28476 29652 28532 30046
rect 29036 29988 29092 29998
rect 29148 29988 29204 30940
rect 29484 30884 29540 32620
rect 29820 32564 29876 32574
rect 29820 32470 29876 32508
rect 29708 31780 29764 31790
rect 29708 30996 29764 31724
rect 29708 30930 29764 30940
rect 29820 31220 29876 31230
rect 29820 30994 29876 31164
rect 29820 30942 29822 30994
rect 29874 30942 29876 30994
rect 29372 30828 29540 30884
rect 29596 30884 29652 30894
rect 29260 30772 29316 30782
rect 29260 30678 29316 30716
rect 29092 29932 29204 29988
rect 29036 29894 29092 29932
rect 29372 29764 29428 30828
rect 29596 30772 29652 30828
rect 28812 29652 28868 29662
rect 28476 29538 28532 29596
rect 28700 29596 28812 29652
rect 28476 29486 28478 29538
rect 28530 29486 28532 29538
rect 28476 29474 28532 29486
rect 28588 29540 28644 29550
rect 28476 28756 28532 28766
rect 28588 28756 28644 29484
rect 28700 29538 28756 29596
rect 28812 29586 28868 29596
rect 28700 29486 28702 29538
rect 28754 29486 28756 29538
rect 28700 29474 28756 29486
rect 29148 29428 29204 29438
rect 29148 29334 29204 29372
rect 28812 29316 28868 29326
rect 28812 29222 28868 29260
rect 28588 28700 28756 28756
rect 28364 27972 28420 27982
rect 28364 27858 28420 27916
rect 28364 27806 28366 27858
rect 28418 27806 28420 27858
rect 28364 27794 28420 27806
rect 28476 26908 28532 28700
rect 28588 27076 28644 27114
rect 28588 27010 28644 27020
rect 28700 26908 28756 28700
rect 29148 28418 29204 28430
rect 29148 28366 29150 28418
rect 29202 28366 29204 28418
rect 28924 27860 28980 27870
rect 29148 27860 29204 28366
rect 28924 27858 29204 27860
rect 28924 27806 28926 27858
rect 28978 27806 29204 27858
rect 28924 27804 29204 27806
rect 28924 27794 28980 27804
rect 27356 23996 27636 24052
rect 27692 25228 28084 25284
rect 28140 26460 28308 26516
rect 28364 26852 28532 26908
rect 28588 26852 28756 26908
rect 29036 26908 29092 27804
rect 29260 27188 29316 27198
rect 29372 27188 29428 29708
rect 29484 30716 29652 30772
rect 29484 30210 29540 30716
rect 29708 30324 29764 30334
rect 29708 30230 29764 30268
rect 29484 30158 29486 30210
rect 29538 30158 29540 30210
rect 29484 29652 29540 30158
rect 29484 29596 29764 29652
rect 29596 29426 29652 29438
rect 29596 29374 29598 29426
rect 29650 29374 29652 29426
rect 29596 29316 29652 29374
rect 29596 29250 29652 29260
rect 29708 29092 29764 29596
rect 29484 28980 29540 28990
rect 29484 28866 29540 28924
rect 29484 28814 29486 28866
rect 29538 28814 29540 28866
rect 29484 28802 29540 28814
rect 29708 28754 29764 29036
rect 29820 28868 29876 30942
rect 29932 30772 29988 36652
rect 30044 36642 30100 36652
rect 30044 35698 30100 35710
rect 30044 35646 30046 35698
rect 30098 35646 30100 35698
rect 30044 35588 30100 35646
rect 30044 35522 30100 35532
rect 30156 34916 30212 38110
rect 30268 36708 30324 40572
rect 31052 40516 31108 40526
rect 30380 40404 30436 40414
rect 30380 40310 30436 40348
rect 30380 40180 30436 40190
rect 30380 39172 30436 40124
rect 31052 39618 31108 40460
rect 31052 39566 31054 39618
rect 31106 39566 31108 39618
rect 31052 39554 31108 39566
rect 30380 39058 30436 39116
rect 30380 39006 30382 39058
rect 30434 39006 30436 39058
rect 30380 38994 30436 39006
rect 31276 38724 31332 40910
rect 31836 40740 31892 40750
rect 31836 40514 31892 40684
rect 31836 40462 31838 40514
rect 31890 40462 31892 40514
rect 31836 40450 31892 40462
rect 31388 40402 31444 40414
rect 31388 40350 31390 40402
rect 31442 40350 31444 40402
rect 31388 38948 31444 40350
rect 31500 40404 31556 40414
rect 31500 40310 31556 40348
rect 31724 40290 31780 40302
rect 31724 40238 31726 40290
rect 31778 40238 31780 40290
rect 31724 39732 31780 40238
rect 31724 39676 32004 39732
rect 31948 39620 32004 39676
rect 31948 39526 32004 39564
rect 32060 39730 32116 39742
rect 32060 39678 32062 39730
rect 32114 39678 32116 39730
rect 31500 39508 31556 39518
rect 31500 39506 31892 39508
rect 31500 39454 31502 39506
rect 31554 39454 31892 39506
rect 31500 39452 31892 39454
rect 31500 39442 31556 39452
rect 31500 38948 31556 38958
rect 31388 38946 31556 38948
rect 31388 38894 31502 38946
rect 31554 38894 31556 38946
rect 31388 38892 31556 38894
rect 31500 38882 31556 38892
rect 31836 38836 31892 39452
rect 31724 38834 31892 38836
rect 31724 38782 31838 38834
rect 31890 38782 31892 38834
rect 31724 38780 31892 38782
rect 31612 38724 31668 38734
rect 31276 38722 31668 38724
rect 31276 38670 31614 38722
rect 31666 38670 31668 38722
rect 31276 38668 31668 38670
rect 30940 38052 30996 38062
rect 30492 37492 30548 37502
rect 30492 37398 30548 37436
rect 30940 37492 30996 37996
rect 30940 37398 30996 37436
rect 30268 36642 30324 36652
rect 30828 37380 30884 37390
rect 30828 36482 30884 37324
rect 30828 36430 30830 36482
rect 30882 36430 30884 36482
rect 30828 36418 30884 36430
rect 30156 34850 30212 34860
rect 30268 36370 30324 36382
rect 30268 36318 30270 36370
rect 30322 36318 30324 36370
rect 30268 34132 30324 36318
rect 31052 36260 31108 36270
rect 31052 36166 31108 36204
rect 31612 35924 31668 38668
rect 30940 35868 31668 35924
rect 30492 35698 30548 35710
rect 30492 35646 30494 35698
rect 30546 35646 30548 35698
rect 30492 35588 30548 35646
rect 30492 35522 30548 35532
rect 30380 35476 30436 35486
rect 30380 35026 30436 35420
rect 30380 34974 30382 35026
rect 30434 34974 30436 35026
rect 30380 34962 30436 34974
rect 30380 34132 30436 34142
rect 30268 34130 30436 34132
rect 30268 34078 30382 34130
rect 30434 34078 30436 34130
rect 30268 34076 30436 34078
rect 30380 34020 30436 34076
rect 30828 34132 30884 34142
rect 30828 34038 30884 34076
rect 30380 33954 30436 33964
rect 30604 34018 30660 34030
rect 30604 33966 30606 34018
rect 30658 33966 30660 34018
rect 30380 33122 30436 33134
rect 30380 33070 30382 33122
rect 30434 33070 30436 33122
rect 30044 32562 30100 32574
rect 30044 32510 30046 32562
rect 30098 32510 30100 32562
rect 30044 31892 30100 32510
rect 30380 32564 30436 33070
rect 30380 32498 30436 32508
rect 30604 32004 30660 33966
rect 30940 33796 30996 35868
rect 31164 35700 31220 35710
rect 31612 35700 31668 35710
rect 31164 35698 31668 35700
rect 31164 35646 31166 35698
rect 31218 35646 31614 35698
rect 31666 35646 31668 35698
rect 31164 35644 31668 35646
rect 31164 35634 31220 35644
rect 31612 35634 31668 35644
rect 31276 35474 31332 35486
rect 31276 35422 31278 35474
rect 31330 35422 31332 35474
rect 31276 34914 31332 35422
rect 31276 34862 31278 34914
rect 31330 34862 31332 34914
rect 31276 34692 31332 34862
rect 31500 34916 31556 34954
rect 31500 34850 31556 34860
rect 31276 34626 31332 34636
rect 31500 34690 31556 34702
rect 31500 34638 31502 34690
rect 31554 34638 31556 34690
rect 31500 34580 31556 34638
rect 31724 34692 31780 38780
rect 31836 38770 31892 38780
rect 31948 38722 32004 38734
rect 31948 38670 31950 38722
rect 32002 38670 32004 38722
rect 31948 37716 32004 38670
rect 32060 38668 32116 39678
rect 32172 39620 32228 41132
rect 32508 41186 32564 41356
rect 32956 41580 33348 41636
rect 32956 41410 33012 41580
rect 32956 41358 32958 41410
rect 33010 41358 33012 41410
rect 32956 41346 33012 41358
rect 32508 41134 32510 41186
rect 32562 41134 32564 41186
rect 32508 41122 32564 41134
rect 32396 41074 32452 41086
rect 32396 41022 32398 41074
rect 32450 41022 32452 41074
rect 32396 40964 32452 41022
rect 33404 40964 33460 40974
rect 32396 40962 33460 40964
rect 32396 40910 33406 40962
rect 33458 40910 33460 40962
rect 32396 40908 33460 40910
rect 33068 40404 33124 40414
rect 32844 40402 33124 40404
rect 32844 40350 33070 40402
rect 33122 40350 33124 40402
rect 32844 40348 33124 40350
rect 32284 39844 32340 39854
rect 32844 39844 32900 40348
rect 33068 40338 33124 40348
rect 32284 39842 32900 39844
rect 32284 39790 32286 39842
rect 32338 39790 32846 39842
rect 32898 39790 32900 39842
rect 32284 39788 32900 39790
rect 32284 39778 32340 39788
rect 32844 39778 32900 39788
rect 32620 39620 32676 39630
rect 32172 39564 32340 39620
rect 32284 38668 32340 39564
rect 32620 39526 32676 39564
rect 33180 39396 33236 39406
rect 33068 39394 33236 39396
rect 33068 39342 33182 39394
rect 33234 39342 33236 39394
rect 33068 39340 33236 39342
rect 32060 38612 32228 38668
rect 32284 38612 32452 38668
rect 31948 36484 32004 37660
rect 32060 37492 32116 37502
rect 32060 37398 32116 37436
rect 31948 36428 32116 36484
rect 31948 36260 32004 36270
rect 31836 35810 31892 35822
rect 31836 35758 31838 35810
rect 31890 35758 31892 35810
rect 31836 35476 31892 35758
rect 31836 35410 31892 35420
rect 31948 35698 32004 36204
rect 31948 35646 31950 35698
rect 32002 35646 32004 35698
rect 31948 35252 32004 35646
rect 31948 35186 32004 35196
rect 31836 34916 31892 34926
rect 31836 34914 32004 34916
rect 31836 34862 31838 34914
rect 31890 34862 32004 34914
rect 31836 34860 32004 34862
rect 31836 34850 31892 34860
rect 31948 34804 32004 34860
rect 31948 34738 32004 34748
rect 31724 34636 31892 34692
rect 31500 34524 31780 34580
rect 31500 34356 31556 34366
rect 31052 34354 31556 34356
rect 31052 34302 31502 34354
rect 31554 34302 31556 34354
rect 31052 34300 31556 34302
rect 31052 34242 31108 34300
rect 31500 34290 31556 34300
rect 31052 34190 31054 34242
rect 31106 34190 31108 34242
rect 31052 34178 31108 34190
rect 31388 34130 31444 34142
rect 31388 34078 31390 34130
rect 31442 34078 31444 34130
rect 31388 34020 31444 34078
rect 31612 34132 31668 34142
rect 31612 34038 31668 34076
rect 31388 33954 31444 33964
rect 31052 33796 31108 33806
rect 30940 33740 31052 33796
rect 31052 33730 31108 33740
rect 31052 33572 31108 33582
rect 31052 32786 31108 33516
rect 31724 32900 31780 34524
rect 31836 33460 31892 34636
rect 32060 34356 32116 36428
rect 32172 35140 32228 38612
rect 32396 37380 32452 38612
rect 32732 38050 32788 38062
rect 32732 37998 32734 38050
rect 32786 37998 32788 38050
rect 32396 37286 32452 37324
rect 32508 37492 32564 37502
rect 32508 37378 32564 37436
rect 32508 37326 32510 37378
rect 32562 37326 32564 37378
rect 32508 37314 32564 37326
rect 32396 37044 32452 37054
rect 32732 37044 32788 37998
rect 33068 37268 33124 39340
rect 33180 39330 33236 39340
rect 33404 39284 33460 40908
rect 33404 38052 33460 39228
rect 33516 39394 33572 39406
rect 33516 39342 33518 39394
rect 33570 39342 33572 39394
rect 33516 38276 33572 39342
rect 33740 38668 33796 43652
rect 34188 43650 34468 43652
rect 34188 43598 34414 43650
rect 34466 43598 34468 43650
rect 34188 43596 34468 43598
rect 34188 42754 34244 43596
rect 34412 43586 34468 43596
rect 34300 43428 34356 43438
rect 34300 43334 34356 43372
rect 34636 43316 34692 43326
rect 34412 43260 34636 43316
rect 34412 42980 34468 43260
rect 34636 43222 34692 43260
rect 34412 42886 34468 42924
rect 34748 43092 34804 43102
rect 34748 42978 34804 43036
rect 34748 42926 34750 42978
rect 34802 42926 34804 42978
rect 34188 42702 34190 42754
rect 34242 42702 34244 42754
rect 34188 42420 34244 42702
rect 34188 42354 34244 42364
rect 34076 41860 34132 41870
rect 33852 41858 34132 41860
rect 33852 41806 34078 41858
rect 34130 41806 34132 41858
rect 33852 41804 34132 41806
rect 33852 40290 33908 41804
rect 34076 41794 34132 41804
rect 33964 40404 34020 40414
rect 34020 40348 34132 40404
rect 33964 40310 34020 40348
rect 33852 40238 33854 40290
rect 33906 40238 33908 40290
rect 33852 39842 33908 40238
rect 33852 39790 33854 39842
rect 33906 39790 33908 39842
rect 33852 39778 33908 39790
rect 34076 39730 34132 40348
rect 34076 39678 34078 39730
rect 34130 39678 34132 39730
rect 34076 39666 34132 39678
rect 33516 38210 33572 38220
rect 33628 38612 33796 38668
rect 34748 38724 34804 42926
rect 34972 42754 35028 43652
rect 35644 43652 36708 43708
rect 37324 44098 37380 44110
rect 37324 44046 37326 44098
rect 37378 44046 37380 44098
rect 34972 42702 34974 42754
rect 35026 42702 35028 42754
rect 34972 42690 35028 42702
rect 35084 43426 35140 43438
rect 35084 43374 35086 43426
rect 35138 43374 35140 43426
rect 35084 41972 35140 43374
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 35308 42644 35364 42654
rect 35308 42550 35364 42588
rect 35196 42532 35252 42542
rect 35196 42438 35252 42476
rect 35084 41906 35140 41916
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 35084 40516 35140 40526
rect 35084 40422 35140 40460
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 35196 39396 35252 39406
rect 35196 39060 35252 39340
rect 34972 39004 35252 39060
rect 34748 38722 34916 38724
rect 34748 38670 34750 38722
rect 34802 38670 34916 38722
rect 34748 38668 34916 38670
rect 34748 38658 34804 38668
rect 33628 38052 33684 38612
rect 34524 38610 34580 38622
rect 34524 38558 34526 38610
rect 34578 38558 34580 38610
rect 33404 37986 33460 37996
rect 33516 38050 33684 38052
rect 33516 37998 33630 38050
rect 33682 37998 33684 38050
rect 33516 37996 33684 37998
rect 33292 37940 33348 37950
rect 33292 37846 33348 37884
rect 33180 37826 33236 37838
rect 33180 37774 33182 37826
rect 33234 37774 33236 37826
rect 33180 37380 33236 37774
rect 33404 37826 33460 37838
rect 33404 37774 33406 37826
rect 33458 37774 33460 37826
rect 33292 37380 33348 37390
rect 33180 37324 33292 37380
rect 33292 37314 33348 37324
rect 33404 37268 33460 37774
rect 33068 37212 33236 37268
rect 32396 37042 32732 37044
rect 32396 36990 32398 37042
rect 32450 36990 32732 37042
rect 32396 36988 32732 36990
rect 32396 36482 32452 36988
rect 32732 36950 32788 36988
rect 33068 37042 33124 37054
rect 33068 36990 33070 37042
rect 33122 36990 33124 37042
rect 32396 36430 32398 36482
rect 32450 36430 32452 36482
rect 32396 36418 32452 36430
rect 32732 36484 32788 36494
rect 33068 36484 33124 36990
rect 32732 36482 33124 36484
rect 32732 36430 32734 36482
rect 32786 36430 33124 36482
rect 32732 36428 33124 36430
rect 32732 36418 32788 36428
rect 32396 35586 32452 35598
rect 32396 35534 32398 35586
rect 32450 35534 32452 35586
rect 32396 35476 32452 35534
rect 32396 35410 32452 35420
rect 32172 35074 32228 35084
rect 32396 34916 32452 34926
rect 32396 34822 32452 34860
rect 32732 34914 32788 34926
rect 32732 34862 32734 34914
rect 32786 34862 32788 34914
rect 32284 34804 32340 34814
rect 32284 34710 32340 34748
rect 32172 34692 32228 34702
rect 32172 34598 32228 34636
rect 32060 34300 32228 34356
rect 32060 34130 32116 34142
rect 32060 34078 32062 34130
rect 32114 34078 32116 34130
rect 32060 33572 32116 34078
rect 32060 33506 32116 33516
rect 31836 33366 31892 33404
rect 32060 33348 32116 33358
rect 32172 33348 32228 34300
rect 32732 33572 32788 34862
rect 33180 34914 33236 37212
rect 33404 37174 33460 37212
rect 33516 36482 33572 37996
rect 33628 37986 33684 37996
rect 33740 38164 33796 38174
rect 33628 37380 33684 37390
rect 33628 37286 33684 37324
rect 33740 36932 33796 38108
rect 33964 38050 34020 38062
rect 33964 37998 33966 38050
rect 34018 37998 34020 38050
rect 33964 37940 34020 37998
rect 33964 37874 34020 37884
rect 34300 37940 34356 37950
rect 34300 37938 34468 37940
rect 34300 37886 34302 37938
rect 34354 37886 34468 37938
rect 34300 37884 34468 37886
rect 34300 37874 34356 37884
rect 33852 37828 33908 37838
rect 33852 37734 33908 37772
rect 34412 37490 34468 37884
rect 34412 37438 34414 37490
rect 34466 37438 34468 37490
rect 34412 37426 34468 37438
rect 34300 37380 34356 37390
rect 34300 37266 34356 37324
rect 34300 37214 34302 37266
rect 34354 37214 34356 37266
rect 34300 37202 34356 37214
rect 34524 37268 34580 38558
rect 34860 38050 34916 38668
rect 34860 37998 34862 38050
rect 34914 37998 34916 38050
rect 34860 37986 34916 37998
rect 34972 38052 35028 39004
rect 35084 38834 35140 38846
rect 35084 38782 35086 38834
rect 35138 38782 35140 38834
rect 35084 38668 35140 38782
rect 35196 38834 35252 39004
rect 35196 38782 35198 38834
rect 35250 38782 35252 38834
rect 35196 38770 35252 38782
rect 35644 38668 35700 43652
rect 35868 43540 35924 43550
rect 35868 43446 35924 43484
rect 37212 43538 37268 43550
rect 37212 43486 37214 43538
rect 37266 43486 37268 43538
rect 37100 43426 37156 43438
rect 37100 43374 37102 43426
rect 37154 43374 37156 43426
rect 37100 42978 37156 43374
rect 37100 42926 37102 42978
rect 37154 42926 37156 42978
rect 37100 42914 37156 42926
rect 37212 42980 37268 43486
rect 37212 42914 37268 42924
rect 37324 43540 37380 44046
rect 37212 42756 37268 42766
rect 37100 42530 37156 42542
rect 37100 42478 37102 42530
rect 37154 42478 37156 42530
rect 36540 41860 36596 41870
rect 36540 41300 36596 41804
rect 36204 41188 36260 41198
rect 36204 41094 36260 41132
rect 36428 40964 36484 40974
rect 36428 40870 36484 40908
rect 36540 40740 36596 41244
rect 35756 40684 36372 40740
rect 35756 40402 35812 40684
rect 36316 40626 36372 40684
rect 36316 40574 36318 40626
rect 36370 40574 36372 40626
rect 36316 40562 36372 40574
rect 36428 40684 36596 40740
rect 36764 40964 36820 40974
rect 35756 40350 35758 40402
rect 35810 40350 35812 40402
rect 35756 40338 35812 40350
rect 35868 40290 35924 40302
rect 35868 40238 35870 40290
rect 35922 40238 35924 40290
rect 35868 39842 35924 40238
rect 35868 39790 35870 39842
rect 35922 39790 35924 39842
rect 35868 39778 35924 39790
rect 35980 39620 36036 39630
rect 36428 39620 36484 40684
rect 36540 40514 36596 40526
rect 36540 40462 36542 40514
rect 36594 40462 36596 40514
rect 36540 40292 36596 40462
rect 36652 40516 36708 40526
rect 36764 40516 36820 40908
rect 37100 40628 37156 42478
rect 37212 41188 37268 42700
rect 37324 41972 37380 43484
rect 37436 43316 37492 44942
rect 37548 44996 37604 45614
rect 37548 44930 37604 44940
rect 37660 45666 37940 45668
rect 37660 45614 37886 45666
rect 37938 45614 37940 45666
rect 37660 45612 37940 45614
rect 37660 44436 37716 45612
rect 37884 45602 37940 45612
rect 38668 45668 38724 45838
rect 39004 45780 39060 49200
rect 39676 46228 39732 49200
rect 40348 46340 40404 49200
rect 40348 46284 40628 46340
rect 39676 46172 40516 46228
rect 39004 45714 39060 45724
rect 40012 45890 40068 45902
rect 40012 45838 40014 45890
rect 40066 45838 40068 45890
rect 40012 45780 40068 45838
rect 40012 45714 40068 45724
rect 40460 45890 40516 46172
rect 40460 45838 40462 45890
rect 40514 45838 40516 45890
rect 38892 45668 38948 45678
rect 38668 45602 38724 45612
rect 38780 45666 38948 45668
rect 38780 45614 38894 45666
rect 38946 45614 38948 45666
rect 38780 45612 38948 45614
rect 38220 45106 38276 45118
rect 38220 45054 38222 45106
rect 38274 45054 38276 45106
rect 38108 44996 38164 45006
rect 37548 44380 38052 44436
rect 37548 44212 37604 44380
rect 37548 44118 37604 44156
rect 37660 44210 37716 44222
rect 37660 44158 37662 44210
rect 37714 44158 37716 44210
rect 37660 43540 37716 44158
rect 37660 43474 37716 43484
rect 37772 43650 37828 43662
rect 37772 43598 37774 43650
rect 37826 43598 37828 43650
rect 37436 42756 37492 43260
rect 37548 42756 37604 42766
rect 37436 42754 37604 42756
rect 37436 42702 37550 42754
rect 37602 42702 37604 42754
rect 37436 42700 37604 42702
rect 37548 42690 37604 42700
rect 37772 42756 37828 43598
rect 37772 42690 37828 42700
rect 37660 42532 37716 42542
rect 37548 42530 37716 42532
rect 37548 42478 37662 42530
rect 37714 42478 37716 42530
rect 37548 42476 37716 42478
rect 37548 42420 37604 42476
rect 37660 42466 37716 42476
rect 37884 42530 37940 42542
rect 37884 42478 37886 42530
rect 37938 42478 37940 42530
rect 37548 42082 37604 42364
rect 37548 42030 37550 42082
rect 37602 42030 37604 42082
rect 37548 42018 37604 42030
rect 37436 41972 37492 41982
rect 37324 41970 37492 41972
rect 37324 41918 37438 41970
rect 37490 41918 37492 41970
rect 37324 41916 37492 41918
rect 37436 41906 37492 41916
rect 37660 41970 37716 41982
rect 37660 41918 37662 41970
rect 37714 41918 37716 41970
rect 37660 41298 37716 41918
rect 37884 41636 37940 42478
rect 37884 41570 37940 41580
rect 37660 41246 37662 41298
rect 37714 41246 37716 41298
rect 37660 41234 37716 41246
rect 37772 41300 37828 41310
rect 37324 41188 37380 41198
rect 37212 41132 37324 41188
rect 37324 41094 37380 41132
rect 37772 41186 37828 41244
rect 37772 41134 37774 41186
rect 37826 41134 37828 41186
rect 37772 41122 37828 41134
rect 37548 41076 37604 41086
rect 37436 41020 37548 41076
rect 37324 40628 37380 40638
rect 37436 40628 37492 41020
rect 37548 40982 37604 41020
rect 37884 40964 37940 40974
rect 37884 40740 37940 40908
rect 37100 40626 37492 40628
rect 37100 40574 37326 40626
rect 37378 40574 37492 40626
rect 37100 40572 37492 40574
rect 37548 40684 37940 40740
rect 37324 40562 37380 40572
rect 36988 40516 37044 40526
rect 36652 40514 36932 40516
rect 36652 40462 36654 40514
rect 36706 40462 36932 40514
rect 36652 40460 36932 40462
rect 36652 40450 36708 40460
rect 36876 40292 36932 40460
rect 36988 40514 37156 40516
rect 36988 40462 36990 40514
rect 37042 40462 37156 40514
rect 36988 40460 37156 40462
rect 36988 40450 37044 40460
rect 37100 40292 37156 40460
rect 37548 40404 37604 40684
rect 37996 40628 38052 44380
rect 38108 43650 38164 44940
rect 38220 44212 38276 45054
rect 38220 44146 38276 44156
rect 38108 43598 38110 43650
rect 38162 43598 38164 43650
rect 38108 43586 38164 43598
rect 38444 43650 38500 43662
rect 38444 43598 38446 43650
rect 38498 43598 38500 43650
rect 38332 41188 38388 41198
rect 38332 41094 38388 41132
rect 38444 41076 38500 43598
rect 38780 43538 38836 45612
rect 38892 45602 38948 45612
rect 39788 45666 39844 45678
rect 39788 45614 39790 45666
rect 39842 45614 39844 45666
rect 39564 45108 39620 45118
rect 39564 45014 39620 45052
rect 39116 44994 39172 45006
rect 39116 44942 39118 44994
rect 39170 44942 39172 44994
rect 39116 44548 39172 44942
rect 38892 44492 39508 44548
rect 38892 44322 38948 44492
rect 38892 44270 38894 44322
rect 38946 44270 38948 44322
rect 38892 44258 38948 44270
rect 39116 44322 39172 44334
rect 39116 44270 39118 44322
rect 39170 44270 39172 44322
rect 39116 44212 39172 44270
rect 39340 44212 39396 44222
rect 39116 44146 39172 44156
rect 39228 44210 39396 44212
rect 39228 44158 39342 44210
rect 39394 44158 39396 44210
rect 39228 44156 39396 44158
rect 38780 43486 38782 43538
rect 38834 43486 38836 43538
rect 38780 43316 38836 43486
rect 39116 43316 39172 43326
rect 38780 43260 39116 43316
rect 39116 43250 39172 43260
rect 39004 42980 39060 42990
rect 39004 42754 39060 42924
rect 39228 42756 39284 44156
rect 39340 44146 39396 44156
rect 39340 43764 39396 43774
rect 39452 43764 39508 44492
rect 39676 44324 39732 44334
rect 39676 44230 39732 44268
rect 39340 43762 39508 43764
rect 39340 43710 39342 43762
rect 39394 43710 39508 43762
rect 39340 43708 39508 43710
rect 39788 43708 39844 45614
rect 40236 45218 40292 45230
rect 40236 45166 40238 45218
rect 40290 45166 40292 45218
rect 40236 45108 40292 45166
rect 40236 45042 40292 45052
rect 40348 45106 40404 45118
rect 40348 45054 40350 45106
rect 40402 45054 40404 45106
rect 40348 44996 40404 45054
rect 40348 44930 40404 44940
rect 40236 44884 40292 44894
rect 40236 44790 40292 44828
rect 40348 44772 40404 44782
rect 40348 44322 40404 44716
rect 40348 44270 40350 44322
rect 40402 44270 40404 44322
rect 40348 44258 40404 44270
rect 40236 44212 40292 44222
rect 40012 44098 40068 44110
rect 40012 44046 40014 44098
rect 40066 44046 40068 44098
rect 40012 43708 40068 44046
rect 39340 43698 39396 43708
rect 39004 42702 39006 42754
rect 39058 42702 39060 42754
rect 39004 42690 39060 42702
rect 39116 42700 39284 42756
rect 39564 43652 39844 43708
rect 39900 43652 40068 43708
rect 40124 43652 40180 43662
rect 39564 43650 39620 43652
rect 39564 43598 39566 43650
rect 39618 43598 39620 43650
rect 38556 41970 38612 41982
rect 38556 41918 38558 41970
rect 38610 41918 38612 41970
rect 38556 41410 38612 41918
rect 38556 41358 38558 41410
rect 38610 41358 38612 41410
rect 38556 41346 38612 41358
rect 39004 41186 39060 41198
rect 39004 41134 39006 41186
rect 39058 41134 39060 41186
rect 38556 41076 38612 41086
rect 38444 41020 38556 41076
rect 38556 40982 38612 41020
rect 39004 40964 39060 41134
rect 39004 40898 39060 40908
rect 37772 40626 38052 40628
rect 37772 40574 37998 40626
rect 38050 40574 38052 40626
rect 37772 40572 38052 40574
rect 36540 40236 36708 40292
rect 36876 40236 37044 40292
rect 35980 39618 36484 39620
rect 35980 39566 35982 39618
rect 36034 39566 36430 39618
rect 36482 39566 36484 39618
rect 35980 39564 36484 39566
rect 35980 39554 36036 39564
rect 36428 39554 36484 39564
rect 36540 40068 36596 40078
rect 35868 39508 35924 39518
rect 35868 39414 35924 39452
rect 36540 39508 36596 40012
rect 36540 38948 36596 39452
rect 36428 38892 36596 38948
rect 36652 39732 36708 40236
rect 36652 38948 36708 39676
rect 36988 39620 37044 40236
rect 37100 39844 37156 40236
rect 37100 39778 37156 39788
rect 37324 40348 37604 40404
rect 37660 40514 37716 40526
rect 37660 40462 37662 40514
rect 37714 40462 37716 40514
rect 37660 40404 37716 40462
rect 36988 39554 37044 39564
rect 37324 39506 37380 40348
rect 37660 40338 37716 40348
rect 37772 40180 37828 40572
rect 37996 40562 38052 40572
rect 39116 40404 39172 42700
rect 39340 42644 39396 42654
rect 39340 42550 39396 42588
rect 39228 42530 39284 42542
rect 39228 42478 39230 42530
rect 39282 42478 39284 42530
rect 39228 42420 39284 42478
rect 39564 42420 39620 43598
rect 39228 42364 39620 42420
rect 39452 42082 39508 42094
rect 39452 42030 39454 42082
rect 39506 42030 39508 42082
rect 39452 41300 39508 42030
rect 39564 41972 39620 42364
rect 39676 43538 39732 43550
rect 39676 43486 39678 43538
rect 39730 43486 39732 43538
rect 39676 42420 39732 43486
rect 39788 43428 39844 43438
rect 39788 42532 39844 43372
rect 39900 42756 39956 43652
rect 40124 43558 40180 43596
rect 40012 43538 40068 43550
rect 40012 43486 40014 43538
rect 40066 43486 40068 43538
rect 40012 43316 40068 43486
rect 40012 43250 40068 43260
rect 40124 43316 40180 43326
rect 40236 43316 40292 44156
rect 40124 43314 40292 43316
rect 40124 43262 40126 43314
rect 40178 43262 40292 43314
rect 40124 43260 40292 43262
rect 40348 43652 40404 43662
rect 40124 43250 40180 43260
rect 39900 42700 40068 42756
rect 39900 42532 39956 42542
rect 39788 42530 39956 42532
rect 39788 42478 39902 42530
rect 39954 42478 39956 42530
rect 39788 42476 39956 42478
rect 39676 42354 39732 42364
rect 39900 42308 39956 42476
rect 39900 42242 39956 42252
rect 39676 41972 39732 41982
rect 39564 41970 39732 41972
rect 39564 41918 39678 41970
rect 39730 41918 39732 41970
rect 39564 41916 39732 41918
rect 39676 41906 39732 41916
rect 39788 41636 39844 41646
rect 39844 41580 39956 41636
rect 39788 41570 39844 41580
rect 39452 41188 39508 41244
rect 39788 41188 39844 41198
rect 39452 41186 39844 41188
rect 39452 41134 39790 41186
rect 39842 41134 39844 41186
rect 39452 41132 39844 41134
rect 39788 40628 39844 41132
rect 39788 40562 39844 40572
rect 39116 40348 39620 40404
rect 37436 40124 37828 40180
rect 37436 39618 37492 40124
rect 37436 39566 37438 39618
rect 37490 39566 37492 39618
rect 37436 39554 37492 39566
rect 37324 39454 37326 39506
rect 37378 39454 37380 39506
rect 37324 39442 37380 39454
rect 35084 38612 35588 38668
rect 35644 38612 35924 38668
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 35084 38052 35140 38062
rect 34972 38050 35140 38052
rect 34972 37998 35086 38050
rect 35138 37998 35140 38050
rect 34972 37996 35140 37998
rect 35084 37986 35140 37996
rect 35532 38050 35588 38612
rect 35532 37998 35534 38050
rect 35586 37998 35588 38050
rect 34524 37174 34580 37212
rect 34972 37826 35028 37838
rect 34972 37774 34974 37826
rect 35026 37774 35028 37826
rect 34076 37044 34132 37054
rect 34076 36950 34132 36988
rect 33516 36430 33518 36482
rect 33570 36430 33572 36482
rect 33516 36418 33572 36430
rect 33628 36876 33796 36932
rect 33628 35924 33684 36876
rect 33516 35868 33684 35924
rect 33740 36706 33796 36718
rect 33740 36654 33742 36706
rect 33794 36654 33796 36706
rect 33740 35924 33796 36654
rect 34972 36036 35028 37774
rect 35532 37378 35588 37998
rect 35532 37326 35534 37378
rect 35586 37326 35588 37378
rect 35532 37314 35588 37326
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35644 36820 35700 36830
rect 35196 36810 35460 36820
rect 34972 35970 35028 35980
rect 35532 36764 35644 36820
rect 33740 35922 34244 35924
rect 33740 35870 33742 35922
rect 33794 35870 34244 35922
rect 33740 35868 34244 35870
rect 33404 35140 33460 35150
rect 33404 35046 33460 35084
rect 33180 34862 33182 34914
rect 33234 34862 33236 34914
rect 33180 34850 33236 34862
rect 33516 34804 33572 35868
rect 33740 35858 33796 35868
rect 34188 35812 34244 35868
rect 35420 35812 35476 35822
rect 35532 35812 35588 36764
rect 35644 36754 35700 36764
rect 34188 35810 35140 35812
rect 34188 35758 34190 35810
rect 34242 35758 35140 35810
rect 34188 35756 35140 35758
rect 34188 35746 34244 35756
rect 33628 35698 33684 35710
rect 33628 35646 33630 35698
rect 33682 35646 33684 35698
rect 33628 35588 33684 35646
rect 33964 35700 34020 35710
rect 33964 35698 34132 35700
rect 33964 35646 33966 35698
rect 34018 35646 34132 35698
rect 33964 35644 34132 35646
rect 33964 35634 34020 35644
rect 33628 35522 33684 35532
rect 33964 35140 34020 35150
rect 34076 35140 34132 35644
rect 35084 35698 35140 35756
rect 35084 35646 35086 35698
rect 35138 35646 35140 35698
rect 35084 35634 35140 35646
rect 35420 35810 35588 35812
rect 35420 35758 35422 35810
rect 35474 35758 35588 35810
rect 35420 35756 35588 35758
rect 34412 35588 34468 35598
rect 34412 35494 34468 35532
rect 35420 35588 35476 35756
rect 35420 35522 35476 35532
rect 34748 35474 34804 35486
rect 34748 35422 34750 35474
rect 34802 35422 34804 35474
rect 34076 35084 34580 35140
rect 33628 35028 33684 35038
rect 33628 34934 33684 34972
rect 33740 34804 33796 34814
rect 33516 34748 33684 34804
rect 33628 34244 33684 34748
rect 33740 34802 33908 34804
rect 33740 34750 33742 34802
rect 33794 34750 33908 34802
rect 33740 34748 33908 34750
rect 33740 34738 33796 34748
rect 33740 34244 33796 34254
rect 33628 34188 33740 34244
rect 33740 34150 33796 34188
rect 33628 33796 33684 33806
rect 32732 33506 32788 33516
rect 33516 33572 33572 33582
rect 32844 33460 32900 33470
rect 32060 33346 32788 33348
rect 32060 33294 32062 33346
rect 32114 33294 32788 33346
rect 32060 33292 32788 33294
rect 32060 33282 32116 33292
rect 32396 33122 32452 33134
rect 32396 33070 32398 33122
rect 32450 33070 32452 33122
rect 31724 32844 32228 32900
rect 31052 32734 31054 32786
rect 31106 32734 31108 32786
rect 31052 32722 31108 32734
rect 31724 32732 32116 32788
rect 30604 31938 30660 31948
rect 30716 32562 30772 32574
rect 30716 32510 30718 32562
rect 30770 32510 30772 32562
rect 30044 31826 30100 31836
rect 30044 31556 30100 31566
rect 30380 31556 30436 31566
rect 30716 31556 30772 32510
rect 30100 31554 30772 31556
rect 30100 31502 30382 31554
rect 30434 31502 30772 31554
rect 30100 31500 30772 31502
rect 30940 32452 30996 32462
rect 30940 31778 30996 32396
rect 31724 32452 31780 32732
rect 32060 32674 32116 32732
rect 32060 32622 32062 32674
rect 32114 32622 32116 32674
rect 32060 32610 32116 32622
rect 31724 32358 31780 32396
rect 31836 32564 31892 32574
rect 30940 31726 30942 31778
rect 30994 31726 30996 31778
rect 30044 31218 30100 31500
rect 30380 31490 30436 31500
rect 30044 31166 30046 31218
rect 30098 31166 30100 31218
rect 30044 31154 30100 31166
rect 29932 30322 29988 30716
rect 29932 30270 29934 30322
rect 29986 30270 29988 30322
rect 29932 30100 29988 30270
rect 29932 29652 29988 30044
rect 29932 29586 29988 29596
rect 30044 30996 30100 31006
rect 30044 29650 30100 30940
rect 30492 30882 30548 30894
rect 30492 30830 30494 30882
rect 30546 30830 30548 30882
rect 30492 30436 30548 30830
rect 30492 30342 30548 30380
rect 30268 30100 30324 30110
rect 30268 30006 30324 30044
rect 30828 29988 30884 29998
rect 30044 29598 30046 29650
rect 30098 29598 30100 29650
rect 30044 29586 30100 29598
rect 30380 29986 30884 29988
rect 30380 29934 30830 29986
rect 30882 29934 30884 29986
rect 30380 29932 30884 29934
rect 30380 29650 30436 29932
rect 30380 29598 30382 29650
rect 30434 29598 30436 29650
rect 30380 29586 30436 29598
rect 30716 28980 30772 29932
rect 30828 29922 30884 29932
rect 30828 29540 30884 29550
rect 30940 29540 30996 31726
rect 31388 31778 31444 31790
rect 31388 31726 31390 31778
rect 31442 31726 31444 31778
rect 31388 30996 31444 31726
rect 31388 30930 31444 30940
rect 31836 31778 31892 32508
rect 32060 32452 32116 32462
rect 32060 32358 32116 32396
rect 32172 32228 32228 32844
rect 32284 32562 32340 32574
rect 32284 32510 32286 32562
rect 32338 32510 32340 32562
rect 32284 32340 32340 32510
rect 32396 32340 32452 33070
rect 32620 33122 32676 33134
rect 32620 33070 32622 33122
rect 32674 33070 32676 33122
rect 32620 32562 32676 33070
rect 32732 33012 32788 33292
rect 32844 33234 32900 33404
rect 32844 33182 32846 33234
rect 32898 33182 32900 33234
rect 32844 33170 32900 33182
rect 32956 33234 33012 33246
rect 32956 33182 32958 33234
rect 33010 33182 33012 33234
rect 32956 33012 33012 33182
rect 32732 32956 33012 33012
rect 32620 32510 32622 32562
rect 32674 32510 32676 32562
rect 32620 32498 32676 32510
rect 33180 32452 33236 32462
rect 32732 32450 33236 32452
rect 32732 32398 33182 32450
rect 33234 32398 33236 32450
rect 32732 32396 33236 32398
rect 32732 32340 32788 32396
rect 33180 32386 33236 32396
rect 32284 32284 32788 32340
rect 33516 32340 33572 33516
rect 33628 32562 33684 33740
rect 33628 32510 33630 32562
rect 33682 32510 33684 32562
rect 33628 32498 33684 32510
rect 33628 32340 33684 32350
rect 33516 32284 33628 32340
rect 32172 32172 32452 32228
rect 31836 31726 31838 31778
rect 31890 31726 31892 31778
rect 31836 30882 31892 31726
rect 31836 30830 31838 30882
rect 31890 30830 31892 30882
rect 31836 30772 31892 30830
rect 31388 30716 31892 30772
rect 32284 30996 32340 31006
rect 30884 29484 30996 29540
rect 31276 30212 31332 30222
rect 31388 30212 31444 30716
rect 32284 30436 32340 30940
rect 32284 30370 32340 30380
rect 32396 30434 32452 32172
rect 33292 32004 33348 32014
rect 33180 31890 33236 31902
rect 33180 31838 33182 31890
rect 33234 31838 33236 31890
rect 32508 31108 32564 31118
rect 32508 31014 32564 31052
rect 32396 30382 32398 30434
rect 32450 30382 32452 30434
rect 32396 30370 32452 30382
rect 31612 30324 31668 30334
rect 31612 30230 31668 30268
rect 31276 30210 31444 30212
rect 31276 30158 31278 30210
rect 31330 30158 31444 30210
rect 31276 30156 31444 30158
rect 32060 30212 32116 30222
rect 30828 29474 30884 29484
rect 30044 28868 30100 28878
rect 29820 28866 30100 28868
rect 29820 28814 30046 28866
rect 30098 28814 30100 28866
rect 29820 28812 30100 28814
rect 30044 28802 30100 28812
rect 29708 28702 29710 28754
rect 29762 28702 29764 28754
rect 29708 28690 29764 28702
rect 30380 28644 30436 28654
rect 30268 28588 30380 28644
rect 30156 28420 30212 28430
rect 30156 28326 30212 28364
rect 29260 27186 29428 27188
rect 29260 27134 29262 27186
rect 29314 27134 29428 27186
rect 29260 27132 29428 27134
rect 29484 28308 29540 28318
rect 29484 27188 29540 28252
rect 30268 28196 30324 28588
rect 30380 28550 30436 28588
rect 30716 28530 30772 28924
rect 31052 29092 31108 29102
rect 30828 28644 30884 28654
rect 30828 28550 30884 28588
rect 31052 28642 31108 29036
rect 31052 28590 31054 28642
rect 31106 28590 31108 28642
rect 31052 28578 31108 28590
rect 30716 28478 30718 28530
rect 30770 28478 30772 28530
rect 30716 28466 30772 28478
rect 30156 28140 30324 28196
rect 29260 27122 29316 27132
rect 28924 26852 28980 26862
rect 29036 26852 29428 26908
rect 27244 23940 27300 23950
rect 27244 23846 27300 23884
rect 27020 22540 27188 22596
rect 27244 22932 27300 22942
rect 27020 21812 27076 22540
rect 27244 22370 27300 22876
rect 27244 22318 27246 22370
rect 27298 22318 27300 22370
rect 27244 22306 27300 22318
rect 27356 22148 27412 23996
rect 27692 23828 27748 25228
rect 27804 24948 27860 24958
rect 27804 24612 27860 24892
rect 28028 24948 28084 24958
rect 28028 24834 28084 24892
rect 28028 24782 28030 24834
rect 28082 24782 28084 24834
rect 27916 24724 27972 24734
rect 27916 24630 27972 24668
rect 27804 23938 27860 24556
rect 28028 24164 28084 24782
rect 28028 24098 28084 24108
rect 27804 23886 27806 23938
rect 27858 23886 27860 23938
rect 27804 23874 27860 23886
rect 27468 23772 27692 23828
rect 27468 22258 27524 23772
rect 27692 23762 27748 23772
rect 27468 22206 27470 22258
rect 27522 22206 27524 22258
rect 27468 22194 27524 22206
rect 27020 21746 27076 21756
rect 27132 22092 27412 22148
rect 28140 22148 28196 26460
rect 28364 26402 28420 26852
rect 28588 26740 28644 26852
rect 28364 26350 28366 26402
rect 28418 26350 28420 26402
rect 28252 26290 28308 26302
rect 28252 26238 28254 26290
rect 28306 26238 28308 26290
rect 28252 25956 28308 26238
rect 28252 25890 28308 25900
rect 28252 25396 28308 25406
rect 28252 25302 28308 25340
rect 28364 25284 28420 26350
rect 28364 25218 28420 25228
rect 28476 26684 28644 26740
rect 28476 25060 28532 26684
rect 28924 26514 28980 26796
rect 28924 26462 28926 26514
rect 28978 26462 28980 26514
rect 28588 26404 28644 26414
rect 28588 26310 28644 26348
rect 28924 25620 28980 26462
rect 29148 26516 29204 26526
rect 29148 26422 29204 26460
rect 29260 26404 29316 26414
rect 29260 26310 29316 26348
rect 28924 25554 28980 25564
rect 29036 26068 29092 26078
rect 28588 25284 28644 25322
rect 28588 25218 28644 25228
rect 28252 25004 28532 25060
rect 28588 25060 28644 25070
rect 28252 22372 28308 25004
rect 28588 24722 28644 25004
rect 28812 24836 28868 24846
rect 28812 24742 28868 24780
rect 28588 24670 28590 24722
rect 28642 24670 28644 24722
rect 28588 24658 28644 24670
rect 28588 24052 28644 24062
rect 28364 23714 28420 23726
rect 28364 23662 28366 23714
rect 28418 23662 28420 23714
rect 28364 23604 28420 23662
rect 28364 23538 28420 23548
rect 28588 22708 28644 23996
rect 29036 23604 29092 26012
rect 29372 25506 29428 26852
rect 29372 25454 29374 25506
rect 29426 25454 29428 25506
rect 29372 25442 29428 25454
rect 29484 26402 29540 27132
rect 29932 27970 29988 27982
rect 29932 27918 29934 27970
rect 29986 27918 29988 27970
rect 29596 27076 29652 27086
rect 29596 26982 29652 27020
rect 29932 27076 29988 27918
rect 30156 27858 30212 28140
rect 30940 28084 30996 28094
rect 30156 27806 30158 27858
rect 30210 27806 30212 27858
rect 30156 27794 30212 27806
rect 30604 27858 30660 27870
rect 30604 27806 30606 27858
rect 30658 27806 30660 27858
rect 30380 27636 30436 27646
rect 30156 27188 30212 27198
rect 30156 27094 30212 27132
rect 29932 27010 29988 27020
rect 29484 26350 29486 26402
rect 29538 26350 29540 26402
rect 29484 25508 29540 26350
rect 29820 26964 29876 26974
rect 29708 26178 29764 26190
rect 29708 26126 29710 26178
rect 29762 26126 29764 26178
rect 29484 25442 29540 25452
rect 29596 26068 29652 26078
rect 29148 25284 29204 25294
rect 29148 25190 29204 25228
rect 29484 24722 29540 24734
rect 29484 24670 29486 24722
rect 29538 24670 29540 24722
rect 29484 24612 29540 24670
rect 29484 24546 29540 24556
rect 29148 24500 29204 24510
rect 29148 23938 29204 24444
rect 29596 24388 29652 26012
rect 29708 25732 29764 26126
rect 29708 25666 29764 25676
rect 29596 24322 29652 24332
rect 29708 24724 29764 24734
rect 29708 24162 29764 24668
rect 29708 24110 29710 24162
rect 29762 24110 29764 24162
rect 29708 24098 29764 24110
rect 29148 23886 29150 23938
rect 29202 23886 29204 23938
rect 29148 23874 29204 23886
rect 29372 23716 29428 23726
rect 29372 23622 29428 23660
rect 29596 23714 29652 23726
rect 29596 23662 29598 23714
rect 29650 23662 29652 23714
rect 29036 23548 29316 23604
rect 28252 22370 28420 22372
rect 28252 22318 28254 22370
rect 28306 22318 28420 22370
rect 28252 22316 28420 22318
rect 28252 22306 28308 22316
rect 28140 22092 28308 22148
rect 27020 21028 27076 21038
rect 27020 20934 27076 20972
rect 26908 20748 27076 20804
rect 26124 20514 26180 20524
rect 26908 20580 26964 20590
rect 26908 20486 26964 20524
rect 26012 20178 26068 20188
rect 26236 20468 26292 20478
rect 25676 20078 25678 20130
rect 25730 20078 25732 20130
rect 25676 20066 25732 20078
rect 26124 20132 26180 20142
rect 26012 20020 26068 20030
rect 26012 19926 26068 19964
rect 25788 19796 25844 19806
rect 25788 19458 25844 19740
rect 25788 19406 25790 19458
rect 25842 19406 25844 19458
rect 25788 19394 25844 19406
rect 25452 19346 25620 19348
rect 25452 19294 25454 19346
rect 25506 19294 25620 19346
rect 25452 19292 25620 19294
rect 25452 19282 25508 19292
rect 26124 19234 26180 20076
rect 26236 20130 26292 20412
rect 26236 20078 26238 20130
rect 26290 20078 26292 20130
rect 26236 20066 26292 20078
rect 27020 20132 27076 20748
rect 27020 20066 27076 20076
rect 26124 19182 26126 19234
rect 26178 19182 26180 19234
rect 26124 19170 26180 19182
rect 27020 19906 27076 19918
rect 27020 19854 27022 19906
rect 27074 19854 27076 19906
rect 27020 19234 27076 19854
rect 27132 19796 27188 22092
rect 28140 21474 28196 21486
rect 28140 21422 28142 21474
rect 28194 21422 28196 21474
rect 28140 21252 28196 21422
rect 28140 21186 28196 21196
rect 28140 21028 28196 21038
rect 28140 20934 28196 20972
rect 27244 20860 28084 20916
rect 27244 20802 27300 20860
rect 27244 20750 27246 20802
rect 27298 20750 27300 20802
rect 27244 20738 27300 20750
rect 28028 20804 28084 20860
rect 28252 20804 28308 22092
rect 28028 20748 28308 20804
rect 27580 20692 27636 20702
rect 27580 20598 27636 20636
rect 27804 20692 27860 20702
rect 27804 20598 27860 20636
rect 28252 20580 28308 20590
rect 28252 20486 28308 20524
rect 27692 20132 27748 20142
rect 28364 20132 28420 22316
rect 28588 22036 28644 22652
rect 28924 23044 28980 23054
rect 28700 22148 28756 22158
rect 28700 22054 28756 22092
rect 28476 21980 28644 22036
rect 28476 21026 28532 21980
rect 28812 21700 28868 21710
rect 28812 21586 28868 21644
rect 28812 21534 28814 21586
rect 28866 21534 28868 21586
rect 28812 21522 28868 21534
rect 28476 20974 28478 21026
rect 28530 20974 28532 21026
rect 28476 20962 28532 20974
rect 28924 20580 28980 22988
rect 29260 22484 29316 23548
rect 29596 23044 29652 23662
rect 29596 22978 29652 22988
rect 29820 23266 29876 26908
rect 30044 26516 30100 26526
rect 30044 25618 30100 26460
rect 30380 26402 30436 27580
rect 30492 27076 30548 27086
rect 30604 27076 30660 27806
rect 30548 27020 30660 27076
rect 30492 26982 30548 27020
rect 30940 26908 30996 28028
rect 30828 26852 30996 26908
rect 31052 27074 31108 27086
rect 31052 27022 31054 27074
rect 31106 27022 31108 27074
rect 30380 26350 30382 26402
rect 30434 26350 30436 26402
rect 30380 26338 30436 26350
rect 30716 26404 30772 26414
rect 30716 26290 30772 26348
rect 30716 26238 30718 26290
rect 30770 26238 30772 26290
rect 30716 26226 30772 26238
rect 30044 25566 30046 25618
rect 30098 25566 30100 25618
rect 30044 25554 30100 25566
rect 30268 26178 30324 26190
rect 30268 26126 30270 26178
rect 30322 26126 30324 26178
rect 30044 24946 30100 24958
rect 30044 24894 30046 24946
rect 30098 24894 30100 24946
rect 30044 24388 30100 24894
rect 30044 24322 30100 24332
rect 30044 23938 30100 23950
rect 30268 23940 30324 26126
rect 30492 25618 30548 25630
rect 30492 25566 30494 25618
rect 30546 25566 30548 25618
rect 30492 25508 30548 25566
rect 30492 25442 30548 25452
rect 30716 25396 30772 25406
rect 30044 23886 30046 23938
rect 30098 23886 30100 23938
rect 29820 23214 29822 23266
rect 29874 23214 29876 23266
rect 29372 22484 29428 22494
rect 29260 22482 29652 22484
rect 29260 22430 29374 22482
rect 29426 22430 29652 22482
rect 29260 22428 29652 22430
rect 29372 22418 29428 22428
rect 29596 22370 29652 22428
rect 29596 22318 29598 22370
rect 29650 22318 29652 22370
rect 29596 22306 29652 22318
rect 29820 21700 29876 23214
rect 29820 21634 29876 21644
rect 29932 23828 29988 23838
rect 29484 21474 29540 21486
rect 29484 21422 29486 21474
rect 29538 21422 29540 21474
rect 29260 21252 29316 21262
rect 29036 20692 29092 20702
rect 29036 20598 29092 20636
rect 28924 20514 28980 20524
rect 29148 20580 29204 20590
rect 28476 20132 28532 20142
rect 28364 20130 28532 20132
rect 28364 20078 28478 20130
rect 28530 20078 28532 20130
rect 28364 20076 28532 20078
rect 27692 20038 27748 20076
rect 28476 20066 28532 20076
rect 27244 20020 27300 20030
rect 29036 20020 29092 20030
rect 27244 20018 27412 20020
rect 27244 19966 27246 20018
rect 27298 19966 27412 20018
rect 27244 19964 27412 19966
rect 27244 19954 27300 19964
rect 27132 19740 27300 19796
rect 27244 19460 27300 19740
rect 27356 19572 27412 19964
rect 28812 19906 28868 19918
rect 28812 19854 28814 19906
rect 28866 19854 28868 19906
rect 27356 19516 28308 19572
rect 27244 19404 27524 19460
rect 27020 19182 27022 19234
rect 27074 19182 27076 19234
rect 25228 19124 25284 19134
rect 25228 19030 25284 19068
rect 25900 19124 25956 19134
rect 25900 19030 25956 19068
rect 24444 18676 24500 18686
rect 24220 18674 24500 18676
rect 24220 18622 24446 18674
rect 24498 18622 24500 18674
rect 24220 18620 24500 18622
rect 23996 16996 24052 17006
rect 23996 16884 24052 16940
rect 23996 16882 24164 16884
rect 23996 16830 23998 16882
rect 24050 16830 24164 16882
rect 23996 16828 24164 16830
rect 23996 16818 24052 16828
rect 24108 16098 24164 16828
rect 24108 16046 24110 16098
rect 24162 16046 24164 16098
rect 24108 16034 24164 16046
rect 23996 15988 24052 15998
rect 23996 15876 24052 15932
rect 24220 15876 24276 18620
rect 24444 18610 24500 18620
rect 26572 18564 26628 18574
rect 24332 18450 24388 18462
rect 24332 18398 24334 18450
rect 24386 18398 24388 18450
rect 24332 16996 24388 18398
rect 24668 18450 24724 18462
rect 24668 18398 24670 18450
rect 24722 18398 24724 18450
rect 24668 17556 24724 18398
rect 26572 17890 26628 18508
rect 27020 18228 27076 19182
rect 27132 19348 27188 19358
rect 27132 18450 27188 19292
rect 27244 19124 27300 19134
rect 27356 19124 27412 19134
rect 27244 19122 27356 19124
rect 27244 19070 27246 19122
rect 27298 19070 27356 19122
rect 27244 19068 27356 19070
rect 27244 19058 27300 19068
rect 27132 18398 27134 18450
rect 27186 18398 27188 18450
rect 27132 18386 27188 18398
rect 27244 18452 27300 18462
rect 26572 17838 26574 17890
rect 26626 17838 26628 17890
rect 26572 17826 26628 17838
rect 26908 18172 27076 18228
rect 25116 17666 25172 17678
rect 25116 17614 25118 17666
rect 25170 17614 25172 17666
rect 24668 17490 24724 17500
rect 24780 17554 24836 17566
rect 24780 17502 24782 17554
rect 24834 17502 24836 17554
rect 24668 16996 24724 17006
rect 24332 16994 24724 16996
rect 24332 16942 24670 16994
rect 24722 16942 24724 16994
rect 24332 16940 24724 16942
rect 24668 16930 24724 16940
rect 24780 16996 24836 17502
rect 24780 16930 24836 16940
rect 25004 16324 25060 16334
rect 25116 16324 25172 17614
rect 26796 17668 26852 17678
rect 26460 17554 26516 17566
rect 26460 17502 26462 17554
rect 26514 17502 26516 17554
rect 25564 17444 25620 17454
rect 25564 17350 25620 17388
rect 26460 17444 26516 17502
rect 26460 17378 26516 17388
rect 26572 17556 26628 17566
rect 26572 17106 26628 17500
rect 26572 17054 26574 17106
rect 26626 17054 26628 17106
rect 26572 17042 26628 17054
rect 26796 17106 26852 17612
rect 26796 17054 26798 17106
rect 26850 17054 26852 17106
rect 26796 17042 26852 17054
rect 26012 16994 26068 17006
rect 26012 16942 26014 16994
rect 26066 16942 26068 16994
rect 25788 16660 25844 16670
rect 25060 16268 25172 16324
rect 25452 16658 25844 16660
rect 25452 16606 25790 16658
rect 25842 16606 25844 16658
rect 25452 16604 25844 16606
rect 25004 16098 25060 16268
rect 25004 16046 25006 16098
rect 25058 16046 25060 16098
rect 25004 16034 25060 16046
rect 23996 15820 24276 15876
rect 23884 15708 24164 15764
rect 23884 15540 23940 15550
rect 23884 15446 23940 15484
rect 23660 15374 23662 15426
rect 23714 15374 23716 15426
rect 23660 15362 23716 15374
rect 23996 15428 24052 15438
rect 23996 15334 24052 15372
rect 23100 15316 23156 15326
rect 23436 15316 23492 15326
rect 23100 15314 23492 15316
rect 23100 15262 23102 15314
rect 23154 15262 23438 15314
rect 23490 15262 23492 15314
rect 23100 15260 23492 15262
rect 23100 15250 23156 15260
rect 23436 15250 23492 15260
rect 23548 15316 23604 15326
rect 22204 14642 22484 14644
rect 22204 14590 22206 14642
rect 22258 14590 22484 14642
rect 22204 14588 22484 14590
rect 22540 15092 22708 15148
rect 22204 13972 22260 14588
rect 22428 14420 22484 14430
rect 22428 14326 22484 14364
rect 22540 14196 22596 15092
rect 23548 14530 23604 15260
rect 24108 15148 24164 15708
rect 23548 14478 23550 14530
rect 23602 14478 23604 14530
rect 23548 14466 23604 14478
rect 23996 15092 24164 15148
rect 25452 15148 25508 16604
rect 25788 16594 25844 16604
rect 26012 16100 26068 16942
rect 26460 16882 26516 16894
rect 26460 16830 26462 16882
rect 26514 16830 26516 16882
rect 26124 16660 26180 16670
rect 26124 16658 26404 16660
rect 26124 16606 26126 16658
rect 26178 16606 26404 16658
rect 26124 16604 26404 16606
rect 26124 16594 26180 16604
rect 26236 16210 26292 16222
rect 26236 16158 26238 16210
rect 26290 16158 26292 16210
rect 26012 16044 26180 16100
rect 25676 15988 25732 15998
rect 25676 15894 25732 15932
rect 26124 15876 26180 16044
rect 25900 15820 26180 15876
rect 26236 15988 26292 16158
rect 26348 16098 26404 16604
rect 26348 16046 26350 16098
rect 26402 16046 26404 16098
rect 26348 16034 26404 16046
rect 25900 15540 25956 15820
rect 25900 15446 25956 15484
rect 26124 15540 26180 15550
rect 26236 15540 26292 15932
rect 26124 15538 26292 15540
rect 26124 15486 26126 15538
rect 26178 15486 26292 15538
rect 26124 15484 26292 15486
rect 26124 15474 26180 15484
rect 26460 15428 26516 16830
rect 26908 16322 26964 18172
rect 27020 17668 27076 17678
rect 27020 17574 27076 17612
rect 27244 17668 27300 18396
rect 27244 17574 27300 17612
rect 27356 18338 27412 19068
rect 27356 18286 27358 18338
rect 27410 18286 27412 18338
rect 26908 16270 26910 16322
rect 26962 16270 26964 16322
rect 26908 16258 26964 16270
rect 26236 15372 26516 15428
rect 25676 15316 25732 15326
rect 26236 15316 26292 15372
rect 25564 15314 25732 15316
rect 25564 15262 25678 15314
rect 25730 15262 25732 15314
rect 25564 15260 25732 15262
rect 25564 15148 25620 15260
rect 25676 15250 25732 15260
rect 26124 15260 26292 15316
rect 25452 15092 25620 15148
rect 25788 15202 25844 15214
rect 25788 15150 25790 15202
rect 25842 15150 25844 15202
rect 25788 15148 25844 15150
rect 26124 15148 26180 15260
rect 26348 15204 26404 15214
rect 25788 15092 26180 15148
rect 26236 15092 26404 15148
rect 27356 15204 27412 18286
rect 27468 18338 27524 19404
rect 27692 19348 27748 19358
rect 27692 19122 27748 19292
rect 28140 19236 28196 19246
rect 28140 19142 28196 19180
rect 28252 19234 28308 19516
rect 28252 19182 28254 19234
rect 28306 19182 28308 19234
rect 28252 19170 28308 19182
rect 28476 19348 28532 19358
rect 27692 19070 27694 19122
rect 27746 19070 27748 19122
rect 27692 19058 27748 19070
rect 28476 19122 28532 19292
rect 28476 19070 28478 19122
rect 28530 19070 28532 19122
rect 28476 19058 28532 19070
rect 28588 19124 28644 19134
rect 28588 19030 28644 19068
rect 28812 19012 28868 19854
rect 29036 19236 29092 19964
rect 29148 19346 29204 20524
rect 29148 19294 29150 19346
rect 29202 19294 29204 19346
rect 29148 19282 29204 19294
rect 29260 20578 29316 21196
rect 29372 20692 29428 20702
rect 29372 20598 29428 20636
rect 29260 20526 29262 20578
rect 29314 20526 29316 20578
rect 29036 19170 29092 19180
rect 29260 19012 29316 20526
rect 29484 20580 29540 21422
rect 29820 20802 29876 20814
rect 29820 20750 29822 20802
rect 29874 20750 29876 20802
rect 29708 20580 29764 20590
rect 29484 20578 29764 20580
rect 29484 20526 29710 20578
rect 29762 20526 29764 20578
rect 29484 20524 29764 20526
rect 29708 20514 29764 20524
rect 29820 20356 29876 20750
rect 29820 20290 29876 20300
rect 29932 20188 29988 23772
rect 30044 23716 30100 23886
rect 30044 23650 30100 23660
rect 30156 23884 30324 23940
rect 30380 25060 30436 25070
rect 30156 23492 30212 23884
rect 30268 23716 30324 23726
rect 30380 23716 30436 25004
rect 30716 24722 30772 25340
rect 30828 24836 30884 26852
rect 31052 26402 31108 27022
rect 31052 26350 31054 26402
rect 31106 26350 31108 26402
rect 30828 24770 30884 24780
rect 30940 25284 30996 25294
rect 30716 24670 30718 24722
rect 30770 24670 30772 24722
rect 30716 24658 30772 24670
rect 30268 23714 30436 23716
rect 30268 23662 30270 23714
rect 30322 23662 30436 23714
rect 30268 23660 30436 23662
rect 30604 23940 30660 23950
rect 30268 23650 30324 23660
rect 30044 23436 30212 23492
rect 30044 21026 30100 23436
rect 30604 21812 30660 23884
rect 30828 23940 30884 23950
rect 30828 23714 30884 23884
rect 30828 23662 30830 23714
rect 30882 23662 30884 23714
rect 30828 22372 30884 23662
rect 30940 23716 30996 25228
rect 30940 23650 30996 23660
rect 31052 23492 31108 26350
rect 31164 26740 31220 26750
rect 31164 26292 31220 26684
rect 31276 26516 31332 30156
rect 31500 30100 31556 30110
rect 31500 30006 31556 30044
rect 31948 30100 32004 30110
rect 31948 30006 32004 30044
rect 32060 29650 32116 30156
rect 32508 30212 32564 30222
rect 32508 30118 32564 30156
rect 33068 30212 33124 30222
rect 32172 30100 32228 30110
rect 32172 30006 32228 30044
rect 32732 29988 32788 29998
rect 32732 29986 33012 29988
rect 32732 29934 32734 29986
rect 32786 29934 33012 29986
rect 32732 29932 33012 29934
rect 32732 29922 32788 29932
rect 32060 29598 32062 29650
rect 32114 29598 32116 29650
rect 32060 29586 32116 29598
rect 31724 29538 31780 29550
rect 31724 29486 31726 29538
rect 31778 29486 31780 29538
rect 31388 29426 31444 29438
rect 31388 29374 31390 29426
rect 31442 29374 31444 29426
rect 31388 29316 31444 29374
rect 31388 29250 31444 29260
rect 31724 28756 31780 29486
rect 32284 29428 32340 29438
rect 31724 28690 31780 28700
rect 31836 29316 31892 29326
rect 31500 27746 31556 27758
rect 31500 27694 31502 27746
rect 31554 27694 31556 27746
rect 31500 27076 31556 27694
rect 31612 27076 31668 27086
rect 31500 27074 31668 27076
rect 31500 27022 31614 27074
rect 31666 27022 31668 27074
rect 31500 27020 31668 27022
rect 31612 26964 31668 27020
rect 31612 26898 31668 26908
rect 31836 26628 31892 29260
rect 32060 29204 32116 29214
rect 31836 26562 31892 26572
rect 31948 28420 32004 28430
rect 31276 26450 31332 26460
rect 31612 26292 31668 26302
rect 31164 26290 31444 26292
rect 31164 26238 31166 26290
rect 31218 26238 31444 26290
rect 31164 26236 31444 26238
rect 31164 26226 31220 26236
rect 31388 25618 31444 26236
rect 31388 25566 31390 25618
rect 31442 25566 31444 25618
rect 31388 25554 31444 25566
rect 31612 25396 31668 26236
rect 31948 25618 32004 28364
rect 32060 26292 32116 29148
rect 32284 28754 32340 29372
rect 32284 28702 32286 28754
rect 32338 28702 32340 28754
rect 32284 26908 32340 28702
rect 32396 29426 32452 29438
rect 32396 29374 32398 29426
rect 32450 29374 32452 29426
rect 32396 28868 32452 29374
rect 32956 28980 33012 29932
rect 33068 29426 33124 30156
rect 33068 29374 33070 29426
rect 33122 29374 33124 29426
rect 33068 29362 33124 29374
rect 33180 29204 33236 31838
rect 33180 29138 33236 29148
rect 33292 29202 33348 31948
rect 33516 31778 33572 32284
rect 33628 32274 33684 32284
rect 33516 31726 33518 31778
rect 33570 31726 33572 31778
rect 33516 31714 33572 31726
rect 33852 31220 33908 34748
rect 33964 34132 34020 35084
rect 34412 34916 34468 34926
rect 34300 34914 34468 34916
rect 34300 34862 34414 34914
rect 34466 34862 34468 34914
rect 34300 34860 34468 34862
rect 34300 34354 34356 34860
rect 34412 34850 34468 34860
rect 34524 34804 34580 35084
rect 34748 34916 34804 35422
rect 35084 35474 35140 35486
rect 35084 35422 35086 35474
rect 35138 35422 35140 35474
rect 35084 35140 35140 35422
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35084 35084 35364 35140
rect 34748 34850 34804 34860
rect 34972 35026 35028 35038
rect 34972 34974 34974 35026
rect 35026 34974 35028 35026
rect 34524 34710 34580 34748
rect 34300 34302 34302 34354
rect 34354 34302 34356 34354
rect 34300 34290 34356 34302
rect 34860 34354 34916 34366
rect 34860 34302 34862 34354
rect 34914 34302 34916 34354
rect 34748 34244 34804 34254
rect 34860 34244 34916 34302
rect 34804 34188 34916 34244
rect 34748 34178 34804 34188
rect 33964 34038 34020 34076
rect 34636 34132 34692 34142
rect 34636 34038 34692 34076
rect 34748 34018 34804 34030
rect 34748 33966 34750 34018
rect 34802 33966 34804 34018
rect 34748 33460 34804 33966
rect 34972 33572 35028 34974
rect 35308 34914 35364 35084
rect 35308 34862 35310 34914
rect 35362 34862 35364 34914
rect 35308 34850 35364 34862
rect 35756 34690 35812 34702
rect 35756 34638 35758 34690
rect 35810 34638 35812 34690
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 34300 33348 34356 33358
rect 34300 33254 34356 33292
rect 34636 33348 34692 33358
rect 34748 33348 34804 33404
rect 34636 33346 34804 33348
rect 34636 33294 34638 33346
rect 34690 33294 34804 33346
rect 34636 33292 34804 33294
rect 34860 33516 35028 33572
rect 34636 33282 34692 33292
rect 34748 33122 34804 33134
rect 34748 33070 34750 33122
rect 34802 33070 34804 33122
rect 34076 32450 34132 32462
rect 34076 32398 34078 32450
rect 34130 32398 34132 32450
rect 34076 31332 34132 32398
rect 34524 31892 34580 31902
rect 34524 31798 34580 31836
rect 34748 31668 34804 33070
rect 34748 31602 34804 31612
rect 34860 31890 34916 33516
rect 35532 33460 35588 33470
rect 34972 33346 35028 33358
rect 34972 33294 34974 33346
rect 35026 33294 35028 33346
rect 34972 33236 35028 33294
rect 34972 33170 35028 33180
rect 35084 33346 35140 33358
rect 35084 33294 35086 33346
rect 35138 33294 35140 33346
rect 35084 32340 35140 33294
rect 35532 33346 35588 33404
rect 35532 33294 35534 33346
rect 35586 33294 35588 33346
rect 35532 33282 35588 33294
rect 35644 33348 35700 33358
rect 35644 33254 35700 33292
rect 35756 33346 35812 34638
rect 35756 33294 35758 33346
rect 35810 33294 35812 33346
rect 35756 33236 35812 33294
rect 35756 33170 35812 33180
rect 35084 32274 35140 32284
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 34860 31838 34862 31890
rect 34914 31838 34916 31890
rect 34860 31556 34916 31838
rect 35196 31892 35252 31902
rect 35196 31778 35252 31836
rect 35196 31726 35198 31778
rect 35250 31726 35252 31778
rect 35196 31714 35252 31726
rect 34972 31556 35028 31566
rect 34860 31500 34972 31556
rect 34972 31490 35028 31500
rect 34076 31276 35140 31332
rect 33852 31164 34580 31220
rect 34188 30996 34244 31006
rect 34076 30210 34132 30222
rect 34076 30158 34078 30210
rect 34130 30158 34132 30210
rect 33740 29986 33796 29998
rect 33740 29934 33742 29986
rect 33794 29934 33796 29986
rect 33740 29764 33796 29934
rect 33740 29698 33796 29708
rect 33292 29150 33294 29202
rect 33346 29150 33348 29202
rect 33292 29138 33348 29150
rect 33516 29650 33572 29662
rect 33516 29598 33518 29650
rect 33570 29598 33572 29650
rect 32956 28924 33348 28980
rect 32396 28084 32452 28812
rect 32732 28756 32788 28766
rect 32732 28642 32788 28700
rect 32732 28590 32734 28642
rect 32786 28590 32788 28642
rect 32732 28578 32788 28590
rect 32732 28084 32788 28094
rect 33180 28084 33236 28094
rect 32396 28018 32452 28028
rect 32508 28028 32732 28084
rect 32396 27188 32452 27198
rect 32508 27188 32564 28028
rect 32732 28018 32788 28028
rect 32844 28028 33124 28084
rect 32396 27186 32564 27188
rect 32396 27134 32398 27186
rect 32450 27134 32564 27186
rect 32396 27132 32564 27134
rect 32396 27122 32452 27132
rect 32284 26852 32452 26908
rect 32060 26198 32116 26236
rect 32396 26404 32452 26852
rect 31948 25566 31950 25618
rect 32002 25566 32004 25618
rect 31948 25554 32004 25566
rect 31276 24722 31332 24734
rect 31276 24670 31278 24722
rect 31330 24670 31332 24722
rect 31276 24052 31332 24670
rect 31276 23986 31332 23996
rect 31612 23938 31668 25340
rect 31836 25282 31892 25294
rect 31836 25230 31838 25282
rect 31890 25230 31892 25282
rect 31836 24948 31892 25230
rect 32060 25282 32116 25294
rect 32060 25230 32062 25282
rect 32114 25230 32116 25282
rect 32060 25060 32116 25230
rect 32060 24994 32116 25004
rect 32284 25284 32340 25294
rect 31836 24882 31892 24892
rect 31612 23886 31614 23938
rect 31666 23886 31668 23938
rect 31612 23874 31668 23886
rect 31724 24834 31780 24846
rect 31724 24782 31726 24834
rect 31778 24782 31780 24834
rect 31612 23716 31668 23726
rect 31164 23492 31220 23502
rect 31052 23436 31164 23492
rect 31164 23426 31220 23436
rect 31612 23378 31668 23660
rect 31724 23492 31780 24782
rect 32060 24834 32116 24846
rect 32060 24782 32062 24834
rect 32114 24782 32116 24834
rect 31836 24722 31892 24734
rect 31836 24670 31838 24722
rect 31890 24670 31892 24722
rect 31836 23716 31892 24670
rect 31836 23650 31892 23660
rect 32060 24052 32116 24782
rect 31724 23426 31780 23436
rect 31612 23326 31614 23378
rect 31666 23326 31668 23378
rect 31612 23314 31668 23326
rect 31948 23266 32004 23278
rect 31948 23214 31950 23266
rect 32002 23214 32004 23266
rect 31948 23044 32004 23214
rect 31948 22978 32004 22988
rect 32060 22820 32116 23996
rect 32172 23940 32228 23950
rect 32172 23846 32228 23884
rect 32172 23268 32228 23278
rect 32284 23268 32340 25228
rect 32396 24722 32452 26348
rect 32508 25508 32564 25518
rect 32508 25506 32788 25508
rect 32508 25454 32510 25506
rect 32562 25454 32788 25506
rect 32508 25452 32788 25454
rect 32508 25442 32564 25452
rect 32732 25394 32788 25452
rect 32732 25342 32734 25394
rect 32786 25342 32788 25394
rect 32732 24948 32788 25342
rect 32844 24948 32900 28028
rect 33068 27970 33124 28028
rect 33180 27990 33236 28028
rect 33292 28082 33348 28924
rect 33516 28532 33572 29598
rect 33628 29428 33684 29438
rect 33628 29334 33684 29372
rect 33852 29428 33908 29438
rect 33852 29334 33908 29372
rect 34076 29204 34132 30158
rect 34076 29138 34132 29148
rect 34188 28980 34244 30940
rect 34524 30548 34580 31164
rect 34860 30772 34916 30782
rect 34860 30770 35028 30772
rect 34860 30718 34862 30770
rect 34914 30718 35028 30770
rect 34860 30716 35028 30718
rect 34860 30706 34916 30716
rect 34524 30492 34916 30548
rect 33516 28466 33572 28476
rect 34076 28924 34244 28980
rect 34748 29426 34804 29438
rect 34748 29374 34750 29426
rect 34802 29374 34804 29426
rect 33292 28030 33294 28082
rect 33346 28030 33348 28082
rect 33292 28018 33348 28030
rect 33628 28308 33684 28318
rect 33068 27918 33070 27970
rect 33122 27918 33124 27970
rect 33068 27906 33124 27918
rect 33404 26628 33460 26638
rect 33404 26178 33460 26572
rect 33404 26126 33406 26178
rect 33458 26126 33460 26178
rect 32956 26066 33012 26078
rect 32956 26014 32958 26066
rect 33010 26014 33012 26066
rect 32956 25506 33012 26014
rect 33404 26066 33460 26126
rect 33404 26014 33406 26066
rect 33458 26014 33460 26066
rect 33404 26002 33460 26014
rect 33628 25732 33684 28252
rect 34076 28082 34132 28924
rect 34748 28644 34804 29374
rect 34860 29426 34916 30492
rect 34860 29374 34862 29426
rect 34914 29374 34916 29426
rect 34860 29362 34916 29374
rect 34972 29426 35028 30716
rect 35084 30210 35140 31276
rect 35868 30996 35924 38612
rect 36316 37268 36372 37278
rect 36316 37174 36372 37212
rect 36428 36482 36484 38892
rect 36652 38882 36708 38892
rect 37100 39394 37156 39406
rect 37100 39342 37102 39394
rect 37154 39342 37156 39394
rect 37100 38948 37156 39342
rect 39116 39396 39172 39406
rect 39116 39302 39172 39340
rect 37100 38946 37380 38948
rect 37100 38894 37102 38946
rect 37154 38894 37380 38946
rect 37100 38892 37380 38894
rect 37100 38882 37156 38892
rect 36540 38724 36596 38734
rect 36540 38630 36596 38668
rect 36428 36430 36430 36482
rect 36482 36430 36484 36482
rect 36428 36418 36484 36430
rect 37100 38164 37156 38174
rect 37100 37268 37156 38108
rect 37100 36482 37156 37212
rect 37100 36430 37102 36482
rect 37154 36430 37156 36482
rect 37100 36418 37156 36430
rect 37212 37828 37268 37838
rect 36988 36372 37044 36382
rect 36876 36370 37044 36372
rect 36876 36318 36990 36370
rect 37042 36318 37044 36370
rect 36876 36316 37044 36318
rect 36092 36258 36148 36270
rect 36092 36206 36094 36258
rect 36146 36206 36148 36258
rect 36092 35812 36148 36206
rect 36092 35746 36148 35756
rect 36316 35810 36372 35822
rect 36316 35758 36318 35810
rect 36370 35758 36372 35810
rect 36316 35588 36372 35758
rect 36540 35812 36596 35822
rect 36540 35718 36596 35756
rect 36876 35700 36932 36316
rect 36988 36306 37044 36316
rect 36876 35606 36932 35644
rect 37100 35698 37156 35710
rect 37100 35646 37102 35698
rect 37154 35646 37156 35698
rect 36204 35532 36316 35588
rect 36092 34916 36148 34926
rect 36092 34822 36148 34860
rect 35980 34804 36036 34814
rect 35980 34710 36036 34748
rect 35980 34356 36036 34366
rect 36204 34356 36260 35532
rect 36316 35522 36372 35532
rect 37100 35588 37156 35646
rect 36652 35476 36708 35486
rect 36652 35382 36708 35420
rect 35980 34354 36260 34356
rect 35980 34302 35982 34354
rect 36034 34302 36260 34354
rect 35980 34300 36260 34302
rect 35980 34290 36036 34300
rect 36204 34242 36260 34300
rect 36204 34190 36206 34242
rect 36258 34190 36260 34242
rect 36204 34178 36260 34190
rect 36316 35140 36372 35150
rect 36316 34242 36372 35084
rect 37100 35026 37156 35532
rect 37100 34974 37102 35026
rect 37154 34974 37156 35026
rect 37100 34962 37156 34974
rect 37212 34356 37268 37772
rect 37324 37266 37380 38892
rect 38444 38946 38500 38958
rect 38444 38894 38446 38946
rect 38498 38894 38500 38946
rect 37324 37214 37326 37266
rect 37378 37214 37380 37266
rect 37324 37202 37380 37214
rect 37772 38724 37828 38734
rect 37772 37154 37828 38668
rect 38444 38164 38500 38894
rect 38668 38836 38724 38846
rect 39004 38836 39060 38846
rect 38668 38834 39060 38836
rect 38668 38782 38670 38834
rect 38722 38782 39006 38834
rect 39058 38782 39060 38834
rect 38668 38780 39060 38782
rect 38668 38770 38724 38780
rect 39004 38770 39060 38780
rect 39228 38668 39284 40348
rect 39564 39618 39620 40348
rect 39564 39566 39566 39618
rect 39618 39566 39620 39618
rect 39564 39554 39620 39566
rect 39676 39620 39732 39630
rect 39676 39526 39732 39564
rect 39788 39506 39844 39518
rect 39788 39454 39790 39506
rect 39842 39454 39844 39506
rect 39788 39396 39844 39454
rect 39676 38946 39732 38958
rect 39676 38894 39678 38946
rect 39730 38894 39732 38946
rect 38444 38098 38500 38108
rect 39116 38612 39284 38668
rect 39452 38722 39508 38734
rect 39452 38670 39454 38722
rect 39506 38670 39508 38722
rect 39116 38050 39172 38612
rect 39116 37998 39118 38050
rect 39170 37998 39172 38050
rect 39116 37986 39172 37998
rect 39340 38276 39396 38286
rect 39340 38050 39396 38220
rect 39340 37998 39342 38050
rect 39394 37998 39396 38050
rect 39340 37986 39396 37998
rect 37772 37102 37774 37154
rect 37826 37102 37828 37154
rect 37772 36932 37828 37102
rect 37660 36876 37772 36932
rect 37660 36482 37716 36876
rect 37772 36866 37828 36876
rect 38332 37380 38388 37390
rect 37660 36430 37662 36482
rect 37714 36430 37716 36482
rect 37660 36418 37716 36430
rect 38332 36482 38388 37324
rect 39452 37380 39508 38670
rect 39676 38274 39732 38894
rect 39676 38222 39678 38274
rect 39730 38222 39732 38274
rect 39676 38210 39732 38222
rect 39564 37940 39620 37950
rect 39788 37940 39844 39340
rect 39900 38834 39956 41580
rect 39900 38782 39902 38834
rect 39954 38782 39956 38834
rect 39900 38770 39956 38782
rect 40012 38836 40068 42700
rect 40348 42644 40404 43596
rect 40348 42578 40404 42588
rect 40236 42530 40292 42542
rect 40236 42478 40238 42530
rect 40290 42478 40292 42530
rect 40124 42420 40180 42430
rect 40124 41412 40180 42364
rect 40236 42196 40292 42478
rect 40236 42130 40292 42140
rect 40348 41972 40404 41982
rect 40460 41972 40516 45838
rect 40572 44324 40628 46284
rect 41020 45892 41076 49200
rect 41020 45826 41076 45836
rect 41356 46116 41412 46126
rect 41356 45892 41412 46060
rect 41356 45890 41524 45892
rect 41356 45838 41358 45890
rect 41410 45838 41524 45890
rect 41356 45836 41524 45838
rect 41356 45826 41412 45836
rect 40796 45666 40852 45678
rect 40796 45614 40798 45666
rect 40850 45614 40852 45666
rect 40572 42868 40628 44268
rect 40684 45220 40740 45230
rect 40684 44210 40740 45164
rect 40684 44158 40686 44210
rect 40738 44158 40740 44210
rect 40684 43764 40740 44158
rect 40684 43698 40740 43708
rect 40684 42868 40740 42878
rect 40572 42866 40740 42868
rect 40572 42814 40686 42866
rect 40738 42814 40740 42866
rect 40572 42812 40740 42814
rect 40684 42802 40740 42812
rect 40348 41970 40516 41972
rect 40348 41918 40350 41970
rect 40402 41918 40516 41970
rect 40348 41916 40516 41918
rect 40348 41906 40404 41916
rect 40124 41356 40292 41412
rect 40124 40964 40180 40974
rect 40124 40870 40180 40908
rect 40012 38770 40068 38780
rect 40124 39844 40180 39854
rect 40124 38668 40180 39788
rect 40012 38612 40180 38668
rect 39564 37938 39844 37940
rect 39564 37886 39566 37938
rect 39618 37886 39844 37938
rect 39564 37884 39844 37886
rect 39900 38276 39956 38286
rect 39564 37874 39620 37884
rect 39788 37492 39844 37502
rect 39900 37492 39956 38220
rect 39844 37436 39956 37492
rect 40012 38052 40068 38612
rect 40236 38388 40292 41356
rect 40460 41188 40516 41198
rect 40796 41188 40852 45614
rect 41020 45332 41076 45342
rect 41020 45106 41076 45276
rect 41020 45054 41022 45106
rect 41074 45054 41076 45106
rect 41020 44772 41076 45054
rect 41020 44706 41076 44716
rect 41356 44996 41412 45006
rect 41356 44100 41412 44940
rect 41356 44034 41412 44044
rect 41468 44322 41524 45836
rect 41468 44270 41470 44322
rect 41522 44270 41524 44322
rect 40908 43764 40964 43774
rect 40908 42756 40964 43708
rect 41020 43652 41076 43662
rect 41244 43652 41300 43662
rect 41020 43650 41244 43652
rect 41020 43598 41022 43650
rect 41074 43598 41244 43650
rect 41020 43596 41244 43598
rect 41020 43586 41076 43596
rect 41132 42980 41188 42990
rect 41132 42886 41188 42924
rect 41020 42756 41076 42766
rect 40908 42754 41076 42756
rect 40908 42702 41022 42754
rect 41074 42702 41076 42754
rect 40908 42700 41076 42702
rect 41020 42084 41076 42700
rect 41020 42018 41076 42028
rect 41132 42644 41188 42654
rect 41132 42530 41188 42588
rect 41132 42478 41134 42530
rect 41186 42478 41188 42530
rect 40460 41186 40852 41188
rect 40460 41134 40462 41186
rect 40514 41134 40798 41186
rect 40850 41134 40852 41186
rect 40460 41132 40852 41134
rect 40460 41122 40516 41132
rect 40796 41122 40852 41132
rect 41132 40962 41188 42478
rect 41244 42196 41300 43596
rect 41356 43540 41412 43550
rect 41356 43446 41412 43484
rect 41468 42308 41524 44270
rect 41580 45108 41636 45118
rect 41580 43708 41636 45052
rect 41692 44660 41748 49200
rect 42364 46450 42420 49200
rect 42364 46398 42366 46450
rect 42418 46398 42420 46450
rect 42364 46386 42420 46398
rect 42252 46228 42308 46238
rect 43036 46228 43092 49200
rect 43708 46676 43764 49200
rect 44380 46900 44436 49200
rect 44380 46834 44436 46844
rect 43708 46620 44436 46676
rect 43036 46172 43540 46228
rect 41804 45890 41860 45902
rect 41804 45838 41806 45890
rect 41858 45838 41860 45890
rect 41804 45108 41860 45838
rect 42252 45890 42308 46172
rect 42252 45838 42254 45890
rect 42306 45838 42308 45890
rect 42252 45444 42308 45838
rect 42588 46116 42644 46126
rect 43484 46116 43540 46172
rect 43484 46060 43764 46116
rect 42364 45780 42420 45790
rect 42364 45686 42420 45724
rect 42588 45778 42644 46060
rect 42588 45726 42590 45778
rect 42642 45726 42644 45778
rect 42588 45714 42644 45726
rect 42812 45890 42868 45902
rect 42812 45838 42814 45890
rect 42866 45838 42868 45890
rect 42252 45388 42756 45444
rect 42252 45220 42308 45230
rect 42252 45126 42308 45164
rect 41804 45042 41860 45052
rect 42028 45106 42084 45118
rect 42028 45054 42030 45106
rect 42082 45054 42084 45106
rect 41692 44594 41748 44604
rect 41916 44210 41972 44222
rect 41916 44158 41918 44210
rect 41970 44158 41972 44210
rect 41916 44100 41972 44158
rect 41916 44034 41972 44044
rect 42028 43988 42084 45054
rect 42028 43922 42084 43932
rect 42588 45108 42644 45118
rect 41580 43652 41972 43708
rect 41244 42130 41300 42140
rect 41356 42252 41524 42308
rect 41580 43540 41636 43550
rect 41356 42082 41412 42252
rect 41356 42030 41358 42082
rect 41410 42030 41412 42082
rect 41356 42018 41412 42030
rect 41468 42084 41524 42094
rect 41580 42084 41636 43484
rect 41804 43540 41860 43550
rect 41804 43446 41860 43484
rect 41804 42756 41860 42766
rect 41804 42662 41860 42700
rect 41916 42642 41972 43652
rect 41916 42590 41918 42642
rect 41970 42590 41972 42642
rect 41916 42578 41972 42590
rect 42028 43650 42084 43662
rect 42028 43598 42030 43650
rect 42082 43598 42084 43650
rect 42028 42644 42084 43598
rect 42588 43540 42644 45052
rect 42700 43708 42756 45388
rect 42812 44884 42868 45838
rect 43596 45890 43652 45902
rect 43596 45838 43598 45890
rect 43650 45838 43652 45890
rect 43036 45780 43092 45790
rect 43036 45218 43092 45724
rect 43596 45780 43652 45838
rect 43596 45714 43652 45724
rect 43148 45668 43204 45678
rect 43708 45668 43764 46060
rect 44156 45668 44212 45678
rect 43708 45666 44212 45668
rect 43708 45614 44158 45666
rect 44210 45614 44212 45666
rect 43708 45612 44212 45614
rect 43148 45574 43204 45612
rect 44156 45332 44212 45612
rect 44156 45276 44324 45332
rect 43036 45166 43038 45218
rect 43090 45166 43092 45218
rect 42924 45108 42980 45118
rect 42924 45014 42980 45052
rect 42812 44828 42980 44884
rect 42812 44212 42868 44222
rect 42812 44118 42868 44156
rect 42700 43642 42756 43652
rect 42924 44100 42980 44828
rect 42924 43650 42980 44044
rect 43036 43764 43092 45166
rect 43820 45218 43876 45230
rect 43820 45166 43822 45218
rect 43874 45166 43876 45218
rect 43372 44996 43428 45006
rect 43372 44902 43428 44940
rect 43036 43698 43092 43708
rect 43708 44548 43764 44558
rect 42924 43598 42926 43650
rect 42978 43598 42980 43650
rect 42924 43586 42980 43598
rect 43708 43540 43764 44492
rect 43820 43652 43876 45166
rect 44268 45220 44324 45276
rect 44268 45154 44324 45164
rect 44156 45108 44212 45118
rect 44156 44212 44212 45052
rect 44380 44884 44436 46620
rect 44940 46450 44996 46462
rect 44940 46398 44942 46450
rect 44994 46398 44996 46450
rect 44604 46116 44660 46126
rect 44604 46002 44660 46060
rect 44604 45950 44606 46002
rect 44658 45950 44660 46002
rect 44604 45938 44660 45950
rect 44940 45892 44996 46398
rect 45052 46228 45108 49200
rect 45052 46172 45556 46228
rect 45052 45892 45108 45902
rect 44940 45890 45108 45892
rect 44940 45838 45054 45890
rect 45106 45838 45108 45890
rect 44940 45836 45108 45838
rect 44716 45220 44772 45230
rect 44380 44818 44436 44828
rect 44492 45218 44772 45220
rect 44492 45166 44718 45218
rect 44770 45166 44772 45218
rect 44492 45164 44772 45166
rect 44380 44436 44436 44446
rect 44492 44436 44548 45164
rect 44716 45154 44772 45164
rect 44940 45220 44996 45230
rect 44380 44434 44548 44436
rect 44380 44382 44382 44434
rect 44434 44382 44548 44434
rect 44380 44380 44548 44382
rect 44380 44370 44436 44380
rect 44156 44146 44212 44156
rect 44268 44322 44324 44334
rect 44268 44270 44270 44322
rect 44322 44270 44324 44322
rect 44156 43708 44212 43718
rect 43820 43596 43988 43652
rect 42588 43538 42868 43540
rect 42588 43486 42590 43538
rect 42642 43486 42868 43538
rect 42588 43484 42868 43486
rect 43708 43484 43876 43540
rect 42588 43474 42644 43484
rect 42140 43092 42196 43102
rect 42140 42754 42196 43036
rect 42140 42702 42142 42754
rect 42194 42702 42196 42754
rect 42140 42690 42196 42702
rect 42812 42756 42868 43484
rect 43036 42756 43092 42766
rect 42868 42754 43092 42756
rect 42868 42702 43038 42754
rect 43090 42702 43092 42754
rect 42868 42700 43092 42702
rect 42812 42662 42868 42700
rect 43036 42690 43092 42700
rect 41468 42082 41636 42084
rect 41468 42030 41470 42082
rect 41522 42030 41636 42082
rect 41468 42028 41636 42030
rect 41692 42532 41748 42542
rect 41468 42018 41524 42028
rect 41692 41970 41748 42476
rect 42028 42196 42084 42588
rect 42700 42644 42756 42654
rect 42364 42530 42420 42542
rect 42364 42478 42366 42530
rect 42418 42478 42420 42530
rect 42028 42140 42196 42196
rect 41804 42084 41860 42094
rect 41860 42028 42084 42084
rect 41804 42018 41860 42028
rect 41692 41918 41694 41970
rect 41746 41918 41748 41970
rect 41692 41906 41748 41918
rect 42028 41970 42084 42028
rect 42028 41918 42030 41970
rect 42082 41918 42084 41970
rect 42028 41906 42084 41918
rect 42140 41186 42196 42140
rect 42140 41134 42142 41186
rect 42194 41134 42196 41186
rect 41692 41074 41748 41086
rect 41692 41022 41694 41074
rect 41746 41022 41748 41074
rect 41132 40910 41134 40962
rect 41186 40910 41188 40962
rect 40348 40740 40404 40750
rect 40348 40292 40404 40684
rect 40348 40226 40404 40236
rect 40460 40628 40516 40638
rect 40348 39618 40404 39630
rect 40348 39566 40350 39618
rect 40402 39566 40404 39618
rect 40348 39284 40404 39566
rect 40460 39284 40516 40572
rect 41020 40404 41076 40414
rect 41132 40404 41188 40910
rect 41356 40964 41412 40974
rect 41356 40870 41412 40908
rect 41580 40962 41636 40974
rect 41580 40910 41582 40962
rect 41634 40910 41636 40962
rect 41580 40852 41636 40910
rect 41580 40786 41636 40796
rect 41692 40740 41748 41022
rect 41692 40674 41748 40684
rect 41020 40402 41188 40404
rect 41020 40350 41022 40402
rect 41074 40350 41188 40402
rect 41020 40348 41188 40350
rect 41244 40514 41300 40526
rect 41244 40462 41246 40514
rect 41298 40462 41300 40514
rect 41020 40338 41076 40348
rect 41132 40180 41188 40190
rect 40684 39732 40740 39742
rect 40684 39638 40740 39676
rect 41132 39506 41188 40124
rect 41244 39956 41300 40462
rect 42140 40180 42196 41134
rect 42252 42082 42308 42094
rect 42252 42030 42254 42082
rect 42306 42030 42308 42082
rect 42252 41188 42308 42030
rect 42364 41860 42420 42478
rect 42700 42420 42756 42588
rect 43372 42532 43428 42542
rect 43708 42532 43764 42542
rect 42700 42354 42756 42364
rect 43148 42530 43428 42532
rect 43148 42478 43374 42530
rect 43426 42478 43428 42530
rect 43148 42476 43428 42478
rect 42476 42084 42532 42094
rect 42812 42084 42868 42094
rect 42532 42028 42756 42084
rect 42476 42018 42532 42028
rect 42700 41970 42756 42028
rect 42700 41918 42702 41970
rect 42754 41918 42756 41970
rect 42700 41906 42756 41918
rect 42364 41412 42420 41804
rect 42476 41748 42532 41758
rect 42476 41654 42532 41692
rect 42812 41524 42868 42028
rect 43148 41972 43204 42476
rect 43372 42466 43428 42476
rect 43484 42530 43764 42532
rect 43484 42478 43710 42530
rect 43762 42478 43764 42530
rect 43484 42476 43764 42478
rect 43372 42084 43428 42094
rect 43484 42084 43540 42476
rect 43708 42466 43764 42476
rect 43820 42532 43876 43484
rect 43820 42466 43876 42476
rect 43932 42308 43988 43596
rect 44156 43650 44212 43652
rect 44156 43598 44158 43650
rect 44210 43598 44212 43650
rect 44156 43586 44212 43598
rect 44268 43540 44324 44270
rect 44044 42756 44100 42766
rect 44268 42756 44324 43484
rect 44492 43708 44548 44380
rect 44940 44434 44996 45164
rect 44940 44382 44942 44434
rect 44994 44382 44996 44434
rect 44940 44370 44996 44382
rect 45052 43988 45108 45836
rect 45500 45890 45556 46172
rect 45500 45838 45502 45890
rect 45554 45838 45556 45890
rect 45388 45106 45444 45118
rect 45388 45054 45390 45106
rect 45442 45054 45444 45106
rect 45276 44994 45332 45006
rect 45276 44942 45278 44994
rect 45330 44942 45332 44994
rect 45276 44436 45332 44942
rect 45276 44370 45332 44380
rect 44940 43932 45108 43988
rect 44604 43764 44660 43774
rect 44492 43652 44660 43708
rect 44044 42754 44324 42756
rect 44044 42702 44046 42754
rect 44098 42702 44324 42754
rect 44044 42700 44324 42702
rect 44380 42980 44436 42990
rect 44044 42690 44100 42700
rect 43428 42028 43540 42084
rect 43708 42252 43988 42308
rect 43372 41990 43428 42028
rect 43708 41972 43764 42252
rect 44156 42082 44212 42094
rect 44156 42030 44158 42082
rect 44210 42030 44212 42082
rect 43148 41636 43204 41916
rect 43484 41916 43764 41972
rect 43484 41858 43540 41916
rect 43484 41806 43486 41858
rect 43538 41806 43540 41858
rect 43148 41580 43316 41636
rect 42364 41346 42420 41356
rect 42476 41468 42868 41524
rect 42252 41186 42420 41188
rect 42252 41134 42254 41186
rect 42306 41134 42420 41186
rect 42252 41132 42420 41134
rect 42252 41122 42308 41132
rect 42140 40114 42196 40124
rect 42364 40404 42420 41132
rect 42476 41186 42532 41468
rect 42588 41300 42644 41310
rect 43148 41300 43204 41310
rect 42588 41298 43204 41300
rect 42588 41246 42590 41298
rect 42642 41246 43150 41298
rect 43202 41246 43204 41298
rect 42588 41244 43204 41246
rect 42588 41234 42644 41244
rect 43148 41234 43204 41244
rect 42476 41134 42478 41186
rect 42530 41134 42532 41186
rect 42476 40516 42532 41134
rect 42588 40964 42644 40974
rect 42588 40870 42644 40908
rect 43036 40740 43092 40750
rect 43260 40740 43316 41580
rect 43092 40684 43316 40740
rect 43372 40740 43428 40750
rect 42812 40516 42868 40526
rect 42476 40514 42868 40516
rect 42476 40462 42814 40514
rect 42866 40462 42868 40514
rect 42476 40460 42868 40462
rect 41244 39900 41412 39956
rect 41132 39454 41134 39506
rect 41186 39454 41188 39506
rect 40348 39228 41076 39284
rect 41020 38946 41076 39228
rect 41020 38894 41022 38946
rect 41074 38894 41076 38946
rect 41020 38882 41076 38894
rect 40908 38836 40964 38846
rect 40908 38742 40964 38780
rect 41132 38668 41188 39454
rect 40236 38276 40292 38332
rect 39788 37398 39844 37436
rect 40012 37380 40068 37996
rect 40124 38220 40292 38276
rect 40572 38612 41188 38668
rect 41244 39732 41300 39742
rect 40124 37604 40180 38220
rect 40348 38164 40404 38174
rect 40236 38050 40292 38062
rect 40236 37998 40238 38050
rect 40290 37998 40292 38050
rect 40236 37940 40292 37998
rect 40236 37874 40292 37884
rect 40348 37826 40404 38108
rect 40348 37774 40350 37826
rect 40402 37774 40404 37826
rect 40348 37762 40404 37774
rect 40460 37940 40516 37950
rect 40124 37548 40292 37604
rect 40124 37380 40180 37390
rect 40012 37378 40180 37380
rect 40012 37326 40126 37378
rect 40178 37326 40180 37378
rect 40012 37324 40180 37326
rect 39452 37314 39508 37324
rect 40124 37314 40180 37324
rect 40236 37378 40292 37548
rect 40460 37490 40516 37884
rect 40460 37438 40462 37490
rect 40514 37438 40516 37490
rect 40460 37426 40516 37438
rect 40236 37326 40238 37378
rect 40290 37326 40292 37378
rect 40236 37314 40292 37326
rect 38332 36430 38334 36482
rect 38386 36430 38388 36482
rect 38332 36418 38388 36430
rect 38444 36484 38500 36494
rect 39004 36484 39060 36494
rect 38444 36482 38724 36484
rect 38444 36430 38446 36482
rect 38498 36430 38724 36482
rect 38444 36428 38724 36430
rect 38444 36418 38500 36428
rect 38556 36260 38612 36270
rect 38444 36258 38612 36260
rect 38444 36206 38558 36258
rect 38610 36206 38612 36258
rect 38444 36204 38612 36206
rect 37660 36036 37716 36046
rect 38444 36036 38500 36204
rect 38556 36194 38612 36204
rect 37324 35812 37380 35822
rect 37324 35718 37380 35756
rect 37436 35700 37492 35710
rect 37436 35606 37492 35644
rect 37436 35476 37492 35486
rect 37436 34802 37492 35420
rect 37660 34914 37716 35980
rect 37884 35980 38500 36036
rect 37884 35922 37940 35980
rect 37884 35870 37886 35922
rect 37938 35870 37940 35922
rect 37884 35858 37940 35870
rect 38108 35812 38164 35822
rect 37660 34862 37662 34914
rect 37714 34862 37716 34914
rect 37660 34850 37716 34862
rect 37996 35700 38052 35710
rect 37996 34914 38052 35644
rect 38108 35698 38164 35756
rect 38108 35646 38110 35698
rect 38162 35646 38164 35698
rect 38108 35634 38164 35646
rect 38444 35698 38500 35710
rect 38444 35646 38446 35698
rect 38498 35646 38500 35698
rect 37996 34862 37998 34914
rect 38050 34862 38052 34914
rect 37996 34850 38052 34862
rect 38332 35586 38388 35598
rect 38332 35534 38334 35586
rect 38386 35534 38388 35586
rect 38332 34916 38388 35534
rect 38444 35476 38500 35646
rect 38444 35410 38500 35420
rect 38556 35588 38612 35598
rect 38332 34850 38388 34860
rect 37436 34750 37438 34802
rect 37490 34750 37492 34802
rect 37436 34738 37492 34750
rect 36316 34190 36318 34242
rect 36370 34190 36372 34242
rect 36316 33908 36372 34190
rect 36988 34300 37268 34356
rect 37324 34690 37380 34702
rect 37324 34638 37326 34690
rect 37378 34638 37380 34690
rect 36316 33842 36372 33852
rect 36540 34130 36596 34142
rect 36540 34078 36542 34130
rect 36594 34078 36596 34130
rect 36540 33460 36596 34078
rect 36876 34132 36932 34142
rect 36876 34038 36932 34076
rect 36540 33394 36596 33404
rect 36988 33236 37044 34300
rect 37324 34244 37380 34638
rect 38332 34692 38388 34702
rect 38556 34692 38612 35532
rect 38332 34690 38612 34692
rect 38332 34638 38334 34690
rect 38386 34638 38612 34690
rect 38332 34636 38612 34638
rect 38332 34626 38388 34636
rect 38668 34356 38724 36428
rect 39004 36482 39620 36484
rect 39004 36430 39006 36482
rect 39058 36430 39620 36482
rect 39004 36428 39620 36430
rect 39004 36418 39060 36428
rect 38780 35700 38836 35710
rect 38780 35606 38836 35644
rect 39228 35700 39284 35710
rect 39228 35606 39284 35644
rect 39564 35026 39620 36428
rect 40572 36370 40628 38612
rect 41132 38050 41188 38062
rect 41132 37998 41134 38050
rect 41186 37998 41188 38050
rect 41132 37716 41188 37998
rect 41244 37938 41300 39676
rect 41244 37886 41246 37938
rect 41298 37886 41300 37938
rect 41244 37874 41300 37886
rect 41356 37716 41412 39900
rect 42364 39620 42420 40348
rect 42476 39620 42532 39630
rect 42364 39618 42532 39620
rect 42364 39566 42478 39618
rect 42530 39566 42532 39618
rect 42364 39564 42532 39566
rect 42476 39554 42532 39564
rect 42252 39508 42308 39518
rect 41468 39396 41524 39406
rect 41524 39340 41636 39396
rect 41468 39302 41524 39340
rect 41132 37660 41412 37716
rect 41468 38722 41524 38734
rect 41468 38670 41470 38722
rect 41522 38670 41524 38722
rect 41132 36932 41188 37660
rect 41468 37604 41524 38670
rect 41580 38724 41636 39340
rect 42252 39394 42308 39452
rect 42252 39342 42254 39394
rect 42306 39342 42308 39394
rect 42252 39172 42308 39342
rect 42588 39172 42644 40460
rect 42812 40450 42868 40460
rect 43036 40514 43092 40684
rect 43036 40462 43038 40514
rect 43090 40462 43092 40514
rect 43036 40450 43092 40462
rect 43260 40404 43316 40414
rect 43260 40310 43316 40348
rect 42700 40290 42756 40302
rect 42700 40238 42702 40290
rect 42754 40238 42756 40290
rect 42700 40180 42756 40238
rect 42700 40114 42756 40124
rect 43372 39620 43428 40684
rect 43484 40404 43540 41806
rect 43708 41860 43764 41916
rect 43820 41972 43876 41982
rect 43820 41878 43876 41916
rect 43708 41794 43764 41804
rect 43596 41748 43652 41758
rect 43596 41186 43652 41692
rect 44156 41636 44212 42030
rect 44380 42084 44436 42924
rect 44492 42196 44548 43652
rect 44604 42196 44660 42206
rect 44492 42194 44660 42196
rect 44492 42142 44606 42194
rect 44658 42142 44660 42194
rect 44492 42140 44660 42142
rect 44604 42130 44660 42140
rect 44828 42196 44884 42206
rect 44828 42102 44884 42140
rect 44380 42028 44548 42084
rect 44492 41970 44548 42028
rect 44492 41918 44494 41970
rect 44546 41918 44548 41970
rect 44492 41906 44548 41918
rect 44716 41636 44772 41646
rect 44156 41580 44324 41636
rect 44156 41412 44212 41422
rect 44156 41318 44212 41356
rect 43596 41134 43598 41186
rect 43650 41134 43652 41186
rect 43596 40628 43652 41134
rect 43932 41186 43988 41198
rect 43932 41134 43934 41186
rect 43986 41134 43988 41186
rect 43596 40562 43652 40572
rect 43708 40628 43764 40638
rect 43932 40628 43988 41134
rect 44268 40852 44324 41580
rect 43708 40626 43988 40628
rect 43708 40574 43710 40626
rect 43762 40574 43988 40626
rect 43708 40572 43988 40574
rect 44156 40628 44212 40638
rect 43708 40562 43764 40572
rect 44156 40534 44212 40572
rect 43484 40348 43652 40404
rect 43372 39564 43540 39620
rect 43148 39508 43204 39518
rect 43148 39414 43204 39452
rect 42812 39396 42868 39406
rect 42812 39394 43092 39396
rect 42812 39342 42814 39394
rect 42866 39342 43092 39394
rect 42812 39340 43092 39342
rect 42812 39330 42868 39340
rect 43036 39284 43092 39340
rect 43372 39394 43428 39406
rect 43372 39342 43374 39394
rect 43426 39342 43428 39394
rect 43372 39284 43428 39342
rect 43484 39396 43540 39564
rect 43596 39618 43652 40348
rect 44044 40292 44100 40302
rect 44044 40198 44100 40236
rect 43932 40180 43988 40190
rect 43820 40178 43988 40180
rect 43820 40126 43934 40178
rect 43986 40126 43988 40178
rect 43820 40124 43988 40126
rect 43708 39732 43764 39742
rect 43820 39732 43876 40124
rect 43932 40114 43988 40124
rect 43708 39730 43876 39732
rect 43708 39678 43710 39730
rect 43762 39678 43876 39730
rect 43708 39676 43876 39678
rect 43708 39666 43764 39676
rect 43596 39566 43598 39618
rect 43650 39566 43652 39618
rect 43596 39554 43652 39566
rect 43484 39340 43652 39396
rect 43036 39228 43428 39284
rect 42588 39116 42868 39172
rect 42252 39106 42308 39116
rect 42252 38948 42308 38958
rect 42028 38946 42308 38948
rect 42028 38894 42254 38946
rect 42306 38894 42308 38946
rect 42028 38892 42308 38894
rect 41916 38836 41972 38846
rect 41916 38742 41972 38780
rect 42028 38668 42084 38892
rect 42252 38882 42308 38892
rect 42812 38836 42868 39116
rect 42924 39060 42980 39070
rect 42924 38966 42980 39004
rect 43148 38836 43204 38846
rect 42812 38834 43204 38836
rect 42812 38782 43150 38834
rect 43202 38782 43204 38834
rect 42812 38780 43204 38782
rect 43148 38770 43204 38780
rect 41580 38658 41636 38668
rect 41804 38612 42084 38668
rect 42252 38724 42308 38734
rect 41804 38274 41860 38612
rect 41804 38222 41806 38274
rect 41858 38222 41860 38274
rect 41580 38052 41636 38062
rect 41580 37958 41636 37996
rect 41804 38052 41860 38222
rect 41804 37986 41860 37996
rect 42140 37828 42196 37838
rect 41804 37826 42196 37828
rect 41804 37774 42142 37826
rect 42194 37774 42196 37826
rect 41804 37772 42196 37774
rect 41468 37548 41636 37604
rect 41468 37378 41524 37390
rect 41468 37326 41470 37378
rect 41522 37326 41524 37378
rect 41132 36876 41412 36932
rect 41132 36708 41188 36718
rect 40684 36484 40740 36494
rect 41132 36484 41188 36652
rect 40684 36482 41188 36484
rect 40684 36430 40686 36482
rect 40738 36430 41188 36482
rect 40684 36428 41188 36430
rect 40684 36418 40740 36428
rect 40572 36318 40574 36370
rect 40626 36318 40628 36370
rect 40572 36306 40628 36318
rect 41132 36370 41188 36428
rect 41132 36318 41134 36370
rect 41186 36318 41188 36370
rect 41132 36306 41188 36318
rect 40348 36260 40404 36270
rect 40124 36258 40404 36260
rect 40124 36206 40350 36258
rect 40402 36206 40404 36258
rect 40124 36204 40404 36206
rect 39564 34974 39566 35026
rect 39618 34974 39620 35026
rect 39564 34962 39620 34974
rect 40012 35812 40068 35822
rect 40012 35586 40068 35756
rect 40012 35534 40014 35586
rect 40066 35534 40068 35586
rect 40012 35026 40068 35534
rect 40012 34974 40014 35026
rect 40066 34974 40068 35026
rect 40012 34962 40068 34974
rect 40124 35700 40180 36204
rect 40348 36194 40404 36204
rect 41356 36258 41412 36876
rect 41468 36596 41524 37326
rect 41468 36502 41524 36540
rect 41580 36932 41636 37548
rect 41804 37268 41860 37772
rect 42140 37762 42196 37772
rect 41804 37266 41972 37268
rect 41804 37214 41806 37266
rect 41858 37214 41972 37266
rect 41804 37212 41972 37214
rect 41804 37202 41860 37212
rect 41580 36482 41636 36876
rect 41580 36430 41582 36482
rect 41634 36430 41636 36482
rect 41580 36418 41636 36430
rect 41692 37154 41748 37166
rect 41692 37102 41694 37154
rect 41746 37102 41748 37154
rect 41356 36206 41358 36258
rect 41410 36206 41412 36258
rect 41356 36148 41412 36206
rect 41356 36082 41412 36092
rect 41692 35924 41748 37102
rect 41916 36482 41972 37212
rect 42252 36820 42308 38668
rect 42700 38052 42756 38062
rect 42476 37940 42532 37950
rect 42476 37846 42532 37884
rect 42700 37938 42756 37996
rect 42700 37886 42702 37938
rect 42754 37886 42756 37938
rect 42700 37874 42756 37886
rect 42588 37826 42644 37838
rect 42588 37774 42590 37826
rect 42642 37774 42644 37826
rect 42588 37604 42644 37774
rect 42364 37548 42644 37604
rect 43260 37826 43316 37838
rect 43260 37774 43262 37826
rect 43314 37774 43316 37826
rect 42364 37266 42420 37548
rect 42364 37214 42366 37266
rect 42418 37214 42420 37266
rect 42364 37202 42420 37214
rect 42252 36764 42532 36820
rect 41916 36430 41918 36482
rect 41970 36430 41972 36482
rect 41916 36418 41972 36430
rect 42028 36596 42084 36606
rect 42028 36370 42084 36540
rect 42028 36318 42030 36370
rect 42082 36318 42084 36370
rect 42028 36306 42084 36318
rect 42476 36484 42532 36764
rect 43260 36708 43316 37774
rect 43372 37604 43428 39228
rect 43596 38388 43652 39340
rect 43708 39394 43764 39406
rect 43708 39342 43710 39394
rect 43762 39342 43764 39394
rect 43708 38836 43764 39342
rect 44268 38836 44324 40796
rect 44716 40740 44772 41580
rect 44940 41298 44996 43932
rect 45052 43764 45108 43774
rect 45052 42754 45108 43708
rect 45388 43426 45444 45054
rect 45388 43374 45390 43426
rect 45442 43374 45444 43426
rect 45388 42980 45444 43374
rect 45388 42886 45444 42924
rect 45052 42702 45054 42754
rect 45106 42702 45108 42754
rect 45052 42690 45108 42702
rect 45164 42532 45220 42542
rect 44940 41246 44942 41298
rect 44994 41246 44996 41298
rect 44940 41234 44996 41246
rect 45052 41860 45108 41870
rect 44716 40626 44772 40684
rect 44716 40574 44718 40626
rect 44770 40574 44772 40626
rect 44716 40562 44772 40574
rect 44604 40404 44660 40414
rect 44604 40310 44660 40348
rect 44940 40402 44996 40414
rect 44940 40350 44942 40402
rect 44994 40350 44996 40402
rect 44940 40292 44996 40350
rect 44940 40226 44996 40236
rect 44828 39060 44884 39070
rect 45052 39060 45108 41804
rect 45164 41748 45220 42476
rect 45276 42530 45332 42542
rect 45276 42478 45278 42530
rect 45330 42478 45332 42530
rect 45276 41972 45332 42478
rect 45276 41906 45332 41916
rect 45276 41748 45332 41758
rect 45164 41746 45332 41748
rect 45164 41694 45278 41746
rect 45330 41694 45332 41746
rect 45164 41692 45332 41694
rect 45276 41682 45332 41692
rect 45500 41636 45556 45838
rect 45724 45220 45780 49200
rect 46396 45892 46452 49200
rect 51436 46900 51492 46910
rect 46396 45826 46452 45836
rect 47404 46228 47460 46238
rect 45724 45154 45780 45164
rect 46060 45778 46116 45790
rect 46060 45726 46062 45778
rect 46114 45726 46116 45778
rect 45836 44210 45892 44222
rect 45836 44158 45838 44210
rect 45890 44158 45892 44210
rect 45836 43708 45892 44158
rect 45724 43652 45892 43708
rect 45612 43540 45668 43550
rect 45612 43446 45668 43484
rect 45724 42196 45780 43652
rect 45836 43586 45892 43596
rect 46060 43650 46116 45726
rect 46732 45780 46788 45790
rect 46732 45686 46788 45724
rect 47404 45778 47460 46172
rect 49868 46172 50260 46228
rect 47404 45726 47406 45778
rect 47458 45726 47460 45778
rect 47404 45714 47460 45726
rect 47740 45778 47796 45790
rect 47740 45726 47742 45778
rect 47794 45726 47796 45778
rect 46284 45668 46340 45678
rect 46284 45106 46340 45612
rect 46396 45666 46452 45678
rect 46396 45614 46398 45666
rect 46450 45614 46452 45666
rect 46396 45332 46452 45614
rect 46396 45266 46452 45276
rect 46284 45054 46286 45106
rect 46338 45054 46340 45106
rect 46284 45042 46340 45054
rect 47628 45106 47684 45118
rect 47628 45054 47630 45106
rect 47682 45054 47684 45106
rect 47628 44996 47684 45054
rect 46060 43598 46062 43650
rect 46114 43598 46116 43650
rect 46060 43540 46116 43598
rect 46060 43474 46116 43484
rect 46284 44322 46340 44334
rect 46284 44270 46286 44322
rect 46338 44270 46340 44322
rect 46284 43762 46340 44270
rect 46284 43710 46286 43762
rect 46338 43710 46340 43762
rect 45948 43428 46004 43438
rect 45836 42532 45892 42542
rect 45836 42438 45892 42476
rect 45948 42196 46004 43372
rect 46284 43204 46340 43710
rect 47292 44322 47348 44334
rect 47292 44270 47294 44322
rect 47346 44270 47348 44322
rect 46956 43652 47012 43662
rect 46508 43538 46564 43550
rect 46508 43486 46510 43538
rect 46562 43486 46564 43538
rect 46508 43428 46564 43486
rect 46956 43538 47012 43596
rect 47292 43652 47348 44270
rect 47292 43650 47572 43652
rect 47292 43598 47294 43650
rect 47346 43598 47572 43650
rect 47292 43596 47572 43598
rect 47292 43586 47348 43596
rect 46956 43486 46958 43538
rect 47010 43486 47012 43538
rect 46956 43474 47012 43486
rect 46284 43138 46340 43148
rect 46396 43372 46508 43428
rect 46396 42980 46452 43372
rect 46508 43362 46564 43372
rect 47180 43426 47236 43438
rect 47180 43374 47182 43426
rect 47234 43374 47236 43426
rect 46172 42924 46452 42980
rect 46172 42754 46228 42924
rect 46172 42702 46174 42754
rect 46226 42702 46228 42754
rect 46172 42690 46228 42702
rect 47068 42866 47124 42878
rect 47068 42814 47070 42866
rect 47122 42814 47124 42866
rect 45948 42140 46228 42196
rect 45724 42130 45780 42140
rect 45388 41580 45556 41636
rect 45612 41972 45668 41982
rect 45836 41972 45892 41982
rect 45612 41970 45892 41972
rect 45612 41918 45614 41970
rect 45666 41918 45838 41970
rect 45890 41918 45892 41970
rect 45612 41916 45892 41918
rect 45388 40626 45444 41580
rect 45500 41300 45556 41310
rect 45612 41300 45668 41916
rect 45836 41906 45892 41916
rect 45948 41972 46004 41982
rect 45724 41412 45780 41422
rect 45724 41318 45780 41356
rect 45948 41410 46004 41916
rect 45948 41358 45950 41410
rect 46002 41358 46004 41410
rect 45948 41346 46004 41358
rect 45500 41298 45668 41300
rect 45500 41246 45502 41298
rect 45554 41246 45668 41298
rect 45500 41244 45668 41246
rect 45836 41300 45892 41310
rect 45500 41234 45556 41244
rect 45388 40574 45390 40626
rect 45442 40574 45444 40626
rect 45388 40562 45444 40574
rect 45836 40628 45892 41244
rect 45948 40628 46004 40638
rect 45836 40572 45948 40628
rect 45948 40534 46004 40572
rect 45724 39396 45780 39406
rect 45164 39060 45220 39070
rect 45052 39058 45220 39060
rect 45052 39006 45166 39058
rect 45218 39006 45220 39058
rect 45052 39004 45220 39006
rect 44828 38966 44884 39004
rect 45164 38994 45220 39004
rect 43708 38780 44324 38836
rect 44268 38668 44324 38780
rect 45500 38946 45556 38958
rect 45500 38894 45502 38946
rect 45554 38894 45556 38946
rect 44268 38612 44436 38668
rect 43372 37378 43428 37548
rect 43484 38052 43540 38062
rect 43484 37492 43540 37996
rect 43596 38050 43652 38332
rect 43596 37998 43598 38050
rect 43650 37998 43652 38050
rect 43596 37986 43652 37998
rect 44156 37938 44212 37950
rect 44156 37886 44158 37938
rect 44210 37886 44212 37938
rect 43820 37828 43876 37838
rect 43820 37734 43876 37772
rect 44044 37828 44100 37838
rect 43932 37492 43988 37502
rect 43484 37490 43988 37492
rect 43484 37438 43486 37490
rect 43538 37438 43934 37490
rect 43986 37438 43988 37490
rect 43484 37436 43988 37438
rect 43484 37426 43540 37436
rect 43932 37426 43988 37436
rect 43372 37326 43374 37378
rect 43426 37326 43428 37378
rect 43372 37314 43428 37326
rect 43708 37266 43764 37278
rect 43708 37214 43710 37266
rect 43762 37214 43764 37266
rect 43708 37156 43764 37214
rect 44044 37156 44100 37772
rect 44156 37604 44212 37886
rect 44156 37538 44212 37548
rect 43708 37090 43764 37100
rect 43820 37100 44100 37156
rect 44268 37378 44324 37390
rect 44268 37326 44270 37378
rect 44322 37326 44324 37378
rect 43260 36642 43316 36652
rect 42476 36428 43540 36484
rect 41244 35868 41748 35924
rect 42252 36258 42308 36270
rect 42252 36206 42254 36258
rect 42306 36206 42308 36258
rect 41244 35812 41300 35868
rect 39900 34916 39956 34926
rect 39900 34692 39956 34860
rect 40124 34914 40180 35644
rect 40908 35700 40964 35738
rect 41244 35718 41300 35756
rect 40908 35634 40964 35644
rect 41132 35586 41188 35598
rect 41132 35534 41134 35586
rect 41186 35534 41188 35586
rect 41132 34916 41188 35534
rect 42252 35364 42308 36206
rect 42476 35810 42532 36428
rect 43484 36370 43540 36428
rect 43484 36318 43486 36370
rect 43538 36318 43540 36370
rect 43484 36306 43540 36318
rect 43596 36372 43652 36382
rect 43596 36278 43652 36316
rect 43260 36260 43316 36270
rect 43260 36258 43428 36260
rect 43260 36206 43262 36258
rect 43314 36206 43428 36258
rect 43260 36204 43428 36206
rect 43260 36194 43316 36204
rect 42476 35758 42478 35810
rect 42530 35758 42532 35810
rect 42476 35746 42532 35758
rect 42588 35812 42644 35822
rect 42588 35810 43316 35812
rect 42588 35758 42590 35810
rect 42642 35758 43316 35810
rect 42588 35756 43316 35758
rect 42588 35746 42644 35756
rect 43260 35698 43316 35756
rect 43260 35646 43262 35698
rect 43314 35646 43316 35698
rect 43260 35634 43316 35646
rect 43148 35586 43204 35598
rect 43148 35534 43150 35586
rect 43202 35534 43204 35586
rect 43148 35364 43204 35534
rect 42252 35308 43204 35364
rect 41356 34916 41412 34926
rect 40124 34862 40126 34914
rect 40178 34862 40180 34914
rect 40124 34850 40180 34862
rect 40908 34914 41412 34916
rect 40908 34862 41358 34914
rect 41410 34862 41412 34914
rect 40908 34860 41412 34862
rect 38780 34356 38836 34366
rect 38668 34354 38836 34356
rect 38668 34302 38782 34354
rect 38834 34302 38836 34354
rect 38668 34300 38836 34302
rect 37324 34242 37940 34244
rect 37324 34190 37326 34242
rect 37378 34190 37940 34242
rect 37324 34188 37940 34190
rect 37324 34178 37380 34188
rect 37100 34130 37156 34142
rect 37100 34078 37102 34130
rect 37154 34078 37156 34130
rect 37100 34020 37156 34078
rect 37884 34132 37940 34188
rect 38444 34132 38500 34142
rect 37884 34130 38500 34132
rect 37884 34078 37886 34130
rect 37938 34078 38446 34130
rect 38498 34078 38500 34130
rect 37884 34076 38500 34078
rect 37884 34066 37940 34076
rect 38444 34066 38500 34076
rect 37100 33954 37156 33964
rect 37212 34018 37268 34030
rect 37212 33966 37214 34018
rect 37266 33966 37268 34018
rect 37100 33460 37156 33470
rect 37212 33460 37268 33966
rect 37660 34020 37716 34030
rect 37660 33926 37716 33964
rect 38780 34020 38836 34300
rect 38780 33954 38836 33964
rect 39004 34242 39060 34254
rect 39004 34190 39006 34242
rect 39058 34190 39060 34242
rect 39004 34132 39060 34190
rect 39900 34244 39956 34636
rect 40012 34244 40068 34254
rect 39900 34242 40068 34244
rect 39900 34190 40014 34242
rect 40066 34190 40068 34242
rect 39900 34188 40068 34190
rect 40012 34178 40068 34188
rect 38220 33908 38276 33918
rect 38220 33906 38612 33908
rect 38220 33854 38222 33906
rect 38274 33854 38612 33906
rect 38220 33852 38612 33854
rect 38220 33842 38276 33852
rect 38220 33684 38276 33694
rect 37212 33404 37604 33460
rect 37100 33366 37156 33404
rect 37324 33236 37380 33246
rect 36988 33234 37380 33236
rect 36988 33182 37326 33234
rect 37378 33182 37380 33234
rect 36988 33180 37380 33182
rect 37324 32340 37380 33180
rect 37548 32786 37604 33404
rect 37548 32734 37550 32786
rect 37602 32734 37604 32786
rect 37548 32722 37604 32734
rect 37660 32564 37716 32574
rect 37660 32470 37716 32508
rect 37772 32562 37828 32574
rect 37772 32510 37774 32562
rect 37826 32510 37828 32562
rect 37772 32340 37828 32510
rect 38220 32562 38276 33628
rect 38556 33348 38612 33852
rect 38668 33906 38724 33918
rect 38668 33854 38670 33906
rect 38722 33854 38724 33906
rect 38668 33684 38724 33854
rect 38668 33618 38724 33628
rect 39004 33572 39060 34076
rect 40348 34132 40404 34142
rect 40908 34132 40964 34860
rect 41356 34850 41412 34860
rect 40348 34130 40964 34132
rect 40348 34078 40350 34130
rect 40402 34078 40910 34130
rect 40962 34078 40964 34130
rect 40348 34076 40964 34078
rect 40348 34066 40404 34076
rect 40908 34066 40964 34076
rect 41132 34692 41188 34702
rect 41132 34130 41188 34636
rect 41132 34078 41134 34130
rect 41186 34078 41188 34130
rect 41132 34066 41188 34078
rect 41244 34690 41300 34702
rect 41244 34638 41246 34690
rect 41298 34638 41300 34690
rect 41244 34132 41300 34638
rect 41580 34690 41636 34702
rect 41580 34638 41582 34690
rect 41634 34638 41636 34690
rect 41580 34356 41636 34638
rect 43148 34692 43204 35308
rect 43260 34916 43316 34926
rect 43372 34916 43428 36204
rect 43820 36148 43876 37100
rect 44268 37044 44324 37326
rect 43932 36988 44324 37044
rect 43932 36372 43988 36988
rect 44380 36932 44436 38612
rect 44940 37828 44996 37838
rect 44940 37734 44996 37772
rect 45500 37828 45556 38894
rect 45724 38276 45780 39340
rect 45948 39396 46004 39406
rect 45948 39302 46004 39340
rect 46060 39060 46116 39070
rect 45836 38836 45892 38846
rect 45836 38742 45892 38780
rect 46060 38834 46116 39004
rect 46060 38782 46062 38834
rect 46114 38782 46116 38834
rect 46060 38770 46116 38782
rect 46172 38668 46228 42140
rect 47068 42082 47124 42814
rect 47180 42756 47236 43374
rect 47516 43428 47572 43596
rect 47628 43650 47684 44940
rect 47740 44660 47796 45726
rect 49644 45780 49700 45790
rect 49868 45780 49924 46172
rect 49644 45778 49924 45780
rect 49644 45726 49646 45778
rect 49698 45726 49924 45778
rect 49644 45724 49924 45726
rect 49644 45714 49700 45724
rect 48076 45668 48132 45678
rect 48076 45666 48356 45668
rect 48076 45614 48078 45666
rect 48130 45614 48356 45666
rect 48076 45612 48356 45614
rect 48076 45602 48132 45612
rect 47740 44594 47796 44604
rect 48188 44660 48244 44670
rect 48076 44210 48132 44222
rect 48076 44158 48078 44210
rect 48130 44158 48132 44210
rect 48076 43708 48132 44158
rect 47628 43598 47630 43650
rect 47682 43598 47684 43650
rect 47628 43586 47684 43598
rect 47852 43652 48132 43708
rect 47740 43428 47796 43438
rect 47516 43426 47796 43428
rect 47516 43374 47742 43426
rect 47794 43374 47796 43426
rect 47516 43372 47796 43374
rect 47740 43362 47796 43372
rect 47852 42756 47908 43652
rect 47964 43540 48020 43550
rect 47964 43446 48020 43484
rect 47180 42690 47236 42700
rect 47516 42754 47908 42756
rect 47516 42702 47854 42754
rect 47906 42702 47908 42754
rect 47516 42700 47908 42702
rect 47068 42030 47070 42082
rect 47122 42030 47124 42082
rect 46508 41972 46564 41982
rect 46508 41858 46564 41916
rect 46508 41806 46510 41858
rect 46562 41806 46564 41858
rect 46508 41794 46564 41806
rect 46620 41970 46676 41982
rect 46620 41918 46622 41970
rect 46674 41918 46676 41970
rect 46620 41412 46676 41918
rect 46620 41346 46676 41356
rect 47068 41188 47124 42030
rect 47516 41298 47572 42700
rect 47852 42690 47908 42700
rect 47964 42532 48020 42542
rect 47964 42082 48020 42476
rect 47964 42030 47966 42082
rect 48018 42030 48020 42082
rect 47964 42018 48020 42030
rect 48076 42084 48132 42094
rect 48076 41990 48132 42028
rect 47516 41246 47518 41298
rect 47570 41246 47572 41298
rect 47516 41234 47572 41246
rect 48076 41300 48132 41310
rect 48188 41300 48244 44604
rect 48300 43708 48356 45612
rect 48412 45666 48468 45678
rect 48412 45614 48414 45666
rect 48466 45614 48468 45666
rect 48412 44884 48468 45614
rect 48748 45668 48804 45678
rect 48748 45574 48804 45612
rect 49084 45666 49140 45678
rect 49084 45614 49086 45666
rect 49138 45614 49140 45666
rect 49084 45332 49140 45614
rect 48412 44818 48468 44828
rect 48972 45276 49084 45332
rect 48860 44436 48916 44446
rect 48860 44322 48916 44380
rect 48860 44270 48862 44322
rect 48914 44270 48916 44322
rect 48860 44258 48916 44270
rect 48972 44324 49028 45276
rect 49084 45266 49140 45276
rect 49868 45106 49924 45724
rect 49868 45054 49870 45106
rect 49922 45054 49924 45106
rect 49868 45042 49924 45054
rect 49980 46002 50036 46014
rect 49980 45950 49982 46002
rect 50034 45950 50036 46002
rect 49084 44996 49140 45006
rect 49084 44994 49476 44996
rect 49084 44942 49086 44994
rect 49138 44942 49476 44994
rect 49084 44940 49476 44942
rect 49084 44930 49140 44940
rect 49420 44772 49476 44940
rect 49980 44772 50036 45950
rect 49420 44716 49924 44772
rect 49532 44436 49588 44446
rect 49084 44324 49140 44334
rect 48972 44322 49364 44324
rect 48972 44270 49086 44322
rect 49138 44270 49364 44322
rect 48972 44268 49364 44270
rect 49084 44258 49140 44268
rect 49084 44100 49140 44110
rect 48300 43652 48468 43708
rect 48300 41972 48356 41982
rect 48300 41878 48356 41916
rect 48412 41636 48468 43652
rect 48860 43652 48916 43662
rect 48860 43650 49028 43652
rect 48860 43598 48862 43650
rect 48914 43598 49028 43650
rect 48860 43596 49028 43598
rect 48860 43586 48916 43596
rect 48748 43538 48804 43550
rect 48748 43486 48750 43538
rect 48802 43486 48804 43538
rect 48748 43428 48804 43486
rect 48748 43362 48804 43372
rect 48748 43204 48804 43214
rect 48748 42754 48804 43148
rect 48748 42702 48750 42754
rect 48802 42702 48804 42754
rect 48748 42690 48804 42702
rect 48860 42532 48916 42542
rect 48860 41972 48916 42476
rect 48972 42420 49028 43596
rect 49084 43650 49140 44044
rect 49084 43598 49086 43650
rect 49138 43598 49140 43650
rect 49084 43586 49140 43598
rect 49308 43540 49364 44268
rect 49308 43446 49364 43484
rect 49532 43764 49588 44380
rect 49532 43538 49588 43708
rect 49532 43486 49534 43538
rect 49586 43486 49588 43538
rect 49532 43474 49588 43486
rect 49756 44324 49812 44334
rect 49756 43538 49812 44268
rect 49756 43486 49758 43538
rect 49810 43486 49812 43538
rect 49756 43474 49812 43486
rect 49196 42868 49252 42878
rect 49196 42866 49476 42868
rect 49196 42814 49198 42866
rect 49250 42814 49476 42866
rect 49196 42812 49476 42814
rect 49196 42802 49252 42812
rect 48972 42354 49028 42364
rect 49420 42196 49476 42812
rect 49532 42756 49588 42766
rect 49532 42662 49588 42700
rect 49868 42308 49924 44716
rect 49980 44706 50036 44716
rect 50092 45890 50148 45902
rect 50092 45838 50094 45890
rect 50146 45838 50148 45890
rect 50092 44548 50148 45838
rect 50092 44482 50148 44492
rect 49980 44434 50036 44446
rect 49980 44382 49982 44434
rect 50034 44382 50036 44434
rect 49980 43652 50036 44382
rect 50204 44324 50260 46172
rect 51436 46004 51492 46844
rect 51436 45890 51492 45948
rect 53788 46004 53844 46014
rect 53788 45910 53844 45948
rect 51436 45838 51438 45890
rect 51490 45838 51492 45890
rect 51436 45826 51492 45838
rect 52108 45890 52164 45902
rect 52108 45838 52110 45890
rect 52162 45838 52164 45890
rect 51212 45666 51268 45678
rect 51212 45614 51214 45666
rect 51266 45614 51268 45666
rect 50556 45500 50820 45510
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50556 45434 50820 45444
rect 50988 45218 51044 45230
rect 50988 45166 50990 45218
rect 51042 45166 51044 45218
rect 50876 44434 50932 44446
rect 50876 44382 50878 44434
rect 50930 44382 50932 44434
rect 50204 44230 50260 44268
rect 50652 44322 50708 44334
rect 50652 44270 50654 44322
rect 50706 44270 50708 44322
rect 50652 44212 50708 44270
rect 50428 44156 50708 44212
rect 49980 42644 50036 43596
rect 50092 43764 50148 43774
rect 50092 42866 50148 43708
rect 50092 42814 50094 42866
rect 50146 42814 50148 42866
rect 50092 42802 50148 42814
rect 50204 43314 50260 43326
rect 50204 43262 50206 43314
rect 50258 43262 50260 43314
rect 49980 42588 50148 42644
rect 49868 42252 50036 42308
rect 49420 42140 49812 42196
rect 48412 41570 48468 41580
rect 48748 41970 48916 41972
rect 48748 41918 48862 41970
rect 48914 41918 48916 41970
rect 48748 41916 48916 41918
rect 48076 41298 48244 41300
rect 48076 41246 48078 41298
rect 48130 41246 48244 41298
rect 48076 41244 48244 41246
rect 48076 41234 48132 41244
rect 46844 41186 47124 41188
rect 46844 41134 47070 41186
rect 47122 41134 47124 41186
rect 46844 41132 47124 41134
rect 46620 41074 46676 41086
rect 46620 41022 46622 41074
rect 46674 41022 46676 41074
rect 46396 40964 46452 40974
rect 46396 40962 46564 40964
rect 46396 40910 46398 40962
rect 46450 40910 46564 40962
rect 46396 40908 46564 40910
rect 46396 40898 46452 40908
rect 46284 40516 46340 40526
rect 46284 40422 46340 40460
rect 46508 40404 46564 40908
rect 46620 40628 46676 41022
rect 46620 40572 46788 40628
rect 46620 40404 46676 40414
rect 46508 40402 46676 40404
rect 46508 40350 46622 40402
rect 46674 40350 46676 40402
rect 46508 40348 46676 40350
rect 46620 40338 46676 40348
rect 46284 39620 46340 39630
rect 46732 39620 46788 40572
rect 46844 40402 46900 41132
rect 47068 41122 47124 41132
rect 48748 41186 48804 41916
rect 48860 41906 48916 41916
rect 49196 42082 49252 42094
rect 49196 42030 49198 42082
rect 49250 42030 49252 42082
rect 49196 41412 49252 42030
rect 49756 42082 49812 42140
rect 49756 42030 49758 42082
rect 49810 42030 49812 42082
rect 49644 41860 49700 41870
rect 49196 41356 49476 41412
rect 48748 41134 48750 41186
rect 48802 41134 48804 41186
rect 48748 41122 48804 41134
rect 49308 41186 49364 41198
rect 49308 41134 49310 41186
rect 49362 41134 49364 41186
rect 49308 41076 49364 41134
rect 48860 40962 48916 40974
rect 48860 40910 48862 40962
rect 48914 40910 48916 40962
rect 47404 40628 47460 40638
rect 46844 40350 46846 40402
rect 46898 40350 46900 40402
rect 46844 40338 46900 40350
rect 47180 40514 47236 40526
rect 47180 40462 47182 40514
rect 47234 40462 47236 40514
rect 46956 39956 47012 39966
rect 46732 39564 46900 39620
rect 46284 39526 46340 39564
rect 46620 39508 46676 39518
rect 46508 39506 46676 39508
rect 46508 39454 46622 39506
rect 46674 39454 46676 39506
rect 46508 39452 46676 39454
rect 46508 38948 46564 39452
rect 46620 39442 46676 39452
rect 46732 39394 46788 39406
rect 46732 39342 46734 39394
rect 46786 39342 46788 39394
rect 46732 39284 46788 39342
rect 46732 39218 46788 39228
rect 46396 38722 46452 38734
rect 46396 38670 46398 38722
rect 46450 38670 46452 38722
rect 45724 38210 45780 38220
rect 45948 38612 46340 38668
rect 45948 38162 46004 38612
rect 45948 38110 45950 38162
rect 46002 38110 46004 38162
rect 45948 38098 46004 38110
rect 46284 38164 46340 38612
rect 46396 38500 46452 38670
rect 46396 38434 46452 38444
rect 46284 38108 46452 38164
rect 45500 37762 45556 37772
rect 46284 37938 46340 37950
rect 46284 37886 46286 37938
rect 46338 37886 46340 37938
rect 46284 37716 46340 37886
rect 46396 37938 46452 38108
rect 46396 37886 46398 37938
rect 46450 37886 46452 37938
rect 46396 37874 46452 37886
rect 46508 37716 46564 38892
rect 46732 39060 46788 39070
rect 46732 38946 46788 39004
rect 46732 38894 46734 38946
rect 46786 38894 46788 38946
rect 46732 38836 46788 38894
rect 46732 38770 46788 38780
rect 46844 38668 46900 39564
rect 46956 39618 47012 39900
rect 46956 39566 46958 39618
rect 47010 39566 47012 39618
rect 46956 39554 47012 39566
rect 47180 39396 47236 40462
rect 47404 40402 47460 40572
rect 47404 40350 47406 40402
rect 47458 40350 47460 40402
rect 47404 40338 47460 40350
rect 48860 39620 48916 40910
rect 49084 40964 49140 40974
rect 49084 40870 49140 40908
rect 49308 40628 49364 41020
rect 49308 40562 49364 40572
rect 49420 41074 49476 41356
rect 49644 41186 49700 41804
rect 49644 41134 49646 41186
rect 49698 41134 49700 41186
rect 49644 41122 49700 41134
rect 49420 41022 49422 41074
rect 49474 41022 49476 41074
rect 49308 40292 49364 40302
rect 49308 40198 49364 40236
rect 48860 39554 48916 39564
rect 47292 39396 47348 39406
rect 47180 39394 47348 39396
rect 47180 39342 47294 39394
rect 47346 39342 47348 39394
rect 47180 39340 47348 39342
rect 47292 39284 47348 39340
rect 47292 39218 47348 39228
rect 47068 38948 47124 38958
rect 47068 38854 47124 38892
rect 49420 38948 49476 41022
rect 49532 40852 49588 40862
rect 49532 40404 49588 40796
rect 49532 40402 49700 40404
rect 49532 40350 49534 40402
rect 49586 40350 49700 40402
rect 49532 40348 49700 40350
rect 49532 40338 49588 40348
rect 49644 39730 49700 40348
rect 49644 39678 49646 39730
rect 49698 39678 49700 39730
rect 49644 39666 49700 39678
rect 49420 38882 49476 38892
rect 49196 38834 49252 38846
rect 49196 38782 49198 38834
rect 49250 38782 49252 38834
rect 47740 38724 47796 38734
rect 46844 38612 47124 38668
rect 46620 38388 46676 38398
rect 46620 38050 46676 38332
rect 46620 37998 46622 38050
rect 46674 37998 46676 38050
rect 46620 37986 46676 37998
rect 46284 37660 46564 37716
rect 47068 37938 47124 38612
rect 47068 37886 47070 37938
rect 47122 37886 47124 37938
rect 44828 37604 44884 37614
rect 44716 37156 44772 37166
rect 44716 37062 44772 37100
rect 44044 36876 44772 36932
rect 44044 36482 44100 36876
rect 44044 36430 44046 36482
rect 44098 36430 44100 36482
rect 44044 36418 44100 36430
rect 44156 36708 44212 36718
rect 43932 36306 43988 36316
rect 44156 36258 44212 36652
rect 44380 36484 44436 36494
rect 44380 36390 44436 36428
rect 44156 36206 44158 36258
rect 44210 36206 44212 36258
rect 43820 36092 44100 36148
rect 43932 35700 43988 35710
rect 43596 35698 43988 35700
rect 43596 35646 43934 35698
rect 43986 35646 43988 35698
rect 43596 35644 43988 35646
rect 43260 34914 43428 34916
rect 43260 34862 43262 34914
rect 43314 34862 43428 34914
rect 43260 34860 43428 34862
rect 43484 35474 43540 35486
rect 43484 35422 43486 35474
rect 43538 35422 43540 35474
rect 43260 34850 43316 34860
rect 43372 34692 43428 34702
rect 43148 34690 43428 34692
rect 43148 34638 43374 34690
rect 43426 34638 43428 34690
rect 43148 34636 43428 34638
rect 43372 34626 43428 34636
rect 41244 34066 41300 34076
rect 41356 34300 41580 34356
rect 41356 34130 41412 34300
rect 41580 34290 41636 34300
rect 42252 34356 42308 34366
rect 42812 34356 42868 34366
rect 43260 34356 43316 34366
rect 43484 34356 43540 35422
rect 42252 34354 42532 34356
rect 42252 34302 42254 34354
rect 42306 34302 42532 34354
rect 42252 34300 42532 34302
rect 42252 34290 42308 34300
rect 41356 34078 41358 34130
rect 41410 34078 41412 34130
rect 41356 34066 41412 34078
rect 41804 34132 41860 34142
rect 42028 34132 42084 34142
rect 41804 34130 42084 34132
rect 41804 34078 41806 34130
rect 41858 34078 42030 34130
rect 42082 34078 42084 34130
rect 41804 34076 42084 34078
rect 41804 34066 41860 34076
rect 42028 34066 42084 34076
rect 42252 34132 42308 34142
rect 42252 34038 42308 34076
rect 40124 34018 40180 34030
rect 40124 33966 40126 34018
rect 40178 33966 40180 34018
rect 40124 33796 40180 33966
rect 40124 33730 40180 33740
rect 41020 33796 41076 33806
rect 39564 33572 39620 33582
rect 39004 33570 39620 33572
rect 39004 33518 39566 33570
rect 39618 33518 39620 33570
rect 39004 33516 39620 33518
rect 39564 33506 39620 33516
rect 39676 33460 39732 33470
rect 39676 33366 39732 33404
rect 38668 33348 38724 33358
rect 38556 33346 38724 33348
rect 38556 33294 38670 33346
rect 38722 33294 38724 33346
rect 38556 33292 38724 33294
rect 38668 33282 38724 33292
rect 41020 33346 41076 33740
rect 41132 33572 41188 33582
rect 41132 33570 41636 33572
rect 41132 33518 41134 33570
rect 41186 33518 41636 33570
rect 41132 33516 41636 33518
rect 41132 33506 41188 33516
rect 41020 33294 41022 33346
rect 41074 33294 41076 33346
rect 41020 33282 41076 33294
rect 39004 33122 39060 33134
rect 39004 33070 39006 33122
rect 39058 33070 39060 33122
rect 38220 32510 38222 32562
rect 38274 32510 38276 32562
rect 38220 32498 38276 32510
rect 38892 32900 38948 32910
rect 38892 32562 38948 32844
rect 38892 32510 38894 32562
rect 38946 32510 38948 32562
rect 38892 32498 38948 32510
rect 37324 32284 37828 32340
rect 37884 32452 37940 32462
rect 36092 31892 36148 31902
rect 36092 31798 36148 31836
rect 36988 31890 37044 31902
rect 36988 31838 36990 31890
rect 37042 31838 37044 31890
rect 36204 31780 36260 31790
rect 36204 31666 36260 31724
rect 36204 31614 36206 31666
rect 36258 31614 36260 31666
rect 36204 31602 36260 31614
rect 36428 31668 36484 31678
rect 36428 31574 36484 31612
rect 35868 30930 35924 30940
rect 36092 31108 36148 31118
rect 36092 30996 36148 31052
rect 36988 31106 37044 31838
rect 37100 31780 37156 31790
rect 37100 31666 37156 31724
rect 37100 31614 37102 31666
rect 37154 31614 37156 31666
rect 37100 31602 37156 31614
rect 37212 31668 37268 31678
rect 37212 31220 37268 31612
rect 37324 31666 37380 31678
rect 37324 31614 37326 31666
rect 37378 31614 37380 31666
rect 37324 31556 37380 31614
rect 37324 31490 37380 31500
rect 37212 31126 37268 31164
rect 36988 31054 36990 31106
rect 37042 31054 37044 31106
rect 36988 31042 37044 31054
rect 36092 30994 36372 30996
rect 36092 30942 36094 30994
rect 36146 30942 36372 30994
rect 36092 30940 36372 30942
rect 36092 30930 36148 30940
rect 35420 30882 35476 30894
rect 35420 30830 35422 30882
rect 35474 30830 35476 30882
rect 35196 30772 35252 30810
rect 35420 30772 35476 30830
rect 35756 30772 35812 30782
rect 35420 30770 35812 30772
rect 35420 30718 35758 30770
rect 35810 30718 35812 30770
rect 35420 30716 35812 30718
rect 35196 30706 35252 30716
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35084 30158 35086 30210
rect 35138 30158 35140 30210
rect 35084 30146 35140 30158
rect 35308 30100 35364 30110
rect 35196 29988 35252 29998
rect 34972 29374 34974 29426
rect 35026 29374 35028 29426
rect 34972 29362 35028 29374
rect 35084 29986 35252 29988
rect 35084 29934 35198 29986
rect 35250 29934 35252 29986
rect 35084 29932 35252 29934
rect 34748 28578 34804 28588
rect 34524 28532 34580 28542
rect 34524 28438 34580 28476
rect 34300 28420 34356 28430
rect 34300 28326 34356 28364
rect 34412 28418 34468 28430
rect 34412 28366 34414 28418
rect 34466 28366 34468 28418
rect 34076 28030 34078 28082
rect 34130 28030 34132 28082
rect 33852 27972 33908 27982
rect 33740 27970 33908 27972
rect 33740 27918 33854 27970
rect 33906 27918 33908 27970
rect 33740 27916 33908 27918
rect 33740 27858 33796 27916
rect 33852 27906 33908 27916
rect 33740 27806 33742 27858
rect 33794 27806 33796 27858
rect 33740 27794 33796 27806
rect 34076 27748 34132 28030
rect 34188 27972 34244 27982
rect 34188 27878 34244 27916
rect 34412 27972 34468 28366
rect 34748 28420 34804 28430
rect 35084 28420 35140 29932
rect 35196 29922 35252 29932
rect 35196 29764 35252 29774
rect 35308 29764 35364 30044
rect 35756 29988 35812 30716
rect 35756 29922 35812 29932
rect 35868 30772 35924 30782
rect 35252 29708 35364 29764
rect 35868 29764 35924 30716
rect 36092 30770 36148 30782
rect 36092 30718 36094 30770
rect 36146 30718 36148 30770
rect 36092 30098 36148 30718
rect 36204 30212 36260 30222
rect 36204 30118 36260 30156
rect 36092 30046 36094 30098
rect 36146 30046 36148 30098
rect 36092 30034 36148 30046
rect 36204 29988 36260 29998
rect 35980 29764 36036 29774
rect 35868 29708 35980 29764
rect 35196 29698 35252 29708
rect 35756 29652 35812 29662
rect 35308 29650 35812 29652
rect 35308 29598 35758 29650
rect 35810 29598 35812 29650
rect 35308 29596 35812 29598
rect 35308 29538 35364 29596
rect 35756 29586 35812 29596
rect 35308 29486 35310 29538
rect 35362 29486 35364 29538
rect 35308 29474 35364 29486
rect 35644 29428 35700 29438
rect 35868 29428 35924 29708
rect 35980 29698 36036 29708
rect 36204 29652 36260 29932
rect 36092 29596 36204 29652
rect 35980 29540 36036 29550
rect 36092 29540 36148 29596
rect 36204 29586 36260 29596
rect 35980 29538 36148 29540
rect 35980 29486 35982 29538
rect 36034 29486 36148 29538
rect 35980 29484 36148 29486
rect 35980 29474 36036 29484
rect 35644 29426 35924 29428
rect 35644 29374 35646 29426
rect 35698 29374 35924 29426
rect 35644 29372 35924 29374
rect 36204 29428 36260 29438
rect 36316 29428 36372 30940
rect 37324 30772 37380 30782
rect 37324 30770 37716 30772
rect 37324 30718 37326 30770
rect 37378 30718 37716 30770
rect 37324 30716 37716 30718
rect 37324 30706 37380 30716
rect 36988 30212 37044 30222
rect 36988 30118 37044 30156
rect 37660 30210 37716 30716
rect 37884 30436 37940 32396
rect 39004 32450 39060 33070
rect 39676 32900 39732 32910
rect 39676 32786 39732 32844
rect 39676 32734 39678 32786
rect 39730 32734 39732 32786
rect 39676 32722 39732 32734
rect 40236 32900 40292 32910
rect 39004 32398 39006 32450
rect 39058 32398 39060 32450
rect 38556 32338 38612 32350
rect 38556 32286 38558 32338
rect 38610 32286 38612 32338
rect 38108 31778 38164 31790
rect 38108 31726 38110 31778
rect 38162 31726 38164 31778
rect 38108 31556 38164 31726
rect 38556 31780 38612 32286
rect 38556 31686 38612 31724
rect 39004 31668 39060 32398
rect 39788 32002 39844 32014
rect 39788 31950 39790 32002
rect 39842 31950 39844 32002
rect 39228 31892 39284 31902
rect 39788 31892 39844 31950
rect 40236 31892 40292 32844
rect 41580 32676 41636 33516
rect 42476 33124 42532 34300
rect 42868 34354 43540 34356
rect 42868 34302 43262 34354
rect 43314 34302 43540 34354
rect 42868 34300 43540 34302
rect 43596 34914 43652 35644
rect 43932 35634 43988 35644
rect 44044 35364 44100 36092
rect 44156 35924 44212 36206
rect 44716 36148 44772 36876
rect 44828 36482 44884 37548
rect 44828 36430 44830 36482
rect 44882 36430 44884 36482
rect 44828 36418 44884 36430
rect 45052 37266 45108 37278
rect 45052 37214 45054 37266
rect 45106 37214 45108 37266
rect 45052 36484 45108 37214
rect 45612 37154 45668 37166
rect 45612 37102 45614 37154
rect 45666 37102 45668 37154
rect 45612 36820 45668 37102
rect 45612 36754 45668 36764
rect 45052 36418 45108 36428
rect 45724 36484 45780 36522
rect 45724 36418 45780 36428
rect 46284 36484 46340 37660
rect 46732 37268 46788 37278
rect 46396 37044 46452 37054
rect 46396 36950 46452 36988
rect 46284 36390 46340 36428
rect 46620 36484 46676 36494
rect 46732 36484 46788 37212
rect 47068 37154 47124 37886
rect 47404 37940 47460 37950
rect 47404 37846 47460 37884
rect 47180 37826 47236 37838
rect 47180 37774 47182 37826
rect 47234 37774 47236 37826
rect 47180 37268 47236 37774
rect 47180 37202 47236 37212
rect 47292 37380 47348 37390
rect 47068 37102 47070 37154
rect 47122 37102 47124 37154
rect 47068 37090 47124 37102
rect 47292 36708 47348 37324
rect 46620 36482 46788 36484
rect 46620 36430 46622 36482
rect 46674 36430 46788 36482
rect 46620 36428 46788 36430
rect 46844 36652 47348 36708
rect 46620 36418 46676 36428
rect 45276 36372 45332 36382
rect 45332 36316 45444 36372
rect 45276 36278 45332 36316
rect 44716 36092 45332 36148
rect 44604 35924 44660 35934
rect 44156 35922 44660 35924
rect 44156 35870 44606 35922
rect 44658 35870 44660 35922
rect 44156 35868 44660 35870
rect 44604 35858 44660 35868
rect 44044 35298 44100 35308
rect 44940 35810 44996 35822
rect 44940 35758 44942 35810
rect 44994 35758 44996 35810
rect 43596 34862 43598 34914
rect 43650 34862 43652 34914
rect 42588 34244 42644 34254
rect 42588 33346 42644 34188
rect 42812 33458 42868 34300
rect 43260 34290 43316 34300
rect 43036 34130 43092 34142
rect 43036 34078 43038 34130
rect 43090 34078 43092 34130
rect 43036 33796 43092 34078
rect 43148 34132 43204 34142
rect 43148 34038 43204 34076
rect 43596 34130 43652 34862
rect 44940 34916 44996 35758
rect 45276 35810 45332 36092
rect 45276 35758 45278 35810
rect 45330 35758 45332 35810
rect 45276 35746 45332 35758
rect 45388 35810 45444 36316
rect 45836 36260 45892 36270
rect 45836 36166 45892 36204
rect 46396 36258 46452 36270
rect 46396 36206 46398 36258
rect 46450 36206 46452 36258
rect 45388 35758 45390 35810
rect 45442 35758 45444 35810
rect 45388 35588 45444 35758
rect 45612 35700 45668 35710
rect 45612 35606 45668 35644
rect 44940 34850 44996 34860
rect 45276 35532 45444 35588
rect 45948 35588 46004 35598
rect 46396 35588 46452 36206
rect 45948 35586 46452 35588
rect 45948 35534 45950 35586
rect 46002 35534 46452 35586
rect 45948 35532 46452 35534
rect 45276 34914 45332 35532
rect 45836 35364 45892 35374
rect 45948 35364 46004 35532
rect 45892 35308 46004 35364
rect 45836 35298 45892 35308
rect 45276 34862 45278 34914
rect 45330 34862 45332 34914
rect 45276 34850 45332 34862
rect 45836 34916 45892 34926
rect 45052 34692 45108 34702
rect 43596 34078 43598 34130
rect 43650 34078 43652 34130
rect 43596 34066 43652 34078
rect 44940 34690 45108 34692
rect 44940 34638 45054 34690
rect 45106 34638 45108 34690
rect 44940 34636 45108 34638
rect 43932 33908 43988 33918
rect 43988 33852 44100 33908
rect 43932 33842 43988 33852
rect 43036 33730 43092 33740
rect 42812 33406 42814 33458
rect 42866 33406 42868 33458
rect 42812 33394 42868 33406
rect 42588 33294 42590 33346
rect 42642 33294 42644 33346
rect 42588 33282 42644 33294
rect 44044 33236 44100 33852
rect 44156 33572 44212 33582
rect 44380 33572 44436 33582
rect 44156 33570 44380 33572
rect 44156 33518 44158 33570
rect 44210 33518 44380 33570
rect 44156 33516 44380 33518
rect 44156 33506 44212 33516
rect 44380 33506 44436 33516
rect 44156 33236 44212 33246
rect 44044 33234 44212 33236
rect 44044 33182 44158 33234
rect 44210 33182 44212 33234
rect 44044 33180 44212 33182
rect 44156 33170 44212 33180
rect 44268 33236 44324 33246
rect 44940 33236 44996 34636
rect 45052 34626 45108 34636
rect 45836 34356 45892 34860
rect 45164 34244 45220 34254
rect 45500 34244 45556 34254
rect 45164 34242 45332 34244
rect 45164 34190 45166 34242
rect 45218 34190 45332 34242
rect 45164 34188 45332 34190
rect 45164 34178 45220 34188
rect 45052 34132 45108 34142
rect 45052 34038 45108 34076
rect 45164 33906 45220 33918
rect 45164 33854 45166 33906
rect 45218 33854 45220 33906
rect 45052 33236 45108 33246
rect 44940 33180 45052 33236
rect 44268 33142 44324 33180
rect 45052 33170 45108 33180
rect 42476 33068 42756 33124
rect 41468 32564 41524 32574
rect 41468 32470 41524 32508
rect 41580 32450 41636 32620
rect 42700 32674 42756 33068
rect 45164 32788 45220 33854
rect 45276 33572 45332 34188
rect 45500 34150 45556 34188
rect 45724 34242 45780 34254
rect 45724 34190 45726 34242
rect 45778 34190 45780 34242
rect 45276 33346 45332 33516
rect 45388 34132 45444 34142
rect 45388 33458 45444 34076
rect 45724 33908 45780 34190
rect 45836 34242 45892 34300
rect 45836 34190 45838 34242
rect 45890 34190 45892 34242
rect 45836 34178 45892 34190
rect 46732 33908 46788 33918
rect 45724 33842 45780 33852
rect 46620 33852 46732 33908
rect 45388 33406 45390 33458
rect 45442 33406 45444 33458
rect 45388 33394 45444 33406
rect 45836 33458 45892 33470
rect 45836 33406 45838 33458
rect 45890 33406 45892 33458
rect 45276 33294 45278 33346
rect 45330 33294 45332 33346
rect 45276 33282 45332 33294
rect 45164 32722 45220 32732
rect 45836 32788 45892 33406
rect 46284 32788 46340 32798
rect 45836 32786 46340 32788
rect 45836 32734 46286 32786
rect 46338 32734 46340 32786
rect 45836 32732 46340 32734
rect 42700 32622 42702 32674
rect 42754 32622 42756 32674
rect 42700 32610 42756 32622
rect 43260 32676 43316 32686
rect 43260 32582 43316 32620
rect 43596 32676 43652 32686
rect 42364 32564 42420 32574
rect 42924 32564 42980 32574
rect 42364 32562 42532 32564
rect 42364 32510 42366 32562
rect 42418 32510 42532 32562
rect 42364 32508 42532 32510
rect 42364 32498 42420 32508
rect 41580 32398 41582 32450
rect 41634 32398 41636 32450
rect 41580 32386 41636 32398
rect 42476 32004 42532 32508
rect 42924 32470 42980 32508
rect 43148 32564 43204 32574
rect 43148 32470 43204 32508
rect 42476 31948 43428 32004
rect 40348 31892 40404 31902
rect 39228 31798 39284 31836
rect 39564 31836 39844 31892
rect 39900 31890 40404 31892
rect 39900 31838 40350 31890
rect 40402 31838 40404 31890
rect 39900 31836 40404 31838
rect 39452 31780 39508 31790
rect 39564 31780 39620 31836
rect 39452 31778 39620 31780
rect 39452 31726 39454 31778
rect 39506 31726 39620 31778
rect 39452 31724 39620 31726
rect 39452 31714 39508 31724
rect 38108 31490 38164 31500
rect 38780 31612 39004 31668
rect 38780 31444 38836 31612
rect 39004 31602 39060 31612
rect 39676 31668 39732 31678
rect 39676 31574 39732 31612
rect 39788 31668 39844 31678
rect 39900 31668 39956 31836
rect 40348 31826 40404 31836
rect 41356 31892 41412 31902
rect 39788 31666 39956 31668
rect 39788 31614 39790 31666
rect 39842 31614 39956 31666
rect 39788 31612 39956 31614
rect 38444 31388 38836 31444
rect 38108 31220 38164 31230
rect 38108 31126 38164 31164
rect 38444 30994 38500 31388
rect 38444 30942 38446 30994
rect 38498 30942 38500 30994
rect 38444 30930 38500 30942
rect 38668 31220 38724 31230
rect 38668 30994 38724 31164
rect 39788 31220 39844 31612
rect 39900 31332 39956 31342
rect 39956 31276 40068 31332
rect 39900 31266 39956 31276
rect 39788 31126 39844 31164
rect 38668 30942 38670 30994
rect 38722 30942 38724 30994
rect 38668 30930 38724 30942
rect 39340 30882 39396 30894
rect 39340 30830 39342 30882
rect 39394 30830 39396 30882
rect 37884 30370 37940 30380
rect 38668 30548 38724 30558
rect 37660 30158 37662 30210
rect 37714 30158 37716 30210
rect 37100 30100 37156 30110
rect 36764 29988 36820 29998
rect 36764 29538 36820 29932
rect 37100 29764 37156 30044
rect 37324 30100 37380 30110
rect 37324 30006 37380 30044
rect 36764 29486 36766 29538
rect 36818 29486 36820 29538
rect 36764 29474 36820 29486
rect 36988 29708 37156 29764
rect 37212 29986 37268 29998
rect 37212 29934 37214 29986
rect 37266 29934 37268 29986
rect 36204 29426 36372 29428
rect 36204 29374 36206 29426
rect 36258 29374 36372 29426
rect 36204 29372 36372 29374
rect 35644 29362 35700 29372
rect 36204 29362 36260 29372
rect 35196 29314 35252 29326
rect 35196 29262 35198 29314
rect 35250 29262 35252 29314
rect 35196 29204 35252 29262
rect 36876 29316 36932 29326
rect 36876 29222 36932 29260
rect 36204 29204 36260 29214
rect 35196 29148 35700 29204
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 34748 28326 34804 28364
rect 34972 28364 35140 28420
rect 35308 28868 35364 28878
rect 35308 28642 35364 28812
rect 35308 28590 35310 28642
rect 35362 28590 35364 28642
rect 34412 27906 34468 27916
rect 34748 27858 34804 27870
rect 34748 27806 34750 27858
rect 34802 27806 34804 27858
rect 34076 27692 34580 27748
rect 32956 25454 32958 25506
rect 33010 25454 33012 25506
rect 32956 25284 33012 25454
rect 33516 25676 33684 25732
rect 33740 27188 33796 27198
rect 33516 25284 33572 25676
rect 33628 25508 33684 25518
rect 33740 25508 33796 27132
rect 34524 27186 34580 27692
rect 34524 27134 34526 27186
rect 34578 27134 34580 27186
rect 34524 26852 34580 27134
rect 34748 27188 34804 27806
rect 34748 27122 34804 27132
rect 34524 26786 34580 26796
rect 34860 26516 34916 26526
rect 34972 26516 35028 28364
rect 35308 27748 35364 28590
rect 35532 28644 35588 28654
rect 35532 28530 35588 28588
rect 35532 28478 35534 28530
rect 35586 28478 35588 28530
rect 35532 28466 35588 28478
rect 35532 27972 35588 27982
rect 35532 27878 35588 27916
rect 35308 27692 35588 27748
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 35084 26852 35140 26862
rect 35084 26758 35140 26796
rect 34860 26514 35028 26516
rect 34860 26462 34862 26514
rect 34914 26462 35028 26514
rect 34860 26460 35028 26462
rect 34860 26450 34916 26460
rect 34636 26292 34692 26302
rect 33628 25506 33796 25508
rect 33628 25454 33630 25506
rect 33682 25454 33796 25506
rect 33628 25452 33796 25454
rect 33628 25442 33684 25452
rect 33516 25228 33684 25284
rect 32956 25218 33012 25228
rect 33404 25060 33460 25070
rect 33180 24948 33236 24958
rect 32844 24946 33236 24948
rect 32844 24894 33182 24946
rect 33234 24894 33236 24946
rect 32844 24892 33236 24894
rect 32732 24882 32788 24892
rect 33180 24882 33236 24892
rect 32396 24670 32398 24722
rect 32450 24670 32452 24722
rect 32396 24500 32452 24670
rect 33068 24724 33124 24734
rect 33292 24724 33348 24734
rect 33404 24724 33460 25004
rect 33068 24722 33236 24724
rect 33068 24670 33070 24722
rect 33122 24670 33236 24722
rect 33068 24668 33236 24670
rect 33068 24658 33124 24668
rect 32396 24444 33124 24500
rect 33068 23938 33124 24444
rect 33068 23886 33070 23938
rect 33122 23886 33124 23938
rect 33068 23874 33124 23886
rect 32620 23826 32676 23838
rect 32620 23774 32622 23826
rect 32674 23774 32676 23826
rect 32620 23492 32676 23774
rect 32956 23828 33012 23838
rect 32956 23734 33012 23772
rect 32620 23426 32676 23436
rect 32228 23212 32340 23268
rect 32396 23268 32452 23278
rect 32172 23202 32228 23212
rect 32396 23174 32452 23212
rect 30828 22306 30884 22316
rect 31948 22764 32116 22820
rect 30604 21746 30660 21756
rect 30044 20974 30046 21026
rect 30098 20974 30100 21026
rect 30044 20962 30100 20974
rect 30156 21700 30212 21710
rect 29708 20132 29988 20188
rect 29708 20130 29764 20132
rect 29708 20078 29710 20130
rect 29762 20078 29764 20130
rect 29708 20066 29764 20078
rect 29932 20020 29988 20030
rect 29820 20018 29988 20020
rect 29820 19966 29934 20018
rect 29986 19966 29988 20018
rect 29820 19964 29988 19966
rect 29820 19348 29876 19964
rect 29932 19954 29988 19964
rect 29596 19292 29876 19348
rect 28812 18900 28868 18956
rect 28364 18844 28868 18900
rect 28924 18956 29316 19012
rect 29484 19122 29540 19134
rect 29484 19070 29486 19122
rect 29538 19070 29540 19122
rect 28252 18676 28308 18686
rect 27916 18564 27972 18574
rect 27916 18470 27972 18508
rect 28028 18562 28084 18574
rect 28028 18510 28030 18562
rect 28082 18510 28084 18562
rect 28028 18452 28084 18510
rect 28028 18386 28084 18396
rect 28252 18450 28308 18620
rect 28252 18398 28254 18450
rect 28306 18398 28308 18450
rect 28252 18386 28308 18398
rect 27468 18286 27470 18338
rect 27522 18286 27524 18338
rect 27468 18274 27524 18286
rect 27916 17780 27972 17790
rect 28364 17780 28420 18844
rect 27916 17778 28420 17780
rect 27916 17726 27918 17778
rect 27970 17726 28420 17778
rect 27916 17724 28420 17726
rect 28588 18452 28644 18462
rect 27916 17714 27972 17724
rect 28476 16884 28532 16894
rect 28588 16884 28644 18396
rect 28476 16882 28644 16884
rect 28476 16830 28478 16882
rect 28530 16830 28644 16882
rect 28476 16828 28644 16830
rect 28476 16818 28532 16828
rect 28588 15314 28644 15326
rect 28588 15262 28590 15314
rect 28642 15262 28644 15314
rect 27356 15138 27412 15148
rect 28140 15202 28196 15214
rect 28140 15150 28142 15202
rect 28194 15150 28196 15202
rect 22204 13906 22260 13916
rect 22428 14140 22596 14196
rect 22204 13746 22260 13758
rect 22204 13694 22206 13746
rect 22258 13694 22260 13746
rect 22204 12292 22260 13694
rect 22316 13746 22372 13758
rect 22316 13694 22318 13746
rect 22370 13694 22372 13746
rect 22316 13636 22372 13694
rect 22316 13570 22372 13580
rect 22428 13748 22484 14140
rect 22540 13972 22596 13982
rect 22540 13970 23156 13972
rect 22540 13918 22542 13970
rect 22594 13918 23156 13970
rect 22540 13916 23156 13918
rect 22540 13906 22596 13916
rect 23100 13860 23156 13916
rect 23100 13766 23156 13804
rect 23436 13860 23492 13870
rect 22652 13748 22708 13758
rect 22428 13746 22708 13748
rect 22428 13694 22654 13746
rect 22706 13694 22708 13746
rect 22428 13692 22708 13694
rect 22316 13076 22372 13086
rect 22428 13076 22484 13692
rect 22652 13682 22708 13692
rect 23324 13522 23380 13534
rect 23324 13470 23326 13522
rect 23378 13470 23380 13522
rect 22316 13074 22484 13076
rect 22316 13022 22318 13074
rect 22370 13022 22484 13074
rect 22316 13020 22484 13022
rect 23100 13076 23156 13086
rect 22316 13010 22372 13020
rect 23100 12982 23156 13020
rect 23212 12964 23268 12974
rect 23212 12870 23268 12908
rect 22316 12292 22372 12302
rect 23324 12292 23380 13470
rect 23436 12402 23492 13804
rect 23436 12350 23438 12402
rect 23490 12350 23492 12402
rect 23436 12338 23492 12350
rect 23548 13748 23604 13758
rect 22204 12290 22372 12292
rect 22204 12238 22318 12290
rect 22370 12238 22372 12290
rect 22204 12236 22372 12238
rect 22316 12226 22372 12236
rect 23212 12236 23380 12292
rect 23212 12178 23268 12236
rect 23548 12180 23604 13692
rect 23660 13522 23716 13534
rect 23660 13470 23662 13522
rect 23714 13470 23716 13522
rect 23660 12962 23716 13470
rect 23660 12910 23662 12962
rect 23714 12910 23716 12962
rect 23660 12898 23716 12910
rect 23772 12964 23828 12974
rect 23212 12126 23214 12178
rect 23266 12126 23268 12178
rect 23212 11788 23268 12126
rect 23436 12124 23604 12180
rect 23772 12178 23828 12908
rect 23772 12126 23774 12178
rect 23826 12126 23828 12178
rect 23324 12068 23380 12078
rect 23436 12068 23492 12124
rect 23772 12114 23828 12126
rect 23324 12066 23492 12068
rect 23324 12014 23326 12066
rect 23378 12014 23492 12066
rect 23324 12012 23492 12014
rect 23324 12002 23380 12012
rect 23212 11732 23380 11788
rect 22876 11508 22932 11518
rect 22876 11394 22932 11452
rect 22876 11342 22878 11394
rect 22930 11342 22932 11394
rect 22876 11330 22932 11342
rect 23212 11172 23268 11182
rect 22092 11116 22708 11172
rect 20412 10782 20414 10834
rect 20466 10782 20468 10834
rect 20412 10770 20468 10782
rect 19180 10518 19236 10556
rect 20188 10556 20356 10612
rect 22316 10610 22372 10622
rect 22316 10558 22318 10610
rect 22370 10558 22372 10610
rect 18284 9762 18340 9772
rect 19068 9826 19124 9838
rect 19740 9828 19796 9838
rect 19068 9774 19070 9826
rect 19122 9774 19124 9826
rect 17724 9662 17726 9714
rect 17778 9662 17780 9714
rect 17724 9650 17780 9662
rect 18732 9714 18788 9726
rect 18732 9662 18734 9714
rect 18786 9662 18788 9714
rect 17948 9604 18004 9614
rect 17948 9510 18004 9548
rect 18732 9604 18788 9662
rect 18732 9156 18788 9548
rect 18844 9156 18900 9166
rect 18732 9100 18844 9156
rect 18844 9090 18900 9100
rect 15708 8930 16212 8932
rect 15708 8878 15710 8930
rect 15762 8878 16212 8930
rect 15708 8876 16212 8878
rect 16268 9042 16324 9054
rect 16268 8990 16270 9042
rect 16322 8990 16324 9042
rect 15708 7812 15764 8876
rect 15820 8148 15876 8158
rect 15820 7924 15876 8092
rect 16268 7924 16324 8990
rect 15820 7868 16212 7924
rect 15708 7756 15988 7812
rect 15484 7634 15540 7644
rect 15932 7474 15988 7756
rect 15932 7422 15934 7474
rect 15986 7422 15988 7474
rect 15932 7410 15988 7422
rect 16156 7474 16212 7868
rect 16268 7858 16324 7868
rect 16492 9044 16548 9054
rect 16492 7698 16548 8988
rect 17948 9044 18004 9054
rect 19068 9044 19124 9774
rect 19628 9826 19796 9828
rect 19628 9774 19742 9826
rect 19794 9774 19796 9826
rect 19628 9772 19796 9774
rect 19628 9268 19684 9772
rect 19740 9762 19796 9772
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 20188 9268 20244 10556
rect 20412 9828 20468 9838
rect 21420 9828 21476 9838
rect 20412 9826 21476 9828
rect 20412 9774 20414 9826
rect 20466 9774 21422 9826
rect 21474 9774 21476 9826
rect 20412 9772 21476 9774
rect 20412 9762 20468 9772
rect 19404 9212 19908 9268
rect 19292 9044 19348 9054
rect 19068 9042 19348 9044
rect 19068 8990 19294 9042
rect 19346 8990 19348 9042
rect 19068 8988 19348 8990
rect 17948 8950 18004 8988
rect 18172 8372 18228 8382
rect 18172 8278 18228 8316
rect 16828 8258 16884 8270
rect 16828 8206 16830 8258
rect 16882 8206 16884 8258
rect 16828 7924 16884 8206
rect 16828 7858 16884 7868
rect 18844 8260 18900 8270
rect 19292 8260 19348 8988
rect 18844 8258 19348 8260
rect 18844 8206 18846 8258
rect 18898 8206 19348 8258
rect 18844 8204 19348 8206
rect 19404 8372 19460 9212
rect 19852 9154 19908 9212
rect 20076 9212 20244 9268
rect 19852 9102 19854 9154
rect 19906 9102 19908 9154
rect 19852 9090 19908 9102
rect 19964 9156 20020 9166
rect 19404 8258 19460 8316
rect 19404 8206 19406 8258
rect 19458 8206 19460 8258
rect 16492 7646 16494 7698
rect 16546 7646 16548 7698
rect 16492 7634 16548 7646
rect 16156 7422 16158 7474
rect 16210 7422 16212 7474
rect 16156 7410 16212 7422
rect 15708 7364 15764 7374
rect 15708 7270 15764 7308
rect 18844 7252 18900 8204
rect 19404 8194 19460 8206
rect 19516 8148 19572 8158
rect 19852 8148 19908 8158
rect 19516 8146 19908 8148
rect 19516 8094 19518 8146
rect 19570 8094 19854 8146
rect 19906 8094 19908 8146
rect 19516 8092 19908 8094
rect 19516 8082 19572 8092
rect 19852 8082 19908 8092
rect 19964 8146 20020 9100
rect 20076 8930 20132 9212
rect 20860 9154 20916 9772
rect 21420 9762 21476 9772
rect 21532 9826 21588 9838
rect 21532 9774 21534 9826
rect 21586 9774 21588 9826
rect 21532 9716 21588 9774
rect 21532 9650 21588 9660
rect 22092 9716 22148 9726
rect 20972 9604 21028 9614
rect 20972 9266 21028 9548
rect 22092 9380 22148 9660
rect 20972 9214 20974 9266
rect 21026 9214 21028 9266
rect 20972 9202 21028 9214
rect 21980 9324 22148 9380
rect 20860 9102 20862 9154
rect 20914 9102 20916 9154
rect 20860 9090 20916 9102
rect 21196 9156 21252 9166
rect 21196 9062 21252 9100
rect 21980 9156 22036 9324
rect 22316 9266 22372 10558
rect 22652 9604 22708 11116
rect 22764 11170 23268 11172
rect 22764 11118 23214 11170
rect 23266 11118 23268 11170
rect 22764 11116 23268 11118
rect 22764 10498 22820 11116
rect 23212 11106 23268 11116
rect 22764 10446 22766 10498
rect 22818 10446 22820 10498
rect 22764 9828 22820 10446
rect 23324 9938 23380 11732
rect 23996 11396 24052 15092
rect 24220 14532 24276 14542
rect 24220 14438 24276 14476
rect 25004 14532 25060 14542
rect 25452 14532 25508 14542
rect 25004 14530 25508 14532
rect 25004 14478 25006 14530
rect 25058 14478 25454 14530
rect 25506 14478 25508 14530
rect 25004 14476 25508 14478
rect 25004 14466 25060 14476
rect 25452 14466 25508 14476
rect 24668 14418 24724 14430
rect 24668 14366 24670 14418
rect 24722 14366 24724 14418
rect 24668 13748 24724 14366
rect 24780 14308 24836 14318
rect 24780 14214 24836 14252
rect 25340 14308 25396 14318
rect 24668 13682 24724 13692
rect 25116 13748 25172 13758
rect 25340 13748 25396 14252
rect 25452 13972 25508 13982
rect 25564 13972 25620 15092
rect 26236 14754 26292 15092
rect 26236 14702 26238 14754
rect 26290 14702 26292 14754
rect 26236 14690 26292 14702
rect 25452 13970 25620 13972
rect 25452 13918 25454 13970
rect 25506 13918 25620 13970
rect 25452 13916 25620 13918
rect 25676 14642 25732 14654
rect 25676 14590 25678 14642
rect 25730 14590 25732 14642
rect 25676 14532 25732 14590
rect 27916 14642 27972 14654
rect 27916 14590 27918 14642
rect 27970 14590 27972 14642
rect 26012 14532 26068 14542
rect 25452 13906 25508 13916
rect 25452 13748 25508 13758
rect 25340 13746 25508 13748
rect 25340 13694 25454 13746
rect 25506 13694 25508 13746
rect 25340 13692 25508 13694
rect 25116 13654 25172 13692
rect 25452 13682 25508 13692
rect 25676 13746 25732 14476
rect 25676 13694 25678 13746
rect 25730 13694 25732 13746
rect 25676 13682 25732 13694
rect 25900 14476 26012 14532
rect 25900 13186 25956 14476
rect 26012 14466 26068 14476
rect 27020 14530 27076 14542
rect 27020 14478 27022 14530
rect 27074 14478 27076 14530
rect 25900 13134 25902 13186
rect 25954 13134 25956 13186
rect 25900 13122 25956 13134
rect 26572 13076 26628 13086
rect 26012 13074 26740 13076
rect 26012 13022 26574 13074
rect 26626 13022 26740 13074
rect 26012 13020 26740 13022
rect 25788 12964 25844 12974
rect 26012 12964 26068 13020
rect 26572 13010 26628 13020
rect 25788 12962 26068 12964
rect 25788 12910 25790 12962
rect 25842 12910 26068 12962
rect 25788 12908 26068 12910
rect 25788 12898 25844 12908
rect 25900 12740 25956 12750
rect 25900 12646 25956 12684
rect 26684 11956 26740 13020
rect 26908 12852 26964 12862
rect 26908 12758 26964 12796
rect 27020 12628 27076 14478
rect 27580 14532 27636 14542
rect 27580 14438 27636 14476
rect 27356 13746 27412 13758
rect 27356 13694 27358 13746
rect 27410 13694 27412 13746
rect 26908 12572 27076 12628
rect 27132 12740 27188 12750
rect 26908 12402 26964 12572
rect 26908 12350 26910 12402
rect 26962 12350 26964 12402
rect 26908 12338 26964 12350
rect 26908 12180 26964 12190
rect 26796 11956 26852 11966
rect 26684 11954 26852 11956
rect 26684 11902 26798 11954
rect 26850 11902 26852 11954
rect 26684 11900 26852 11902
rect 23548 11340 24052 11396
rect 25452 11396 25508 11406
rect 25452 11394 25732 11396
rect 25452 11342 25454 11394
rect 25506 11342 25732 11394
rect 25452 11340 25732 11342
rect 23548 10834 23604 11340
rect 25452 11330 25508 11340
rect 25116 11284 25172 11294
rect 25116 11190 25172 11228
rect 23548 10782 23550 10834
rect 23602 10782 23604 10834
rect 23548 10770 23604 10782
rect 25676 10612 25732 11340
rect 26572 11282 26628 11294
rect 26572 11230 26574 11282
rect 26626 11230 26628 11282
rect 26572 10836 26628 11230
rect 26572 10770 26628 10780
rect 23324 9886 23326 9938
rect 23378 9886 23380 9938
rect 23324 9874 23380 9886
rect 25564 10610 25732 10612
rect 25564 10558 25678 10610
rect 25730 10558 25732 10610
rect 25564 10556 25732 10558
rect 25564 9940 25620 10556
rect 25676 10546 25732 10556
rect 25788 10612 25844 10622
rect 25564 9846 25620 9884
rect 22764 9762 22820 9772
rect 23772 9828 23828 9838
rect 23772 9734 23828 9772
rect 25788 9826 25844 10556
rect 26460 10612 26516 10650
rect 26460 10546 26516 10556
rect 26348 10500 26404 10510
rect 25788 9774 25790 9826
rect 25842 9774 25844 9826
rect 23212 9716 23268 9726
rect 23212 9622 23268 9660
rect 23548 9714 23604 9726
rect 23548 9662 23550 9714
rect 23602 9662 23604 9714
rect 22764 9604 22820 9614
rect 22652 9602 22820 9604
rect 22652 9550 22766 9602
rect 22818 9550 22820 9602
rect 22652 9548 22820 9550
rect 22764 9538 22820 9548
rect 23548 9492 23604 9662
rect 22316 9214 22318 9266
rect 22370 9214 22372 9266
rect 22316 9202 22372 9214
rect 23436 9436 23604 9492
rect 21980 9062 22036 9100
rect 22092 9154 22148 9166
rect 22092 9102 22094 9154
rect 22146 9102 22148 9154
rect 20076 8878 20078 8930
rect 20130 8878 20132 8930
rect 20076 8866 20132 8878
rect 22092 9044 22148 9102
rect 20188 8484 20244 8494
rect 20188 8258 20244 8428
rect 22092 8484 22148 8988
rect 23436 9044 23492 9436
rect 23436 8978 23492 8988
rect 25564 8930 25620 8942
rect 25564 8878 25566 8930
rect 25618 8878 25620 8930
rect 22092 8418 22148 8428
rect 24668 8484 24724 8494
rect 24668 8390 24724 8428
rect 25004 8372 25060 8382
rect 25004 8278 25060 8316
rect 20188 8206 20190 8258
rect 20242 8206 20244 8258
rect 20188 8194 20244 8206
rect 24668 8258 24724 8270
rect 24668 8206 24670 8258
rect 24722 8206 24724 8258
rect 19964 8094 19966 8146
rect 20018 8094 20020 8146
rect 19964 8082 20020 8094
rect 24332 8146 24388 8158
rect 24332 8094 24334 8146
rect 24386 8094 24388 8146
rect 22876 8036 22932 8046
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 22876 7474 22932 7980
rect 22876 7422 22878 7474
rect 22930 7422 22932 7474
rect 22876 7410 22932 7422
rect 23212 7476 23268 7486
rect 23212 7382 23268 7420
rect 24220 7474 24276 7486
rect 24220 7422 24222 7474
rect 24274 7422 24276 7474
rect 18844 7186 18900 7196
rect 15148 6860 15428 6916
rect 15148 6804 15204 6860
rect 15036 6748 15204 6804
rect 15036 6690 15092 6748
rect 15036 6638 15038 6690
rect 15090 6638 15092 6690
rect 15036 6626 15092 6638
rect 24220 6692 24276 7422
rect 24332 6914 24388 8094
rect 24668 8036 24724 8206
rect 24668 7970 24724 7980
rect 25228 8260 25284 8270
rect 25564 8260 25620 8878
rect 25788 8484 25844 9774
rect 26012 9828 26068 9838
rect 26348 9828 26404 10444
rect 26460 10388 26516 10398
rect 26460 10050 26516 10332
rect 26460 9998 26462 10050
rect 26514 9998 26516 10050
rect 26460 9986 26516 9998
rect 26012 9826 26404 9828
rect 26012 9774 26014 9826
rect 26066 9774 26404 9826
rect 26012 9772 26404 9774
rect 25788 8418 25844 8428
rect 25900 9042 25956 9054
rect 25900 8990 25902 9042
rect 25954 8990 25956 9042
rect 25900 8372 25956 8990
rect 25900 8306 25956 8316
rect 25228 8258 25620 8260
rect 25228 8206 25230 8258
rect 25282 8206 25620 8258
rect 25228 8204 25620 8206
rect 24668 7588 24724 7598
rect 25228 7588 25284 8204
rect 25564 8036 25620 8046
rect 26012 8036 26068 9772
rect 26348 9156 26404 9166
rect 26684 9156 26740 11900
rect 26796 11890 26852 11900
rect 26908 11788 26964 12124
rect 27132 12178 27188 12684
rect 27132 12126 27134 12178
rect 27186 12126 27188 12178
rect 27132 11956 27188 12126
rect 27356 12180 27412 13694
rect 27916 13634 27972 14590
rect 27916 13582 27918 13634
rect 27970 13582 27972 13634
rect 27916 13300 27972 13582
rect 28028 14418 28084 14430
rect 28028 14366 28030 14418
rect 28082 14366 28084 14418
rect 28028 13412 28084 14366
rect 28140 14420 28196 15150
rect 28140 13858 28196 14364
rect 28140 13806 28142 13858
rect 28194 13806 28196 13858
rect 28140 13794 28196 13806
rect 28476 14532 28532 14542
rect 28028 13356 28420 13412
rect 27916 13244 28196 13300
rect 27356 12114 27412 12124
rect 27468 12178 27524 12190
rect 27468 12126 27470 12178
rect 27522 12126 27524 12178
rect 27132 11890 27188 11900
rect 26796 11732 26964 11788
rect 26796 11506 26852 11732
rect 27468 11618 27524 12126
rect 28140 12066 28196 13244
rect 28364 12850 28420 13356
rect 28364 12798 28366 12850
rect 28418 12798 28420 12850
rect 28364 12404 28420 12798
rect 28476 12738 28532 14476
rect 28588 14308 28644 15262
rect 28812 14308 28868 14318
rect 28588 14306 28812 14308
rect 28588 14254 28590 14306
rect 28642 14254 28812 14306
rect 28588 14252 28812 14254
rect 28588 14242 28644 14252
rect 28812 14242 28868 14252
rect 28476 12686 28478 12738
rect 28530 12686 28532 12738
rect 28476 12674 28532 12686
rect 28364 12338 28420 12348
rect 28476 12290 28532 12302
rect 28476 12238 28478 12290
rect 28530 12238 28532 12290
rect 28252 12180 28308 12190
rect 28252 12086 28308 12124
rect 28476 12180 28532 12238
rect 28476 12114 28532 12124
rect 28140 12014 28142 12066
rect 28194 12014 28196 12066
rect 28140 12002 28196 12014
rect 27468 11566 27470 11618
rect 27522 11566 27524 11618
rect 27468 11554 27524 11566
rect 28252 11956 28308 11966
rect 26796 11454 26798 11506
rect 26850 11454 26852 11506
rect 26796 11442 26852 11454
rect 27132 11396 27188 11406
rect 27020 11394 27188 11396
rect 27020 11342 27134 11394
rect 27186 11342 27188 11394
rect 27020 11340 27188 11342
rect 27020 10388 27076 11340
rect 27132 11330 27188 11340
rect 27804 11396 27860 11406
rect 27804 11302 27860 11340
rect 27356 11282 27412 11294
rect 27356 11230 27358 11282
rect 27410 11230 27412 11282
rect 27356 11172 27412 11230
rect 27132 10724 27188 10734
rect 27356 10724 27412 11116
rect 28028 10836 28084 10846
rect 28028 10742 28084 10780
rect 28252 10834 28308 11900
rect 28588 11732 28644 11742
rect 28588 11396 28644 11676
rect 28588 11394 28756 11396
rect 28588 11342 28590 11394
rect 28642 11342 28756 11394
rect 28588 11340 28756 11342
rect 28588 11330 28644 11340
rect 28252 10782 28254 10834
rect 28306 10782 28308 10834
rect 28252 10770 28308 10782
rect 28476 10836 28532 10846
rect 28476 10742 28532 10780
rect 27132 10722 27412 10724
rect 27132 10670 27134 10722
rect 27186 10670 27412 10722
rect 27132 10668 27412 10670
rect 27132 10658 27188 10668
rect 27468 10612 27524 10622
rect 27468 10518 27524 10556
rect 28588 10610 28644 10622
rect 28588 10558 28590 10610
rect 28642 10558 28644 10610
rect 27692 10500 27748 10510
rect 27692 10406 27748 10444
rect 28588 10388 28644 10558
rect 28700 10500 28756 11340
rect 28924 10724 28980 18956
rect 29484 18788 29540 19070
rect 29484 18722 29540 18732
rect 29596 19122 29652 19292
rect 30156 19236 30212 21644
rect 31612 21474 31668 21486
rect 31612 21422 31614 21474
rect 31666 21422 31668 21474
rect 30380 20804 30436 20814
rect 30380 20710 30436 20748
rect 30604 20692 30660 20702
rect 30828 20692 30884 20702
rect 30604 20690 30884 20692
rect 30604 20638 30606 20690
rect 30658 20638 30830 20690
rect 30882 20638 30884 20690
rect 30604 20636 30884 20638
rect 30604 20626 30660 20636
rect 30828 20626 30884 20636
rect 31164 20692 31220 20702
rect 31164 20598 31220 20636
rect 31052 20578 31108 20590
rect 31052 20526 31054 20578
rect 31106 20526 31108 20578
rect 31052 20468 31108 20526
rect 31612 20578 31668 21422
rect 31612 20526 31614 20578
rect 31666 20526 31668 20578
rect 31612 20468 31668 20526
rect 31052 20412 31668 20468
rect 31612 20356 31668 20412
rect 31612 20300 31892 20356
rect 31052 20244 31108 20254
rect 30380 20020 30436 20030
rect 30380 19926 30436 19964
rect 30604 20020 30660 20030
rect 30604 20018 30772 20020
rect 30604 19966 30606 20018
rect 30658 19966 30772 20018
rect 30604 19964 30772 19966
rect 30604 19954 30660 19964
rect 30492 19908 30548 19918
rect 30492 19814 30548 19852
rect 30492 19236 30548 19246
rect 30156 19234 30660 19236
rect 30156 19182 30494 19234
rect 30546 19182 30660 19234
rect 30156 19180 30660 19182
rect 30492 19170 30548 19180
rect 29596 19070 29598 19122
rect 29650 19070 29652 19122
rect 29596 18676 29652 19070
rect 29708 19124 29764 19134
rect 29708 19030 29764 19068
rect 29932 19012 29988 19022
rect 29932 18918 29988 18956
rect 29596 18610 29652 18620
rect 30268 18676 30324 18686
rect 30268 18450 30324 18620
rect 30268 18398 30270 18450
rect 30322 18398 30324 18450
rect 30268 18386 30324 18398
rect 30604 18674 30660 19180
rect 30716 19012 30772 19964
rect 30716 18946 30772 18956
rect 30604 18622 30606 18674
rect 30658 18622 30660 18674
rect 30604 18452 30660 18622
rect 31052 18676 31108 20188
rect 31724 20132 31780 20142
rect 31276 20130 31780 20132
rect 31276 20078 31726 20130
rect 31778 20078 31780 20130
rect 31276 20076 31780 20078
rect 31276 19346 31332 20076
rect 31724 20066 31780 20076
rect 31276 19294 31278 19346
rect 31330 19294 31332 19346
rect 31276 19282 31332 19294
rect 31052 18610 31108 18620
rect 29708 17892 29764 17902
rect 29596 17444 29652 17454
rect 29148 17442 29652 17444
rect 29148 17390 29598 17442
rect 29650 17390 29652 17442
rect 29148 17388 29652 17390
rect 29148 16994 29204 17388
rect 29596 17378 29652 17388
rect 29708 17108 29764 17836
rect 29932 17556 29988 17566
rect 30380 17556 30436 17566
rect 29932 17554 30436 17556
rect 29932 17502 29934 17554
rect 29986 17502 30382 17554
rect 30434 17502 30436 17554
rect 29932 17500 30436 17502
rect 29932 17490 29988 17500
rect 30380 17490 30436 17500
rect 29148 16942 29150 16994
rect 29202 16942 29204 16994
rect 29148 16930 29204 16942
rect 29260 17052 29764 17108
rect 29148 15874 29204 15886
rect 29148 15822 29150 15874
rect 29202 15822 29204 15874
rect 29148 15652 29204 15822
rect 29260 15874 29316 17052
rect 30604 16772 30660 18396
rect 30716 17668 30772 17678
rect 30716 17666 30884 17668
rect 30716 17614 30718 17666
rect 30770 17614 30884 17666
rect 30716 17612 30884 17614
rect 30716 17602 30772 17612
rect 30828 16884 30884 17612
rect 31388 17666 31444 17678
rect 31388 17614 31390 17666
rect 31442 17614 31444 17666
rect 31388 17556 31444 17614
rect 31388 17490 31444 17500
rect 31500 17554 31556 17566
rect 31500 17502 31502 17554
rect 31554 17502 31556 17554
rect 30828 16828 31332 16884
rect 30604 16716 31220 16772
rect 30156 16212 30212 16222
rect 29820 16210 30212 16212
rect 29820 16158 30158 16210
rect 30210 16158 30212 16210
rect 29820 16156 30212 16158
rect 29820 16098 29876 16156
rect 30156 16146 30212 16156
rect 31164 16210 31220 16716
rect 31164 16158 31166 16210
rect 31218 16158 31220 16210
rect 31164 16146 31220 16158
rect 31276 16770 31332 16828
rect 31276 16718 31278 16770
rect 31330 16718 31332 16770
rect 29820 16046 29822 16098
rect 29874 16046 29876 16098
rect 29820 16034 29876 16046
rect 30044 15986 30100 15998
rect 30044 15934 30046 15986
rect 30098 15934 30100 15986
rect 29260 15822 29262 15874
rect 29314 15822 29316 15874
rect 29260 15810 29316 15822
rect 29372 15876 29428 15886
rect 29372 15782 29428 15820
rect 30044 15764 30100 15934
rect 29484 15708 30100 15764
rect 30380 15986 30436 15998
rect 30380 15934 30382 15986
rect 30434 15934 30436 15986
rect 30380 15876 30436 15934
rect 29484 15652 29540 15708
rect 29036 15596 29540 15652
rect 29036 15426 29092 15596
rect 29036 15374 29038 15426
rect 29090 15374 29092 15426
rect 29036 15362 29092 15374
rect 30044 15428 30100 15438
rect 29484 15314 29540 15326
rect 29484 15262 29486 15314
rect 29538 15262 29540 15314
rect 29484 14754 29540 15262
rect 30044 15202 30100 15372
rect 30044 15150 30046 15202
rect 30098 15150 30100 15202
rect 30044 15138 30100 15150
rect 30156 15426 30212 15438
rect 30156 15374 30158 15426
rect 30210 15374 30212 15426
rect 29484 14702 29486 14754
rect 29538 14702 29540 14754
rect 29484 14690 29540 14702
rect 29484 14532 29540 14542
rect 29484 14530 29764 14532
rect 29484 14478 29486 14530
rect 29538 14478 29764 14530
rect 29484 14476 29764 14478
rect 29148 14420 29204 14430
rect 29148 14326 29204 14364
rect 29484 14308 29540 14476
rect 29484 14242 29540 14252
rect 29708 13636 29764 14476
rect 30156 14530 30212 15374
rect 30380 15428 30436 15820
rect 30604 15986 30660 15998
rect 30604 15934 30606 15986
rect 30658 15934 30660 15986
rect 30604 15652 30660 15934
rect 30604 15586 30660 15596
rect 31276 15540 31332 16718
rect 31388 16324 31444 16334
rect 31388 16098 31444 16268
rect 31500 16212 31556 17502
rect 31836 16884 31892 20300
rect 31948 20132 32004 22764
rect 33180 22484 33236 24668
rect 33292 24722 33460 24724
rect 33292 24670 33294 24722
rect 33346 24670 33460 24722
rect 33292 24668 33460 24670
rect 33516 24948 33572 24958
rect 33292 24164 33348 24668
rect 33516 24276 33572 24892
rect 33516 24210 33572 24220
rect 33292 24098 33348 24108
rect 33180 22418 33236 22428
rect 33404 24050 33460 24062
rect 33404 23998 33406 24050
rect 33458 23998 33460 24050
rect 32060 21700 32116 21710
rect 32060 21606 32116 21644
rect 32508 21700 32564 21710
rect 32508 21606 32564 21644
rect 33068 21700 33124 21710
rect 33068 21586 33124 21644
rect 33068 21534 33070 21586
rect 33122 21534 33124 21586
rect 33068 21522 33124 21534
rect 32060 21252 32116 21262
rect 32060 20914 32116 21196
rect 33404 21028 33460 23998
rect 33516 23940 33572 23950
rect 33516 23268 33572 23884
rect 33516 22482 33572 23212
rect 33516 22430 33518 22482
rect 33570 22430 33572 22482
rect 33516 22418 33572 22430
rect 33516 21028 33572 21038
rect 33404 21026 33572 21028
rect 33404 20974 33518 21026
rect 33570 20974 33572 21026
rect 33404 20972 33572 20974
rect 33516 20962 33572 20972
rect 32060 20862 32062 20914
rect 32114 20862 32116 20914
rect 32060 20244 32116 20862
rect 33292 20804 33348 20814
rect 33292 20710 33348 20748
rect 32060 20178 32116 20188
rect 31948 20066 32004 20076
rect 32060 20020 32116 20030
rect 33180 20020 33236 20030
rect 32060 20018 33236 20020
rect 32060 19966 32062 20018
rect 32114 19966 33182 20018
rect 33234 19966 33236 20018
rect 32060 19964 33236 19966
rect 32060 19954 32116 19964
rect 33180 19954 33236 19964
rect 33516 19796 33572 19806
rect 33404 19794 33572 19796
rect 33404 19742 33518 19794
rect 33570 19742 33572 19794
rect 33404 19740 33572 19742
rect 33404 19346 33460 19740
rect 33516 19730 33572 19740
rect 33404 19294 33406 19346
rect 33458 19294 33460 19346
rect 33404 18564 33460 19294
rect 33628 18788 33684 25228
rect 33740 25060 33796 25452
rect 33740 24994 33796 25004
rect 33852 26290 34692 26292
rect 33852 26238 34638 26290
rect 34690 26238 34692 26290
rect 33852 26236 34692 26238
rect 33740 24052 33796 24062
rect 33740 23938 33796 23996
rect 33852 24050 33908 26236
rect 34636 26226 34692 26236
rect 35196 26292 35252 26302
rect 35196 26198 35252 26236
rect 34748 26178 34804 26190
rect 34748 26126 34750 26178
rect 34802 26126 34804 26178
rect 34748 25844 34804 26126
rect 34300 25788 34804 25844
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 34300 25618 34356 25788
rect 34300 25566 34302 25618
rect 34354 25566 34356 25618
rect 34300 25554 34356 25566
rect 34076 25172 34132 25182
rect 33852 23998 33854 24050
rect 33906 23998 33908 24050
rect 33852 23986 33908 23998
rect 33964 24164 34020 24174
rect 33740 23886 33742 23938
rect 33794 23886 33796 23938
rect 33740 23874 33796 23886
rect 33964 23938 34020 24108
rect 33964 23886 33966 23938
rect 34018 23886 34020 23938
rect 33964 23874 34020 23886
rect 34076 22372 34132 25116
rect 34188 25060 34244 25070
rect 34188 24722 34244 25004
rect 35532 24948 35588 27692
rect 35644 26908 35700 29148
rect 35868 28644 35924 28654
rect 35644 26852 35812 26908
rect 35532 24882 35588 24892
rect 34188 24670 34190 24722
rect 34242 24670 34244 24722
rect 34188 24658 34244 24670
rect 34972 24610 35028 24622
rect 34972 24558 34974 24610
rect 35026 24558 35028 24610
rect 34636 24388 34692 24398
rect 34188 24276 34244 24286
rect 34188 23940 34244 24220
rect 34524 23940 34580 23950
rect 34188 23938 34580 23940
rect 34188 23886 34526 23938
rect 34578 23886 34580 23938
rect 34188 23884 34580 23886
rect 34188 23826 34244 23884
rect 34524 23874 34580 23884
rect 34188 23774 34190 23826
rect 34242 23774 34244 23826
rect 34188 23762 34244 23774
rect 34636 23156 34692 24332
rect 34748 24164 34804 24174
rect 34804 24108 34916 24164
rect 34748 24098 34804 24108
rect 34748 23828 34804 23838
rect 34860 23828 34916 24108
rect 34972 24052 35028 24558
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 34972 23986 35028 23996
rect 35644 24052 35700 24062
rect 35644 23958 35700 23996
rect 35084 23940 35140 23950
rect 35532 23940 35588 23950
rect 35084 23938 35588 23940
rect 35084 23886 35086 23938
rect 35138 23886 35534 23938
rect 35586 23886 35588 23938
rect 35084 23884 35588 23886
rect 35084 23874 35140 23884
rect 35532 23874 35588 23884
rect 35756 23938 35812 26852
rect 35756 23886 35758 23938
rect 35810 23886 35812 23938
rect 35756 23874 35812 23886
rect 34972 23828 35028 23838
rect 34860 23826 35028 23828
rect 34860 23774 34974 23826
rect 35026 23774 35028 23826
rect 34860 23772 35028 23774
rect 34748 23604 34804 23772
rect 34972 23762 35028 23772
rect 35196 23714 35252 23726
rect 35196 23662 35198 23714
rect 35250 23662 35252 23714
rect 35196 23604 35252 23662
rect 34748 23548 35252 23604
rect 34636 23090 34692 23100
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 35420 22596 35476 22606
rect 33964 22316 34132 22372
rect 35196 22372 35252 22382
rect 33852 21474 33908 21486
rect 33852 21422 33854 21474
rect 33906 21422 33908 21474
rect 33852 20914 33908 21422
rect 33964 21252 34020 22316
rect 33964 21186 34020 21196
rect 34076 22148 34132 22158
rect 35196 22148 35252 22316
rect 34076 21026 34132 22092
rect 34972 22146 35252 22148
rect 34972 22094 35198 22146
rect 35250 22094 35252 22146
rect 34972 22092 35252 22094
rect 34076 20974 34078 21026
rect 34130 20974 34132 21026
rect 34076 20962 34132 20974
rect 34188 22036 34244 22046
rect 33852 20862 33854 20914
rect 33906 20862 33908 20914
rect 33852 20850 33908 20862
rect 33964 20916 34020 20926
rect 33964 20802 34020 20860
rect 33964 20750 33966 20802
rect 34018 20750 34020 20802
rect 33964 20738 34020 20750
rect 34188 20018 34244 21980
rect 34412 21812 34468 21822
rect 34412 20802 34468 21756
rect 34972 21028 35028 22092
rect 35196 22082 35252 22092
rect 35420 22370 35476 22540
rect 35420 22318 35422 22370
rect 35474 22318 35476 22370
rect 35420 22036 35476 22318
rect 35756 22148 35812 22158
rect 35756 22054 35812 22092
rect 35420 21970 35476 21980
rect 35196 21924 35252 21934
rect 34972 20962 35028 20972
rect 35084 21868 35196 21924
rect 34412 20750 34414 20802
rect 34466 20750 34468 20802
rect 34412 20738 34468 20750
rect 34860 20916 34916 20926
rect 34860 20802 34916 20860
rect 34860 20750 34862 20802
rect 34914 20750 34916 20802
rect 34860 20738 34916 20750
rect 34636 20580 34692 20590
rect 34636 20486 34692 20524
rect 34748 20578 34804 20590
rect 34748 20526 34750 20578
rect 34802 20526 34804 20578
rect 34748 20356 34804 20526
rect 34972 20580 35028 20590
rect 34972 20486 35028 20524
rect 34300 20300 34804 20356
rect 34300 20130 34356 20300
rect 34300 20078 34302 20130
rect 34354 20078 34356 20130
rect 34300 20066 34356 20078
rect 34188 19966 34190 20018
rect 34242 19966 34244 20018
rect 34188 19954 34244 19966
rect 34748 19796 34804 19806
rect 33628 18732 33796 18788
rect 33404 18508 33684 18564
rect 31948 17780 32004 17790
rect 31948 17686 32004 17724
rect 33516 17108 33572 17118
rect 33516 17014 33572 17052
rect 32060 16994 32116 17006
rect 32060 16942 32062 16994
rect 32114 16942 32116 16994
rect 31836 16828 32004 16884
rect 31836 16660 31892 16670
rect 31500 16146 31556 16156
rect 31612 16658 31892 16660
rect 31612 16606 31838 16658
rect 31890 16606 31892 16658
rect 31612 16604 31892 16606
rect 31612 16322 31668 16604
rect 31836 16594 31892 16604
rect 31948 16436 32004 16828
rect 31612 16270 31614 16322
rect 31666 16270 31668 16322
rect 31388 16046 31390 16098
rect 31442 16046 31444 16098
rect 31388 15876 31444 16046
rect 31388 15820 31556 15876
rect 31276 15484 31444 15540
rect 30940 15428 30996 15438
rect 30380 15426 30996 15428
rect 30380 15374 30942 15426
rect 30994 15374 30996 15426
rect 30380 15372 30996 15374
rect 30492 15314 30548 15372
rect 30940 15362 30996 15372
rect 30492 15262 30494 15314
rect 30546 15262 30548 15314
rect 30492 15250 30548 15262
rect 30156 14478 30158 14530
rect 30210 14478 30212 14530
rect 30156 14466 30212 14478
rect 30828 14532 30884 14542
rect 30828 14438 30884 14476
rect 31276 14532 31332 14542
rect 29820 14420 29876 14430
rect 29820 14326 29876 14364
rect 29932 14306 29988 14318
rect 29932 14254 29934 14306
rect 29986 14254 29988 14306
rect 29932 13636 29988 14254
rect 30940 13746 30996 13758
rect 30940 13694 30942 13746
rect 30994 13694 30996 13746
rect 30156 13636 30212 13646
rect 30604 13636 30660 13646
rect 29708 13634 30212 13636
rect 29708 13582 29710 13634
rect 29762 13582 30158 13634
rect 30210 13582 30212 13634
rect 29708 13580 30212 13582
rect 29708 13570 29764 13580
rect 29596 12292 29652 12302
rect 29596 12180 29652 12236
rect 29260 12178 29652 12180
rect 29260 12126 29598 12178
rect 29650 12126 29652 12178
rect 29260 12124 29652 12126
rect 29036 11284 29092 11294
rect 29036 11190 29092 11228
rect 29260 11282 29316 12124
rect 29260 11230 29262 11282
rect 29314 11230 29316 11282
rect 29260 11218 29316 11230
rect 29372 11284 29428 11294
rect 29372 11190 29428 11228
rect 29596 10836 29652 12124
rect 29820 12290 29876 12302
rect 29820 12238 29822 12290
rect 29874 12238 29876 12290
rect 29820 11956 29876 12238
rect 29820 11890 29876 11900
rect 30044 11396 30100 13580
rect 30156 13570 30212 13580
rect 30380 13580 30604 13636
rect 30156 12404 30212 12414
rect 30156 12310 30212 12348
rect 30380 11732 30436 13580
rect 30604 13542 30660 13580
rect 30380 11666 30436 11676
rect 30492 12962 30548 12974
rect 30492 12910 30494 12962
rect 30546 12910 30548 12962
rect 30492 12180 30548 12910
rect 30716 12740 30772 12750
rect 30716 12290 30772 12684
rect 30716 12238 30718 12290
rect 30770 12238 30772 12290
rect 30604 12180 30660 12190
rect 30492 12178 30660 12180
rect 30492 12126 30606 12178
rect 30658 12126 30660 12178
rect 30492 12124 30660 12126
rect 30044 11340 30436 11396
rect 29596 10742 29652 10780
rect 29708 11284 29764 11294
rect 29708 11172 29764 11228
rect 29820 11172 29876 11182
rect 30268 11172 30324 11182
rect 29708 11170 30324 11172
rect 29708 11118 29822 11170
rect 29874 11118 30270 11170
rect 30322 11118 30324 11170
rect 29708 11116 30324 11118
rect 28924 10668 29540 10724
rect 29148 10500 29204 10510
rect 28700 10498 29204 10500
rect 28700 10446 29150 10498
rect 29202 10446 29204 10498
rect 28700 10444 29204 10446
rect 29148 10434 29204 10444
rect 28588 10332 28868 10388
rect 27020 10322 27076 10332
rect 26348 9154 26740 9156
rect 26348 9102 26350 9154
rect 26402 9102 26740 9154
rect 26348 9100 26740 9102
rect 26796 9940 26852 9950
rect 26796 9154 26852 9884
rect 28588 9828 28644 9838
rect 28476 9716 28532 9726
rect 27916 9602 27972 9614
rect 27916 9550 27918 9602
rect 27970 9550 27972 9602
rect 26796 9102 26798 9154
rect 26850 9102 26852 9154
rect 26348 9090 26404 9100
rect 26796 9090 26852 9102
rect 27580 9156 27636 9166
rect 27468 9044 27524 9054
rect 26908 8820 26964 8830
rect 25564 8034 26068 8036
rect 25564 7982 25566 8034
rect 25618 7982 26068 8034
rect 25564 7980 26068 7982
rect 26236 8036 26292 8046
rect 25564 7970 25620 7980
rect 26236 7698 26292 7980
rect 26236 7646 26238 7698
rect 26290 7646 26292 7698
rect 26236 7634 26292 7646
rect 26908 8034 26964 8764
rect 26908 7982 26910 8034
rect 26962 7982 26964 8034
rect 24668 7586 25284 7588
rect 24668 7534 24670 7586
rect 24722 7534 25284 7586
rect 24668 7532 25284 7534
rect 26460 7586 26516 7598
rect 26460 7534 26462 7586
rect 26514 7534 26516 7586
rect 24668 7522 24724 7532
rect 24332 6862 24334 6914
rect 24386 6862 24388 6914
rect 24332 6850 24388 6862
rect 24444 7476 24500 7486
rect 24220 6626 24276 6636
rect 24444 6690 24500 7420
rect 26460 7140 26516 7534
rect 26908 7586 26964 7982
rect 26908 7534 26910 7586
rect 26962 7534 26964 7586
rect 26908 7522 26964 7534
rect 27020 8316 27300 8372
rect 27020 7586 27076 8316
rect 27244 8260 27300 8316
rect 27020 7534 27022 7586
rect 27074 7534 27076 7586
rect 26460 7074 26516 7084
rect 26572 7474 26628 7486
rect 26572 7422 26574 7474
rect 26626 7422 26628 7474
rect 24444 6638 24446 6690
rect 24498 6638 24500 6690
rect 24444 6626 24500 6638
rect 24668 6802 24724 6814
rect 24668 6750 24670 6802
rect 24722 6750 24724 6802
rect 24668 6692 24724 6750
rect 24668 6626 24724 6636
rect 25340 6692 25396 6702
rect 14812 6526 14814 6578
rect 14866 6526 14868 6578
rect 14812 6514 14868 6526
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 25340 6130 25396 6636
rect 26124 6692 26180 6702
rect 26124 6578 26180 6636
rect 26124 6526 26126 6578
rect 26178 6526 26180 6578
rect 26124 6514 26180 6526
rect 25788 6466 25844 6478
rect 25788 6414 25790 6466
rect 25842 6414 25844 6466
rect 25340 6078 25342 6130
rect 25394 6078 25396 6130
rect 25340 6066 25396 6078
rect 25564 6132 25620 6142
rect 25788 6132 25844 6414
rect 25564 6130 25844 6132
rect 25564 6078 25566 6130
rect 25618 6078 25844 6130
rect 25564 6076 25844 6078
rect 25564 6066 25620 6076
rect 25676 5908 25732 5918
rect 14364 5852 14756 5908
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 14140 3444 14196 3454
rect 14364 3444 14420 3454
rect 14140 3442 14420 3444
rect 14140 3390 14142 3442
rect 14194 3390 14366 3442
rect 14418 3390 14420 3442
rect 14140 3388 14420 3390
rect 14140 800 14196 3388
rect 14364 3378 14420 3388
rect 14700 3442 14756 5852
rect 25676 5814 25732 5852
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 14700 3390 14702 3442
rect 14754 3390 14756 3442
rect 14700 3378 14756 3390
rect 25116 3556 25172 3566
rect 25116 3388 25172 3500
rect 25564 3442 25620 3454
rect 25564 3390 25566 3442
rect 25618 3390 25620 3442
rect 21756 3332 21812 3342
rect 25116 3332 25284 3388
rect 21532 3330 21812 3332
rect 21532 3278 21758 3330
rect 21810 3278 21812 3330
rect 21532 3276 21812 3278
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 21532 800 21588 3276
rect 21756 3266 21812 3276
rect 25228 3108 25284 3332
rect 25564 3220 25620 3390
rect 25788 3442 25844 6076
rect 26460 6466 26516 6478
rect 26460 6414 26462 6466
rect 26514 6414 26516 6466
rect 26460 6132 26516 6414
rect 26460 5908 26516 6076
rect 26572 6244 26628 7422
rect 27020 7252 27076 7534
rect 27020 7186 27076 7196
rect 27132 8146 27188 8158
rect 27132 8094 27134 8146
rect 27186 8094 27188 8146
rect 27132 6916 27188 8094
rect 27244 8146 27300 8204
rect 27468 8258 27524 8988
rect 27580 9042 27636 9100
rect 27580 8990 27582 9042
rect 27634 8990 27636 9042
rect 27580 8978 27636 8990
rect 27916 8820 27972 9550
rect 27916 8754 27972 8764
rect 28252 9602 28308 9614
rect 28252 9550 28254 9602
rect 28306 9550 28308 9602
rect 28140 8372 28196 8382
rect 28140 8278 28196 8316
rect 27468 8206 27470 8258
rect 27522 8206 27524 8258
rect 27468 8194 27524 8206
rect 28252 8260 28308 9550
rect 28252 8194 28308 8204
rect 27244 8094 27246 8146
rect 27298 8094 27300 8146
rect 27244 8082 27300 8094
rect 27468 8036 27524 8046
rect 27356 7980 27468 8036
rect 27244 7700 27300 7710
rect 27356 7700 27412 7980
rect 27468 7970 27524 7980
rect 28028 8036 28084 8046
rect 28028 7942 28084 7980
rect 28252 8034 28308 8046
rect 28252 7982 28254 8034
rect 28306 7982 28308 8034
rect 27244 7698 27412 7700
rect 27244 7646 27246 7698
rect 27298 7646 27412 7698
rect 27244 7644 27412 7646
rect 27244 7634 27300 7644
rect 27692 7474 27748 7486
rect 27692 7422 27694 7474
rect 27746 7422 27748 7474
rect 27580 7364 27636 7374
rect 26796 6860 27132 6916
rect 26796 6578 26852 6860
rect 27132 6822 27188 6860
rect 27244 7362 27636 7364
rect 27244 7310 27582 7362
rect 27634 7310 27636 7362
rect 27244 7308 27636 7310
rect 26796 6526 26798 6578
rect 26850 6526 26852 6578
rect 26796 6468 26852 6526
rect 26796 6402 26852 6412
rect 26908 6692 26964 6702
rect 27244 6692 27300 7308
rect 27580 7298 27636 7308
rect 27580 7140 27636 7150
rect 26572 6020 26628 6188
rect 26796 6132 26852 6142
rect 26908 6132 26964 6636
rect 26796 6130 26964 6132
rect 26796 6078 26798 6130
rect 26850 6078 26964 6130
rect 26796 6076 26964 6078
rect 27020 6636 27300 6692
rect 27468 6804 27524 6814
rect 27020 6130 27076 6636
rect 27468 6578 27524 6748
rect 27468 6526 27470 6578
rect 27522 6526 27524 6578
rect 27468 6514 27524 6526
rect 27020 6078 27022 6130
rect 27074 6078 27076 6130
rect 26796 6066 26852 6076
rect 27020 6066 27076 6078
rect 27132 6466 27188 6478
rect 27132 6414 27134 6466
rect 27186 6414 27188 6466
rect 27132 6244 27188 6414
rect 26684 6020 26740 6030
rect 26572 6018 26740 6020
rect 26572 5966 26686 6018
rect 26738 5966 26740 6018
rect 26572 5964 26740 5966
rect 26684 5954 26740 5964
rect 26460 5460 26516 5852
rect 27132 5684 27188 6188
rect 27244 6468 27300 6478
rect 27244 6018 27300 6412
rect 27580 6356 27636 7084
rect 27468 6300 27636 6356
rect 27356 6244 27412 6254
rect 27356 6130 27412 6188
rect 27356 6078 27358 6130
rect 27410 6078 27412 6130
rect 27356 6066 27412 6078
rect 27244 5966 27246 6018
rect 27298 5966 27300 6018
rect 27244 5954 27300 5966
rect 27244 5684 27300 5694
rect 27132 5628 27244 5684
rect 27244 5618 27300 5628
rect 26460 5404 26628 5460
rect 26012 3556 26068 3566
rect 26012 3462 26068 3500
rect 25788 3390 25790 3442
rect 25842 3390 25844 3442
rect 25788 3378 25844 3390
rect 26460 3442 26516 3454
rect 26460 3390 26462 3442
rect 26514 3390 26516 3442
rect 26460 3388 26516 3390
rect 26572 3444 26628 5404
rect 26908 4226 26964 4238
rect 26908 4174 26910 4226
rect 26962 4174 26964 4226
rect 26796 3444 26852 3454
rect 26572 3442 26852 3444
rect 26572 3390 26798 3442
rect 26850 3390 26852 3442
rect 26572 3388 26852 3390
rect 26236 3332 26516 3388
rect 26796 3378 26852 3388
rect 26908 3332 26964 4174
rect 27132 3442 27188 3454
rect 27132 3390 27134 3442
rect 27186 3390 27188 3442
rect 27132 3332 27188 3390
rect 27468 3442 27524 6300
rect 27580 6132 27636 6142
rect 27692 6132 27748 7422
rect 28028 6804 28084 6814
rect 27916 6690 27972 6702
rect 27916 6638 27918 6690
rect 27970 6638 27972 6690
rect 27916 6580 27972 6638
rect 27916 6514 27972 6524
rect 28028 6466 28084 6748
rect 28252 6802 28308 7982
rect 28252 6750 28254 6802
rect 28306 6750 28308 6802
rect 28252 6738 28308 6750
rect 28364 6916 28420 6926
rect 28364 6690 28420 6860
rect 28364 6638 28366 6690
rect 28418 6638 28420 6690
rect 28364 6626 28420 6638
rect 28476 6692 28532 9660
rect 28588 9714 28644 9772
rect 28588 9662 28590 9714
rect 28642 9662 28644 9714
rect 28588 9650 28644 9662
rect 28588 9044 28644 9054
rect 28588 8950 28644 8988
rect 28812 8820 28868 10332
rect 29260 9826 29316 9838
rect 29260 9774 29262 9826
rect 29314 9774 29316 9826
rect 29260 9716 29316 9774
rect 29260 9650 29316 9660
rect 29036 8932 29092 8942
rect 29036 8838 29092 8876
rect 28812 8754 28868 8764
rect 28700 8260 28756 8270
rect 28700 8258 29316 8260
rect 28700 8206 28702 8258
rect 28754 8206 29316 8258
rect 28700 8204 29316 8206
rect 28700 8194 28756 8204
rect 29036 8036 29092 8046
rect 29036 7474 29092 7980
rect 29036 7422 29038 7474
rect 29090 7422 29092 7474
rect 29036 7410 29092 7422
rect 29260 6914 29316 8204
rect 29260 6862 29262 6914
rect 29314 6862 29316 6914
rect 29260 6850 29316 6862
rect 29372 6916 29428 6926
rect 29148 6692 29204 6702
rect 28476 6690 29204 6692
rect 28476 6638 29150 6690
rect 29202 6638 29204 6690
rect 28476 6636 29204 6638
rect 28028 6414 28030 6466
rect 28082 6414 28084 6466
rect 28028 6244 28084 6414
rect 28252 6468 28308 6478
rect 28252 6374 28308 6412
rect 28476 6244 28532 6636
rect 29148 6626 29204 6636
rect 29372 6690 29428 6860
rect 29372 6638 29374 6690
rect 29426 6638 29428 6690
rect 29372 6626 29428 6638
rect 28028 6188 28532 6244
rect 27580 6130 27748 6132
rect 27580 6078 27582 6130
rect 27634 6078 27748 6130
rect 27580 6076 27748 6078
rect 27580 6066 27636 6076
rect 29484 5908 29540 10668
rect 29708 9826 29764 11116
rect 29820 11106 29876 11116
rect 30268 11106 30324 11116
rect 30380 10948 30436 11340
rect 30380 10882 30436 10892
rect 29932 10610 29988 10622
rect 29932 10558 29934 10610
rect 29986 10558 29988 10610
rect 29708 9774 29710 9826
rect 29762 9774 29764 9826
rect 29708 9380 29764 9774
rect 29708 9314 29764 9324
rect 29820 10052 29876 10062
rect 29820 7586 29876 9996
rect 29932 9156 29988 10558
rect 30492 10052 30548 12124
rect 30604 12114 30660 12124
rect 30716 11284 30772 12238
rect 30940 12178 30996 13694
rect 31276 13186 31332 14476
rect 31276 13134 31278 13186
rect 31330 13134 31332 13186
rect 31276 13122 31332 13134
rect 31164 12962 31220 12974
rect 31164 12910 31166 12962
rect 31218 12910 31220 12962
rect 31164 12402 31220 12910
rect 31388 12516 31444 15484
rect 31500 15316 31556 15820
rect 31500 15250 31556 15260
rect 31612 15202 31668 16270
rect 31612 15150 31614 15202
rect 31666 15150 31668 15202
rect 31612 14754 31668 15150
rect 31612 14702 31614 14754
rect 31666 14702 31668 14754
rect 31612 14690 31668 14702
rect 31836 16380 32004 16436
rect 31500 14530 31556 14542
rect 31500 14478 31502 14530
rect 31554 14478 31556 14530
rect 31500 14308 31556 14478
rect 31500 14242 31556 14252
rect 31164 12350 31166 12402
rect 31218 12350 31220 12402
rect 31164 12338 31220 12350
rect 31276 12460 31444 12516
rect 31276 12180 31332 12460
rect 31388 12292 31444 12302
rect 31388 12198 31444 12236
rect 30940 12126 30942 12178
rect 30994 12126 30996 12178
rect 30940 11956 30996 12126
rect 30940 11890 30996 11900
rect 31164 12124 31332 12180
rect 31500 12178 31556 12190
rect 31500 12126 31502 12178
rect 31554 12126 31556 12178
rect 30940 11284 30996 11294
rect 30716 11282 30996 11284
rect 30716 11230 30942 11282
rect 30994 11230 30996 11282
rect 30716 11228 30996 11230
rect 30940 11218 30996 11228
rect 31164 10948 31220 12124
rect 31276 11172 31332 11182
rect 31500 11172 31556 12126
rect 31276 11170 31556 11172
rect 31276 11118 31278 11170
rect 31330 11118 31556 11170
rect 31276 11116 31556 11118
rect 31276 11106 31332 11116
rect 31164 10892 31332 10948
rect 30492 9986 30548 9996
rect 30604 10722 30660 10734
rect 30604 10670 30606 10722
rect 30658 10670 30660 10722
rect 30604 10050 30660 10670
rect 30604 9998 30606 10050
rect 30658 9998 30660 10050
rect 30604 9986 30660 9998
rect 31164 10610 31220 10622
rect 31164 10558 31166 10610
rect 31218 10558 31220 10610
rect 31164 10050 31220 10558
rect 31164 9998 31166 10050
rect 31218 9998 31220 10050
rect 31164 9986 31220 9998
rect 30716 9714 30772 9726
rect 30716 9662 30718 9714
rect 30770 9662 30772 9714
rect 30604 9602 30660 9614
rect 30604 9550 30606 9602
rect 30658 9550 30660 9602
rect 30604 9156 30660 9550
rect 30716 9268 30772 9662
rect 31052 9716 31108 9726
rect 31052 9622 31108 9660
rect 30716 9202 30772 9212
rect 31164 9602 31220 9614
rect 31164 9550 31166 9602
rect 31218 9550 31220 9602
rect 29932 9100 30660 9156
rect 29820 7534 29822 7586
rect 29874 7534 29876 7586
rect 29820 7522 29876 7534
rect 29820 7364 29876 7374
rect 29596 6692 29652 6702
rect 29596 6468 29652 6636
rect 29820 6690 29876 7308
rect 29820 6638 29822 6690
rect 29874 6638 29876 6690
rect 29820 6626 29876 6638
rect 29596 6402 29652 6412
rect 29932 5908 29988 5918
rect 29484 5906 29988 5908
rect 29484 5854 29934 5906
rect 29986 5854 29988 5906
rect 29484 5852 29988 5854
rect 29932 5842 29988 5852
rect 27468 3390 27470 3442
rect 27522 3390 27524 3442
rect 27468 3378 27524 3390
rect 28028 5682 28084 5694
rect 28028 5630 28030 5682
rect 28082 5630 28084 5682
rect 28028 3388 28084 5630
rect 28700 5236 28756 5246
rect 28700 5234 29876 5236
rect 28700 5182 28702 5234
rect 28754 5182 29876 5234
rect 28700 5180 29876 5182
rect 28700 5170 28756 5180
rect 28812 5012 28868 5022
rect 28252 4226 28308 4238
rect 28252 4174 28254 4226
rect 28306 4174 28308 4226
rect 28252 3444 28308 4174
rect 28700 4116 28756 4126
rect 28476 4114 28756 4116
rect 28476 4062 28702 4114
rect 28754 4062 28756 4114
rect 28476 4060 28756 4062
rect 28364 3444 28420 3482
rect 28252 3388 28364 3444
rect 26236 3220 26292 3332
rect 25564 3164 26292 3220
rect 25228 3052 25620 3108
rect 25564 800 25620 3052
rect 26236 800 26292 3164
rect 26908 3276 27188 3332
rect 27692 3332 28084 3388
rect 28364 3378 28420 3388
rect 26908 800 26964 3276
rect 27692 980 27748 3332
rect 28476 2100 28532 4060
rect 28700 4050 28756 4060
rect 28700 3444 28756 3454
rect 28812 3444 28868 4956
rect 29372 5012 29428 5022
rect 29372 4918 29428 4956
rect 29484 5010 29540 5022
rect 29484 4958 29486 5010
rect 29538 4958 29540 5010
rect 29148 4898 29204 4910
rect 29148 4846 29150 4898
rect 29202 4846 29204 4898
rect 29148 3892 29204 4846
rect 29484 4564 29540 4958
rect 29484 4498 29540 4508
rect 29148 3836 29428 3892
rect 28700 3442 28868 3444
rect 28700 3390 28702 3442
rect 28754 3390 28868 3442
rect 28700 3388 28868 3390
rect 29260 3666 29316 3678
rect 29260 3614 29262 3666
rect 29314 3614 29316 3666
rect 29260 3388 29316 3614
rect 28700 3378 28756 3388
rect 27580 924 27748 980
rect 28252 2044 28532 2100
rect 29148 3332 29316 3388
rect 27580 800 27636 924
rect 28252 800 28308 2044
rect 29148 980 29204 3332
rect 29372 3220 29428 3836
rect 29372 3154 29428 3164
rect 28924 924 29204 980
rect 28924 800 28980 924
rect 29596 800 29652 5180
rect 29820 5122 29876 5180
rect 29820 5070 29822 5122
rect 29874 5070 29876 5122
rect 29820 5058 29876 5070
rect 30156 5010 30212 9100
rect 31164 9044 31220 9550
rect 30268 8932 30324 8942
rect 30268 8484 30324 8876
rect 30380 8484 30436 8494
rect 30268 8482 30436 8484
rect 30268 8430 30382 8482
rect 30434 8430 30436 8482
rect 30268 8428 30436 8430
rect 30380 8418 30436 8428
rect 30492 8148 30548 8158
rect 30492 8054 30548 8092
rect 30940 8148 30996 8158
rect 30380 8036 30436 8046
rect 30380 7942 30436 7980
rect 30828 8036 30884 8046
rect 30940 8036 30996 8092
rect 31164 8146 31220 8988
rect 31164 8094 31166 8146
rect 31218 8094 31220 8146
rect 31164 8082 31220 8094
rect 30828 8034 30996 8036
rect 30828 7982 30830 8034
rect 30882 7982 30996 8034
rect 30828 7980 30996 7982
rect 30604 7588 30660 7598
rect 30604 7494 30660 7532
rect 30380 7476 30436 7486
rect 30380 7382 30436 7420
rect 30716 7476 30772 7486
rect 30828 7476 30884 7980
rect 31164 7476 31220 7486
rect 30716 7474 31220 7476
rect 30716 7422 30718 7474
rect 30770 7422 31166 7474
rect 31218 7422 31220 7474
rect 30716 7420 31220 7422
rect 30716 7410 30772 7420
rect 30940 6468 30996 6478
rect 30940 6466 31108 6468
rect 30940 6414 30942 6466
rect 30994 6414 31108 6466
rect 30940 6412 31108 6414
rect 30940 6402 30996 6412
rect 31052 5908 31108 6412
rect 31164 6130 31220 7420
rect 31164 6078 31166 6130
rect 31218 6078 31220 6130
rect 31164 6066 31220 6078
rect 31052 5842 31108 5852
rect 30940 5796 30996 5806
rect 31276 5796 31332 10892
rect 31388 9716 31444 11116
rect 31836 10052 31892 16380
rect 32060 16324 32116 16942
rect 33292 16884 33348 16894
rect 33292 16790 33348 16828
rect 33068 16772 33124 16782
rect 32172 16660 32228 16670
rect 32172 16658 32564 16660
rect 32172 16606 32174 16658
rect 32226 16606 32564 16658
rect 32172 16604 32564 16606
rect 32172 16594 32228 16604
rect 32060 16258 32116 16268
rect 32508 16322 32564 16604
rect 32508 16270 32510 16322
rect 32562 16270 32564 16322
rect 32508 16258 32564 16270
rect 32956 16212 33012 16222
rect 32956 16118 33012 16156
rect 31948 16100 32004 16110
rect 32284 16100 32340 16110
rect 31948 16098 32340 16100
rect 31948 16046 31950 16098
rect 32002 16046 32286 16098
rect 32338 16046 32340 16098
rect 31948 16044 32340 16046
rect 31948 16034 32004 16044
rect 32284 16034 32340 16044
rect 32844 16098 32900 16110
rect 32844 16046 32846 16098
rect 32898 16046 32900 16098
rect 32844 15652 32900 16046
rect 32844 15586 32900 15596
rect 32956 15876 33012 15886
rect 33068 15876 33124 16716
rect 33180 16100 33236 16110
rect 33180 16006 33236 16044
rect 32956 15874 33124 15876
rect 32956 15822 32958 15874
rect 33010 15822 33124 15874
rect 32956 15820 33124 15822
rect 32060 15314 32116 15326
rect 32060 15262 32062 15314
rect 32114 15262 32116 15314
rect 32060 14756 32116 15262
rect 32956 15204 33012 15820
rect 33292 15426 33348 15438
rect 33292 15374 33294 15426
rect 33346 15374 33348 15426
rect 32956 15138 33012 15148
rect 33180 15316 33236 15326
rect 33180 15202 33236 15260
rect 33180 15150 33182 15202
rect 33234 15150 33236 15202
rect 33180 15138 33236 15150
rect 32172 14756 32228 14766
rect 32060 14754 32228 14756
rect 32060 14702 32174 14754
rect 32226 14702 32228 14754
rect 32060 14700 32228 14702
rect 32172 14690 32228 14700
rect 33180 14532 33236 14542
rect 33292 14532 33348 15374
rect 33236 14476 33348 14532
rect 33516 15314 33572 15326
rect 33516 15262 33518 15314
rect 33570 15262 33572 15314
rect 33516 14642 33572 15262
rect 33628 15148 33684 18508
rect 33740 18340 33796 18732
rect 33740 18274 33796 18284
rect 34412 17780 34468 17790
rect 34076 17554 34132 17566
rect 34076 17502 34078 17554
rect 34130 17502 34132 17554
rect 34076 17108 34132 17502
rect 34076 17042 34132 17052
rect 34412 16996 34468 17724
rect 34076 16884 34132 16894
rect 34076 16790 34132 16828
rect 34412 16770 34468 16940
rect 34412 16718 34414 16770
rect 34466 16718 34468 16770
rect 34412 16706 34468 16718
rect 34748 17108 34804 19740
rect 35084 18452 35140 21868
rect 35196 21858 35252 21868
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 35868 20916 35924 28588
rect 36092 28644 36148 28654
rect 36092 28530 36148 28588
rect 36092 28478 36094 28530
rect 36146 28478 36148 28530
rect 36092 28466 36148 28478
rect 36204 28530 36260 29148
rect 36988 28868 37044 29708
rect 37100 29540 37156 29550
rect 37100 29446 37156 29484
rect 37212 29316 37268 29934
rect 37660 29988 37716 30158
rect 38668 30210 38724 30492
rect 38892 30548 38948 30558
rect 39340 30548 39396 30830
rect 38668 30158 38670 30210
rect 38722 30158 38724 30210
rect 38668 30146 38724 30158
rect 38780 30436 38836 30446
rect 37660 29922 37716 29932
rect 37772 29986 37828 29998
rect 37772 29934 37774 29986
rect 37826 29934 37828 29986
rect 37772 29652 37828 29934
rect 37324 29596 37828 29652
rect 37884 29988 37940 29998
rect 38108 29988 38164 29998
rect 37324 29538 37380 29596
rect 37324 29486 37326 29538
rect 37378 29486 37380 29538
rect 37324 29474 37380 29486
rect 37884 29540 37940 29932
rect 37884 29474 37940 29484
rect 37996 29986 38164 29988
rect 37996 29934 38110 29986
rect 38162 29934 38164 29986
rect 37996 29932 38164 29934
rect 37212 29250 37268 29260
rect 37996 28980 38052 29932
rect 38108 29922 38164 29932
rect 38444 29652 38500 29662
rect 38444 29202 38500 29596
rect 38668 29426 38724 29438
rect 38668 29374 38670 29426
rect 38722 29374 38724 29426
rect 38668 29316 38724 29374
rect 38780 29428 38836 30380
rect 38892 30434 38948 30492
rect 38892 30382 38894 30434
rect 38946 30382 38948 30434
rect 38892 30370 38948 30382
rect 39004 30492 39396 30548
rect 39004 30212 39060 30492
rect 39900 30436 39956 30446
rect 39228 30434 39956 30436
rect 39228 30382 39902 30434
rect 39954 30382 39956 30434
rect 39228 30380 39956 30382
rect 39228 30322 39284 30380
rect 39900 30370 39956 30380
rect 39228 30270 39230 30322
rect 39282 30270 39284 30322
rect 39228 30258 39284 30270
rect 38780 29372 38948 29428
rect 38724 29260 38836 29316
rect 38668 29250 38724 29260
rect 38444 29150 38446 29202
rect 38498 29150 38500 29202
rect 38444 29138 38500 29150
rect 37660 28924 38052 28980
rect 36988 28812 37604 28868
rect 37548 28756 37604 28812
rect 37100 28644 37156 28654
rect 36204 28478 36206 28530
rect 36258 28478 36260 28530
rect 36204 28466 36260 28478
rect 36988 28642 37156 28644
rect 36988 28590 37102 28642
rect 37154 28590 37156 28642
rect 36988 28588 37156 28590
rect 36428 28418 36484 28430
rect 36428 28366 36430 28418
rect 36482 28366 36484 28418
rect 36428 26908 36484 28366
rect 36316 26852 36484 26908
rect 36988 27972 37044 28588
rect 37100 28578 37156 28588
rect 36204 24500 36260 24510
rect 36204 23938 36260 24444
rect 36204 23886 36206 23938
rect 36258 23886 36260 23938
rect 36204 23874 36260 23886
rect 35980 22708 36036 22718
rect 35980 22258 36036 22652
rect 35980 22206 35982 22258
rect 36034 22206 36036 22258
rect 35980 21474 36036 22206
rect 36092 22258 36148 22270
rect 36092 22206 36094 22258
rect 36146 22206 36148 22258
rect 36092 22148 36148 22206
rect 36092 22082 36148 22092
rect 36316 21924 36372 26852
rect 36988 26516 37044 27916
rect 37436 27860 37492 27870
rect 36876 26460 37044 26516
rect 37100 27188 37156 27198
rect 37100 26514 37156 27132
rect 37436 26962 37492 27804
rect 37548 27524 37604 28700
rect 37660 28644 37716 28924
rect 37660 28550 37716 28588
rect 38108 28644 38164 28654
rect 38108 28084 38164 28588
rect 38220 28420 38276 28430
rect 38276 28364 38388 28420
rect 38220 28354 38276 28364
rect 37660 28082 38164 28084
rect 37660 28030 38110 28082
rect 38162 28030 38164 28082
rect 37660 28028 38164 28030
rect 37660 27746 37716 28028
rect 38108 28018 38164 28028
rect 38332 28082 38388 28364
rect 38332 28030 38334 28082
rect 38386 28030 38388 28082
rect 38332 28018 38388 28030
rect 38444 28418 38500 28430
rect 38444 28366 38446 28418
rect 38498 28366 38500 28418
rect 38444 28082 38500 28366
rect 38668 28420 38724 28430
rect 38668 28326 38724 28364
rect 38444 28030 38446 28082
rect 38498 28030 38500 28082
rect 38444 28018 38500 28030
rect 38668 27972 38724 27982
rect 38668 27878 38724 27916
rect 38780 27970 38836 29260
rect 38892 28642 38948 29372
rect 39004 28756 39060 30156
rect 39788 30212 39844 30222
rect 40012 30212 40068 31276
rect 41356 30996 41412 31836
rect 42364 31892 42420 31902
rect 42364 31798 42420 31836
rect 42476 31778 42532 31948
rect 42476 31726 42478 31778
rect 42530 31726 42532 31778
rect 42476 31714 42532 31726
rect 43372 31666 43428 31948
rect 43372 31614 43374 31666
rect 43426 31614 43428 31666
rect 43372 31602 43428 31614
rect 42588 31556 42644 31566
rect 42588 31554 43092 31556
rect 42588 31502 42590 31554
rect 42642 31502 43092 31554
rect 42588 31500 43092 31502
rect 41916 31220 41972 31230
rect 41356 30994 41524 30996
rect 41356 30942 41358 30994
rect 41410 30942 41524 30994
rect 41356 30940 41524 30942
rect 41356 30930 41412 30940
rect 40460 30772 40516 30782
rect 39788 30210 40068 30212
rect 39788 30158 39790 30210
rect 39842 30158 40068 30210
rect 39788 30156 40068 30158
rect 40124 30322 40180 30334
rect 40124 30270 40126 30322
rect 40178 30270 40180 30322
rect 40124 30212 40180 30270
rect 39788 30146 39844 30156
rect 40124 30146 40180 30156
rect 39116 30098 39172 30110
rect 39116 30046 39118 30098
rect 39170 30046 39172 30098
rect 39116 29652 39172 30046
rect 39116 29586 39172 29596
rect 39228 30100 39284 30110
rect 39116 29428 39172 29438
rect 39228 29428 39284 30044
rect 39340 30098 39396 30110
rect 39340 30046 39342 30098
rect 39394 30046 39396 30098
rect 39340 29764 39396 30046
rect 39340 29698 39396 29708
rect 40236 30098 40292 30110
rect 40236 30046 40238 30098
rect 40290 30046 40292 30098
rect 39116 29426 39284 29428
rect 39116 29374 39118 29426
rect 39170 29374 39284 29426
rect 39116 29372 39284 29374
rect 39116 29362 39172 29372
rect 39004 28690 39060 28700
rect 39116 28924 39732 28980
rect 38892 28590 38894 28642
rect 38946 28590 38948 28642
rect 38892 28578 38948 28590
rect 38780 27918 38782 27970
rect 38834 27918 38836 27970
rect 38780 27906 38836 27918
rect 39004 28532 39060 28542
rect 39116 28532 39172 28924
rect 39228 28756 39284 28766
rect 39564 28756 39620 28766
rect 39228 28754 39508 28756
rect 39228 28702 39230 28754
rect 39282 28702 39508 28754
rect 39228 28700 39508 28702
rect 39228 28690 39284 28700
rect 39004 28530 39172 28532
rect 39004 28478 39006 28530
rect 39058 28478 39172 28530
rect 39004 28476 39172 28478
rect 37996 27860 38052 27870
rect 37996 27766 38052 27804
rect 37660 27694 37662 27746
rect 37714 27694 37716 27746
rect 37660 27682 37716 27694
rect 37548 27468 37940 27524
rect 37436 26910 37438 26962
rect 37490 26910 37492 26962
rect 37436 26898 37492 26910
rect 37772 26852 37828 26862
rect 37772 26758 37828 26796
rect 37100 26462 37102 26514
rect 37154 26462 37156 26514
rect 36764 26178 36820 26190
rect 36764 26126 36766 26178
rect 36818 26126 36820 26178
rect 36428 25620 36484 25630
rect 36428 25526 36484 25564
rect 36764 25620 36820 26126
rect 36764 25554 36820 25564
rect 36876 25172 36932 26460
rect 37100 26450 37156 26462
rect 36988 26292 37044 26302
rect 36988 25732 37044 26236
rect 37100 25732 37156 25742
rect 36988 25730 37156 25732
rect 36988 25678 37102 25730
rect 37154 25678 37156 25730
rect 36988 25676 37156 25678
rect 37100 25666 37156 25676
rect 37212 25620 37268 25630
rect 37212 25508 37268 25564
rect 37100 25452 37268 25508
rect 37100 25394 37156 25452
rect 37100 25342 37102 25394
rect 37154 25342 37156 25394
rect 37100 25330 37156 25342
rect 37212 25338 37268 25350
rect 37212 25286 37214 25338
rect 37266 25286 37268 25338
rect 37212 25284 37268 25286
rect 37772 25284 37828 25294
rect 37212 25282 37828 25284
rect 37212 25230 37774 25282
rect 37826 25230 37828 25282
rect 37212 25228 37828 25230
rect 36876 25106 36932 25116
rect 37548 24836 37604 24846
rect 37436 24834 37604 24836
rect 37436 24782 37550 24834
rect 37602 24782 37604 24834
rect 37436 24780 37604 24782
rect 37100 24612 37156 24622
rect 37436 24612 37492 24780
rect 37548 24770 37604 24780
rect 37100 24610 37492 24612
rect 37100 24558 37102 24610
rect 37154 24558 37492 24610
rect 37100 24556 37492 24558
rect 37100 24546 37156 24556
rect 37436 24388 37492 24556
rect 37660 24722 37716 25228
rect 37772 25218 37828 25228
rect 37660 24670 37662 24722
rect 37714 24670 37716 24722
rect 37548 24500 37604 24510
rect 37548 24406 37604 24444
rect 37436 24322 37492 24332
rect 37660 23940 37716 24670
rect 37436 23884 37716 23940
rect 37324 23044 37380 23054
rect 37100 22594 37156 22606
rect 37100 22542 37102 22594
rect 37154 22542 37156 22594
rect 36988 22484 37044 22494
rect 36988 22390 37044 22428
rect 36316 21858 36372 21868
rect 37100 21698 37156 22542
rect 37212 22372 37268 22382
rect 37212 22278 37268 22316
rect 37100 21646 37102 21698
rect 37154 21646 37156 21698
rect 37100 21634 37156 21646
rect 35980 21422 35982 21474
rect 36034 21422 36036 21474
rect 35980 21410 36036 21422
rect 36316 21586 36372 21598
rect 36316 21534 36318 21586
rect 36370 21534 36372 21586
rect 35980 20916 36036 20926
rect 35868 20860 35980 20916
rect 35980 20822 36036 20860
rect 35420 20804 35476 20814
rect 35420 20710 35476 20748
rect 35756 20802 35812 20814
rect 35756 20750 35758 20802
rect 35810 20750 35812 20802
rect 35644 20132 35700 20142
rect 35644 20020 35700 20076
rect 35532 20018 35700 20020
rect 35532 19966 35646 20018
rect 35698 19966 35700 20018
rect 35532 19964 35700 19966
rect 35196 19906 35252 19918
rect 35196 19854 35198 19906
rect 35250 19854 35252 19906
rect 35196 19796 35252 19854
rect 35196 19730 35252 19740
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 35084 18386 35140 18396
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 35532 17892 35588 19964
rect 35644 19954 35700 19964
rect 35756 19796 35812 20750
rect 36316 20132 36372 21534
rect 36988 20916 37044 20926
rect 36988 20822 37044 20860
rect 37212 20802 37268 20814
rect 37212 20750 37214 20802
rect 37266 20750 37268 20802
rect 36540 20580 36596 20590
rect 36540 20486 36596 20524
rect 36316 20066 36372 20076
rect 36316 19908 36372 19918
rect 35756 19730 35812 19740
rect 36092 19906 36372 19908
rect 36092 19854 36318 19906
rect 36370 19854 36372 19906
rect 36092 19852 36372 19854
rect 36092 19122 36148 19852
rect 36316 19842 36372 19852
rect 37212 19908 37268 20750
rect 37324 20804 37380 22988
rect 37436 22148 37492 23884
rect 37884 23828 37940 27468
rect 38220 27188 38276 27198
rect 38108 26852 38164 26862
rect 38108 25508 38164 26796
rect 38108 25414 38164 25452
rect 38220 26850 38276 27132
rect 39004 26908 39060 28476
rect 39228 27972 39284 27982
rect 39228 27878 39284 27916
rect 39228 27076 39284 27086
rect 39228 26982 39284 27020
rect 38220 26798 38222 26850
rect 38274 26798 38276 26850
rect 37660 23772 37940 23828
rect 38108 24612 38164 24622
rect 38220 24612 38276 26798
rect 38444 26852 38500 26862
rect 38444 26514 38500 26796
rect 38444 26462 38446 26514
rect 38498 26462 38500 26514
rect 38444 26450 38500 26462
rect 38892 26852 39060 26908
rect 38780 26404 38836 26414
rect 38780 25394 38836 26348
rect 38780 25342 38782 25394
rect 38834 25342 38836 25394
rect 38780 25330 38836 25342
rect 38892 25396 38948 26852
rect 39004 26292 39060 26302
rect 39452 26292 39508 28700
rect 39564 28420 39620 28700
rect 39676 28754 39732 28924
rect 39676 28702 39678 28754
rect 39730 28702 39732 28754
rect 39676 28690 39732 28702
rect 39564 28354 39620 28364
rect 39676 27972 39732 27982
rect 39676 27878 39732 27916
rect 39564 27858 39620 27870
rect 39564 27806 39566 27858
rect 39618 27806 39620 27858
rect 39564 26908 39620 27806
rect 39900 27858 39956 27870
rect 39900 27806 39902 27858
rect 39954 27806 39956 27858
rect 39900 27188 39956 27806
rect 40012 27188 40068 27198
rect 39900 27186 40068 27188
rect 39900 27134 40014 27186
rect 40066 27134 40068 27186
rect 39900 27132 40068 27134
rect 40012 27122 40068 27132
rect 39564 26852 39844 26908
rect 39564 26292 39620 26302
rect 39452 26290 39620 26292
rect 39452 26238 39566 26290
rect 39618 26238 39620 26290
rect 39452 26236 39620 26238
rect 39004 26068 39060 26236
rect 39564 26226 39620 26236
rect 39788 26178 39844 26852
rect 40124 26402 40180 26414
rect 40124 26350 40126 26402
rect 40178 26350 40180 26402
rect 39900 26292 39956 26302
rect 39900 26290 40068 26292
rect 39900 26238 39902 26290
rect 39954 26238 40068 26290
rect 39900 26236 40068 26238
rect 39900 26226 39956 26236
rect 39788 26126 39790 26178
rect 39842 26126 39844 26178
rect 39788 26114 39844 26126
rect 39004 26002 39060 26012
rect 39004 25508 39060 25518
rect 39060 25452 39508 25508
rect 39004 25414 39060 25452
rect 38892 25330 38948 25340
rect 39452 25394 39508 25452
rect 40012 25506 40068 26236
rect 40124 25732 40180 26350
rect 40124 25666 40180 25676
rect 40236 25508 40292 30046
rect 40460 30100 40516 30716
rect 40460 30034 40516 30044
rect 41132 30324 41188 30334
rect 41132 30098 41188 30268
rect 41468 30210 41524 30940
rect 41468 30158 41470 30210
rect 41522 30158 41524 30210
rect 41468 30146 41524 30158
rect 41916 30324 41972 31164
rect 42588 30324 42644 31500
rect 42812 31220 42868 31230
rect 42812 30994 42868 31164
rect 42812 30942 42814 30994
rect 42866 30942 42868 30994
rect 42812 30930 42868 30942
rect 43036 30996 43092 31500
rect 43148 31554 43204 31566
rect 43148 31502 43150 31554
rect 43202 31502 43204 31554
rect 43148 31220 43204 31502
rect 43148 31154 43204 31164
rect 43372 31108 43428 31118
rect 43260 31052 43372 31108
rect 43148 30996 43204 31006
rect 43036 30994 43204 30996
rect 43036 30942 43150 30994
rect 43202 30942 43204 30994
rect 43036 30940 43204 30942
rect 43148 30930 43204 30940
rect 41916 30210 41972 30268
rect 41916 30158 41918 30210
rect 41970 30158 41972 30210
rect 41916 30146 41972 30158
rect 42140 30322 42644 30324
rect 42140 30270 42590 30322
rect 42642 30270 42644 30322
rect 42140 30268 42644 30270
rect 42140 30210 42196 30268
rect 42588 30258 42644 30268
rect 42140 30158 42142 30210
rect 42194 30158 42196 30210
rect 42140 30146 42196 30158
rect 41132 30046 41134 30098
rect 41186 30046 41188 30098
rect 41132 30034 41188 30046
rect 41244 30100 41300 30110
rect 41244 30006 41300 30044
rect 42476 30100 42532 30110
rect 43036 30100 43092 30110
rect 42476 30006 42532 30044
rect 42924 30098 43092 30100
rect 42924 30046 43038 30098
rect 43090 30046 43092 30098
rect 42924 30044 43092 30046
rect 40908 29988 40964 29998
rect 40908 29894 40964 29932
rect 41692 29986 41748 29998
rect 41692 29934 41694 29986
rect 41746 29934 41748 29986
rect 40908 29428 40964 29438
rect 40908 29334 40964 29372
rect 41692 29426 41748 29934
rect 41692 29374 41694 29426
rect 41746 29374 41748 29426
rect 41692 29362 41748 29374
rect 42924 29428 42980 30044
rect 43036 30034 43092 30044
rect 43260 30098 43316 31052
rect 43372 31042 43428 31052
rect 43372 30324 43428 30334
rect 43372 30230 43428 30268
rect 43260 30046 43262 30098
rect 43314 30046 43316 30098
rect 42924 29314 42980 29372
rect 43036 29428 43092 29438
rect 43260 29428 43316 30046
rect 43036 29426 43316 29428
rect 43036 29374 43038 29426
rect 43090 29374 43316 29426
rect 43036 29372 43316 29374
rect 43036 29362 43092 29372
rect 42924 29262 42926 29314
rect 42978 29262 42980 29314
rect 42924 29250 42980 29262
rect 43596 28756 43652 32620
rect 45388 32564 45444 32574
rect 45388 32470 45444 32508
rect 45836 32562 45892 32732
rect 46284 32722 46340 32732
rect 45836 32510 45838 32562
rect 45890 32510 45892 32562
rect 45836 32498 45892 32510
rect 46396 32562 46452 32574
rect 46396 32510 46398 32562
rect 46450 32510 46452 32562
rect 43708 32450 43764 32462
rect 43708 32398 43710 32450
rect 43762 32398 43764 32450
rect 43708 31892 43764 32398
rect 44380 32452 44436 32462
rect 44380 32450 44660 32452
rect 44380 32398 44382 32450
rect 44434 32398 44660 32450
rect 44380 32396 44660 32398
rect 44380 32386 44436 32396
rect 43708 31778 43764 31836
rect 43708 31726 43710 31778
rect 43762 31726 43764 31778
rect 43708 31714 43764 31726
rect 44156 31556 44212 31566
rect 43820 31108 43876 31118
rect 43820 31106 44100 31108
rect 43820 31054 43822 31106
rect 43874 31054 44100 31106
rect 43820 31052 44100 31054
rect 43820 31042 43876 31052
rect 44044 30436 44100 31052
rect 43820 30324 43876 30334
rect 43876 30268 43988 30324
rect 43820 30230 43876 30268
rect 43708 30212 43764 30222
rect 43708 30118 43764 30156
rect 43820 29876 43876 29886
rect 43820 29650 43876 29820
rect 43820 29598 43822 29650
rect 43874 29598 43876 29650
rect 43820 29586 43876 29598
rect 43932 29650 43988 30268
rect 43932 29598 43934 29650
rect 43986 29598 43988 29650
rect 43932 29586 43988 29598
rect 43708 29428 43764 29438
rect 44044 29428 44100 30380
rect 43708 29426 44100 29428
rect 43708 29374 43710 29426
rect 43762 29374 44100 29426
rect 43708 29372 44100 29374
rect 44156 29428 44212 31500
rect 44604 31108 44660 32396
rect 45500 31948 46228 32004
rect 44940 31780 44996 31790
rect 44940 31666 44996 31724
rect 45500 31778 45556 31948
rect 45500 31726 45502 31778
rect 45554 31726 45556 31778
rect 45500 31714 45556 31726
rect 45836 31780 45892 31790
rect 44940 31614 44942 31666
rect 44994 31614 44996 31666
rect 44940 31602 44996 31614
rect 45164 31668 45220 31678
rect 45164 31574 45220 31612
rect 44604 31014 44660 31052
rect 44828 31554 44884 31566
rect 44828 31502 44830 31554
rect 44882 31502 44884 31554
rect 44828 30434 44884 31502
rect 44828 30382 44830 30434
rect 44882 30382 44884 30434
rect 44828 30370 44884 30382
rect 45276 31556 45332 31566
rect 45276 30994 45332 31500
rect 45724 31332 45780 31342
rect 45276 30942 45278 30994
rect 45330 30942 45332 30994
rect 44940 30324 44996 30334
rect 43708 29362 43764 29372
rect 43036 28754 43652 28756
rect 43036 28702 43598 28754
rect 43650 28702 43652 28754
rect 43036 28700 43652 28702
rect 41020 28420 41076 28430
rect 41020 28082 41076 28364
rect 41020 28030 41022 28082
rect 41074 28030 41076 28082
rect 41020 28018 41076 28030
rect 42140 28420 42196 28430
rect 40796 27972 40852 27982
rect 40796 27878 40852 27916
rect 41132 27858 41188 27870
rect 41132 27806 41134 27858
rect 41186 27806 41188 27858
rect 41132 27748 41188 27806
rect 41580 27748 41636 27758
rect 41132 27746 41636 27748
rect 41132 27694 41582 27746
rect 41634 27694 41636 27746
rect 41132 27692 41636 27694
rect 40012 25454 40014 25506
rect 40066 25454 40068 25506
rect 40012 25442 40068 25454
rect 40124 25452 40292 25508
rect 40348 26516 40404 26526
rect 40348 25620 40404 26460
rect 41132 26404 41188 27692
rect 41580 27682 41636 27692
rect 42140 27186 42196 28364
rect 43036 28082 43092 28700
rect 43596 28690 43652 28700
rect 43708 28756 43764 28766
rect 43036 28030 43038 28082
rect 43090 28030 43092 28082
rect 43036 28018 43092 28030
rect 43260 28084 43316 28094
rect 43260 27990 43316 28028
rect 42700 27860 42756 27870
rect 42924 27860 42980 27870
rect 42700 27858 42924 27860
rect 42700 27806 42702 27858
rect 42754 27806 42924 27858
rect 42700 27804 42924 27806
rect 42700 27794 42756 27804
rect 42924 27766 42980 27804
rect 42140 27134 42142 27186
rect 42194 27134 42196 27186
rect 42140 27122 42196 27134
rect 43372 27634 43428 27646
rect 43372 27582 43374 27634
rect 43426 27582 43428 27634
rect 41132 26338 41188 26348
rect 42588 26962 42644 26974
rect 42588 26910 42590 26962
rect 42642 26910 42644 26962
rect 41020 26292 41076 26302
rect 40796 25620 40852 25630
rect 40348 25618 40852 25620
rect 40348 25566 40798 25618
rect 40850 25566 40852 25618
rect 40348 25564 40852 25566
rect 40348 25506 40404 25564
rect 40796 25554 40852 25564
rect 40348 25454 40350 25506
rect 40402 25454 40404 25506
rect 39788 25396 39844 25406
rect 39452 25342 39454 25394
rect 39506 25342 39508 25394
rect 39452 25330 39508 25342
rect 39676 25340 39788 25396
rect 38892 24948 38948 24958
rect 38892 24854 38948 24892
rect 39228 24836 39284 24846
rect 38108 24610 38276 24612
rect 38108 24558 38110 24610
rect 38162 24558 38276 24610
rect 38108 24556 38276 24558
rect 39116 24780 39228 24836
rect 37548 23716 37604 23726
rect 37548 22594 37604 23660
rect 37660 23380 37716 23772
rect 38108 23604 38164 24556
rect 38556 23940 38612 23950
rect 38556 23846 38612 23884
rect 38108 23548 38724 23604
rect 38668 23492 38724 23548
rect 38668 23436 38836 23492
rect 37660 23286 37716 23324
rect 38332 23380 38388 23390
rect 37548 22542 37550 22594
rect 37602 22542 37604 22594
rect 37548 22530 37604 22542
rect 37884 23154 37940 23166
rect 37884 23102 37886 23154
rect 37938 23102 37940 23154
rect 37884 23044 37940 23102
rect 37884 22596 37940 22988
rect 38108 23156 38164 23166
rect 38108 22930 38164 23100
rect 38332 23154 38388 23324
rect 38556 23380 38612 23390
rect 38556 23286 38612 23324
rect 38332 23102 38334 23154
rect 38386 23102 38388 23154
rect 38332 23090 38388 23102
rect 38668 23154 38724 23166
rect 38668 23102 38670 23154
rect 38722 23102 38724 23154
rect 38108 22878 38110 22930
rect 38162 22878 38164 22930
rect 38108 22866 38164 22878
rect 37884 22530 37940 22540
rect 38332 22594 38388 22606
rect 38332 22542 38334 22594
rect 38386 22542 38388 22594
rect 38108 22484 38164 22494
rect 38332 22484 38388 22542
rect 38164 22428 38388 22484
rect 38668 22484 38724 23102
rect 38108 22418 38164 22428
rect 38668 22418 38724 22428
rect 38780 23156 38836 23436
rect 37660 22372 37716 22382
rect 37548 22148 37604 22158
rect 37436 22092 37548 22148
rect 37548 22082 37604 22092
rect 37548 21028 37604 21038
rect 37660 21028 37716 22316
rect 37772 22372 37828 22382
rect 37772 22370 38052 22372
rect 37772 22318 37774 22370
rect 37826 22318 38052 22370
rect 37772 22316 38052 22318
rect 37772 22306 37828 22316
rect 37996 21476 38052 22316
rect 38220 22258 38276 22270
rect 38220 22206 38222 22258
rect 38274 22206 38276 22258
rect 38220 22148 38276 22206
rect 38220 22082 38276 22092
rect 38332 22148 38388 22158
rect 38332 22146 38724 22148
rect 38332 22094 38334 22146
rect 38386 22094 38724 22146
rect 38332 22092 38724 22094
rect 38332 22082 38388 22092
rect 38668 21700 38724 22092
rect 38668 21634 38724 21644
rect 37996 21420 38388 21476
rect 37548 21026 37716 21028
rect 37548 20974 37550 21026
rect 37602 20974 37716 21026
rect 37548 20972 37716 20974
rect 37548 20962 37604 20972
rect 38332 20914 38388 21420
rect 38332 20862 38334 20914
rect 38386 20862 38388 20914
rect 38332 20850 38388 20862
rect 37884 20804 37940 20814
rect 37324 20802 37940 20804
rect 37324 20750 37886 20802
rect 37938 20750 37940 20802
rect 37324 20748 37940 20750
rect 37884 20738 37940 20748
rect 38220 20804 38276 20814
rect 38108 20690 38164 20702
rect 38108 20638 38110 20690
rect 38162 20638 38164 20690
rect 37212 19842 37268 19852
rect 37996 20580 38052 20590
rect 36988 19684 37044 19694
rect 36092 19070 36094 19122
rect 36146 19070 36148 19122
rect 36092 19058 36148 19070
rect 36428 19124 36484 19134
rect 36428 19030 36484 19068
rect 35308 17836 35588 17892
rect 35756 18340 35812 18350
rect 35308 17780 35364 17836
rect 34860 17778 35364 17780
rect 34860 17726 35310 17778
rect 35362 17726 35364 17778
rect 34860 17724 35364 17726
rect 34860 17666 34916 17724
rect 35308 17714 35364 17724
rect 35756 17780 35812 18284
rect 36316 17780 36372 17790
rect 35756 17778 36316 17780
rect 35756 17726 35758 17778
rect 35810 17726 36316 17778
rect 35756 17724 36316 17726
rect 35756 17714 35812 17724
rect 34860 17614 34862 17666
rect 34914 17614 34916 17666
rect 34860 17602 34916 17614
rect 36316 17666 36372 17724
rect 36988 17668 37044 19628
rect 37996 19460 38052 20524
rect 38108 19684 38164 20638
rect 38108 19618 38164 19628
rect 37996 19404 38164 19460
rect 37436 19234 37492 19246
rect 37436 19182 37438 19234
rect 37490 19182 37492 19234
rect 37100 19124 37156 19134
rect 37100 19030 37156 19068
rect 37212 18452 37268 18462
rect 36316 17614 36318 17666
rect 36370 17614 36372 17666
rect 36316 17602 36372 17614
rect 36876 17612 37044 17668
rect 37100 17668 37156 17678
rect 34748 16772 34804 17052
rect 35196 17556 35252 17566
rect 34748 16706 34804 16716
rect 35084 16994 35140 17006
rect 35084 16942 35086 16994
rect 35138 16942 35140 16994
rect 34188 16212 34244 16222
rect 34524 16212 34580 16222
rect 34188 16210 34580 16212
rect 34188 16158 34190 16210
rect 34242 16158 34526 16210
rect 34578 16158 34580 16210
rect 34188 16156 34580 16158
rect 35084 16212 35140 16942
rect 35196 16882 35252 17500
rect 36092 17442 36148 17454
rect 36092 17390 36094 17442
rect 36146 17390 36148 17442
rect 35756 16996 35812 17006
rect 35644 16884 35700 16894
rect 35196 16830 35198 16882
rect 35250 16830 35252 16882
rect 35196 16818 35252 16830
rect 35532 16828 35644 16884
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 35532 16324 35588 16828
rect 35644 16818 35700 16828
rect 35756 16772 35812 16940
rect 35756 16706 35812 16716
rect 35308 16268 35588 16324
rect 35196 16212 35252 16222
rect 35084 16210 35252 16212
rect 35084 16158 35198 16210
rect 35250 16158 35252 16210
rect 35084 16156 35252 16158
rect 34188 16146 34244 16156
rect 34524 16146 34580 16156
rect 35196 16146 35252 16156
rect 34748 16100 34804 16110
rect 34636 16098 34804 16100
rect 34636 16046 34750 16098
rect 34802 16046 34804 16098
rect 34636 16044 34804 16046
rect 33852 15986 33908 15998
rect 33852 15934 33854 15986
rect 33906 15934 33908 15986
rect 33628 15092 33796 15148
rect 33516 14590 33518 14642
rect 33570 14590 33572 14642
rect 33180 14438 33236 14476
rect 32172 14420 32228 14430
rect 32172 14326 32228 14364
rect 32284 14418 32340 14430
rect 32284 14366 32286 14418
rect 32338 14366 32340 14418
rect 32284 14308 32340 14366
rect 32284 13748 32340 14252
rect 32284 13682 32340 13692
rect 33068 13074 33124 13086
rect 33068 13022 33070 13074
rect 33122 13022 33124 13074
rect 31948 12740 32004 12750
rect 31948 12402 32004 12684
rect 31948 12350 31950 12402
rect 32002 12350 32004 12402
rect 31948 12338 32004 12350
rect 33068 12402 33124 13022
rect 33516 13076 33572 14590
rect 33516 13010 33572 13020
rect 33068 12350 33070 12402
rect 33122 12350 33124 12402
rect 33068 12338 33124 12350
rect 33516 12850 33572 12862
rect 33516 12798 33518 12850
rect 33570 12798 33572 12850
rect 33292 12290 33348 12302
rect 33292 12238 33294 12290
rect 33346 12238 33348 12290
rect 33068 11956 33124 11966
rect 32508 11396 32564 11406
rect 32508 10722 32564 11340
rect 33068 10948 33124 11900
rect 33292 11844 33348 12238
rect 33404 12178 33460 12190
rect 33404 12126 33406 12178
rect 33458 12126 33460 12178
rect 33404 12068 33460 12126
rect 33404 12002 33460 12012
rect 33292 11778 33348 11788
rect 33180 11508 33236 11518
rect 33180 11414 33236 11452
rect 33292 11396 33348 11406
rect 33516 11396 33572 12798
rect 33292 11394 33572 11396
rect 33292 11342 33294 11394
rect 33346 11342 33572 11394
rect 33292 11340 33572 11342
rect 33628 11508 33684 11518
rect 33292 11330 33348 11340
rect 33404 11284 33460 11340
rect 33404 11218 33460 11228
rect 33628 11282 33684 11452
rect 33628 11230 33630 11282
rect 33682 11230 33684 11282
rect 33516 11170 33572 11182
rect 33516 11118 33518 11170
rect 33570 11118 33572 11170
rect 33516 10948 33572 11118
rect 33068 10892 33572 10948
rect 33628 10836 33684 11230
rect 33628 10770 33684 10780
rect 32508 10670 32510 10722
rect 32562 10670 32564 10722
rect 32508 10658 32564 10670
rect 31836 9986 31892 9996
rect 32060 10610 32116 10622
rect 32060 10558 32062 10610
rect 32114 10558 32116 10610
rect 31836 9828 31892 9838
rect 31724 9716 31780 9726
rect 31388 9714 31780 9716
rect 31388 9662 31726 9714
rect 31778 9662 31780 9714
rect 31388 9660 31780 9662
rect 31724 9492 31780 9660
rect 31836 9714 31892 9772
rect 32060 9826 32116 10558
rect 32060 9774 32062 9826
rect 32114 9774 32116 9826
rect 32060 9762 32116 9774
rect 32284 10612 32340 10622
rect 31836 9662 31838 9714
rect 31890 9662 31892 9714
rect 31836 9650 31892 9662
rect 31724 9436 31892 9492
rect 31388 9156 31444 9166
rect 31388 9042 31444 9100
rect 31388 8990 31390 9042
rect 31442 8990 31444 9042
rect 31388 8978 31444 8990
rect 31612 9042 31668 9054
rect 31612 8990 31614 9042
rect 31666 8990 31668 9042
rect 31612 8932 31668 8990
rect 31612 8866 31668 8876
rect 31836 8484 31892 9436
rect 31836 8418 31892 8428
rect 31948 9156 32004 9166
rect 31948 8370 32004 9100
rect 32284 9154 32340 10556
rect 33628 10612 33684 10622
rect 33628 10518 33684 10556
rect 32284 9102 32286 9154
rect 32338 9102 32340 9154
rect 32284 9090 32340 9102
rect 33516 8484 33572 8494
rect 33404 8428 33516 8484
rect 31948 8318 31950 8370
rect 32002 8318 32004 8370
rect 31948 8306 32004 8318
rect 33292 8372 33348 8382
rect 31836 8258 31892 8270
rect 31836 8206 31838 8258
rect 31890 8206 31892 8258
rect 31612 8146 31668 8158
rect 31612 8094 31614 8146
rect 31666 8094 31668 8146
rect 31612 7812 31668 8094
rect 31388 7756 31668 7812
rect 31836 8148 31892 8206
rect 31388 7698 31444 7756
rect 31388 7646 31390 7698
rect 31442 7646 31444 7698
rect 31388 6692 31444 7646
rect 31724 7586 31780 7598
rect 31724 7534 31726 7586
rect 31778 7534 31780 7586
rect 31724 7364 31780 7534
rect 31724 7298 31780 7308
rect 31388 6626 31444 6636
rect 31836 6578 31892 8092
rect 32508 8258 32564 8270
rect 32508 8206 32510 8258
rect 32562 8206 32564 8258
rect 32284 7588 32340 7598
rect 32060 7476 32116 7486
rect 32060 7474 32228 7476
rect 32060 7422 32062 7474
rect 32114 7422 32228 7474
rect 32060 7420 32228 7422
rect 32060 7410 32116 7420
rect 31836 6526 31838 6578
rect 31890 6526 31892 6578
rect 31836 6514 31892 6526
rect 32172 6690 32228 7420
rect 32172 6638 32174 6690
rect 32226 6638 32228 6690
rect 32172 6580 32228 6638
rect 32172 6514 32228 6524
rect 32284 6578 32340 7532
rect 32508 7364 32564 8206
rect 32508 6690 32564 7308
rect 33068 8258 33124 8270
rect 33068 8206 33070 8258
rect 33122 8206 33124 8258
rect 33068 8036 33124 8206
rect 33292 8146 33348 8316
rect 33292 8094 33294 8146
rect 33346 8094 33348 8146
rect 33292 8082 33348 8094
rect 33068 7140 33124 7980
rect 33068 7074 33124 7084
rect 33180 7362 33236 7374
rect 33180 7310 33182 7362
rect 33234 7310 33236 7362
rect 32508 6638 32510 6690
rect 32562 6638 32564 6690
rect 32508 6626 32564 6638
rect 32284 6526 32286 6578
rect 32338 6526 32340 6578
rect 32284 6514 32340 6526
rect 32732 6578 32788 6590
rect 32732 6526 32734 6578
rect 32786 6526 32788 6578
rect 31500 6466 31556 6478
rect 31500 6414 31502 6466
rect 31554 6414 31556 6466
rect 31500 6132 31556 6414
rect 31500 6066 31556 6076
rect 32284 6244 32340 6254
rect 32172 6020 32228 6030
rect 32060 6018 32228 6020
rect 32060 5966 32174 6018
rect 32226 5966 32228 6018
rect 32060 5964 32228 5966
rect 30940 5702 30996 5740
rect 31164 5740 31332 5796
rect 31500 5908 31556 5918
rect 31836 5908 31892 5918
rect 30156 4958 30158 5010
rect 30210 4958 30212 5010
rect 30156 4946 30212 4958
rect 30604 5236 30660 5246
rect 30604 4338 30660 5180
rect 30940 5124 30996 5134
rect 30940 5030 30996 5068
rect 30604 4286 30606 4338
rect 30658 4286 30660 4338
rect 30604 4274 30660 4286
rect 31164 3554 31220 5740
rect 31388 5684 31444 5694
rect 31276 5628 31388 5684
rect 31276 5010 31332 5628
rect 31388 5618 31444 5628
rect 31276 4958 31278 5010
rect 31330 4958 31332 5010
rect 31276 4946 31332 4958
rect 31388 4564 31444 4574
rect 31388 4470 31444 4508
rect 31164 3502 31166 3554
rect 31218 3502 31220 3554
rect 31164 3490 31220 3502
rect 30268 3444 30324 3454
rect 30268 800 30324 3388
rect 31500 3332 31556 5852
rect 30940 3276 31556 3332
rect 31612 5906 31892 5908
rect 31612 5854 31838 5906
rect 31890 5854 31892 5906
rect 31612 5852 31892 5854
rect 31612 5796 31668 5852
rect 31836 5842 31892 5852
rect 30940 800 30996 3276
rect 31612 800 31668 5740
rect 31948 5796 32004 5806
rect 31724 5348 31780 5358
rect 31724 4562 31780 5292
rect 31724 4510 31726 4562
rect 31778 4510 31780 4562
rect 31724 4498 31780 4510
rect 31948 5122 32004 5740
rect 31948 5070 31950 5122
rect 32002 5070 32004 5122
rect 31948 4340 32004 5070
rect 32060 4564 32116 5964
rect 32172 5954 32228 5964
rect 32284 5796 32340 6188
rect 32172 5740 32340 5796
rect 32172 5010 32228 5740
rect 32732 5348 32788 6526
rect 32844 6466 32900 6478
rect 32844 6414 32846 6466
rect 32898 6414 32900 6466
rect 32844 6132 32900 6414
rect 33068 6468 33124 6478
rect 33068 6374 33124 6412
rect 32844 6066 32900 6076
rect 33068 6018 33124 6030
rect 33068 5966 33070 6018
rect 33122 5966 33124 6018
rect 32956 5460 33012 5470
rect 32732 5282 32788 5292
rect 32844 5404 32956 5460
rect 32620 5124 32676 5134
rect 32620 5030 32676 5068
rect 32844 5122 32900 5404
rect 32956 5394 33012 5404
rect 33068 5124 33124 5966
rect 33180 5908 33236 7310
rect 33404 6914 33460 8428
rect 33516 8418 33572 8428
rect 33628 8260 33684 8270
rect 33628 8036 33684 8204
rect 33628 7970 33684 7980
rect 33628 7364 33684 7374
rect 33740 7364 33796 15092
rect 33852 14420 33908 15934
rect 34076 15874 34132 15886
rect 34076 15822 34078 15874
rect 34130 15822 34132 15874
rect 34076 15540 34132 15822
rect 34524 15540 34580 15550
rect 34636 15540 34692 16044
rect 34748 16034 34804 16044
rect 34972 16098 35028 16110
rect 34972 16046 34974 16098
rect 35026 16046 35028 16098
rect 34076 15474 34132 15484
rect 34188 15538 34692 15540
rect 34188 15486 34526 15538
rect 34578 15486 34692 15538
rect 34188 15484 34692 15486
rect 34972 15652 35028 16046
rect 35196 15988 35252 15998
rect 35308 15988 35364 16268
rect 35420 16100 35476 16110
rect 35420 16006 35476 16044
rect 35196 15986 35364 15988
rect 35196 15934 35198 15986
rect 35250 15934 35364 15986
rect 35196 15932 35364 15934
rect 35196 15922 35252 15932
rect 34188 15314 34244 15484
rect 34524 15474 34580 15484
rect 34188 15262 34190 15314
rect 34242 15262 34244 15314
rect 34188 15250 34244 15262
rect 34972 15316 35028 15596
rect 34972 15250 35028 15260
rect 35084 15540 35140 15550
rect 35084 15314 35140 15484
rect 35084 15262 35086 15314
rect 35138 15262 35140 15314
rect 35084 15250 35140 15262
rect 35980 15426 36036 15438
rect 35980 15374 35982 15426
rect 36034 15374 36036 15426
rect 34412 15092 34468 15102
rect 34860 15092 34916 15102
rect 34412 14642 34468 15036
rect 34412 14590 34414 14642
rect 34466 14590 34468 14642
rect 34412 14578 34468 14590
rect 34524 15090 34916 15092
rect 34524 15038 34862 15090
rect 34914 15038 34916 15090
rect 34524 15036 34916 15038
rect 34524 14420 34580 15036
rect 34860 15026 34916 15036
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35980 14644 36036 15374
rect 36092 15316 36148 17390
rect 36428 17108 36484 17118
rect 36876 17108 36932 17612
rect 36988 17444 37044 17454
rect 37100 17444 37156 17612
rect 37212 17668 37268 18396
rect 37324 18450 37380 18462
rect 37324 18398 37326 18450
rect 37378 18398 37380 18450
rect 37324 17892 37380 18398
rect 37436 18452 37492 19182
rect 37996 19122 38052 19134
rect 37996 19070 37998 19122
rect 38050 19070 38052 19122
rect 37884 18676 37940 18686
rect 37996 18676 38052 19070
rect 37884 18674 38052 18676
rect 37884 18622 37886 18674
rect 37938 18622 38052 18674
rect 37884 18620 38052 18622
rect 37884 18610 37940 18620
rect 38108 18564 38164 19404
rect 37996 18508 38108 18564
rect 37436 18386 37492 18396
rect 37772 18452 37828 18462
rect 37772 18450 37940 18452
rect 37772 18398 37774 18450
rect 37826 18398 37940 18450
rect 37772 18396 37940 18398
rect 37772 18386 37828 18396
rect 37324 17826 37380 17836
rect 37660 17668 37716 17678
rect 37212 17666 37716 17668
rect 37212 17614 37214 17666
rect 37266 17614 37662 17666
rect 37714 17614 37716 17666
rect 37212 17612 37716 17614
rect 37212 17602 37268 17612
rect 37660 17602 37716 17612
rect 37884 17556 37940 18396
rect 37996 18450 38052 18508
rect 38108 18470 38164 18508
rect 38220 19234 38276 20748
rect 38780 20802 38836 23100
rect 39004 23154 39060 23166
rect 39004 23102 39006 23154
rect 39058 23102 39060 23154
rect 39004 23044 39060 23102
rect 39004 22596 39060 22988
rect 39004 22530 39060 22540
rect 38780 20750 38782 20802
rect 38834 20750 38836 20802
rect 38780 20738 38836 20750
rect 38892 22258 38948 22270
rect 38892 22206 38894 22258
rect 38946 22206 38948 22258
rect 38444 20690 38500 20702
rect 38444 20638 38446 20690
rect 38498 20638 38500 20690
rect 38444 20188 38500 20638
rect 38444 20132 38724 20188
rect 38668 20020 38724 20132
rect 38220 19182 38222 19234
rect 38274 19182 38276 19234
rect 37996 18398 37998 18450
rect 38050 18398 38052 18450
rect 37996 18386 38052 18398
rect 37996 17556 38052 17566
rect 37884 17554 38052 17556
rect 37884 17502 37998 17554
rect 38050 17502 38052 17554
rect 37884 17500 38052 17502
rect 36988 17442 37156 17444
rect 36988 17390 36990 17442
rect 37042 17390 37156 17442
rect 36988 17388 37156 17390
rect 36988 17378 37044 17388
rect 36988 17108 37044 17118
rect 36428 17106 37044 17108
rect 36428 17054 36430 17106
rect 36482 17054 36990 17106
rect 37042 17054 37044 17106
rect 36428 17052 37044 17054
rect 36428 17042 36484 17052
rect 36988 17042 37044 17052
rect 36204 16884 36260 16894
rect 36204 16790 36260 16828
rect 36540 16884 36596 16894
rect 36540 16790 36596 16828
rect 37100 16100 37156 17388
rect 37548 17332 37604 17342
rect 37436 16884 37492 16894
rect 37100 16034 37156 16044
rect 37324 16772 37380 16782
rect 36988 15428 37044 15438
rect 36092 15250 36148 15260
rect 36316 15314 36372 15326
rect 36316 15262 36318 15314
rect 36370 15262 36372 15314
rect 33852 14418 34580 14420
rect 33852 14366 33854 14418
rect 33906 14366 34580 14418
rect 33852 14364 34580 14366
rect 35532 14588 36036 14644
rect 35532 14418 35588 14588
rect 35980 14530 36036 14588
rect 35980 14478 35982 14530
rect 36034 14478 36036 14530
rect 35980 14466 36036 14478
rect 36204 14532 36260 14542
rect 36204 14438 36260 14476
rect 35532 14366 35534 14418
rect 35586 14366 35588 14418
rect 33852 14354 33908 14364
rect 35308 14308 35364 14318
rect 35308 14214 35364 14252
rect 35532 13860 35588 14366
rect 35644 14420 35700 14430
rect 35644 14326 35700 14364
rect 36316 14420 36372 15262
rect 36988 15314 37044 15372
rect 36988 15262 36990 15314
rect 37042 15262 37044 15314
rect 36988 15250 37044 15262
rect 37324 15148 37380 16716
rect 37436 16436 37492 16828
rect 37436 16370 37492 16380
rect 37548 15538 37604 17276
rect 37996 17108 38052 17500
rect 38220 17556 38276 19182
rect 38444 19906 38500 19918
rect 38444 19854 38446 19906
rect 38498 19854 38500 19906
rect 38444 18452 38500 19854
rect 38668 19124 38724 19964
rect 38780 20132 38836 20142
rect 38892 20132 38948 22206
rect 39004 22148 39060 22158
rect 39116 22148 39172 24780
rect 39228 24742 39284 24780
rect 39340 24052 39396 24062
rect 39228 23604 39284 23614
rect 39228 22930 39284 23548
rect 39228 22878 39230 22930
rect 39282 22878 39284 22930
rect 39228 22866 39284 22878
rect 39228 22372 39284 22382
rect 39340 22372 39396 23996
rect 39676 23548 39732 25340
rect 39788 25302 39844 25340
rect 40124 24612 40180 25452
rect 40348 25442 40404 25454
rect 40236 25282 40292 25294
rect 40236 25230 40238 25282
rect 40290 25230 40292 25282
rect 40236 24836 40292 25230
rect 40236 24770 40292 24780
rect 40908 24722 40964 24734
rect 40908 24670 40910 24722
rect 40962 24670 40964 24722
rect 39564 23492 39732 23548
rect 39788 24556 40180 24612
rect 40460 24612 40516 24622
rect 40684 24612 40740 24622
rect 40460 24610 40684 24612
rect 40460 24558 40462 24610
rect 40514 24558 40684 24610
rect 40460 24556 40684 24558
rect 39788 23548 39844 24556
rect 40460 24546 40516 24556
rect 40684 24546 40740 24556
rect 40908 24052 40964 24670
rect 40908 23986 40964 23996
rect 40236 23940 40292 23950
rect 40292 23884 40404 23940
rect 40236 23846 40292 23884
rect 39788 23492 39956 23548
rect 39452 23268 39508 23278
rect 39452 23154 39508 23212
rect 39452 23102 39454 23154
rect 39506 23102 39508 23154
rect 39452 23090 39508 23102
rect 39564 22820 39620 23492
rect 39788 23154 39844 23166
rect 39788 23102 39790 23154
rect 39842 23102 39844 23154
rect 39676 23044 39732 23054
rect 39676 22950 39732 22988
rect 39788 22820 39844 23102
rect 39564 22754 39620 22764
rect 39676 22764 39844 22820
rect 39228 22370 39396 22372
rect 39228 22318 39230 22370
rect 39282 22318 39396 22370
rect 39228 22316 39396 22318
rect 39564 22372 39620 22382
rect 39228 22306 39284 22316
rect 39564 22278 39620 22316
rect 39060 22092 39172 22148
rect 39452 22146 39508 22158
rect 39452 22094 39454 22146
rect 39506 22094 39508 22146
rect 39004 22054 39060 22092
rect 39228 21700 39284 21710
rect 39228 21474 39284 21644
rect 39228 21422 39230 21474
rect 39282 21422 39284 21474
rect 39228 21410 39284 21422
rect 39452 20916 39508 22094
rect 39676 21924 39732 22764
rect 39788 22596 39844 22606
rect 39900 22596 39956 23492
rect 40012 22820 40068 22830
rect 40068 22764 40180 22820
rect 40012 22754 40068 22764
rect 39788 22594 39956 22596
rect 39788 22542 39790 22594
rect 39842 22542 39956 22594
rect 39788 22540 39956 22542
rect 40012 22596 40068 22606
rect 39788 22530 39844 22540
rect 39900 22372 39956 22382
rect 39900 21924 39956 22316
rect 39676 21868 39844 21924
rect 39676 21700 39732 21710
rect 39676 21606 39732 21644
rect 39564 20916 39620 20926
rect 39452 20914 39620 20916
rect 39452 20862 39566 20914
rect 39618 20862 39620 20914
rect 39452 20860 39620 20862
rect 39564 20850 39620 20860
rect 39452 20132 39508 20142
rect 38892 20076 39396 20132
rect 38780 19346 38836 20076
rect 38892 19906 38948 19918
rect 38892 19854 38894 19906
rect 38946 19854 38948 19906
rect 38892 19684 38948 19854
rect 38892 19618 38948 19628
rect 38780 19294 38782 19346
rect 38834 19294 38836 19346
rect 38780 19282 38836 19294
rect 38668 19068 38836 19124
rect 38444 18340 38500 18396
rect 38556 18340 38612 18350
rect 38444 18338 38612 18340
rect 38444 18286 38558 18338
rect 38610 18286 38612 18338
rect 38444 18284 38612 18286
rect 38556 17892 38612 18284
rect 38556 17826 38612 17836
rect 38220 17490 38276 17500
rect 38332 17780 38388 17790
rect 38332 17666 38388 17724
rect 38332 17614 38334 17666
rect 38386 17614 38388 17666
rect 38332 17332 38388 17614
rect 38668 17444 38724 17454
rect 38668 17350 38724 17388
rect 37996 17042 38052 17052
rect 38108 17276 38388 17332
rect 38108 17106 38164 17276
rect 38108 17054 38110 17106
rect 38162 17054 38164 17106
rect 38108 17042 38164 17054
rect 38780 16436 38836 19068
rect 39228 18564 39284 18574
rect 39004 18338 39060 18350
rect 39004 18286 39006 18338
rect 39058 18286 39060 18338
rect 39004 18228 39060 18286
rect 39004 18162 39060 18172
rect 39228 17778 39284 18508
rect 39228 17726 39230 17778
rect 39282 17726 39284 17778
rect 39228 17714 39284 17726
rect 39340 17668 39396 20076
rect 39452 19348 39508 20076
rect 39452 19234 39508 19292
rect 39452 19182 39454 19234
rect 39506 19182 39508 19234
rect 39452 19170 39508 19182
rect 39788 18116 39844 21868
rect 39900 21858 39956 21868
rect 40012 21810 40068 22540
rect 40012 21758 40014 21810
rect 40066 21758 40068 21810
rect 40012 21746 40068 21758
rect 40124 21588 40180 22764
rect 40348 22484 40404 23884
rect 41020 23828 41076 26236
rect 42588 26292 42644 26910
rect 42588 26226 42644 26236
rect 43036 26850 43092 26862
rect 43036 26798 43038 26850
rect 43090 26798 43092 26850
rect 41692 26180 41748 26190
rect 41692 26178 42084 26180
rect 41692 26126 41694 26178
rect 41746 26126 42084 26178
rect 41692 26124 42084 26126
rect 41692 26114 41748 26124
rect 41356 25844 41412 25854
rect 41132 25732 41188 25742
rect 41132 25282 41188 25676
rect 41356 25506 41412 25788
rect 42028 25730 42084 26124
rect 42700 26068 42756 26078
rect 43036 26068 43092 26798
rect 42756 26012 43092 26068
rect 43372 26404 43428 27582
rect 43596 27300 43652 27310
rect 43708 27300 43764 28700
rect 44156 28754 44212 29372
rect 44268 30210 44324 30222
rect 44268 30158 44270 30210
rect 44322 30158 44324 30210
rect 44268 29988 44324 30158
rect 44268 29426 44324 29932
rect 44268 29374 44270 29426
rect 44322 29374 44324 29426
rect 44268 29362 44324 29374
rect 44380 30212 44436 30222
rect 44156 28702 44158 28754
rect 44210 28702 44212 28754
rect 44156 28690 44212 28702
rect 43820 27972 43876 27982
rect 43820 27858 43876 27916
rect 44268 27972 44324 27982
rect 44380 27972 44436 30156
rect 44940 30210 44996 30268
rect 44940 30158 44942 30210
rect 44994 30158 44996 30210
rect 44940 30146 44996 30158
rect 45276 30212 45332 30942
rect 45612 31276 45724 31332
rect 45388 30436 45444 30446
rect 45388 30342 45444 30380
rect 45612 30436 45668 31276
rect 45724 31266 45780 31276
rect 45836 30994 45892 31724
rect 45948 31668 46004 31678
rect 45948 31108 46004 31612
rect 46060 31554 46116 31566
rect 46060 31502 46062 31554
rect 46114 31502 46116 31554
rect 46060 31332 46116 31502
rect 46060 31266 46116 31276
rect 46172 31556 46228 31948
rect 46396 31780 46452 32510
rect 46508 32564 46564 32574
rect 46508 32470 46564 32508
rect 46396 31714 46452 31724
rect 46284 31666 46340 31678
rect 46284 31614 46286 31666
rect 46338 31614 46340 31666
rect 46284 31556 46340 31614
rect 46620 31556 46676 33852
rect 46732 33842 46788 33852
rect 46732 32788 46788 32798
rect 46732 32694 46788 32732
rect 46172 31500 46676 31556
rect 46732 32116 46788 32126
rect 45948 31052 46116 31108
rect 45836 30942 45838 30994
rect 45890 30942 45892 30994
rect 45836 30930 45892 30942
rect 46060 30994 46116 31052
rect 46172 31106 46228 31500
rect 46172 31054 46174 31106
rect 46226 31054 46228 31106
rect 46172 31042 46228 31054
rect 46060 30942 46062 30994
rect 46114 30942 46116 30994
rect 46060 30930 46116 30942
rect 46620 30772 46676 30782
rect 46396 30770 46676 30772
rect 46396 30718 46622 30770
rect 46674 30718 46676 30770
rect 46396 30716 46676 30718
rect 45612 30434 46340 30436
rect 45612 30382 45614 30434
rect 45666 30382 46340 30434
rect 45612 30380 46340 30382
rect 45612 30370 45668 30380
rect 46284 30212 46340 30380
rect 46396 30434 46452 30716
rect 46620 30706 46676 30716
rect 46396 30382 46398 30434
rect 46450 30382 46452 30434
rect 46396 30370 46452 30382
rect 46620 30212 46676 30222
rect 45276 30156 45444 30212
rect 46284 30210 46676 30212
rect 46284 30158 46622 30210
rect 46674 30158 46676 30210
rect 46284 30156 46676 30158
rect 45164 30100 45220 30110
rect 45164 30098 45332 30100
rect 45164 30046 45166 30098
rect 45218 30046 45332 30098
rect 45164 30044 45332 30046
rect 45164 30034 45220 30044
rect 44716 29652 44772 29662
rect 45276 29652 45332 30044
rect 45388 29876 45444 30156
rect 46620 30146 46676 30156
rect 45388 29810 45444 29820
rect 45500 30100 45556 30110
rect 45388 29652 45444 29662
rect 44716 29650 45444 29652
rect 44716 29598 44718 29650
rect 44770 29598 45390 29650
rect 45442 29598 45444 29650
rect 44716 29596 45444 29598
rect 44716 29586 44772 29596
rect 45388 29586 45444 29596
rect 45500 29538 45556 30044
rect 46060 29988 46116 29998
rect 46060 29894 46116 29932
rect 46284 29988 46340 29998
rect 45948 29876 46004 29886
rect 45500 29486 45502 29538
rect 45554 29486 45556 29538
rect 44940 29428 44996 29438
rect 45500 29428 45556 29486
rect 44940 29426 45556 29428
rect 44940 29374 44942 29426
rect 44994 29374 45556 29426
rect 44940 29372 45556 29374
rect 45612 29652 45668 29662
rect 44940 29362 44996 29372
rect 44604 29202 44660 29214
rect 44604 29150 44606 29202
rect 44658 29150 44660 29202
rect 44604 28868 44660 29150
rect 45388 29204 45444 29214
rect 45388 29110 45444 29148
rect 44604 28802 44660 28812
rect 44940 28756 44996 28766
rect 44940 28662 44996 28700
rect 44268 27970 44436 27972
rect 44268 27918 44270 27970
rect 44322 27918 44436 27970
rect 44268 27916 44436 27918
rect 44716 28084 44772 28094
rect 44716 27970 44772 28028
rect 45052 28084 45108 28094
rect 44716 27918 44718 27970
rect 44770 27918 44772 27970
rect 44268 27906 44324 27916
rect 44716 27906 44772 27918
rect 44828 27972 44884 27982
rect 44828 27878 44884 27916
rect 43820 27806 43822 27858
rect 43874 27806 43876 27858
rect 43820 27794 43876 27806
rect 44044 27858 44100 27870
rect 44044 27806 44046 27858
rect 44098 27806 44100 27858
rect 43932 27636 43988 27646
rect 43596 27298 43764 27300
rect 43596 27246 43598 27298
rect 43650 27246 43764 27298
rect 43596 27244 43764 27246
rect 43820 27524 43876 27534
rect 43820 27298 43876 27468
rect 43820 27246 43822 27298
rect 43874 27246 43876 27298
rect 43596 27234 43652 27244
rect 43820 27234 43876 27246
rect 43932 27298 43988 27580
rect 43932 27246 43934 27298
rect 43986 27246 43988 27298
rect 43932 27234 43988 27246
rect 44044 26908 44100 27806
rect 45052 27858 45108 28028
rect 45052 27806 45054 27858
rect 45106 27806 45108 27858
rect 45052 27794 45108 27806
rect 45500 28084 45556 28094
rect 45612 28084 45668 29596
rect 45948 29650 46004 29820
rect 45948 29598 45950 29650
rect 46002 29598 46004 29650
rect 45948 29586 46004 29598
rect 45500 28082 45668 28084
rect 45500 28030 45502 28082
rect 45554 28030 45668 28082
rect 45500 28028 45668 28030
rect 45948 28532 46004 28542
rect 44380 27748 44436 27758
rect 44380 27654 44436 27692
rect 45500 27748 45556 28028
rect 45500 27682 45556 27692
rect 45612 27636 45668 27646
rect 43932 26852 44100 26908
rect 45052 27524 45108 27534
rect 44716 26852 44772 26862
rect 43932 26850 43988 26852
rect 43932 26798 43934 26850
rect 43986 26798 43988 26850
rect 43932 26786 43988 26798
rect 44380 26850 44772 26852
rect 44380 26798 44718 26850
rect 44770 26798 44772 26850
rect 44380 26796 44772 26798
rect 42028 25678 42030 25730
rect 42082 25678 42084 25730
rect 42028 25666 42084 25678
rect 42588 25956 42644 25966
rect 41468 25620 41524 25630
rect 41468 25618 41972 25620
rect 41468 25566 41470 25618
rect 41522 25566 41972 25618
rect 41468 25564 41972 25566
rect 41468 25554 41524 25564
rect 41356 25454 41358 25506
rect 41410 25454 41412 25506
rect 41356 25442 41412 25454
rect 41916 25506 41972 25564
rect 42364 25508 42420 25518
rect 41916 25454 41918 25506
rect 41970 25454 41972 25506
rect 41916 25442 41972 25454
rect 42028 25506 42420 25508
rect 42028 25454 42366 25506
rect 42418 25454 42420 25506
rect 42028 25452 42420 25454
rect 41132 25230 41134 25282
rect 41186 25230 41188 25282
rect 41132 25172 41188 25230
rect 41580 25394 41636 25406
rect 41580 25342 41582 25394
rect 41634 25342 41636 25394
rect 41356 25172 41412 25182
rect 41132 25116 41356 25172
rect 41356 24946 41412 25116
rect 41356 24894 41358 24946
rect 41410 24894 41412 24946
rect 41356 24882 41412 24894
rect 41580 24946 41636 25342
rect 42028 25394 42084 25452
rect 42364 25442 42420 25452
rect 42028 25342 42030 25394
rect 42082 25342 42084 25394
rect 42028 25330 42084 25342
rect 42588 25394 42644 25900
rect 42700 25506 42756 26012
rect 42700 25454 42702 25506
rect 42754 25454 42756 25506
rect 42700 25442 42756 25454
rect 42588 25342 42590 25394
rect 42642 25342 42644 25394
rect 42588 25330 42644 25342
rect 43036 25396 43092 25406
rect 43036 25302 43092 25340
rect 43372 25394 43428 26348
rect 44156 26404 44212 26414
rect 44156 26290 44212 26348
rect 44156 26238 44158 26290
rect 44210 26238 44212 26290
rect 44156 26226 44212 26238
rect 44380 26402 44436 26796
rect 44716 26786 44772 26796
rect 44380 26350 44382 26402
rect 44434 26350 44436 26402
rect 43820 26178 43876 26190
rect 43820 26126 43822 26178
rect 43874 26126 43876 26178
rect 43820 25956 43876 26126
rect 44380 26068 44436 26350
rect 44940 26628 44996 26638
rect 44940 26514 44996 26572
rect 44940 26462 44942 26514
rect 44994 26462 44996 26514
rect 43820 25890 43876 25900
rect 44156 26012 44436 26068
rect 44492 26290 44548 26302
rect 44492 26238 44494 26290
rect 44546 26238 44548 26290
rect 43372 25342 43374 25394
rect 43426 25342 43428 25394
rect 43372 25330 43428 25342
rect 43932 25396 43988 25406
rect 43988 25340 44100 25396
rect 43932 25330 43988 25340
rect 41580 24894 41582 24946
rect 41634 24894 41636 24946
rect 41580 24882 41636 24894
rect 41804 24834 41860 24846
rect 41804 24782 41806 24834
rect 41858 24782 41860 24834
rect 41132 24724 41188 24734
rect 41132 24630 41188 24668
rect 41468 24498 41524 24510
rect 41468 24446 41470 24498
rect 41522 24446 41524 24498
rect 41468 23940 41524 24446
rect 41468 23874 41524 23884
rect 41244 23828 41300 23838
rect 41804 23828 41860 24782
rect 43932 24836 43988 24846
rect 43932 24742 43988 24780
rect 41020 23826 41300 23828
rect 41020 23774 41246 23826
rect 41298 23774 41300 23826
rect 41020 23772 41300 23774
rect 41244 23156 41300 23772
rect 41244 23062 41300 23100
rect 41580 23772 41860 23828
rect 41916 24722 41972 24734
rect 41916 24670 41918 24722
rect 41970 24670 41972 24722
rect 41916 24612 41972 24670
rect 40908 22484 40964 22494
rect 40348 22428 40740 22484
rect 40236 22372 40292 22382
rect 40236 22278 40292 22316
rect 40348 22260 40404 22270
rect 40572 22260 40628 22270
rect 40348 22258 40628 22260
rect 40348 22206 40350 22258
rect 40402 22206 40574 22258
rect 40626 22206 40628 22258
rect 40348 22204 40628 22206
rect 40348 22194 40404 22204
rect 40572 22194 40628 22204
rect 40348 21812 40404 21822
rect 40236 21588 40292 21598
rect 40124 21586 40292 21588
rect 40124 21534 40238 21586
rect 40290 21534 40292 21586
rect 40124 21532 40292 21534
rect 40236 21522 40292 21532
rect 40236 20132 40292 20142
rect 39900 20020 39956 20030
rect 39900 19926 39956 19964
rect 40236 19346 40292 20076
rect 40236 19294 40238 19346
rect 40290 19294 40292 19346
rect 40236 19282 40292 19294
rect 39788 18050 39844 18060
rect 39452 17668 39508 17678
rect 39340 17666 39508 17668
rect 39340 17614 39454 17666
rect 39506 17614 39508 17666
rect 39340 17612 39508 17614
rect 38780 16370 38836 16380
rect 39116 17442 39172 17454
rect 39116 17390 39118 17442
rect 39170 17390 39172 17442
rect 37548 15486 37550 15538
rect 37602 15486 37604 15538
rect 37548 15474 37604 15486
rect 38556 16324 38612 16334
rect 38556 15540 38612 16268
rect 38556 15446 38612 15484
rect 38780 16100 38836 16110
rect 38780 15986 38836 16044
rect 39116 16098 39172 17390
rect 39340 17444 39396 17454
rect 39340 17350 39396 17388
rect 39452 17332 39508 17612
rect 39788 17668 39844 17678
rect 40124 17668 40180 17678
rect 39844 17666 40180 17668
rect 39844 17614 40126 17666
rect 40178 17614 40180 17666
rect 39844 17612 40180 17614
rect 39788 17574 39844 17612
rect 40124 17602 40180 17612
rect 40348 17666 40404 21756
rect 40684 21588 40740 22428
rect 40908 22370 40964 22428
rect 41244 22484 41300 22494
rect 41300 22428 41412 22484
rect 41244 22418 41300 22428
rect 40908 22318 40910 22370
rect 40962 22318 40964 22370
rect 40908 22306 40964 22318
rect 41244 22260 41300 22270
rect 41244 22166 41300 22204
rect 40796 22146 40852 22158
rect 40796 22094 40798 22146
rect 40850 22094 40852 22146
rect 40796 21812 40852 22094
rect 40796 21756 41076 21812
rect 40908 21588 40964 21598
rect 40460 21586 40964 21588
rect 40460 21534 40910 21586
rect 40962 21534 40964 21586
rect 40460 21532 40964 21534
rect 40460 20242 40516 21532
rect 40908 21522 40964 21532
rect 41020 20916 41076 21756
rect 41132 20916 41188 20926
rect 41020 20860 41132 20916
rect 41132 20850 41188 20860
rect 40460 20190 40462 20242
rect 40514 20190 40516 20242
rect 40460 20178 40516 20190
rect 41356 20468 41412 22428
rect 41468 22260 41524 22270
rect 41580 22260 41636 23772
rect 41468 22258 41636 22260
rect 41468 22206 41470 22258
rect 41522 22206 41636 22258
rect 41468 22204 41636 22206
rect 41804 22260 41860 22270
rect 41468 22148 41524 22204
rect 41804 22166 41860 22204
rect 41468 22082 41524 22092
rect 41692 22146 41748 22158
rect 41692 22094 41694 22146
rect 41746 22094 41748 22146
rect 41692 21364 41748 22094
rect 41692 21298 41748 21308
rect 41692 20916 41748 20926
rect 41692 20822 41748 20860
rect 40908 20132 40964 20142
rect 40908 20038 40964 20076
rect 41244 20018 41300 20030
rect 41244 19966 41246 20018
rect 41298 19966 41300 20018
rect 41132 18564 41188 18574
rect 41132 18470 41188 18508
rect 41244 18452 41300 19966
rect 41244 18386 41300 18396
rect 41356 18450 41412 20412
rect 41356 18398 41358 18450
rect 41410 18398 41412 18450
rect 41356 18386 41412 18398
rect 41804 18340 41860 18350
rect 41804 18226 41860 18284
rect 41804 18174 41806 18226
rect 41858 18174 41860 18226
rect 40348 17614 40350 17666
rect 40402 17614 40404 17666
rect 39452 17266 39508 17276
rect 40348 17220 40404 17614
rect 41020 18116 41076 18126
rect 40572 17554 40628 17566
rect 40572 17502 40574 17554
rect 40626 17502 40628 17554
rect 40460 17444 40516 17454
rect 40572 17444 40628 17502
rect 40516 17388 40628 17444
rect 40684 17444 40740 17454
rect 40460 17378 40516 17388
rect 40684 17350 40740 17388
rect 40796 17442 40852 17454
rect 40796 17390 40798 17442
rect 40850 17390 40852 17442
rect 40460 17220 40516 17230
rect 40348 17164 40460 17220
rect 40460 17154 40516 17164
rect 39676 17108 39732 17118
rect 39116 16046 39118 16098
rect 39170 16046 39172 16098
rect 39116 16034 39172 16046
rect 39340 17106 39732 17108
rect 39340 17054 39678 17106
rect 39730 17054 39732 17106
rect 39340 17052 39732 17054
rect 39340 16100 39396 17052
rect 39676 17042 39732 17052
rect 40796 16996 40852 17390
rect 40684 16940 40852 16996
rect 39340 16034 39396 16044
rect 39452 16882 39508 16894
rect 39452 16830 39454 16882
rect 39506 16830 39508 16882
rect 39452 16098 39508 16830
rect 39900 16882 39956 16894
rect 39900 16830 39902 16882
rect 39954 16830 39956 16882
rect 39788 16772 39844 16782
rect 39788 16678 39844 16716
rect 39900 16436 39956 16830
rect 39452 16046 39454 16098
rect 39506 16046 39508 16098
rect 39004 15988 39060 15998
rect 38780 15934 38782 15986
rect 38834 15934 38836 15986
rect 37772 15428 37828 15438
rect 37324 15092 37492 15148
rect 35644 13860 35700 13870
rect 35532 13858 35700 13860
rect 35532 13806 35646 13858
rect 35698 13806 35700 13858
rect 35532 13804 35700 13806
rect 35644 13794 35700 13804
rect 35084 13746 35140 13758
rect 35084 13694 35086 13746
rect 35138 13694 35140 13746
rect 34748 13634 34804 13646
rect 34748 13582 34750 13634
rect 34802 13582 34804 13634
rect 34636 12962 34692 12974
rect 34636 12910 34638 12962
rect 34690 12910 34692 12962
rect 33852 12178 33908 12190
rect 33852 12126 33854 12178
rect 33906 12126 33908 12178
rect 33852 11844 33908 12126
rect 33852 11778 33908 11788
rect 33964 12178 34020 12190
rect 33964 12126 33966 12178
rect 34018 12126 34020 12178
rect 33964 12068 34020 12126
rect 34076 12180 34132 12190
rect 34636 12180 34692 12910
rect 34076 12178 34692 12180
rect 34076 12126 34078 12178
rect 34130 12126 34692 12178
rect 34076 12124 34692 12126
rect 34748 12738 34804 13582
rect 34748 12686 34750 12738
rect 34802 12686 34804 12738
rect 34748 12180 34804 12686
rect 35084 12292 35140 13694
rect 36316 13524 36372 14364
rect 36876 14530 36932 14542
rect 36876 14478 36878 14530
rect 36930 14478 36932 14530
rect 36876 14308 36932 14478
rect 36876 14242 36932 14252
rect 36316 13458 36372 13468
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 37100 13076 37156 13086
rect 35980 12404 36036 12442
rect 35980 12338 36036 12348
rect 35084 12198 35140 12236
rect 34972 12180 35028 12190
rect 34748 12178 35028 12180
rect 34748 12126 34974 12178
rect 35026 12126 35028 12178
rect 34748 12124 35028 12126
rect 34076 12114 34132 12124
rect 33964 11394 34020 12012
rect 34524 11954 34580 11966
rect 34524 11902 34526 11954
rect 34578 11902 34580 11954
rect 33964 11342 33966 11394
rect 34018 11342 34020 11394
rect 33964 11172 34020 11342
rect 33964 11106 34020 11116
rect 34188 11844 34244 11854
rect 34188 11282 34244 11788
rect 34524 11620 34580 11902
rect 34636 11732 34692 12124
rect 34972 12114 35028 12124
rect 35980 12178 36036 12190
rect 35980 12126 35982 12178
rect 36034 12126 36036 12178
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 34636 11676 35140 11732
rect 35196 11722 35460 11732
rect 34524 11554 34580 11564
rect 34188 11230 34190 11282
rect 34242 11230 34244 11282
rect 33964 10836 34020 10846
rect 33964 10722 34020 10780
rect 34188 10834 34244 11230
rect 34972 11508 35028 11518
rect 34972 11170 35028 11452
rect 34972 11118 34974 11170
rect 35026 11118 35028 11170
rect 34972 11106 35028 11118
rect 35084 11394 35140 11676
rect 35084 11342 35086 11394
rect 35138 11342 35140 11394
rect 34188 10782 34190 10834
rect 34242 10782 34244 10834
rect 34188 10770 34244 10782
rect 34860 10836 34916 10846
rect 33964 10670 33966 10722
rect 34018 10670 34020 10722
rect 33964 9604 34020 10670
rect 34524 10724 34580 10734
rect 34524 10630 34580 10668
rect 34748 9716 34804 9726
rect 34636 9714 34804 9716
rect 34636 9662 34750 9714
rect 34802 9662 34804 9714
rect 34636 9660 34804 9662
rect 33964 9538 34020 9548
rect 34412 9604 34468 9614
rect 34468 9548 34580 9604
rect 34412 9510 34468 9548
rect 34188 8932 34244 8942
rect 33852 8930 34244 8932
rect 33852 8878 34190 8930
rect 34242 8878 34244 8930
rect 33852 8876 34244 8878
rect 33852 8372 33908 8876
rect 34188 8866 34244 8876
rect 34412 8818 34468 8830
rect 34412 8766 34414 8818
rect 34466 8766 34468 8818
rect 33852 7698 33908 8316
rect 33852 7646 33854 7698
rect 33906 7646 33908 7698
rect 33852 7634 33908 7646
rect 33964 8596 34020 8606
rect 33740 7308 33908 7364
rect 33628 7270 33684 7308
rect 33404 6862 33406 6914
rect 33458 6862 33460 6914
rect 33404 6850 33460 6862
rect 33740 7140 33796 7150
rect 33292 6578 33348 6590
rect 33292 6526 33294 6578
rect 33346 6526 33348 6578
rect 33292 6244 33348 6526
rect 33292 6178 33348 6188
rect 33404 6466 33460 6478
rect 33404 6414 33406 6466
rect 33458 6414 33460 6466
rect 33292 5908 33348 5918
rect 33180 5906 33348 5908
rect 33180 5854 33294 5906
rect 33346 5854 33348 5906
rect 33180 5852 33348 5854
rect 32844 5070 32846 5122
rect 32898 5070 32900 5122
rect 32844 5058 32900 5070
rect 32956 5068 33124 5124
rect 33180 5572 33236 5582
rect 33180 5122 33236 5516
rect 33180 5070 33182 5122
rect 33234 5070 33236 5122
rect 32172 4958 32174 5010
rect 32226 4958 32228 5010
rect 32172 4946 32228 4958
rect 32732 5012 32788 5022
rect 32732 4788 32788 4956
rect 32060 4470 32116 4508
rect 32396 4732 32788 4788
rect 32396 4562 32452 4732
rect 32396 4510 32398 4562
rect 32450 4510 32452 4562
rect 32396 4498 32452 4510
rect 31948 4284 32228 4340
rect 32172 3442 32228 4284
rect 32508 3556 32564 3566
rect 32956 3556 33012 5068
rect 33068 4900 33124 4910
rect 33068 4562 33124 4844
rect 33180 4676 33236 5070
rect 33180 4610 33236 4620
rect 33068 4510 33070 4562
rect 33122 4510 33124 4562
rect 33068 4498 33124 4510
rect 33292 4228 33348 5852
rect 33404 5684 33460 6414
rect 33740 6130 33796 7084
rect 33740 6078 33742 6130
rect 33794 6078 33796 6130
rect 33740 6066 33796 6078
rect 33740 5908 33796 5918
rect 33404 5618 33460 5628
rect 33628 5684 33684 5694
rect 33516 5460 33572 5470
rect 33404 5404 33516 5460
rect 33404 4676 33460 5404
rect 33516 5394 33572 5404
rect 33516 5236 33572 5246
rect 33516 5142 33572 5180
rect 33628 4900 33684 5628
rect 33740 5122 33796 5852
rect 33740 5070 33742 5122
rect 33794 5070 33796 5122
rect 33740 5058 33796 5070
rect 33628 4834 33684 4844
rect 33404 4620 33796 4676
rect 33404 4562 33460 4620
rect 33404 4510 33406 4562
rect 33458 4510 33460 4562
rect 33404 4498 33460 4510
rect 32508 3554 33012 3556
rect 32508 3502 32510 3554
rect 32562 3502 32958 3554
rect 33010 3502 33012 3554
rect 32508 3500 33012 3502
rect 32508 3490 32564 3500
rect 32956 3490 33012 3500
rect 33068 4172 33348 4228
rect 32172 3390 32174 3442
rect 32226 3390 32228 3442
rect 32172 3378 32228 3390
rect 33068 3332 33124 4172
rect 33628 4116 33684 4126
rect 33516 3556 33572 3566
rect 33180 3500 33516 3556
rect 33180 3442 33236 3500
rect 33516 3462 33572 3500
rect 33180 3390 33182 3442
rect 33234 3390 33236 3442
rect 33180 3378 33236 3390
rect 32284 3276 33124 3332
rect 33292 3332 33348 3342
rect 32284 800 32340 3276
rect 33292 3220 33348 3276
rect 32956 3164 33348 3220
rect 32956 800 33012 3164
rect 33628 800 33684 4060
rect 33740 3442 33796 4620
rect 33852 4338 33908 7308
rect 33964 7362 34020 8540
rect 34412 8260 34468 8766
rect 34188 8204 34412 8260
rect 34524 8260 34580 9548
rect 34636 8596 34692 9660
rect 34748 9650 34804 9660
rect 34748 9492 34804 9502
rect 34748 9266 34804 9436
rect 34748 9214 34750 9266
rect 34802 9214 34804 9266
rect 34748 9202 34804 9214
rect 34636 8530 34692 8540
rect 34636 8260 34692 8270
rect 34524 8258 34692 8260
rect 34524 8206 34638 8258
rect 34690 8206 34692 8258
rect 34524 8204 34692 8206
rect 34076 8148 34132 8158
rect 34076 8054 34132 8092
rect 34188 7476 34244 8204
rect 34412 8166 34468 8204
rect 34188 7410 34244 7420
rect 34300 8036 34356 8046
rect 34300 7586 34356 7980
rect 34636 7812 34692 8204
rect 34748 8260 34804 8270
rect 34860 8260 34916 10780
rect 35084 10722 35140 11342
rect 35420 11620 35476 11630
rect 35420 11394 35476 11564
rect 35644 11620 35700 11630
rect 35644 11526 35700 11564
rect 35980 11618 36036 12126
rect 35980 11566 35982 11618
rect 36034 11566 36036 11618
rect 35980 11554 36036 11566
rect 36428 12178 36484 12190
rect 36428 12126 36430 12178
rect 36482 12126 36484 12178
rect 36428 11620 36484 12126
rect 36428 11554 36484 11564
rect 36652 12178 36708 12190
rect 36652 12126 36654 12178
rect 36706 12126 36708 12178
rect 35420 11342 35422 11394
rect 35474 11342 35476 11394
rect 35420 11330 35476 11342
rect 35868 11394 35924 11406
rect 35868 11342 35870 11394
rect 35922 11342 35924 11394
rect 35868 11284 35924 11342
rect 35868 11218 35924 11228
rect 36652 10834 36708 12126
rect 36652 10782 36654 10834
rect 36706 10782 36708 10834
rect 36652 10770 36708 10782
rect 35084 10670 35086 10722
rect 35138 10670 35140 10722
rect 35084 10658 35140 10670
rect 36764 10722 36820 10734
rect 36764 10670 36766 10722
rect 36818 10670 36820 10722
rect 35644 10612 35700 10622
rect 35084 10388 35140 10398
rect 34972 9716 35028 9726
rect 34972 9268 35028 9660
rect 35084 9602 35140 10332
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35644 9828 35700 10556
rect 35980 10612 36036 10622
rect 36764 10612 36820 10670
rect 35980 10610 36820 10612
rect 35980 10558 35982 10610
rect 36034 10558 36820 10610
rect 35980 10556 36820 10558
rect 35868 10498 35924 10510
rect 35868 10446 35870 10498
rect 35922 10446 35924 10498
rect 35868 10388 35924 10446
rect 35868 10322 35924 10332
rect 35644 9734 35700 9772
rect 35980 9826 36036 10556
rect 36540 10388 36596 10398
rect 36540 10294 36596 10332
rect 36652 10276 36708 10286
rect 35980 9774 35982 9826
rect 36034 9774 36036 9826
rect 35980 9762 36036 9774
rect 36540 9828 36596 9838
rect 36652 9828 36708 10220
rect 37100 9938 37156 13020
rect 37212 12180 37268 12190
rect 37212 12086 37268 12124
rect 37100 9886 37102 9938
rect 37154 9886 37156 9938
rect 37100 9874 37156 9886
rect 36540 9826 36708 9828
rect 36540 9774 36542 9826
rect 36594 9774 36708 9826
rect 36540 9772 36708 9774
rect 36540 9762 36596 9772
rect 35084 9550 35086 9602
rect 35138 9550 35140 9602
rect 35084 9538 35140 9550
rect 35308 9714 35364 9726
rect 35308 9662 35310 9714
rect 35362 9662 35364 9714
rect 35308 9492 35364 9662
rect 36204 9714 36260 9726
rect 36204 9662 36206 9714
rect 36258 9662 36260 9714
rect 35756 9604 35812 9614
rect 35308 9426 35364 9436
rect 35532 9548 35756 9604
rect 35196 9268 35252 9278
rect 34972 9266 35252 9268
rect 34972 9214 35198 9266
rect 35250 9214 35252 9266
rect 34972 9212 35252 9214
rect 35196 9202 35252 9212
rect 35532 9266 35588 9548
rect 35756 9510 35812 9548
rect 36204 9492 36260 9662
rect 36316 9716 36372 9726
rect 36316 9622 36372 9660
rect 36204 9426 36260 9436
rect 36876 9492 36932 9502
rect 35532 9214 35534 9266
rect 35586 9214 35588 9266
rect 35308 9156 35364 9166
rect 35308 9062 35364 9100
rect 34804 8204 34916 8260
rect 35084 9042 35140 9054
rect 35084 8990 35086 9042
rect 35138 8990 35140 9042
rect 34748 8194 34804 8204
rect 35084 8148 35140 8990
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 35308 8260 35364 8270
rect 35308 8258 35476 8260
rect 35308 8206 35310 8258
rect 35362 8206 35476 8258
rect 35308 8204 35476 8206
rect 35308 8194 35364 8204
rect 35084 8082 35140 8092
rect 34636 7746 34692 7756
rect 35308 7700 35364 7710
rect 35308 7606 35364 7644
rect 34300 7534 34302 7586
rect 34354 7534 34356 7586
rect 33964 7310 33966 7362
rect 34018 7310 34020 7362
rect 33964 7298 34020 7310
rect 34300 6916 34356 7534
rect 35420 7588 35476 8204
rect 35532 8146 35588 9214
rect 36428 9268 36484 9278
rect 36484 9212 36596 9268
rect 35980 9156 36036 9166
rect 35980 9062 36036 9100
rect 36316 9156 36372 9166
rect 36092 9044 36148 9054
rect 36092 8950 36148 8988
rect 35868 8148 35924 8158
rect 35532 8094 35534 8146
rect 35586 8094 35588 8146
rect 35532 8082 35588 8094
rect 35756 8146 35924 8148
rect 35756 8094 35870 8146
rect 35922 8094 35924 8146
rect 35756 8092 35924 8094
rect 35420 7522 35476 7532
rect 34636 7474 34692 7486
rect 34636 7422 34638 7474
rect 34690 7422 34692 7474
rect 34300 6850 34356 6860
rect 34412 7364 34468 7374
rect 34412 6578 34468 7308
rect 34412 6526 34414 6578
rect 34466 6526 34468 6578
rect 34412 6514 34468 6526
rect 34076 6468 34132 6478
rect 33964 6466 34132 6468
rect 33964 6414 34078 6466
rect 34130 6414 34132 6466
rect 33964 6412 34132 6414
rect 33964 5572 34020 6412
rect 34076 6402 34132 6412
rect 34636 6468 34692 7422
rect 35084 7474 35140 7486
rect 35756 7476 35812 8092
rect 35868 8082 35924 8092
rect 35980 8148 36036 8158
rect 35980 8054 36036 8092
rect 36204 8036 36260 8046
rect 36204 7942 36260 7980
rect 35084 7422 35086 7474
rect 35138 7422 35140 7474
rect 34636 6402 34692 6412
rect 34860 6466 34916 6478
rect 34860 6414 34862 6466
rect 34914 6414 34916 6466
rect 34860 6132 34916 6414
rect 34300 6076 34916 6132
rect 33964 5506 34020 5516
rect 34076 5908 34132 5918
rect 34300 5908 34356 6076
rect 34076 5906 34356 5908
rect 34076 5854 34078 5906
rect 34130 5854 34356 5906
rect 34076 5852 34356 5854
rect 34524 5908 34580 5918
rect 33964 5348 34020 5358
rect 33964 5010 34020 5292
rect 33964 4958 33966 5010
rect 34018 4958 34020 5010
rect 33964 4946 34020 4958
rect 33852 4286 33854 4338
rect 33906 4286 33908 4338
rect 33852 4274 33908 4286
rect 33740 3390 33742 3442
rect 33794 3390 33796 3442
rect 33740 3378 33796 3390
rect 33964 3444 34020 3454
rect 34076 3444 34132 5852
rect 34524 5814 34580 5852
rect 34636 5906 34692 5918
rect 34636 5854 34638 5906
rect 34690 5854 34692 5906
rect 34636 5124 34692 5854
rect 34748 5906 34804 5918
rect 34748 5854 34750 5906
rect 34802 5854 34804 5906
rect 34748 5684 34804 5854
rect 35084 5684 35140 7422
rect 35644 7474 35812 7476
rect 35644 7422 35758 7474
rect 35810 7422 35812 7474
rect 35644 7420 35812 7422
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35644 6916 35700 7420
rect 35756 7410 35812 7420
rect 35868 7700 35924 7710
rect 35308 6860 35700 6916
rect 35196 6580 35252 6590
rect 35308 6580 35364 6860
rect 35756 6804 35812 6814
rect 35756 6710 35812 6748
rect 35868 6690 35924 7644
rect 36316 7474 36372 9100
rect 36316 7422 36318 7474
rect 36370 7422 36372 7474
rect 36316 7410 36372 7422
rect 35868 6638 35870 6690
rect 35922 6638 35924 6690
rect 35868 6626 35924 6638
rect 35196 6578 35364 6580
rect 35196 6526 35198 6578
rect 35250 6526 35364 6578
rect 35196 6524 35364 6526
rect 35420 6580 35476 6590
rect 35196 6244 35252 6524
rect 35420 6356 35476 6524
rect 36204 6578 36260 6590
rect 36204 6526 36206 6578
rect 36258 6526 36260 6578
rect 35644 6468 35700 6478
rect 35196 6178 35252 6188
rect 35308 6300 35476 6356
rect 35532 6356 35588 6366
rect 34748 5628 35140 5684
rect 35196 5908 35252 5918
rect 35308 5908 35364 6300
rect 35420 6132 35476 6142
rect 35532 6132 35588 6300
rect 35420 6130 35588 6132
rect 35420 6078 35422 6130
rect 35474 6078 35588 6130
rect 35420 6076 35588 6078
rect 35420 6066 35476 6076
rect 35196 5906 35364 5908
rect 35196 5854 35198 5906
rect 35250 5854 35364 5906
rect 35196 5852 35364 5854
rect 35644 5908 35700 6412
rect 36204 6356 36260 6526
rect 36428 6580 36484 9212
rect 36540 9154 36596 9212
rect 36876 9266 36932 9436
rect 36876 9214 36878 9266
rect 36930 9214 36932 9266
rect 36876 9202 36932 9214
rect 36540 9102 36542 9154
rect 36594 9102 36596 9154
rect 36540 9090 36596 9102
rect 36652 8260 36708 8270
rect 36652 7700 36708 8204
rect 36988 8148 37044 8158
rect 36652 7586 36708 7644
rect 36876 8146 37044 8148
rect 36876 8094 36990 8146
rect 37042 8094 37044 8146
rect 36876 8092 37044 8094
rect 36652 7534 36654 7586
rect 36706 7534 36708 7586
rect 36652 7522 36708 7534
rect 36764 7588 36820 7598
rect 36764 7140 36820 7532
rect 36876 7252 36932 8092
rect 36988 8082 37044 8092
rect 37100 8034 37156 8046
rect 37100 7982 37102 8034
rect 37154 7982 37156 8034
rect 37100 7700 37156 7982
rect 37324 8034 37380 8046
rect 37324 7982 37326 8034
rect 37378 7982 37380 8034
rect 37212 7700 37268 7710
rect 37100 7698 37268 7700
rect 37100 7646 37214 7698
rect 37266 7646 37268 7698
rect 37100 7644 37268 7646
rect 37212 7634 37268 7644
rect 36988 7476 37044 7486
rect 36988 7474 37268 7476
rect 36988 7422 36990 7474
rect 37042 7422 37268 7474
rect 36988 7420 37268 7422
rect 36988 7410 37044 7420
rect 36876 7196 37044 7252
rect 36652 7084 36820 7140
rect 36540 6692 36596 6702
rect 36540 6598 36596 6636
rect 36428 6514 36484 6524
rect 36204 6290 36260 6300
rect 36316 6466 36372 6478
rect 36316 6414 36318 6466
rect 36370 6414 36372 6466
rect 35196 5684 35252 5852
rect 35644 5842 35700 5852
rect 35868 6130 35924 6142
rect 35868 6078 35870 6130
rect 35922 6078 35924 6130
rect 34748 5348 34804 5628
rect 35196 5618 35252 5628
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 34748 5282 34804 5292
rect 34972 5348 35028 5358
rect 34300 5012 34356 5022
rect 34300 3554 34356 4956
rect 34300 3502 34302 3554
rect 34354 3502 34356 3554
rect 34300 3490 34356 3502
rect 34636 3556 34692 5068
rect 34972 5122 35028 5292
rect 34972 5070 34974 5122
rect 35026 5070 35028 5122
rect 34972 5058 35028 5070
rect 35868 5124 35924 6078
rect 36316 6132 36372 6414
rect 36316 6066 36372 6076
rect 35868 5030 35924 5068
rect 36092 5908 36148 5918
rect 36092 5122 36148 5852
rect 36316 5906 36372 5918
rect 36316 5854 36318 5906
rect 36370 5854 36372 5906
rect 36316 5572 36372 5854
rect 36428 5572 36484 5582
rect 36316 5516 36428 5572
rect 36428 5234 36484 5516
rect 36428 5182 36430 5234
rect 36482 5182 36484 5234
rect 36428 5170 36484 5182
rect 36092 5070 36094 5122
rect 36146 5070 36148 5122
rect 36092 5058 36148 5070
rect 36316 5124 36372 5134
rect 35196 5010 35252 5022
rect 35196 4958 35198 5010
rect 35250 4958 35252 5010
rect 34748 4676 34804 4686
rect 34748 3556 34804 4620
rect 35196 4340 35252 4958
rect 35644 5012 35700 5022
rect 35420 4900 35476 4910
rect 35420 4806 35476 4844
rect 35196 4274 35252 4284
rect 34860 4116 34916 4126
rect 34860 4022 34916 4060
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 35084 3780 35140 3790
rect 35084 3686 35140 3724
rect 34972 3668 35028 3678
rect 34860 3556 34916 3566
rect 34748 3500 34860 3556
rect 34636 3490 34692 3500
rect 34860 3462 34916 3500
rect 34020 3388 34132 3444
rect 34412 3444 34468 3454
rect 33964 3378 34020 3388
rect 34412 3332 34468 3388
rect 34300 3276 34468 3332
rect 34300 800 34356 3276
rect 34972 800 35028 3612
rect 35532 3444 35588 3482
rect 35532 3378 35588 3388
rect 35644 800 35700 4956
rect 36316 5010 36372 5068
rect 36316 4958 36318 5010
rect 36370 4958 36372 5010
rect 36316 4946 36372 4958
rect 36652 4788 36708 7084
rect 36988 7028 37044 7196
rect 36764 6972 37044 7028
rect 37100 7250 37156 7262
rect 37100 7198 37102 7250
rect 37154 7198 37156 7250
rect 36764 5908 36820 6972
rect 37100 6916 37156 7198
rect 37212 7252 37268 7420
rect 37212 7186 37268 7196
rect 36764 5814 36820 5852
rect 36876 6860 37156 6916
rect 36876 5572 36932 6860
rect 36988 6692 37044 6702
rect 36988 6690 37156 6692
rect 36988 6638 36990 6690
rect 37042 6638 37156 6690
rect 36988 6636 37156 6638
rect 36988 6626 37044 6636
rect 36876 5506 36932 5516
rect 36988 6468 37044 6478
rect 36988 5010 37044 6412
rect 37100 6132 37156 6636
rect 37212 6690 37268 6702
rect 37212 6638 37214 6690
rect 37266 6638 37268 6690
rect 37212 6356 37268 6638
rect 37212 6290 37268 6300
rect 37324 6244 37380 7982
rect 37436 7028 37492 15092
rect 37772 14642 37828 15372
rect 37772 14590 37774 14642
rect 37826 14590 37828 14642
rect 37772 14578 37828 14590
rect 37660 14532 37716 14542
rect 37660 14438 37716 14476
rect 38332 14420 38388 14430
rect 38780 14420 38836 15934
rect 38892 15932 39004 15988
rect 38892 15874 38948 15932
rect 39004 15922 39060 15932
rect 38892 15822 38894 15874
rect 38946 15822 38948 15874
rect 38892 14644 38948 15822
rect 39004 15314 39060 15326
rect 39004 15262 39006 15314
rect 39058 15262 39060 15314
rect 39004 14980 39060 15262
rect 39004 14914 39060 14924
rect 39116 15314 39172 15326
rect 39116 15262 39118 15314
rect 39170 15262 39172 15314
rect 39116 14756 39172 15262
rect 39340 15316 39396 15326
rect 39340 15222 39396 15260
rect 39452 15148 39508 16046
rect 39564 16380 39956 16436
rect 40012 16882 40068 16894
rect 40012 16830 40014 16882
rect 40066 16830 40068 16882
rect 39564 16098 39620 16380
rect 40012 16324 40068 16830
rect 39564 16046 39566 16098
rect 39618 16046 39620 16098
rect 39564 15988 39620 16046
rect 39564 15922 39620 15932
rect 39788 16268 40068 16324
rect 40124 16660 40180 16670
rect 39788 15986 39844 16268
rect 39900 16100 39956 16110
rect 39900 16006 39956 16044
rect 39788 15934 39790 15986
rect 39842 15934 39844 15986
rect 39676 15314 39732 15326
rect 39676 15262 39678 15314
rect 39730 15262 39732 15314
rect 39452 15092 39620 15148
rect 39116 14700 39284 14756
rect 38892 14588 39172 14644
rect 39004 14420 39060 14430
rect 38780 14418 39060 14420
rect 38780 14366 39006 14418
rect 39058 14366 39060 14418
rect 38780 14364 39060 14366
rect 38332 14326 38388 14364
rect 39004 14354 39060 14364
rect 39116 14196 39172 14588
rect 39004 14140 39172 14196
rect 39228 14530 39284 14700
rect 39228 14478 39230 14530
rect 39282 14478 39284 14530
rect 38556 13858 38612 13870
rect 38556 13806 38558 13858
rect 38610 13806 38612 13858
rect 37660 13748 37716 13758
rect 37548 11396 37604 11406
rect 37548 11302 37604 11340
rect 37660 11172 37716 13692
rect 37996 13748 38052 13758
rect 37996 12404 38052 13692
rect 38444 13748 38500 13758
rect 38444 12964 38500 13692
rect 38556 13300 38612 13806
rect 38892 13746 38948 13758
rect 38892 13694 38894 13746
rect 38946 13694 38948 13746
rect 38556 13244 38836 13300
rect 38556 12964 38612 12974
rect 38444 12962 38612 12964
rect 38444 12910 38558 12962
rect 38610 12910 38612 12962
rect 38444 12908 38612 12910
rect 38556 12898 38612 12908
rect 38780 12962 38836 13244
rect 38780 12910 38782 12962
rect 38834 12910 38836 12962
rect 38780 12898 38836 12910
rect 38332 12852 38388 12862
rect 38108 12740 38164 12750
rect 38108 12646 38164 12684
rect 38220 12738 38276 12750
rect 38220 12686 38222 12738
rect 38274 12686 38276 12738
rect 38220 12628 38276 12686
rect 38220 12562 38276 12572
rect 38220 12404 38276 12414
rect 37996 12402 38276 12404
rect 37996 12350 38222 12402
rect 38274 12350 38276 12402
rect 37996 12348 38276 12350
rect 38220 12338 38276 12348
rect 37996 12178 38052 12190
rect 37996 12126 37998 12178
rect 38050 12126 38052 12178
rect 37548 11116 37716 11172
rect 37884 11394 37940 11406
rect 37884 11342 37886 11394
rect 37938 11342 37940 11394
rect 37548 7362 37604 11116
rect 37884 10834 37940 11342
rect 37884 10782 37886 10834
rect 37938 10782 37940 10834
rect 37884 10770 37940 10782
rect 37996 10500 38052 12126
rect 38332 11508 38388 12796
rect 38444 12740 38500 12750
rect 38444 12738 38612 12740
rect 38444 12686 38446 12738
rect 38498 12686 38612 12738
rect 38444 12684 38612 12686
rect 38444 12674 38500 12684
rect 38444 11508 38500 11518
rect 38332 11506 38500 11508
rect 38332 11454 38446 11506
rect 38498 11454 38500 11506
rect 38332 11452 38500 11454
rect 38444 11442 38500 11452
rect 38444 11284 38500 11294
rect 38332 11228 38444 11284
rect 38108 10836 38164 10846
rect 38108 10742 38164 10780
rect 38220 10724 38276 10734
rect 38332 10724 38388 11228
rect 38444 11218 38500 11228
rect 38220 10722 38388 10724
rect 38220 10670 38222 10722
rect 38274 10670 38388 10722
rect 38220 10668 38388 10670
rect 38444 10724 38500 10734
rect 38556 10724 38612 12684
rect 38892 12628 38948 13694
rect 38892 12562 38948 12572
rect 39004 12850 39060 14140
rect 39228 13748 39284 14478
rect 39228 13682 39284 13692
rect 39564 12964 39620 15092
rect 39676 14980 39732 15262
rect 39676 14914 39732 14924
rect 39788 14196 39844 15934
rect 40124 15538 40180 16604
rect 40124 15486 40126 15538
rect 40178 15486 40180 15538
rect 40124 15474 40180 15486
rect 40236 16100 40292 16110
rect 40236 15426 40292 16044
rect 40348 16100 40404 16110
rect 40572 16100 40628 16110
rect 40348 16098 40628 16100
rect 40348 16046 40350 16098
rect 40402 16046 40574 16098
rect 40626 16046 40628 16098
rect 40348 16044 40628 16046
rect 40348 16034 40404 16044
rect 40572 16034 40628 16044
rect 40236 15374 40238 15426
rect 40290 15374 40292 15426
rect 40236 15362 40292 15374
rect 39900 15316 39956 15326
rect 39956 15260 40180 15316
rect 39900 15222 39956 15260
rect 40012 15092 40068 15102
rect 39900 14196 39956 14206
rect 39788 14140 39900 14196
rect 39788 13746 39844 13758
rect 39788 13694 39790 13746
rect 39842 13694 39844 13746
rect 39788 13186 39844 13694
rect 39788 13134 39790 13186
rect 39842 13134 39844 13186
rect 39788 13122 39844 13134
rect 39228 12908 39844 12964
rect 39004 12798 39006 12850
rect 39058 12798 39060 12850
rect 38892 12404 38948 12414
rect 39004 12404 39060 12798
rect 38892 12402 39060 12404
rect 38892 12350 38894 12402
rect 38946 12350 39060 12402
rect 38892 12348 39060 12350
rect 39116 12850 39172 12862
rect 39116 12798 39118 12850
rect 39170 12798 39172 12850
rect 39116 12740 39172 12798
rect 38892 12338 38948 12348
rect 38668 12178 38724 12190
rect 38668 12126 38670 12178
rect 38722 12126 38724 12178
rect 38668 11508 38724 12126
rect 39116 11844 39172 12684
rect 39004 11788 39172 11844
rect 38668 11452 38948 11508
rect 38892 11396 38948 11452
rect 38780 11282 38836 11294
rect 38780 11230 38782 11282
rect 38834 11230 38836 11282
rect 38500 10668 38612 10724
rect 38668 11060 38724 11070
rect 38220 10658 38276 10668
rect 38444 10658 38500 10668
rect 38668 10612 38724 11004
rect 38780 10836 38836 11230
rect 38780 10770 38836 10780
rect 38780 10612 38836 10622
rect 38668 10610 38836 10612
rect 38668 10558 38782 10610
rect 38834 10558 38836 10610
rect 38668 10556 38836 10558
rect 38780 10546 38836 10556
rect 37996 10434 38052 10444
rect 38668 10388 38724 10398
rect 38332 9938 38388 9950
rect 38332 9886 38334 9938
rect 38386 9886 38388 9938
rect 37548 7310 37550 7362
rect 37602 7310 37604 7362
rect 37548 7298 37604 7310
rect 37660 9826 37716 9838
rect 37660 9774 37662 9826
rect 37714 9774 37716 9826
rect 37436 6972 37604 7028
rect 37436 6804 37492 6814
rect 37436 6710 37492 6748
rect 37548 6580 37604 6972
rect 37548 6514 37604 6524
rect 37324 6178 37380 6188
rect 37100 6066 37156 6076
rect 37660 6132 37716 9774
rect 37884 9828 37940 9838
rect 38332 9828 38388 9886
rect 37884 9826 38388 9828
rect 37884 9774 37886 9826
rect 37938 9774 38388 9826
rect 37884 9772 38388 9774
rect 38444 9828 38500 9838
rect 37884 9762 37940 9772
rect 38332 9604 38388 9614
rect 38220 9602 38388 9604
rect 38220 9550 38334 9602
rect 38386 9550 38388 9602
rect 38220 9548 38388 9550
rect 38220 9492 38276 9548
rect 38332 9538 38388 9548
rect 38220 9426 38276 9436
rect 38444 9266 38500 9772
rect 38444 9214 38446 9266
rect 38498 9214 38500 9266
rect 38444 9202 38500 9214
rect 38668 9826 38724 10332
rect 38892 10276 38948 11340
rect 39004 11060 39060 11788
rect 39116 11284 39172 11294
rect 39228 11284 39284 12908
rect 39788 12850 39844 12908
rect 39788 12798 39790 12850
rect 39842 12798 39844 12850
rect 39788 12786 39844 12798
rect 39900 12850 39956 14140
rect 39900 12798 39902 12850
rect 39954 12798 39956 12850
rect 39900 12628 39956 12798
rect 39116 11282 39284 11284
rect 39116 11230 39118 11282
rect 39170 11230 39284 11282
rect 39116 11228 39284 11230
rect 39116 11218 39172 11228
rect 39228 11172 39284 11228
rect 39228 11106 39284 11116
rect 39452 12572 39956 12628
rect 39116 11060 39172 11070
rect 39004 11004 39116 11060
rect 39116 10994 39172 11004
rect 39452 10836 39508 12572
rect 39564 12178 39620 12190
rect 39564 12126 39566 12178
rect 39618 12126 39620 12178
rect 39564 11618 39620 12126
rect 39564 11566 39566 11618
rect 39618 11566 39620 11618
rect 39564 11554 39620 11566
rect 39788 12066 39844 12078
rect 39788 12014 39790 12066
rect 39842 12014 39844 12066
rect 39564 11396 39620 11406
rect 39788 11396 39844 12014
rect 40012 11954 40068 15036
rect 40124 12292 40180 15260
rect 40684 15148 40740 16940
rect 40796 16772 40852 16782
rect 40796 16322 40852 16716
rect 40908 16660 40964 16670
rect 40908 16566 40964 16604
rect 40796 16270 40798 16322
rect 40850 16270 40852 16322
rect 40796 16258 40852 16270
rect 40908 16436 40964 16446
rect 40348 15092 40740 15148
rect 40236 15036 40404 15092
rect 40236 13858 40292 15036
rect 40908 14868 40964 16380
rect 41020 15876 41076 18060
rect 41804 17668 41860 18174
rect 41916 18228 41972 24556
rect 42364 24612 42420 24622
rect 42364 24610 42644 24612
rect 42364 24558 42366 24610
rect 42418 24558 42644 24610
rect 42364 24556 42644 24558
rect 42364 24546 42420 24556
rect 42252 24500 42308 24510
rect 42028 24498 42308 24500
rect 42028 24446 42254 24498
rect 42306 24446 42308 24498
rect 42028 24444 42308 24446
rect 42028 23266 42084 24444
rect 42252 24434 42308 24444
rect 42028 23214 42030 23266
rect 42082 23214 42084 23266
rect 42028 23202 42084 23214
rect 42252 23156 42308 23166
rect 42140 23044 42196 23054
rect 42140 22370 42196 22988
rect 42140 22318 42142 22370
rect 42194 22318 42196 22370
rect 42140 22306 42196 22318
rect 42028 20692 42084 20702
rect 42028 20598 42084 20636
rect 42028 20132 42084 20142
rect 42252 20132 42308 23100
rect 42028 20130 42308 20132
rect 42028 20078 42030 20130
rect 42082 20078 42308 20130
rect 42028 20076 42308 20078
rect 42476 22596 42532 22606
rect 42476 22370 42532 22540
rect 42588 22482 42644 24556
rect 42588 22430 42590 22482
rect 42642 22430 42644 22482
rect 42588 22418 42644 22430
rect 43036 22484 43092 22494
rect 43036 22390 43092 22428
rect 42476 22318 42478 22370
rect 42530 22318 42532 22370
rect 42028 20066 42084 20076
rect 42476 19908 42532 22318
rect 42700 22372 42756 22382
rect 42700 22278 42756 22316
rect 44044 22370 44100 25340
rect 44156 25394 44212 26012
rect 44156 25342 44158 25394
rect 44210 25342 44212 25394
rect 44156 25330 44212 25342
rect 44268 25508 44324 25518
rect 44492 25508 44548 26238
rect 44268 25506 44548 25508
rect 44268 25454 44270 25506
rect 44322 25454 44548 25506
rect 44268 25452 44548 25454
rect 44268 24946 44324 25452
rect 44940 25396 44996 26462
rect 45052 25618 45108 27468
rect 45500 27412 45556 27422
rect 45500 27074 45556 27356
rect 45500 27022 45502 27074
rect 45554 27022 45556 27074
rect 45500 27010 45556 27022
rect 45612 26908 45668 27580
rect 45948 27186 46004 28476
rect 46284 28420 46340 29932
rect 46284 28354 46340 28364
rect 46060 28084 46116 28094
rect 46060 27990 46116 28028
rect 46732 28084 46788 32060
rect 46844 31892 46900 36652
rect 47068 36484 47124 36494
rect 47068 36390 47124 36428
rect 47292 36260 47348 36270
rect 47292 35700 47348 36204
rect 47404 36258 47460 36270
rect 47404 36206 47406 36258
rect 47458 36206 47460 36258
rect 47404 35924 47460 36206
rect 47404 35858 47460 35868
rect 47628 35812 47684 35822
rect 47404 35700 47460 35710
rect 47292 35698 47460 35700
rect 47292 35646 47406 35698
rect 47458 35646 47460 35698
rect 47292 35644 47460 35646
rect 47404 35634 47460 35644
rect 47516 35700 47572 35710
rect 47516 35026 47572 35644
rect 47628 35698 47684 35756
rect 47628 35646 47630 35698
rect 47682 35646 47684 35698
rect 47628 35634 47684 35646
rect 47740 35028 47796 38668
rect 48748 38724 48804 38734
rect 48748 38630 48804 38668
rect 48300 38500 48356 38510
rect 48300 37938 48356 38444
rect 48300 37886 48302 37938
rect 48354 37886 48356 37938
rect 48300 37268 48356 37886
rect 48524 38050 48580 38062
rect 48524 37998 48526 38050
rect 48578 37998 48580 38050
rect 48524 37828 48580 37998
rect 48524 37762 48580 37772
rect 49196 37940 49252 38782
rect 49756 38836 49812 42030
rect 49980 41970 50036 42252
rect 49980 41918 49982 41970
rect 50034 41918 50036 41970
rect 49868 40292 49924 40302
rect 49868 39842 49924 40236
rect 49980 40180 50036 41918
rect 50092 41860 50148 42588
rect 50092 41794 50148 41804
rect 50092 41188 50148 41198
rect 50204 41188 50260 43262
rect 50428 43316 50484 44156
rect 50556 43932 50820 43942
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50556 43866 50820 43876
rect 50428 43250 50484 43260
rect 50876 43092 50932 44382
rect 50988 44100 51044 45166
rect 51212 45108 51268 45614
rect 51884 45666 51940 45678
rect 51884 45614 51886 45666
rect 51938 45614 51940 45666
rect 51212 45042 51268 45052
rect 51772 45108 51828 45118
rect 51548 44996 51604 45006
rect 51548 44902 51604 44940
rect 51772 44436 51828 45052
rect 51884 44660 51940 45614
rect 52108 45220 52164 45838
rect 52780 45892 52836 45902
rect 52780 45798 52836 45836
rect 54236 45892 54292 45902
rect 54236 45798 54292 45836
rect 53340 45780 53396 45790
rect 53340 45686 53396 45724
rect 52556 45666 52612 45678
rect 52556 45614 52558 45666
rect 52610 45614 52612 45666
rect 52220 45332 52276 45342
rect 52220 45238 52276 45276
rect 52108 45154 52164 45164
rect 51996 45108 52052 45118
rect 51996 45014 52052 45052
rect 52108 44996 52164 45006
rect 52108 44902 52164 44940
rect 51884 44604 52164 44660
rect 51772 44370 51828 44380
rect 50988 44034 51044 44044
rect 51884 44098 51940 44110
rect 51884 44046 51886 44098
rect 51938 44046 51940 44098
rect 51548 43652 51604 43662
rect 51212 43540 51268 43550
rect 51212 43446 51268 43484
rect 51548 43538 51604 43596
rect 51548 43486 51550 43538
rect 51602 43486 51604 43538
rect 51548 43474 51604 43486
rect 51884 43540 51940 44046
rect 51660 43426 51716 43438
rect 51660 43374 51662 43426
rect 51714 43374 51716 43426
rect 51548 43316 51604 43326
rect 50876 43026 50932 43036
rect 51324 43092 51380 43102
rect 51324 42978 51380 43036
rect 51324 42926 51326 42978
rect 51378 42926 51380 42978
rect 51324 42914 51380 42926
rect 51548 42642 51604 43260
rect 51548 42590 51550 42642
rect 51602 42590 51604 42642
rect 51548 42578 51604 42590
rect 51436 42530 51492 42542
rect 51436 42478 51438 42530
rect 51490 42478 51492 42530
rect 50556 42364 50820 42374
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50556 42298 50820 42308
rect 50764 42194 50820 42206
rect 50764 42142 50766 42194
rect 50818 42142 50820 42194
rect 50652 41972 50708 41982
rect 50316 41970 50708 41972
rect 50316 41918 50654 41970
rect 50706 41918 50708 41970
rect 50316 41916 50708 41918
rect 50316 41410 50372 41916
rect 50652 41906 50708 41916
rect 50764 41860 50820 42142
rect 50764 41794 50820 41804
rect 50316 41358 50318 41410
rect 50370 41358 50372 41410
rect 50316 41346 50372 41358
rect 51324 41300 51380 41310
rect 51436 41300 51492 42478
rect 51324 41298 51492 41300
rect 51324 41246 51326 41298
rect 51378 41246 51492 41298
rect 51324 41244 51492 41246
rect 51324 41234 51380 41244
rect 50092 41186 50260 41188
rect 50092 41134 50094 41186
rect 50146 41134 50260 41186
rect 50092 41132 50260 41134
rect 51436 41188 51492 41244
rect 50092 41122 50148 41132
rect 50652 41076 50708 41086
rect 50652 40982 50708 41020
rect 50556 40796 50820 40806
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50556 40730 50820 40740
rect 50204 40404 50260 40414
rect 50204 40310 50260 40348
rect 51100 40404 51156 40414
rect 49980 40124 50372 40180
rect 49868 39790 49870 39842
rect 49922 39790 49924 39842
rect 49868 39778 49924 39790
rect 50204 39394 50260 39406
rect 50204 39342 50206 39394
rect 50258 39342 50260 39394
rect 50092 38836 50148 38846
rect 49756 38834 50148 38836
rect 49756 38782 50094 38834
rect 50146 38782 50148 38834
rect 49756 38780 50148 38782
rect 49532 38722 49588 38734
rect 49532 38670 49534 38722
rect 49586 38670 49588 38722
rect 48300 37202 48356 37212
rect 49196 37266 49252 37884
rect 49196 37214 49198 37266
rect 49250 37214 49252 37266
rect 49196 37202 49252 37214
rect 49420 37940 49476 37950
rect 48300 36370 48356 36382
rect 48300 36318 48302 36370
rect 48354 36318 48356 36370
rect 48188 35924 48244 35934
rect 47852 35700 47908 35710
rect 47852 35606 47908 35644
rect 47516 34974 47518 35026
rect 47570 34974 47572 35026
rect 47516 34962 47572 34974
rect 47628 34972 47796 35028
rect 48188 35588 48244 35868
rect 48300 35812 48356 36318
rect 48300 35746 48356 35756
rect 48412 36258 48468 36270
rect 48412 36206 48414 36258
rect 48466 36206 48468 36258
rect 47516 34244 47572 34254
rect 47516 34150 47572 34188
rect 47404 33908 47460 33918
rect 47180 33906 47460 33908
rect 47180 33854 47406 33906
rect 47458 33854 47460 33906
rect 47180 33852 47460 33854
rect 47180 33460 47236 33852
rect 47404 33842 47460 33852
rect 47180 33346 47236 33404
rect 47180 33294 47182 33346
rect 47234 33294 47236 33346
rect 47180 33282 47236 33294
rect 47404 33346 47460 33358
rect 47404 33294 47406 33346
rect 47458 33294 47460 33346
rect 47404 33236 47460 33294
rect 47404 33170 47460 33180
rect 47516 33122 47572 33134
rect 47516 33070 47518 33122
rect 47570 33070 47572 33122
rect 47516 32228 47572 33070
rect 47628 32900 47684 34972
rect 47740 34802 47796 34814
rect 47740 34750 47742 34802
rect 47794 34750 47796 34802
rect 47740 34354 47796 34750
rect 47740 34302 47742 34354
rect 47794 34302 47796 34354
rect 47740 34290 47796 34302
rect 47852 34356 47908 34366
rect 48076 34356 48132 34366
rect 47908 34300 48020 34356
rect 47852 34290 47908 34300
rect 47964 34242 48020 34300
rect 47964 34190 47966 34242
rect 48018 34190 48020 34242
rect 47964 34178 48020 34190
rect 48076 34242 48132 34300
rect 48076 34190 48078 34242
rect 48130 34190 48132 34242
rect 48076 34020 48132 34190
rect 47740 33964 48132 34020
rect 47740 33346 47796 33964
rect 47740 33294 47742 33346
rect 47794 33294 47796 33346
rect 47740 33282 47796 33294
rect 48188 33346 48244 35532
rect 48300 35474 48356 35486
rect 48300 35422 48302 35474
rect 48354 35422 48356 35474
rect 48300 34132 48356 35422
rect 48412 34916 48468 36206
rect 48524 36260 48580 36270
rect 48524 36166 48580 36204
rect 49084 36260 49140 36270
rect 49084 35922 49140 36204
rect 49084 35870 49086 35922
rect 49138 35870 49140 35922
rect 49084 35858 49140 35870
rect 49308 35812 49364 35822
rect 49308 35718 49364 35756
rect 48636 35700 48692 35710
rect 48636 35606 48692 35644
rect 49196 35586 49252 35598
rect 49196 35534 49198 35586
rect 49250 35534 49252 35586
rect 48972 34916 49028 34926
rect 48412 34914 49028 34916
rect 48412 34862 48974 34914
rect 49026 34862 49028 34914
rect 48412 34860 49028 34862
rect 48972 34850 49028 34860
rect 48300 34066 48356 34076
rect 48748 34468 48804 34478
rect 48748 34132 48804 34412
rect 48972 34356 49028 34366
rect 48972 34242 49028 34300
rect 48972 34190 48974 34242
rect 49026 34190 49028 34242
rect 48972 34178 49028 34190
rect 49196 34244 49252 35534
rect 49196 34150 49252 34188
rect 49308 34132 49364 34142
rect 48748 34130 48916 34132
rect 48748 34078 48750 34130
rect 48802 34078 48916 34130
rect 48748 34076 48916 34078
rect 48748 34066 48804 34076
rect 48860 33684 48916 34076
rect 49308 34038 49364 34076
rect 48860 33628 49140 33684
rect 48748 33460 48804 33470
rect 48748 33366 48804 33404
rect 48188 33294 48190 33346
rect 48242 33294 48244 33346
rect 48188 33124 48244 33294
rect 48972 33348 49028 33358
rect 48972 33254 49028 33292
rect 48412 33236 48468 33246
rect 48412 33142 48468 33180
rect 48188 33058 48244 33068
rect 48524 33122 48580 33134
rect 48524 33070 48526 33122
rect 48578 33070 48580 33122
rect 47628 32834 47684 32844
rect 47516 32172 48020 32228
rect 46844 31798 46900 31836
rect 47068 32004 47124 32014
rect 46732 28018 46788 28028
rect 47068 27412 47124 31948
rect 47964 31892 48020 32172
rect 47964 31778 48020 31836
rect 47964 31726 47966 31778
rect 48018 31726 48020 31778
rect 47964 31714 48020 31726
rect 47964 31444 48020 31454
rect 47292 31108 47348 31118
rect 47292 30994 47348 31052
rect 47964 31106 48020 31388
rect 47964 31054 47966 31106
rect 48018 31054 48020 31106
rect 47964 31042 48020 31054
rect 48524 31108 48580 33070
rect 49084 33124 49140 33628
rect 49420 33348 49476 37884
rect 49532 37826 49588 38670
rect 49644 38164 49700 38174
rect 49644 37938 49700 38108
rect 49644 37886 49646 37938
rect 49698 37886 49700 37938
rect 49644 37874 49700 37886
rect 49532 37774 49534 37826
rect 49586 37774 49588 37826
rect 49532 37266 49588 37774
rect 50092 37828 50148 38780
rect 50204 38276 50260 39342
rect 50204 38210 50260 38220
rect 50316 38834 50372 40124
rect 51100 39618 51156 40348
rect 51100 39566 51102 39618
rect 51154 39566 51156 39618
rect 51100 39554 51156 39566
rect 51436 39618 51492 41132
rect 51548 41412 51604 41422
rect 51660 41412 51716 43374
rect 51884 42756 51940 43484
rect 51884 42690 51940 42700
rect 51548 41410 51660 41412
rect 51548 41358 51550 41410
rect 51602 41358 51660 41410
rect 51548 41356 51660 41358
rect 51548 39730 51604 41356
rect 51660 41318 51716 41356
rect 51772 41186 51828 41198
rect 51772 41134 51774 41186
rect 51826 41134 51828 41186
rect 51660 40964 51716 40974
rect 51660 40514 51716 40908
rect 51660 40462 51662 40514
rect 51714 40462 51716 40514
rect 51660 40450 51716 40462
rect 51772 40404 51828 41134
rect 51772 40338 51828 40348
rect 51996 40964 52052 40974
rect 51996 40402 52052 40908
rect 51996 40350 51998 40402
rect 52050 40350 52052 40402
rect 51996 40338 52052 40350
rect 51548 39678 51550 39730
rect 51602 39678 51604 39730
rect 51548 39666 51604 39678
rect 51436 39566 51438 39618
rect 51490 39566 51492 39618
rect 51436 39554 51492 39566
rect 51772 39506 51828 39518
rect 51772 39454 51774 39506
rect 51826 39454 51828 39506
rect 51100 39396 51156 39406
rect 50556 39228 50820 39238
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50556 39162 50820 39172
rect 50316 38782 50318 38834
rect 50370 38782 50372 38834
rect 50316 38276 50372 38782
rect 51100 39058 51156 39340
rect 51100 39006 51102 39058
rect 51154 39006 51156 39058
rect 51100 38724 51156 39006
rect 51548 38948 51604 38958
rect 51100 38658 51156 38668
rect 51324 38892 51548 38948
rect 50652 38610 50708 38622
rect 50652 38558 50654 38610
rect 50706 38558 50708 38610
rect 50540 38276 50596 38286
rect 50316 38274 50596 38276
rect 50316 38222 50542 38274
rect 50594 38222 50596 38274
rect 50316 38220 50596 38222
rect 50316 38164 50372 38220
rect 50540 38210 50596 38220
rect 50316 38098 50372 38108
rect 50652 37940 50708 38558
rect 51212 38276 51268 38286
rect 51212 38162 51268 38220
rect 51212 38110 51214 38162
rect 51266 38110 51268 38162
rect 50652 37884 50932 37940
rect 50316 37828 50372 37838
rect 50092 37772 50316 37828
rect 50316 37734 50372 37772
rect 50428 37826 50484 37838
rect 50428 37774 50430 37826
rect 50482 37774 50484 37826
rect 49532 37214 49534 37266
rect 49586 37214 49588 37266
rect 49532 37202 49588 37214
rect 50204 37492 50260 37502
rect 49980 36260 50036 36270
rect 49868 36258 50036 36260
rect 49868 36206 49982 36258
rect 50034 36206 50036 36258
rect 49868 36204 50036 36206
rect 49644 35810 49700 35822
rect 49644 35758 49646 35810
rect 49698 35758 49700 35810
rect 49644 34356 49700 35758
rect 49868 35476 49924 36204
rect 49980 36194 50036 36204
rect 49980 35700 50036 35710
rect 49980 35606 50036 35644
rect 49980 35476 50036 35486
rect 49868 35420 49980 35476
rect 49980 35410 50036 35420
rect 49700 34300 49924 34356
rect 49644 34290 49700 34300
rect 49756 34132 49812 34142
rect 49756 34038 49812 34076
rect 49420 33292 49700 33348
rect 49532 33124 49588 33134
rect 49084 33068 49476 33124
rect 49420 32786 49476 33068
rect 49420 32734 49422 32786
rect 49474 32734 49476 32786
rect 49420 32722 49476 32734
rect 48860 32676 48916 32686
rect 48860 32674 49028 32676
rect 48860 32622 48862 32674
rect 48914 32622 49028 32674
rect 48860 32620 49028 32622
rect 48860 32610 48916 32620
rect 48748 32562 48804 32574
rect 48748 32510 48750 32562
rect 48802 32510 48804 32562
rect 48748 32002 48804 32510
rect 48748 31950 48750 32002
rect 48802 31950 48804 32002
rect 48748 31938 48804 31950
rect 48860 32338 48916 32350
rect 48860 32286 48862 32338
rect 48914 32286 48916 32338
rect 48636 31780 48692 31790
rect 48636 31686 48692 31724
rect 48860 31444 48916 32286
rect 48972 32340 49028 32620
rect 49532 32674 49588 33068
rect 49532 32622 49534 32674
rect 49586 32622 49588 32674
rect 49532 32610 49588 32622
rect 49420 32340 49476 32350
rect 48972 32338 49476 32340
rect 48972 32286 49422 32338
rect 49474 32286 49476 32338
rect 48972 32284 49476 32286
rect 49308 31892 49364 31902
rect 49308 31798 49364 31836
rect 49420 31778 49476 32284
rect 49420 31726 49422 31778
rect 49474 31726 49476 31778
rect 49420 31714 49476 31726
rect 48916 31388 49476 31444
rect 48860 31350 48916 31388
rect 48524 31042 48580 31052
rect 48860 31220 48916 31230
rect 47292 30942 47294 30994
rect 47346 30942 47348 30994
rect 47292 30930 47348 30942
rect 48188 30996 48244 31006
rect 48188 30902 48244 30940
rect 47628 30882 47684 30894
rect 47628 30830 47630 30882
rect 47682 30830 47684 30882
rect 47628 30548 47684 30830
rect 47628 30210 47684 30492
rect 48748 30770 48804 30782
rect 48748 30718 48750 30770
rect 48802 30718 48804 30770
rect 47852 30324 47908 30334
rect 47852 30230 47908 30268
rect 48748 30324 48804 30718
rect 48748 30258 48804 30268
rect 47628 30158 47630 30210
rect 47682 30158 47684 30210
rect 47628 30146 47684 30158
rect 47292 30098 47348 30110
rect 47292 30046 47294 30098
rect 47346 30046 47348 30098
rect 47292 29764 47348 30046
rect 47292 29698 47348 29708
rect 45948 27134 45950 27186
rect 46002 27134 46004 27186
rect 45948 27122 46004 27134
rect 46508 27188 46564 27198
rect 46508 27094 46564 27132
rect 47068 27186 47124 27356
rect 47068 27134 47070 27186
rect 47122 27134 47124 27186
rect 47068 27122 47124 27134
rect 47516 27188 47572 27198
rect 47516 27094 47572 27132
rect 45724 27076 45780 27086
rect 45724 26982 45780 27020
rect 48860 26908 48916 31164
rect 49196 31108 49252 31118
rect 49196 31014 49252 31052
rect 49420 31106 49476 31388
rect 49420 31054 49422 31106
rect 49474 31054 49476 31106
rect 49420 31042 49476 31054
rect 49308 30996 49364 31006
rect 49308 30902 49364 30940
rect 49644 27636 49700 33292
rect 49868 33234 49924 34300
rect 49980 33348 50036 33358
rect 49980 33254 50036 33292
rect 49868 33182 49870 33234
rect 49922 33182 49924 33234
rect 49868 33170 49924 33182
rect 50092 33236 50148 33246
rect 50092 33142 50148 33180
rect 50204 32116 50260 37436
rect 50316 37156 50372 37166
rect 50316 37042 50372 37100
rect 50428 37154 50484 37774
rect 50556 37660 50820 37670
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50556 37594 50820 37604
rect 50652 37268 50708 37278
rect 50876 37268 50932 37884
rect 51100 37268 51156 37278
rect 50876 37266 51156 37268
rect 50876 37214 51102 37266
rect 51154 37214 51156 37266
rect 50876 37212 51156 37214
rect 50652 37174 50708 37212
rect 51100 37202 51156 37212
rect 50428 37102 50430 37154
rect 50482 37102 50484 37154
rect 50428 37090 50484 37102
rect 50316 36990 50318 37042
rect 50370 36990 50372 37042
rect 50316 36978 50372 36990
rect 50316 36484 50372 36494
rect 50316 36482 50484 36484
rect 50316 36430 50318 36482
rect 50370 36430 50484 36482
rect 50316 36428 50484 36430
rect 50316 36148 50372 36428
rect 50316 36082 50372 36092
rect 50428 35924 50484 36428
rect 51212 36370 51268 38110
rect 51212 36318 51214 36370
rect 51266 36318 51268 36370
rect 51212 36306 51268 36318
rect 51324 36148 51380 38892
rect 51548 38854 51604 38892
rect 51772 38834 51828 39454
rect 52108 39060 52164 44604
rect 52556 43428 52612 45614
rect 53228 45220 53284 45230
rect 53228 45126 53284 45164
rect 52780 44994 52836 45006
rect 52780 44942 52782 44994
rect 52834 44942 52836 44994
rect 52780 44884 52836 44942
rect 52780 44818 52836 44828
rect 52892 44772 52948 44782
rect 52668 44548 52724 44558
rect 52668 44434 52724 44492
rect 52892 44546 52948 44716
rect 52892 44494 52894 44546
rect 52946 44494 52948 44546
rect 52892 44482 52948 44494
rect 52668 44382 52670 44434
rect 52722 44382 52724 44434
rect 52668 44370 52724 44382
rect 53228 44098 53284 44110
rect 53228 44046 53230 44098
rect 53282 44046 53284 44098
rect 53004 43540 53060 43550
rect 53228 43540 53284 44046
rect 53564 43652 53620 43662
rect 53340 43540 53396 43550
rect 53004 43538 53396 43540
rect 53004 43486 53006 43538
rect 53058 43486 53342 43538
rect 53394 43486 53396 43538
rect 53004 43484 53396 43486
rect 53004 43474 53060 43484
rect 53340 43474 53396 43484
rect 53564 43538 53620 43596
rect 53564 43486 53566 43538
rect 53618 43486 53620 43538
rect 53564 43474 53620 43486
rect 52556 43362 52612 43372
rect 53900 43314 53956 43326
rect 53900 43262 53902 43314
rect 53954 43262 53956 43314
rect 52892 42868 52948 42878
rect 52444 42756 52500 42766
rect 52332 42700 52444 42756
rect 52332 41748 52388 42700
rect 52444 42690 52500 42700
rect 52444 41972 52500 41982
rect 52892 41972 52948 42812
rect 53900 42868 53956 43262
rect 53900 42802 53956 42812
rect 54348 42756 54404 42766
rect 54348 42662 54404 42700
rect 53452 42642 53508 42654
rect 53452 42590 53454 42642
rect 53506 42590 53508 42642
rect 52444 41970 52948 41972
rect 52444 41918 52446 41970
rect 52498 41918 52948 41970
rect 52444 41916 52948 41918
rect 53004 41972 53060 41982
rect 53340 41972 53396 41982
rect 53004 41970 53396 41972
rect 53004 41918 53006 41970
rect 53058 41918 53342 41970
rect 53394 41918 53396 41970
rect 53004 41916 53396 41918
rect 52444 41906 52500 41916
rect 53004 41906 53060 41916
rect 53340 41906 53396 41916
rect 53452 41972 53508 42590
rect 55692 42642 55748 42654
rect 55692 42590 55694 42642
rect 55746 42590 55748 42642
rect 53452 41906 53508 41916
rect 53564 41970 53620 41982
rect 53564 41918 53566 41970
rect 53618 41918 53620 41970
rect 52668 41748 52724 41758
rect 52332 41746 52724 41748
rect 52332 41694 52670 41746
rect 52722 41694 52724 41746
rect 52332 41692 52724 41694
rect 52668 41682 52724 41692
rect 53004 41412 53060 41422
rect 53004 41318 53060 41356
rect 53564 41412 53620 41918
rect 53788 41972 53844 41982
rect 53788 41878 53844 41916
rect 54684 41970 54740 41982
rect 54684 41918 54686 41970
rect 54738 41918 54740 41970
rect 54236 41860 54292 41870
rect 53564 41346 53620 41356
rect 54012 41746 54068 41758
rect 54012 41694 54014 41746
rect 54066 41694 54068 41746
rect 52668 41188 52724 41198
rect 52668 41094 52724 41132
rect 52108 38994 52164 39004
rect 52220 40962 52276 40974
rect 52220 40910 52222 40962
rect 52274 40910 52276 40962
rect 51772 38782 51774 38834
rect 51826 38782 51828 38834
rect 51436 38724 51492 38734
rect 51436 38630 51492 38668
rect 51772 38164 51828 38782
rect 52220 38834 52276 40910
rect 52892 40964 52948 40974
rect 52892 40870 52948 40908
rect 52892 40404 52948 40414
rect 52892 40310 52948 40348
rect 54012 39618 54068 41694
rect 54236 41298 54292 41804
rect 54684 41860 54740 41918
rect 55132 41972 55188 41982
rect 55692 41972 55748 42590
rect 55132 41970 55748 41972
rect 55132 41918 55134 41970
rect 55186 41918 55748 41970
rect 55132 41916 55748 41918
rect 54740 41804 54964 41860
rect 54684 41794 54740 41804
rect 54236 41246 54238 41298
rect 54290 41246 54292 41298
rect 54236 41234 54292 41246
rect 54460 41074 54516 41086
rect 54460 41022 54462 41074
rect 54514 41022 54516 41074
rect 54012 39566 54014 39618
rect 54066 39566 54068 39618
rect 52220 38782 52222 38834
rect 52274 38782 52276 38834
rect 52220 38770 52276 38782
rect 53788 38834 53844 38846
rect 53788 38782 53790 38834
rect 53842 38782 53844 38834
rect 51436 38108 51828 38164
rect 51884 38724 51940 38734
rect 51436 38050 51492 38108
rect 51884 38052 51940 38668
rect 52444 38612 52500 38622
rect 52444 38610 53284 38612
rect 52444 38558 52446 38610
rect 52498 38558 53284 38610
rect 52444 38556 53284 38558
rect 52444 38546 52500 38556
rect 51436 37998 51438 38050
rect 51490 37998 51492 38050
rect 51436 36482 51492 37998
rect 51436 36430 51438 36482
rect 51490 36430 51492 36482
rect 51436 36418 51492 36430
rect 51660 37996 51940 38052
rect 53228 38050 53284 38556
rect 53788 38388 53844 38782
rect 53788 38322 53844 38332
rect 54012 38722 54068 39566
rect 54012 38670 54014 38722
rect 54066 38670 54068 38722
rect 53228 37998 53230 38050
rect 53282 37998 53284 38050
rect 50556 36092 50820 36102
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50556 36026 50820 36036
rect 50876 36092 51380 36148
rect 50764 35924 50820 35934
rect 50428 35922 50820 35924
rect 50428 35870 50766 35922
rect 50818 35870 50820 35922
rect 50428 35868 50820 35870
rect 50764 35858 50820 35868
rect 50652 35700 50708 35710
rect 50876 35700 50932 36092
rect 51660 36036 51716 37996
rect 53228 37986 53284 37998
rect 54012 37938 54068 38670
rect 54236 40178 54292 40190
rect 54236 40126 54238 40178
rect 54290 40126 54292 40178
rect 54236 39730 54292 40126
rect 54236 39678 54238 39730
rect 54290 39678 54292 39730
rect 54236 38836 54292 39678
rect 54460 39956 54516 41022
rect 54908 40402 54964 41804
rect 54908 40350 54910 40402
rect 54962 40350 54964 40402
rect 54908 40338 54964 40350
rect 55132 40290 55188 41916
rect 55692 41186 55748 41916
rect 55692 41134 55694 41186
rect 55746 41134 55748 41186
rect 55692 41122 55748 41134
rect 56028 40962 56084 40974
rect 56028 40910 56030 40962
rect 56082 40910 56084 40962
rect 55580 40292 55636 40302
rect 55132 40238 55134 40290
rect 55186 40238 55188 40290
rect 55132 40226 55188 40238
rect 55356 40290 55636 40292
rect 55356 40238 55582 40290
rect 55634 40238 55636 40290
rect 55356 40236 55636 40238
rect 54460 39396 54516 39900
rect 55356 39618 55412 40236
rect 55580 40226 55636 40236
rect 55356 39566 55358 39618
rect 55410 39566 55412 39618
rect 55356 39554 55412 39566
rect 54572 39508 54628 39518
rect 54572 39506 54964 39508
rect 54572 39454 54574 39506
rect 54626 39454 54964 39506
rect 54572 39452 54964 39454
rect 54572 39442 54628 39452
rect 54460 39330 54516 39340
rect 54236 38050 54292 38780
rect 54684 38388 54740 38398
rect 54684 38162 54740 38332
rect 54908 38274 54964 39452
rect 55468 39396 55524 39406
rect 55468 39302 55524 39340
rect 55692 39396 55748 39406
rect 55692 39394 55972 39396
rect 55692 39342 55694 39394
rect 55746 39342 55972 39394
rect 55692 39340 55972 39342
rect 55692 39330 55748 39340
rect 55132 38836 55188 38846
rect 55132 38742 55188 38780
rect 55804 38612 55860 38622
rect 55804 38518 55860 38556
rect 54908 38222 54910 38274
rect 54962 38222 54964 38274
rect 54908 38210 54964 38222
rect 55132 38276 55188 38286
rect 54684 38110 54686 38162
rect 54738 38110 54740 38162
rect 54684 38098 54740 38110
rect 54236 37998 54238 38050
rect 54290 37998 54292 38050
rect 54236 37986 54292 37998
rect 54012 37886 54014 37938
rect 54066 37886 54068 37938
rect 54012 37874 54068 37886
rect 51772 37826 51828 37838
rect 51772 37774 51774 37826
rect 51826 37774 51828 37826
rect 51772 37044 51828 37774
rect 53452 37826 53508 37838
rect 53452 37774 53454 37826
rect 53506 37774 53508 37826
rect 51772 36978 51828 36988
rect 52220 37378 52276 37390
rect 52220 37326 52222 37378
rect 52274 37326 52276 37378
rect 51884 36820 51940 36830
rect 51884 36482 51940 36764
rect 51884 36430 51886 36482
rect 51938 36430 51940 36482
rect 51884 36418 51940 36430
rect 51324 35980 51716 36036
rect 51996 36258 52052 36270
rect 51996 36206 51998 36258
rect 52050 36206 52052 36258
rect 50988 35924 51044 35934
rect 51324 35924 51380 35980
rect 50988 35830 51044 35868
rect 51100 35922 51380 35924
rect 51100 35870 51326 35922
rect 51378 35870 51380 35922
rect 51100 35868 51380 35870
rect 50708 35644 50932 35700
rect 50652 35606 50708 35644
rect 50988 35028 51044 35038
rect 51100 35028 51156 35868
rect 51324 35858 51380 35868
rect 51996 35812 52052 36206
rect 51212 35698 51268 35710
rect 51212 35646 51214 35698
rect 51266 35646 51268 35698
rect 51212 35588 51268 35646
rect 51212 35522 51268 35532
rect 51548 35698 51604 35710
rect 51548 35646 51550 35698
rect 51602 35646 51604 35698
rect 50988 35026 51156 35028
rect 50988 34974 50990 35026
rect 51042 34974 51156 35026
rect 50988 34972 51156 34974
rect 50988 34962 51044 34972
rect 50316 34802 50372 34814
rect 50316 34750 50318 34802
rect 50370 34750 50372 34802
rect 50316 34244 50372 34750
rect 51548 34804 51604 35646
rect 51996 35698 52052 35756
rect 51996 35646 51998 35698
rect 52050 35646 52052 35698
rect 51996 35634 52052 35646
rect 52220 35924 52276 37326
rect 52444 37266 52500 37278
rect 53228 37268 53284 37278
rect 52444 37214 52446 37266
rect 52498 37214 52500 37266
rect 52444 37044 52500 37214
rect 52444 36978 52500 36988
rect 53116 37266 53284 37268
rect 53116 37214 53230 37266
rect 53282 37214 53284 37266
rect 53116 37212 53284 37214
rect 53004 36820 53060 36830
rect 53116 36820 53172 37212
rect 53228 37202 53284 37212
rect 53060 36764 53172 36820
rect 53228 37044 53284 37054
rect 53004 36706 53060 36764
rect 53004 36654 53006 36706
rect 53058 36654 53060 36706
rect 53004 36642 53060 36654
rect 53228 36594 53284 36988
rect 53228 36542 53230 36594
rect 53282 36542 53284 36594
rect 53228 36530 53284 36542
rect 52220 35698 52276 35868
rect 52220 35646 52222 35698
rect 52274 35646 52276 35698
rect 52220 35634 52276 35646
rect 52668 36258 52724 36270
rect 52668 36206 52670 36258
rect 52722 36206 52724 36258
rect 52668 35586 52724 36206
rect 52668 35534 52670 35586
rect 52722 35534 52724 35586
rect 52668 35522 52724 35534
rect 53452 35586 53508 37774
rect 54460 37492 54516 37502
rect 54236 37156 54292 37166
rect 53788 37154 54292 37156
rect 53788 37102 54238 37154
rect 54290 37102 54292 37154
rect 53788 37100 54292 37102
rect 53676 35700 53732 35710
rect 53788 35700 53844 37100
rect 54236 37090 54292 37100
rect 54348 37156 54404 37166
rect 54348 36372 54404 37100
rect 54460 36706 54516 37436
rect 54572 37380 54628 37390
rect 54572 37044 54628 37324
rect 55132 37268 55188 38220
rect 55916 38052 55972 39340
rect 56028 38276 56084 40910
rect 57820 38724 57876 38734
rect 57708 38722 57876 38724
rect 57708 38670 57822 38722
rect 57874 38670 57876 38722
rect 57708 38668 57876 38670
rect 56028 38210 56084 38220
rect 57036 38612 57092 38622
rect 55916 37996 56868 38052
rect 55804 37938 55860 37950
rect 55804 37886 55806 37938
rect 55858 37886 55860 37938
rect 54572 36978 54628 36988
rect 54684 37266 55188 37268
rect 54684 37214 55134 37266
rect 55186 37214 55188 37266
rect 54684 37212 55188 37214
rect 54460 36654 54462 36706
rect 54514 36654 54516 36706
rect 54460 36642 54516 36654
rect 54572 36484 54628 36494
rect 54684 36484 54740 37212
rect 55132 37202 55188 37212
rect 55244 37826 55300 37838
rect 55244 37774 55246 37826
rect 55298 37774 55300 37826
rect 54572 36482 54740 36484
rect 54572 36430 54574 36482
rect 54626 36430 54740 36482
rect 54572 36428 54740 36430
rect 54908 37044 54964 37054
rect 54572 36418 54628 36428
rect 54460 36372 54516 36382
rect 54348 36370 54516 36372
rect 54348 36318 54462 36370
rect 54514 36318 54516 36370
rect 54348 36316 54516 36318
rect 54460 36306 54516 36316
rect 53676 35698 53788 35700
rect 53676 35646 53678 35698
rect 53730 35646 53788 35698
rect 53676 35644 53788 35646
rect 53676 35634 53732 35644
rect 53788 35606 53844 35644
rect 54236 35700 54292 35710
rect 53452 35534 53454 35586
rect 53506 35534 53508 35586
rect 52332 35476 52388 35486
rect 51548 34738 51604 34748
rect 51772 35474 52388 35476
rect 51772 35422 52334 35474
rect 52386 35422 52388 35474
rect 51772 35420 52388 35422
rect 50556 34524 50820 34534
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50556 34458 50820 34468
rect 50316 34178 50372 34188
rect 50764 34354 50820 34366
rect 50764 34302 50766 34354
rect 50818 34302 50820 34354
rect 50652 34132 50708 34142
rect 50652 34038 50708 34076
rect 50316 33460 50372 33470
rect 50316 33366 50372 33404
rect 50652 33348 50708 33358
rect 50764 33348 50820 34302
rect 50428 33346 50820 33348
rect 50428 33294 50654 33346
rect 50706 33294 50820 33346
rect 50428 33292 50820 33294
rect 51660 34244 51716 34254
rect 51660 34130 51716 34188
rect 51660 34078 51662 34130
rect 51714 34078 51716 34130
rect 51660 33348 51716 34078
rect 50428 32564 50484 33292
rect 50652 33282 50708 33292
rect 51660 33282 51716 33292
rect 51772 34242 51828 35420
rect 52332 35410 52388 35420
rect 52780 35364 52836 35374
rect 51772 34190 51774 34242
rect 51826 34190 51828 34242
rect 51772 33346 51828 34190
rect 52556 34692 52612 34702
rect 51772 33294 51774 33346
rect 51826 33294 51828 33346
rect 51100 33236 51156 33246
rect 50876 33234 51156 33236
rect 50876 33182 51102 33234
rect 51154 33182 51156 33234
rect 50876 33180 51156 33182
rect 50556 32956 50820 32966
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50556 32890 50820 32900
rect 50764 32564 50820 32574
rect 50876 32564 50932 33180
rect 51100 33170 51156 33180
rect 50428 32508 50708 32564
rect 50204 32050 50260 32060
rect 50428 32338 50484 32350
rect 50428 32286 50430 32338
rect 50482 32286 50484 32338
rect 50428 31220 50484 32286
rect 50652 31948 50708 32508
rect 50764 32562 50932 32564
rect 50764 32510 50766 32562
rect 50818 32510 50932 32562
rect 50764 32508 50932 32510
rect 50988 32564 51044 32574
rect 50764 32498 50820 32508
rect 50988 32470 51044 32508
rect 51772 32450 51828 33294
rect 51996 33348 52052 33358
rect 51996 33254 52052 33292
rect 51884 33124 51940 33134
rect 51884 32564 51940 33068
rect 51884 32470 51940 32508
rect 51772 32398 51774 32450
rect 51826 32398 51828 32450
rect 51772 32386 51828 32398
rect 50652 31892 50820 31948
rect 50764 31780 50820 31892
rect 50764 31686 50820 31724
rect 51548 31666 51604 31678
rect 51548 31614 51550 31666
rect 51602 31614 51604 31666
rect 50556 31388 50820 31398
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50556 31322 50820 31332
rect 50428 31164 50596 31220
rect 50092 31106 50148 31118
rect 50092 31054 50094 31106
rect 50146 31054 50148 31106
rect 50092 30996 50148 31054
rect 50092 30930 50148 30940
rect 50204 30996 50260 31006
rect 50428 30996 50484 31006
rect 50204 30994 50484 30996
rect 50204 30942 50206 30994
rect 50258 30942 50430 30994
rect 50482 30942 50484 30994
rect 50204 30940 50484 30942
rect 50204 30930 50260 30940
rect 50428 30930 50484 30940
rect 50092 30772 50148 30782
rect 50092 30678 50148 30716
rect 50540 30772 50596 31164
rect 51548 31108 51604 31614
rect 50876 31052 51604 31108
rect 50876 30994 50932 31052
rect 50876 30942 50878 30994
rect 50930 30942 50932 30994
rect 50876 30930 50932 30942
rect 51548 30994 51604 31052
rect 52444 31108 52500 31118
rect 52444 31014 52500 31052
rect 51548 30942 51550 30994
rect 51602 30942 51604 30994
rect 51548 30930 51604 30942
rect 52332 30994 52388 31006
rect 52332 30942 52334 30994
rect 52386 30942 52388 30994
rect 51100 30884 51156 30894
rect 51100 30790 51156 30828
rect 51324 30882 51380 30894
rect 51324 30830 51326 30882
rect 51378 30830 51380 30882
rect 50540 30706 50596 30716
rect 51324 30772 51380 30830
rect 51324 30706 51380 30716
rect 52332 30772 52388 30942
rect 52332 30706 52388 30716
rect 50556 29820 50820 29830
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50556 29754 50820 29764
rect 52108 29540 52164 29550
rect 52108 28532 52164 29484
rect 52556 28756 52612 34636
rect 52780 33572 52836 35308
rect 53004 35140 53060 35150
rect 53004 35138 53284 35140
rect 53004 35086 53006 35138
rect 53058 35086 53284 35138
rect 53004 35084 53284 35086
rect 53004 35074 53060 35084
rect 53228 34916 53284 35084
rect 53452 35028 53508 35534
rect 53564 35028 53620 35038
rect 53452 35026 53620 35028
rect 53452 34974 53566 35026
rect 53618 34974 53620 35026
rect 53452 34972 53620 34974
rect 53228 34860 53508 34916
rect 53004 34804 53060 34814
rect 53004 34710 53060 34748
rect 53116 34804 53172 34814
rect 53116 34802 53396 34804
rect 53116 34750 53118 34802
rect 53170 34750 53396 34802
rect 53116 34748 53396 34750
rect 53116 34738 53172 34748
rect 53340 34242 53396 34748
rect 53340 34190 53342 34242
rect 53394 34190 53396 34242
rect 53340 34178 53396 34190
rect 52780 33516 53396 33572
rect 52668 33236 52724 33246
rect 52668 33142 52724 33180
rect 52780 33234 52836 33516
rect 53340 33458 53396 33516
rect 53340 33406 53342 33458
rect 53394 33406 53396 33458
rect 53340 33394 53396 33406
rect 52780 33182 52782 33234
rect 52834 33182 52836 33234
rect 52780 33170 52836 33182
rect 52892 33348 52948 33358
rect 52892 32562 52948 33292
rect 53004 33124 53060 33134
rect 53004 33030 53060 33068
rect 52892 32510 52894 32562
rect 52946 32510 52948 32562
rect 52892 32498 52948 32510
rect 53452 31948 53508 34860
rect 53564 34132 53620 34972
rect 53788 34804 53844 34814
rect 53788 34710 53844 34748
rect 53788 34132 53844 34142
rect 53564 34130 53844 34132
rect 53564 34078 53790 34130
rect 53842 34078 53844 34130
rect 53564 34076 53844 34078
rect 53788 34066 53844 34076
rect 54236 34130 54292 35644
rect 54236 34078 54238 34130
rect 54290 34078 54292 34130
rect 54236 34066 54292 34078
rect 54796 33908 54852 33918
rect 54796 33814 54852 33852
rect 53564 32340 53620 32350
rect 53564 32338 53732 32340
rect 53564 32286 53566 32338
rect 53618 32286 53732 32338
rect 53564 32284 53732 32286
rect 53564 32274 53620 32284
rect 53676 31948 53732 32284
rect 53452 31892 53620 31948
rect 53676 31892 53956 31948
rect 53340 31668 53396 31678
rect 53564 31668 53620 31892
rect 53676 31668 53732 31678
rect 53564 31666 53732 31668
rect 53564 31614 53678 31666
rect 53730 31614 53732 31666
rect 53564 31612 53732 31614
rect 53340 31574 53396 31612
rect 53452 31554 53508 31566
rect 53452 31502 53454 31554
rect 53506 31502 53508 31554
rect 52556 28690 52612 28700
rect 52668 31108 52724 31118
rect 53452 31108 53508 31502
rect 53676 31556 53732 31612
rect 53676 31490 53732 31500
rect 53900 31666 53956 31892
rect 54572 31780 54628 31790
rect 54796 31780 54852 31790
rect 54572 31778 54796 31780
rect 54572 31726 54574 31778
rect 54626 31726 54796 31778
rect 54572 31724 54796 31726
rect 54572 31714 54628 31724
rect 54796 31714 54852 31724
rect 53900 31614 53902 31666
rect 53954 31614 53956 31666
rect 52108 28466 52164 28476
rect 50556 28252 50820 28262
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50556 28186 50820 28196
rect 49644 27570 49700 27580
rect 45500 26852 45668 26908
rect 45052 25566 45054 25618
rect 45106 25566 45108 25618
rect 45052 25554 45108 25566
rect 45388 26290 45444 26302
rect 45388 26238 45390 26290
rect 45442 26238 45444 26290
rect 45388 25396 45444 26238
rect 45500 25618 45556 26852
rect 46396 26850 46452 26862
rect 46396 26798 46398 26850
rect 46450 26798 46452 26850
rect 45500 25566 45502 25618
rect 45554 25566 45556 25618
rect 45500 25554 45556 25566
rect 46060 26178 46116 26190
rect 46060 26126 46062 26178
rect 46114 26126 46116 26178
rect 44940 25340 45220 25396
rect 44268 24894 44270 24946
rect 44322 24894 44324 24946
rect 44268 24882 44324 24894
rect 44492 25284 44548 25294
rect 44492 24722 44548 25228
rect 44492 24670 44494 24722
rect 44546 24670 44548 24722
rect 44492 24658 44548 24670
rect 44940 25172 44996 25182
rect 44940 23826 44996 25116
rect 45164 24724 45220 25340
rect 45388 25330 45444 25340
rect 45836 25396 45892 25406
rect 45836 25302 45892 25340
rect 46060 25172 46116 26126
rect 46284 25508 46340 25518
rect 46060 25106 46116 25116
rect 46172 25506 46340 25508
rect 46172 25454 46286 25506
rect 46338 25454 46340 25506
rect 46172 25452 46340 25454
rect 46172 25396 46228 25452
rect 46284 25442 46340 25452
rect 45164 23938 45220 24668
rect 45724 24164 45780 24174
rect 45164 23886 45166 23938
rect 45218 23886 45220 23938
rect 45164 23874 45220 23886
rect 45388 24162 45780 24164
rect 45388 24110 45726 24162
rect 45778 24110 45780 24162
rect 45388 24108 45780 24110
rect 44940 23774 44942 23826
rect 44994 23774 44996 23826
rect 44940 23762 44996 23774
rect 45388 23266 45444 24108
rect 45724 24098 45780 24108
rect 45612 23940 45668 23950
rect 45612 23846 45668 23884
rect 45724 23714 45780 23726
rect 45724 23662 45726 23714
rect 45778 23662 45780 23714
rect 45724 23492 45780 23662
rect 45724 23436 46116 23492
rect 45388 23214 45390 23266
rect 45442 23214 45444 23266
rect 45388 23202 45444 23214
rect 44604 23156 44660 23166
rect 44604 23062 44660 23100
rect 45724 23156 45780 23166
rect 44156 23042 44212 23054
rect 44156 22990 44158 23042
rect 44210 22990 44212 23042
rect 44156 22596 44212 22990
rect 44156 22530 44212 22540
rect 44044 22318 44046 22370
rect 44098 22318 44100 22370
rect 44044 22306 44100 22318
rect 45164 22372 45220 22382
rect 42588 22260 42644 22270
rect 42588 22148 42644 22204
rect 44156 22260 44212 22270
rect 42588 22092 42756 22148
rect 42588 21924 42644 21934
rect 42588 20802 42644 21868
rect 42588 20750 42590 20802
rect 42642 20750 42644 20802
rect 42588 20738 42644 20750
rect 42476 19842 42532 19852
rect 42252 19348 42308 19358
rect 42140 18452 42196 18462
rect 42140 18358 42196 18396
rect 41916 18172 42196 18228
rect 41804 17612 42084 17668
rect 41468 17556 41524 17566
rect 41356 17332 41412 17342
rect 41356 16884 41412 17276
rect 41244 16882 41412 16884
rect 41244 16830 41358 16882
rect 41410 16830 41412 16882
rect 41244 16828 41412 16830
rect 41132 16658 41188 16670
rect 41132 16606 41134 16658
rect 41186 16606 41188 16658
rect 41132 16324 41188 16606
rect 41132 16258 41188 16268
rect 41132 16100 41188 16110
rect 41244 16100 41300 16828
rect 41356 16818 41412 16828
rect 41356 16212 41412 16222
rect 41468 16212 41524 17500
rect 41804 17108 41860 17118
rect 41580 16884 41636 16894
rect 41580 16790 41636 16828
rect 41692 16772 41748 16782
rect 41692 16678 41748 16716
rect 41356 16210 41524 16212
rect 41356 16158 41358 16210
rect 41410 16158 41524 16210
rect 41356 16156 41524 16158
rect 41356 16146 41412 16156
rect 41132 16098 41300 16100
rect 41132 16046 41134 16098
rect 41186 16046 41300 16098
rect 41132 16044 41300 16046
rect 41804 16100 41860 17052
rect 41132 16034 41188 16044
rect 41468 15988 41524 15998
rect 41804 15988 41860 16044
rect 41468 15986 41860 15988
rect 41468 15934 41470 15986
rect 41522 15934 41860 15986
rect 41468 15932 41860 15934
rect 41468 15922 41524 15932
rect 41244 15876 41300 15886
rect 41020 15820 41244 15876
rect 41244 15782 41300 15820
rect 42028 15540 42084 17612
rect 42140 17442 42196 18172
rect 42140 17390 42142 17442
rect 42194 17390 42196 17442
rect 42140 16884 42196 17390
rect 42140 16818 42196 16828
rect 42252 16882 42308 19292
rect 42364 19346 42420 19358
rect 42364 19294 42366 19346
rect 42418 19294 42420 19346
rect 42364 18340 42420 19294
rect 42364 18274 42420 18284
rect 42252 16830 42254 16882
rect 42306 16830 42308 16882
rect 42252 16818 42308 16830
rect 42588 16212 42644 16222
rect 42588 16118 42644 16156
rect 42028 15474 42084 15484
rect 42140 16098 42196 16110
rect 42140 16046 42142 16098
rect 42194 16046 42196 16098
rect 42140 15538 42196 16046
rect 42476 16100 42532 16110
rect 42476 16006 42532 16044
rect 42700 16100 42756 22092
rect 43596 22146 43652 22158
rect 43596 22094 43598 22146
rect 43650 22094 43652 22146
rect 43596 21924 43652 22094
rect 43596 21858 43652 21868
rect 43820 21588 43876 21598
rect 43708 21474 43764 21486
rect 43708 21422 43710 21474
rect 43762 21422 43764 21474
rect 43036 21364 43092 21374
rect 43036 20690 43092 21308
rect 43036 20638 43038 20690
rect 43090 20638 43092 20690
rect 43036 20626 43092 20638
rect 43148 20802 43204 20814
rect 43148 20750 43150 20802
rect 43202 20750 43204 20802
rect 43148 20692 43204 20750
rect 43148 20626 43204 20636
rect 43708 20132 43764 21422
rect 43596 20076 43764 20132
rect 43820 21026 43876 21532
rect 43820 20974 43822 21026
rect 43874 20974 43876 21026
rect 42924 19908 42980 19918
rect 42924 19814 42980 19852
rect 42812 19348 42868 19358
rect 42812 19254 42868 19292
rect 43596 19348 43652 20076
rect 43708 19908 43764 19918
rect 43820 19908 43876 20974
rect 44156 21026 44212 22204
rect 45164 22258 45220 22316
rect 45164 22206 45166 22258
rect 45218 22206 45220 22258
rect 45164 22194 45220 22206
rect 45500 22260 45556 22270
rect 45500 22166 45556 22204
rect 44268 22146 44324 22158
rect 44268 22094 44270 22146
rect 44322 22094 44324 22146
rect 44268 21924 44324 22094
rect 44268 21858 44324 21868
rect 44828 22146 44884 22158
rect 44828 22094 44830 22146
rect 44882 22094 44884 22146
rect 44828 21924 44884 22094
rect 44156 20974 44158 21026
rect 44210 20974 44212 21026
rect 44156 20962 44212 20974
rect 44828 20802 44884 21868
rect 45276 20914 45332 20926
rect 45276 20862 45278 20914
rect 45330 20862 45332 20914
rect 45276 20804 45332 20862
rect 45724 20916 45780 23100
rect 46060 22370 46116 23436
rect 46172 23156 46228 25340
rect 46284 25284 46340 25294
rect 46396 25284 46452 26798
rect 48636 26852 48916 26908
rect 48188 26292 48244 26302
rect 48188 26178 48244 26236
rect 48188 26126 48190 26178
rect 48242 26126 48244 26178
rect 48188 26114 48244 26126
rect 46340 25228 46452 25284
rect 46284 25218 46340 25228
rect 46508 25172 46564 25182
rect 46396 25116 46508 25172
rect 46396 24834 46452 25116
rect 46508 25106 46564 25116
rect 46396 24782 46398 24834
rect 46450 24782 46452 24834
rect 46396 24770 46452 24782
rect 46508 24948 46564 24958
rect 46508 24722 46564 24892
rect 47852 24948 47908 24958
rect 47852 24854 47908 24892
rect 47516 24836 47572 24846
rect 47516 24742 47572 24780
rect 48636 24836 48692 26852
rect 50556 26684 50820 26694
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50556 26618 50820 26628
rect 49084 26516 49140 26526
rect 49084 26422 49140 26460
rect 48860 26292 48916 26302
rect 48860 26198 48916 26236
rect 52108 26292 52164 26302
rect 50556 25116 50820 25126
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50556 25050 50820 25060
rect 48636 24770 48692 24780
rect 46508 24670 46510 24722
rect 46562 24670 46564 24722
rect 46508 24658 46564 24670
rect 46956 24724 47012 24734
rect 46956 24630 47012 24668
rect 46844 24052 46900 24062
rect 47292 24052 47348 24062
rect 46844 24050 47348 24052
rect 46844 23998 46846 24050
rect 46898 23998 47294 24050
rect 47346 23998 47348 24050
rect 46844 23996 47348 23998
rect 46844 23986 46900 23996
rect 47292 23986 47348 23996
rect 46396 23828 46452 23838
rect 46396 23734 46452 23772
rect 46620 23828 46676 23838
rect 46620 23734 46676 23772
rect 46956 23826 47012 23838
rect 46956 23774 46958 23826
rect 47010 23774 47012 23826
rect 46172 23090 46228 23100
rect 46060 22318 46062 22370
rect 46114 22318 46116 22370
rect 46060 22306 46116 22318
rect 46284 23044 46340 23054
rect 46284 22258 46340 22988
rect 46396 22372 46452 22382
rect 46396 22278 46452 22316
rect 46844 22370 46900 22382
rect 46844 22318 46846 22370
rect 46898 22318 46900 22370
rect 46284 22206 46286 22258
rect 46338 22206 46340 22258
rect 46284 22194 46340 22206
rect 45836 22148 45892 22158
rect 45836 22146 46004 22148
rect 45836 22094 45838 22146
rect 45890 22094 46004 22146
rect 45836 22092 46004 22094
rect 45836 22082 45892 22092
rect 45836 20916 45892 20926
rect 45724 20914 45892 20916
rect 45724 20862 45838 20914
rect 45890 20862 45892 20914
rect 45724 20860 45892 20862
rect 45836 20850 45892 20860
rect 44828 20750 44830 20802
rect 44882 20750 44884 20802
rect 44828 20738 44884 20750
rect 45052 20748 45332 20804
rect 43708 19906 43876 19908
rect 43708 19854 43710 19906
rect 43762 19854 43876 19906
rect 43708 19852 43876 19854
rect 43708 19842 43764 19852
rect 43596 19282 43652 19292
rect 44268 19348 44324 19358
rect 44268 19254 44324 19292
rect 44828 19348 44884 19358
rect 44828 19234 44884 19292
rect 44828 19182 44830 19234
rect 44882 19182 44884 19234
rect 44828 19170 44884 19182
rect 43820 18564 43876 18574
rect 43708 18508 43820 18564
rect 43484 17444 43540 17454
rect 43036 17442 43540 17444
rect 43036 17390 43486 17442
rect 43538 17390 43540 17442
rect 43036 17388 43540 17390
rect 43036 16994 43092 17388
rect 43484 17378 43540 17388
rect 43036 16942 43038 16994
rect 43090 16942 43092 16994
rect 43036 16930 43092 16942
rect 43708 16212 43764 18508
rect 43820 18498 43876 18508
rect 44940 18452 44996 18462
rect 44940 18358 44996 18396
rect 45052 18116 45108 20748
rect 45836 20132 45892 20142
rect 45948 20132 46004 22092
rect 46620 21474 46676 21486
rect 46620 21422 46622 21474
rect 46674 21422 46676 21474
rect 46620 20804 46676 21422
rect 46844 20804 46900 22318
rect 46956 22372 47012 23774
rect 49756 23828 49812 23838
rect 47404 23716 47460 23726
rect 47404 23714 47684 23716
rect 47404 23662 47406 23714
rect 47458 23662 47684 23714
rect 47404 23660 47684 23662
rect 47404 23650 47460 23660
rect 47516 23044 47572 23054
rect 47516 22950 47572 22988
rect 47628 22482 47684 23660
rect 47964 23156 48020 23166
rect 47964 23062 48020 23100
rect 47628 22430 47630 22482
rect 47682 22430 47684 22482
rect 47628 22418 47684 22430
rect 49756 22484 49812 23772
rect 50556 23548 50820 23558
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50556 23482 50820 23492
rect 49756 22390 49812 22428
rect 46956 22306 47012 22316
rect 52108 22372 52164 26236
rect 52668 24948 52724 31052
rect 52892 31052 53508 31108
rect 52892 30994 52948 31052
rect 52892 30942 52894 30994
rect 52946 30942 52948 30994
rect 52892 30884 52948 30942
rect 52892 30818 52948 30828
rect 53900 30882 53956 31614
rect 54236 31668 54292 31678
rect 54236 31574 54292 31612
rect 54796 31554 54852 31566
rect 54796 31502 54798 31554
rect 54850 31502 54852 31554
rect 54348 30996 54404 31006
rect 54796 30996 54852 31502
rect 54348 30994 54852 30996
rect 54348 30942 54350 30994
rect 54402 30942 54852 30994
rect 54348 30940 54852 30942
rect 54348 30930 54404 30940
rect 53900 30830 53902 30882
rect 53954 30830 53956 30882
rect 53900 30818 53956 30830
rect 53564 30770 53620 30782
rect 53564 30718 53566 30770
rect 53618 30718 53620 30770
rect 53564 30100 53620 30718
rect 53564 30034 53620 30044
rect 54012 30212 54068 30222
rect 54012 29988 54068 30156
rect 54012 29922 54068 29932
rect 54908 27860 54964 36988
rect 55020 37042 55076 37054
rect 55020 36990 55022 37042
rect 55074 36990 55076 37042
rect 55020 36932 55076 36990
rect 55020 36866 55076 36876
rect 55020 35700 55076 35710
rect 55020 34914 55076 35644
rect 55020 34862 55022 34914
rect 55074 34862 55076 34914
rect 55020 34850 55076 34862
rect 55244 34916 55300 37774
rect 55804 37380 55860 37886
rect 55916 37938 55972 37996
rect 55916 37886 55918 37938
rect 55970 37886 55972 37938
rect 55916 37874 55972 37886
rect 56140 37828 56196 37838
rect 56140 37826 56532 37828
rect 56140 37774 56142 37826
rect 56194 37774 56532 37826
rect 56140 37772 56532 37774
rect 56140 37762 56196 37772
rect 55804 37314 55860 37324
rect 55356 37266 55412 37278
rect 55356 37214 55358 37266
rect 55410 37214 55412 37266
rect 55356 37156 55412 37214
rect 55356 37090 55412 37100
rect 56476 36370 56532 37772
rect 56588 37380 56644 37390
rect 56588 37286 56644 37324
rect 56812 37266 56868 37996
rect 56924 37828 56980 37838
rect 56924 37734 56980 37772
rect 56812 37214 56814 37266
rect 56866 37214 56868 37266
rect 56812 37202 56868 37214
rect 57036 37268 57092 38556
rect 57484 37940 57540 37950
rect 57708 37940 57764 38668
rect 57820 38658 57876 38668
rect 58268 38722 58324 38734
rect 58268 38670 58270 38722
rect 58322 38670 58324 38722
rect 58044 38050 58100 38062
rect 58044 37998 58046 38050
rect 58098 37998 58100 38050
rect 57484 37938 57764 37940
rect 57484 37886 57486 37938
rect 57538 37886 57764 37938
rect 57484 37884 57764 37886
rect 57820 37940 57876 37950
rect 57148 37826 57204 37838
rect 57148 37774 57150 37826
rect 57202 37774 57204 37826
rect 57148 37492 57204 37774
rect 57484 37716 57540 37884
rect 57820 37846 57876 37884
rect 57484 37650 57540 37660
rect 58044 37828 58100 37998
rect 57148 37426 57204 37436
rect 57820 37604 57876 37614
rect 57820 37490 57876 37548
rect 57820 37438 57822 37490
rect 57874 37438 57876 37490
rect 57820 37426 57876 37438
rect 57148 37268 57204 37278
rect 57036 37266 57204 37268
rect 57036 37214 57150 37266
rect 57202 37214 57204 37266
rect 57036 37212 57204 37214
rect 56476 36318 56478 36370
rect 56530 36318 56532 36370
rect 56476 36306 56532 36318
rect 56700 37154 56756 37166
rect 56700 37102 56702 37154
rect 56754 37102 56756 37154
rect 55692 36260 55748 36270
rect 56252 36260 56308 36270
rect 55692 36258 55860 36260
rect 55692 36206 55694 36258
rect 55746 36206 55860 36258
rect 55692 36204 55860 36206
rect 55692 36194 55748 36204
rect 55244 34850 55300 34860
rect 55692 34916 55748 34926
rect 55356 34690 55412 34702
rect 55356 34638 55358 34690
rect 55410 34638 55412 34690
rect 55356 34356 55412 34638
rect 55244 34300 55412 34356
rect 55244 33908 55300 34300
rect 55132 33906 55300 33908
rect 55132 33854 55246 33906
rect 55298 33854 55300 33906
rect 55132 33852 55300 33854
rect 55020 33236 55076 33246
rect 55132 33236 55188 33852
rect 55244 33842 55300 33852
rect 55356 34132 55412 34142
rect 55244 33348 55300 33358
rect 55356 33348 55412 34076
rect 55692 34132 55748 34860
rect 55692 34038 55748 34076
rect 55244 33346 55412 33348
rect 55244 33294 55246 33346
rect 55298 33294 55412 33346
rect 55244 33292 55412 33294
rect 55468 33908 55524 33918
rect 55468 33346 55524 33852
rect 55468 33294 55470 33346
rect 55522 33294 55524 33346
rect 55244 33282 55300 33292
rect 55468 33282 55524 33294
rect 55020 33234 55188 33236
rect 55020 33182 55022 33234
rect 55074 33182 55188 33234
rect 55020 33180 55188 33182
rect 55020 33170 55076 33180
rect 55356 33122 55412 33134
rect 55356 33070 55358 33122
rect 55410 33070 55412 33122
rect 55356 31948 55412 33070
rect 55132 31892 55412 31948
rect 55132 31780 55188 31892
rect 55132 31686 55188 31724
rect 55020 31556 55076 31566
rect 55020 31462 55076 31500
rect 55804 31444 55860 36204
rect 55804 31378 55860 31388
rect 55916 34244 55972 34254
rect 55580 30212 55636 30222
rect 55580 30118 55636 30156
rect 55916 29652 55972 34188
rect 55916 29586 55972 29596
rect 55244 28644 55300 28654
rect 55244 28550 55300 28588
rect 55580 28644 55636 28654
rect 55580 28550 55636 28588
rect 54908 27794 54964 27804
rect 56252 27188 56308 36204
rect 56588 35812 56644 35822
rect 56588 27524 56644 35756
rect 56700 33908 56756 37102
rect 57036 36594 57092 37212
rect 57148 37202 57204 37212
rect 58044 37044 58100 37772
rect 58156 37266 58212 37278
rect 58156 37214 58158 37266
rect 58210 37214 58212 37266
rect 58156 37156 58212 37214
rect 58268 37156 58324 38670
rect 58156 37100 58436 37156
rect 58044 36978 58100 36988
rect 57036 36542 57038 36594
rect 57090 36542 57092 36594
rect 57036 36530 57092 36542
rect 58156 36372 58212 36382
rect 58380 36372 58436 37100
rect 58156 36370 58324 36372
rect 58156 36318 58158 36370
rect 58210 36318 58324 36370
rect 58156 36316 58324 36318
rect 58156 36306 58212 36316
rect 57820 36260 57876 36270
rect 57820 36166 57876 36204
rect 57820 35812 57876 35822
rect 57820 35718 57876 35756
rect 57148 35700 57204 35710
rect 57148 35606 57204 35644
rect 58156 35698 58212 35710
rect 58156 35646 58158 35698
rect 58210 35646 58212 35698
rect 57596 35588 57652 35598
rect 58156 35588 58212 35646
rect 58268 35700 58324 36316
rect 58380 36306 58436 36316
rect 58268 35634 58324 35644
rect 57596 35586 58212 35588
rect 57596 35534 57598 35586
rect 57650 35534 58212 35586
rect 57596 35532 58212 35534
rect 57596 35522 57652 35532
rect 58156 35028 58212 35532
rect 58156 34962 58212 34972
rect 58156 34802 58212 34814
rect 58156 34750 58158 34802
rect 58210 34750 58212 34802
rect 57596 34690 57652 34702
rect 57596 34638 57598 34690
rect 57650 34638 57652 34690
rect 57596 34356 57652 34638
rect 57820 34692 57876 34702
rect 57820 34598 57876 34636
rect 57596 34290 57652 34300
rect 58156 34356 58212 34750
rect 58156 34290 58212 34300
rect 57820 34244 57876 34254
rect 57820 34150 57876 34188
rect 58156 34130 58212 34142
rect 58156 34078 58158 34130
rect 58210 34078 58212 34130
rect 57596 34020 57652 34030
rect 58156 34020 58212 34078
rect 57596 34018 58212 34020
rect 57596 33966 57598 34018
rect 57650 33966 58212 34018
rect 57596 33964 58212 33966
rect 57596 33954 57652 33964
rect 56700 33842 56756 33852
rect 58156 33684 58212 33964
rect 58156 33618 58212 33628
rect 58156 33234 58212 33246
rect 58156 33182 58158 33234
rect 58210 33182 58212 33234
rect 57596 33122 57652 33134
rect 57820 33124 57876 33134
rect 57596 33070 57598 33122
rect 57650 33070 57652 33122
rect 57596 33012 57652 33070
rect 57596 32946 57652 32956
rect 57708 33122 57876 33124
rect 57708 33070 57822 33122
rect 57874 33070 57876 33122
rect 57708 33068 57876 33070
rect 57148 32450 57204 32462
rect 57148 32398 57150 32450
rect 57202 32398 57204 32450
rect 57148 32340 57204 32398
rect 57148 32274 57204 32284
rect 57596 32450 57652 32462
rect 57596 32398 57598 32450
rect 57650 32398 57652 32450
rect 57596 31780 57652 32398
rect 57708 32004 57764 33068
rect 57820 33058 57876 33068
rect 58156 33012 58212 33182
rect 58156 32946 58212 32956
rect 57820 32676 57876 32686
rect 57820 32582 57876 32620
rect 58156 32562 58212 32574
rect 58156 32510 58158 32562
rect 58210 32510 58212 32562
rect 58156 32340 58212 32510
rect 58156 32274 58212 32284
rect 57708 31938 57764 31948
rect 57596 31724 57988 31780
rect 56924 31668 56980 31678
rect 56924 31574 56980 31612
rect 57484 31668 57540 31678
rect 57484 31574 57540 31612
rect 57148 31554 57204 31566
rect 57148 31502 57150 31554
rect 57202 31502 57204 31554
rect 57148 30324 57204 31502
rect 57820 31556 57876 31566
rect 57932 31556 57988 31724
rect 58156 31556 58212 31566
rect 57932 31554 58324 31556
rect 57932 31502 58158 31554
rect 58210 31502 58324 31554
rect 57932 31500 58324 31502
rect 57820 31462 57876 31500
rect 58156 31490 58212 31500
rect 57820 31108 57876 31118
rect 57820 31014 57876 31052
rect 58156 30994 58212 31006
rect 58156 30942 58158 30994
rect 58210 30942 58212 30994
rect 57596 30884 57652 30894
rect 58156 30884 58212 30942
rect 58268 30996 58324 31500
rect 58380 30996 58436 31006
rect 58268 30940 58380 30996
rect 58380 30930 58436 30940
rect 57596 30882 58212 30884
rect 57596 30830 57598 30882
rect 57650 30830 58212 30882
rect 57596 30828 58212 30830
rect 57596 30818 57652 30828
rect 57148 30258 57204 30268
rect 58156 30324 58212 30828
rect 58156 30258 58212 30268
rect 57260 30098 57316 30110
rect 57260 30046 57262 30098
rect 57314 30046 57316 30098
rect 57260 28980 57316 30046
rect 57596 29652 57652 29662
rect 57596 29558 57652 29596
rect 58156 29652 58212 29662
rect 57820 29540 57876 29550
rect 57820 29446 57876 29484
rect 58156 29538 58212 29596
rect 58156 29486 58158 29538
rect 58210 29486 58212 29538
rect 58156 29474 58212 29486
rect 57260 28914 57316 28924
rect 57932 28754 57988 28766
rect 57932 28702 57934 28754
rect 57986 28702 57988 28754
rect 57932 28308 57988 28702
rect 57932 28242 57988 28252
rect 57820 27970 57876 27982
rect 57820 27918 57822 27970
rect 57874 27918 57876 27970
rect 57596 27746 57652 27758
rect 57596 27694 57598 27746
rect 57650 27694 57652 27746
rect 57596 27636 57652 27694
rect 57596 27570 57652 27580
rect 56588 27458 56644 27468
rect 57820 27300 57876 27918
rect 58156 27858 58212 27870
rect 58156 27806 58158 27858
rect 58210 27806 58212 27858
rect 58156 27636 58212 27806
rect 58156 27570 58212 27580
rect 57820 27234 57876 27244
rect 56252 27122 56308 27132
rect 57932 27186 57988 27198
rect 57932 27134 57934 27186
rect 57986 27134 57988 27186
rect 55580 27074 55636 27086
rect 55580 27022 55582 27074
rect 55634 27022 55636 27074
rect 55580 26516 55636 27022
rect 55580 26450 55636 26460
rect 57596 26852 57652 26862
rect 57596 26514 57652 26796
rect 57596 26462 57598 26514
rect 57650 26462 57652 26514
rect 57596 26450 57652 26462
rect 57820 26402 57876 26414
rect 57820 26350 57822 26402
rect 57874 26350 57876 26402
rect 55580 25956 55636 25966
rect 52668 24882 52724 24892
rect 55132 25620 55188 25630
rect 53452 24722 53508 24734
rect 53452 24670 53454 24722
rect 53506 24670 53508 24722
rect 53452 24388 53508 24670
rect 53452 24322 53508 24332
rect 55132 24052 55188 25564
rect 55580 25506 55636 25900
rect 55580 25454 55582 25506
rect 55634 25454 55636 25506
rect 55580 25442 55636 25454
rect 57820 25284 57876 26350
rect 57932 26292 57988 27134
rect 58156 26852 58212 26862
rect 58156 26402 58212 26796
rect 58156 26350 58158 26402
rect 58210 26350 58212 26402
rect 58156 26338 58212 26350
rect 57932 26226 57988 26236
rect 57932 25620 57988 25630
rect 57932 25526 57988 25564
rect 57820 25218 57876 25228
rect 57932 24948 57988 24958
rect 55356 24500 55412 24510
rect 55356 24406 55412 24444
rect 57932 24162 57988 24892
rect 57932 24110 57934 24162
rect 57986 24110 57988 24162
rect 57932 24098 57988 24110
rect 55356 24052 55412 24062
rect 55132 24050 55636 24052
rect 55132 23998 55358 24050
rect 55410 23998 55636 24050
rect 55132 23996 55636 23998
rect 55356 23958 55412 23996
rect 55580 23938 55636 23996
rect 55580 23886 55582 23938
rect 55634 23886 55636 23938
rect 55580 23874 55636 23886
rect 57932 23492 57988 23502
rect 53452 23154 53508 23166
rect 53452 23102 53454 23154
rect 53506 23102 53508 23154
rect 53452 23044 53508 23102
rect 53452 22978 53508 22988
rect 55356 22932 55412 22942
rect 55356 22838 55412 22876
rect 52108 22306 52164 22316
rect 52668 22708 52724 22718
rect 52668 22370 52724 22652
rect 57932 22594 57988 23436
rect 57932 22542 57934 22594
rect 57986 22542 57988 22594
rect 57932 22530 57988 22542
rect 52668 22318 52670 22370
rect 52722 22318 52724 22370
rect 52668 22306 52724 22318
rect 53564 22484 53620 22494
rect 50556 21980 50820 21990
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50556 21914 50820 21924
rect 53452 21588 53508 21598
rect 53452 21494 53508 21532
rect 49756 20916 49812 20926
rect 49644 20914 49812 20916
rect 49644 20862 49758 20914
rect 49810 20862 49812 20914
rect 49644 20860 49812 20862
rect 46620 20802 47012 20804
rect 46620 20750 46846 20802
rect 46898 20750 47012 20802
rect 46620 20748 47012 20750
rect 45836 20130 46004 20132
rect 45836 20078 45838 20130
rect 45890 20078 46004 20130
rect 45836 20076 46004 20078
rect 46508 20580 46564 20590
rect 46620 20580 46676 20748
rect 46844 20738 46900 20748
rect 46508 20578 46676 20580
rect 46508 20526 46510 20578
rect 46562 20526 46676 20578
rect 46508 20524 46676 20526
rect 45836 20066 45892 20076
rect 46508 20018 46564 20524
rect 46508 19966 46510 20018
rect 46562 19966 46564 20018
rect 46508 19348 46564 19966
rect 46508 19282 46564 19292
rect 46956 20132 47012 20748
rect 47628 20690 47684 20702
rect 47628 20638 47630 20690
rect 47682 20638 47684 20690
rect 47628 20242 47684 20638
rect 47628 20190 47630 20242
rect 47682 20190 47684 20242
rect 47628 20178 47684 20190
rect 47068 20132 47124 20142
rect 46956 20130 47124 20132
rect 46956 20078 47070 20130
rect 47122 20078 47124 20130
rect 46956 20076 47124 20078
rect 45612 19124 45668 19134
rect 45164 19122 45668 19124
rect 45164 19070 45614 19122
rect 45666 19070 45668 19122
rect 45164 19068 45668 19070
rect 45164 18674 45220 19068
rect 45612 19058 45668 19068
rect 45164 18622 45166 18674
rect 45218 18622 45220 18674
rect 45164 18610 45220 18622
rect 45724 18562 45780 18574
rect 45724 18510 45726 18562
rect 45778 18510 45780 18562
rect 45164 18116 45220 18126
rect 45052 18060 45164 18116
rect 45164 18050 45220 18060
rect 45612 17780 45668 17790
rect 45276 17668 45332 17678
rect 45164 17612 45276 17668
rect 43820 17556 43876 17566
rect 44940 17556 44996 17566
rect 43820 17554 44996 17556
rect 43820 17502 43822 17554
rect 43874 17502 44942 17554
rect 44994 17502 44996 17554
rect 43820 17500 44996 17502
rect 43820 17490 43876 17500
rect 44940 17490 44996 17500
rect 43820 16884 43876 16894
rect 43820 16660 43876 16828
rect 45164 16770 45220 17612
rect 45276 17574 45332 17612
rect 45612 17106 45668 17724
rect 45612 17054 45614 17106
rect 45666 17054 45668 17106
rect 45612 17042 45668 17054
rect 45164 16718 45166 16770
rect 45218 16718 45220 16770
rect 45164 16706 45220 16718
rect 45724 16772 45780 18510
rect 45948 18450 46004 18462
rect 45948 18398 45950 18450
rect 46002 18398 46004 18450
rect 45948 18116 46004 18398
rect 46732 18452 46788 18462
rect 46732 18358 46788 18396
rect 46396 18340 46452 18350
rect 46396 18246 46452 18284
rect 45948 17666 46004 18060
rect 46956 17780 47012 20076
rect 47068 20066 47124 20076
rect 48972 20130 49028 20142
rect 48972 20078 48974 20130
rect 49026 20078 49028 20130
rect 47964 20020 48020 20030
rect 47964 19926 48020 19964
rect 48860 20018 48916 20030
rect 48860 19966 48862 20018
rect 48914 19966 48916 20018
rect 48188 19908 48244 19918
rect 47740 19346 47796 19358
rect 47740 19294 47742 19346
rect 47794 19294 47796 19346
rect 47740 18452 47796 19294
rect 47740 18386 47796 18396
rect 48076 17780 48132 17790
rect 47012 17724 47348 17780
rect 46956 17686 47012 17724
rect 45948 17614 45950 17666
rect 46002 17614 46004 17666
rect 45948 17602 46004 17614
rect 47292 17666 47348 17724
rect 48076 17686 48132 17724
rect 47292 17614 47294 17666
rect 47346 17614 47348 17666
rect 47292 17602 47348 17614
rect 45836 17556 45892 17566
rect 45836 17462 45892 17500
rect 45724 16706 45780 16716
rect 46508 17220 46564 17230
rect 43820 16594 43876 16604
rect 43708 16146 43764 16156
rect 46508 16210 46564 17164
rect 46508 16158 46510 16210
rect 46562 16158 46564 16210
rect 46508 16146 46564 16158
rect 42700 16006 42756 16044
rect 47068 16098 47124 16110
rect 47068 16046 47070 16098
rect 47122 16046 47124 16098
rect 45276 15986 45332 15998
rect 45276 15934 45278 15986
rect 45330 15934 45332 15986
rect 42140 15486 42142 15538
rect 42194 15486 42196 15538
rect 42140 15474 42196 15486
rect 43708 15876 43764 15886
rect 41132 15428 41188 15438
rect 41132 15334 41188 15372
rect 42476 15426 42532 15438
rect 42476 15374 42478 15426
rect 42530 15374 42532 15426
rect 41356 15314 41412 15326
rect 41356 15262 41358 15314
rect 41410 15262 41412 15314
rect 41356 15204 41412 15262
rect 41580 15316 41636 15326
rect 41580 15222 41636 15260
rect 41804 15316 41860 15326
rect 42028 15316 42084 15326
rect 41804 15314 42084 15316
rect 41804 15262 41806 15314
rect 41858 15262 42030 15314
rect 42082 15262 42084 15314
rect 41804 15260 42084 15262
rect 41804 15250 41860 15260
rect 41356 15138 41412 15148
rect 40908 14802 40964 14812
rect 42028 14754 42084 15260
rect 42252 15314 42308 15326
rect 42252 15262 42254 15314
rect 42306 15262 42308 15314
rect 42252 15204 42308 15262
rect 42476 15316 42532 15374
rect 43708 15426 43764 15820
rect 43708 15374 43710 15426
rect 43762 15374 43764 15426
rect 43708 15362 43764 15374
rect 45052 15874 45108 15886
rect 45052 15822 45054 15874
rect 45106 15822 45108 15874
rect 42476 15250 42532 15260
rect 44380 15314 44436 15326
rect 44380 15262 44382 15314
rect 44434 15262 44436 15314
rect 42252 15138 42308 15148
rect 42028 14702 42030 14754
rect 42082 14702 42084 14754
rect 42028 14690 42084 14702
rect 41468 14642 41524 14654
rect 41468 14590 41470 14642
rect 41522 14590 41524 14642
rect 40908 14532 40964 14542
rect 41356 14532 41412 14542
rect 40908 14530 41412 14532
rect 40908 14478 40910 14530
rect 40962 14478 41358 14530
rect 41410 14478 41412 14530
rect 40908 14476 41412 14478
rect 40908 14466 40964 14476
rect 41356 14466 41412 14476
rect 40572 14418 40628 14430
rect 40572 14366 40574 14418
rect 40626 14366 40628 14418
rect 40572 14196 40628 14366
rect 40572 14130 40628 14140
rect 40684 14306 40740 14318
rect 40684 14254 40686 14306
rect 40738 14254 40740 14306
rect 40236 13806 40238 13858
rect 40290 13806 40292 13858
rect 40236 13794 40292 13806
rect 40124 12236 40292 12292
rect 40012 11902 40014 11954
rect 40066 11902 40068 11954
rect 40012 11890 40068 11902
rect 40236 11732 40292 12236
rect 40684 11956 40740 14254
rect 41244 13972 41300 13982
rect 41468 13972 41524 14590
rect 44380 14532 44436 15262
rect 45052 15316 45108 15822
rect 45052 15250 45108 15260
rect 45164 15874 45220 15886
rect 45164 15822 45166 15874
rect 45218 15822 45220 15874
rect 44380 14466 44436 14476
rect 45164 14530 45220 15822
rect 45276 15204 45332 15934
rect 47068 15540 47124 16046
rect 48076 15988 48132 15998
rect 47964 15986 48132 15988
rect 47964 15934 48078 15986
rect 48130 15934 48132 15986
rect 47964 15932 48132 15934
rect 46956 15484 47124 15540
rect 47180 15540 47236 15550
rect 47964 15540 48020 15932
rect 48076 15922 48132 15932
rect 47180 15538 48020 15540
rect 47180 15486 47182 15538
rect 47234 15486 48020 15538
rect 47180 15484 48020 15486
rect 46396 15426 46452 15438
rect 46396 15374 46398 15426
rect 46450 15374 46452 15426
rect 45276 15138 45332 15148
rect 45388 15316 45444 15326
rect 45388 14980 45444 15260
rect 46172 15314 46228 15326
rect 46172 15262 46174 15314
rect 46226 15262 46228 15314
rect 45164 14478 45166 14530
rect 45218 14478 45220 14530
rect 45164 14466 45220 14478
rect 45276 14924 45444 14980
rect 45724 15204 45780 15214
rect 41244 13970 41524 13972
rect 41244 13918 41246 13970
rect 41298 13918 41524 13970
rect 41244 13916 41524 13918
rect 41244 13906 41300 13916
rect 41020 13858 41076 13870
rect 41020 13806 41022 13858
rect 41074 13806 41076 13858
rect 40908 13748 40964 13758
rect 40908 13654 40964 13692
rect 41020 13636 41076 13806
rect 45052 13860 45108 13870
rect 45276 13860 45332 14924
rect 45612 14532 45668 14542
rect 45612 14438 45668 14476
rect 45052 13858 45332 13860
rect 45052 13806 45054 13858
rect 45106 13806 45332 13858
rect 45052 13804 45332 13806
rect 45052 13794 45108 13804
rect 44604 13746 44660 13758
rect 44604 13694 44606 13746
rect 44658 13694 44660 13746
rect 41020 13570 41076 13580
rect 41580 13636 41636 13646
rect 41580 13542 41636 13580
rect 43036 13634 43092 13646
rect 43036 13582 43038 13634
rect 43090 13582 43092 13634
rect 42700 12964 42756 12974
rect 43036 12964 43092 13582
rect 44268 13634 44324 13646
rect 44268 13582 44270 13634
rect 44322 13582 44324 13634
rect 42700 12962 43036 12964
rect 42700 12910 42702 12962
rect 42754 12910 43036 12962
rect 42700 12908 43036 12910
rect 41692 12850 41748 12862
rect 41692 12798 41694 12850
rect 41746 12798 41748 12850
rect 41356 12738 41412 12750
rect 41356 12686 41358 12738
rect 41410 12686 41412 12738
rect 41356 12628 41412 12686
rect 41580 12738 41636 12750
rect 41580 12686 41582 12738
rect 41634 12686 41636 12738
rect 41468 12628 41524 12638
rect 41356 12572 41468 12628
rect 41468 12562 41524 12572
rect 41580 12068 41636 12686
rect 41580 12002 41636 12012
rect 41692 12292 41748 12798
rect 42476 12850 42532 12862
rect 42476 12798 42478 12850
rect 42530 12798 42532 12850
rect 42476 12628 42532 12798
rect 42476 12562 42532 12572
rect 40012 11676 40292 11732
rect 40572 11900 40740 11956
rect 39900 11396 39956 11406
rect 39788 11394 39956 11396
rect 39788 11342 39902 11394
rect 39954 11342 39956 11394
rect 39788 11340 39956 11342
rect 39564 11282 39620 11340
rect 39900 11330 39956 11340
rect 39564 11230 39566 11282
rect 39618 11230 39620 11282
rect 39564 11218 39620 11230
rect 39676 11284 39732 11294
rect 39676 11190 39732 11228
rect 39900 10836 39956 10846
rect 39452 10834 39956 10836
rect 39452 10782 39902 10834
rect 39954 10782 39956 10834
rect 39452 10780 39956 10782
rect 39900 10770 39956 10780
rect 39116 10724 39172 10734
rect 39116 10630 39172 10668
rect 39340 10612 39396 10622
rect 39340 10518 39396 10556
rect 38668 9774 38670 9826
rect 38722 9774 38724 9826
rect 38220 9042 38276 9054
rect 38220 8990 38222 9042
rect 38274 8990 38276 9042
rect 38220 8260 38276 8990
rect 38220 8194 38276 8204
rect 38444 8820 38500 8830
rect 37772 8146 37828 8158
rect 37772 8094 37774 8146
rect 37826 8094 37828 8146
rect 37772 6692 37828 8094
rect 37884 8034 37940 8046
rect 37884 7982 37886 8034
rect 37938 7982 37940 8034
rect 37884 6916 37940 7982
rect 38108 8034 38164 8046
rect 38108 7982 38110 8034
rect 38162 7982 38164 8034
rect 38108 7474 38164 7982
rect 38108 7422 38110 7474
rect 38162 7422 38164 7474
rect 38108 7410 38164 7422
rect 38332 7476 38388 7486
rect 38332 7362 38388 7420
rect 38332 7310 38334 7362
rect 38386 7310 38388 7362
rect 38332 7298 38388 7310
rect 37884 6914 38276 6916
rect 37884 6862 37886 6914
rect 37938 6862 38276 6914
rect 37884 6860 38276 6862
rect 37884 6850 37940 6860
rect 37772 6626 37828 6636
rect 38108 6692 38164 6702
rect 38108 6598 38164 6636
rect 37660 6066 37716 6076
rect 37996 6580 38052 6590
rect 37212 6020 37268 6030
rect 37100 5794 37156 5806
rect 37100 5742 37102 5794
rect 37154 5742 37156 5794
rect 37100 5348 37156 5742
rect 37100 5282 37156 5292
rect 37212 5124 37268 5964
rect 37548 6018 37604 6030
rect 37548 5966 37550 6018
rect 37602 5966 37604 6018
rect 37548 5460 37604 5966
rect 37772 5908 37828 5918
rect 37548 5394 37604 5404
rect 37660 5572 37716 5582
rect 37212 5030 37268 5068
rect 37660 5124 37716 5516
rect 37660 5030 37716 5068
rect 36988 4958 36990 5010
rect 37042 4958 37044 5010
rect 36988 4946 37044 4958
rect 37772 5012 37828 5852
rect 37772 4946 37828 4956
rect 37884 5348 37940 5358
rect 37548 4900 37604 4910
rect 36764 4788 36820 4798
rect 36652 4732 36764 4788
rect 36764 4722 36820 4732
rect 37212 4450 37268 4462
rect 37212 4398 37214 4450
rect 37266 4398 37268 4450
rect 36988 4340 37044 4350
rect 36988 4246 37044 4284
rect 36316 4004 36372 4014
rect 36204 3668 36260 3678
rect 36204 3574 36260 3612
rect 36316 800 36372 3948
rect 37212 3780 37268 4398
rect 37212 3714 37268 3724
rect 37436 4226 37492 4238
rect 37436 4174 37438 4226
rect 37490 4174 37492 4226
rect 37436 3780 37492 4174
rect 37548 4226 37604 4844
rect 37884 4338 37940 5292
rect 37996 5010 38052 6524
rect 38220 6578 38276 6860
rect 38220 6526 38222 6578
rect 38274 6526 38276 6578
rect 38220 6514 38276 6526
rect 38332 6804 38388 6814
rect 37996 4958 37998 5010
rect 38050 4958 38052 5010
rect 37996 4946 38052 4958
rect 38108 6468 38164 6478
rect 37884 4286 37886 4338
rect 37938 4286 37940 4338
rect 37884 4274 37940 4286
rect 37548 4174 37550 4226
rect 37602 4174 37604 4226
rect 37548 4162 37604 4174
rect 37436 3714 37492 3724
rect 36988 3556 37044 3566
rect 36988 800 37044 3500
rect 38108 3554 38164 6412
rect 38220 5794 38276 5806
rect 38220 5742 38222 5794
rect 38274 5742 38276 5794
rect 38220 5236 38276 5742
rect 38220 4564 38276 5180
rect 38220 4498 38276 4508
rect 38108 3502 38110 3554
rect 38162 3502 38164 3554
rect 38108 3490 38164 3502
rect 37660 924 37940 980
rect 37660 800 37716 924
rect 0 0 112 800
rect 672 0 784 800
rect 1344 0 1456 800
rect 2016 0 2128 800
rect 2688 0 2800 800
rect 3360 0 3472 800
rect 4032 0 4144 800
rect 4704 0 4816 800
rect 5376 0 5488 800
rect 6048 0 6160 800
rect 6720 0 6832 800
rect 7392 0 7504 800
rect 8064 0 8176 800
rect 8736 0 8848 800
rect 9408 0 9520 800
rect 10080 0 10192 800
rect 14112 0 14224 800
rect 21504 0 21616 800
rect 25536 0 25648 800
rect 26208 0 26320 800
rect 26880 0 26992 800
rect 27552 0 27664 800
rect 28224 0 28336 800
rect 28896 0 29008 800
rect 29568 0 29680 800
rect 30240 0 30352 800
rect 30912 0 31024 800
rect 31584 0 31696 800
rect 32256 0 32368 800
rect 32928 0 33040 800
rect 33600 0 33712 800
rect 34272 0 34384 800
rect 34944 0 35056 800
rect 35616 0 35728 800
rect 36288 0 36400 800
rect 36960 0 37072 800
rect 37632 0 37744 800
rect 37884 756 37940 924
rect 38332 756 38388 6748
rect 38444 6580 38500 8764
rect 38668 7364 38724 9774
rect 38780 10220 38948 10276
rect 38780 9044 38836 10220
rect 39452 10052 39508 10062
rect 39340 9996 39452 10052
rect 38892 9714 38948 9726
rect 38892 9662 38894 9714
rect 38946 9662 38948 9714
rect 38892 9268 38948 9662
rect 38892 9174 38948 9212
rect 39340 9602 39396 9996
rect 39452 9986 39508 9996
rect 39900 9828 39956 9838
rect 40012 9828 40068 11676
rect 40236 11394 40292 11406
rect 40236 11342 40238 11394
rect 40290 11342 40292 11394
rect 40124 11172 40180 11182
rect 40124 11078 40180 11116
rect 40236 11060 40292 11342
rect 40236 10994 40292 11004
rect 40572 11282 40628 11900
rect 40684 11508 40740 11518
rect 40684 11506 41188 11508
rect 40684 11454 40686 11506
rect 40738 11454 41188 11506
rect 40684 11452 41188 11454
rect 40684 11442 40740 11452
rect 41132 11396 41188 11452
rect 41580 11506 41636 11518
rect 41580 11454 41582 11506
rect 41634 11454 41636 11506
rect 41356 11396 41412 11406
rect 41132 11394 41412 11396
rect 41132 11342 41358 11394
rect 41410 11342 41412 11394
rect 41132 11340 41412 11342
rect 41356 11330 41412 11340
rect 40572 11230 40574 11282
rect 40626 11230 40628 11282
rect 40572 10724 40628 11230
rect 40572 10658 40628 10668
rect 41020 10722 41076 10734
rect 41020 10670 41022 10722
rect 41074 10670 41076 10722
rect 40236 10610 40292 10622
rect 40236 10558 40238 10610
rect 40290 10558 40292 10610
rect 39956 9772 40068 9828
rect 40124 10388 40180 10398
rect 39900 9734 39956 9772
rect 40124 9716 40180 10332
rect 40236 9828 40292 10558
rect 40908 10610 40964 10622
rect 40908 10558 40910 10610
rect 40962 10558 40964 10610
rect 40908 10388 40964 10558
rect 41020 10612 41076 10670
rect 41580 10722 41636 11454
rect 41580 10670 41582 10722
rect 41634 10670 41636 10722
rect 41020 10546 41076 10556
rect 41244 10612 41300 10622
rect 41468 10612 41524 10622
rect 41244 10610 41524 10612
rect 41244 10558 41246 10610
rect 41298 10558 41470 10610
rect 41522 10558 41524 10610
rect 41244 10556 41524 10558
rect 41244 10546 41300 10556
rect 41468 10546 41524 10556
rect 40908 10322 40964 10332
rect 41580 10276 41636 10670
rect 41580 10210 41636 10220
rect 40908 9940 40964 9950
rect 40796 9828 40852 9838
rect 40236 9772 40404 9828
rect 40012 9714 40180 9716
rect 40012 9662 40126 9714
rect 40178 9662 40180 9714
rect 40012 9660 40180 9662
rect 40012 9604 40068 9660
rect 40124 9650 40180 9660
rect 39340 9550 39342 9602
rect 39394 9550 39396 9602
rect 39340 9268 39396 9550
rect 39340 9202 39396 9212
rect 39788 9548 40068 9604
rect 40236 9604 40292 9614
rect 38780 8978 38836 8988
rect 39228 9042 39284 9054
rect 39228 8990 39230 9042
rect 39282 8990 39284 9042
rect 39228 8428 39284 8990
rect 39788 9042 39844 9548
rect 40124 9268 40180 9278
rect 40124 9154 40180 9212
rect 40236 9266 40292 9548
rect 40348 9492 40404 9772
rect 40348 9426 40404 9436
rect 40460 9826 40852 9828
rect 40460 9774 40798 9826
rect 40850 9774 40852 9826
rect 40460 9772 40852 9774
rect 40236 9214 40238 9266
rect 40290 9214 40292 9266
rect 40236 9202 40292 9214
rect 40460 9266 40516 9772
rect 40796 9762 40852 9772
rect 40908 9602 40964 9884
rect 41692 9714 41748 12236
rect 42028 12178 42084 12190
rect 42028 12126 42030 12178
rect 42082 12126 42084 12178
rect 42028 11396 42084 12126
rect 42476 12180 42532 12190
rect 42476 12066 42532 12124
rect 42476 12014 42478 12066
rect 42530 12014 42532 12066
rect 42476 12002 42532 12014
rect 42588 12180 42644 12190
rect 42700 12180 42756 12908
rect 43036 12870 43092 12908
rect 43148 13524 43204 13534
rect 43148 12740 43204 13468
rect 42588 12178 42756 12180
rect 42588 12126 42590 12178
rect 42642 12126 42756 12178
rect 42588 12124 42756 12126
rect 43036 12684 43204 12740
rect 43260 13522 43316 13534
rect 43260 13470 43262 13522
rect 43314 13470 43316 13522
rect 42588 11844 42644 12124
rect 42924 11956 42980 11966
rect 42924 11862 42980 11900
rect 42252 11788 42644 11844
rect 42252 11618 42308 11788
rect 42252 11566 42254 11618
rect 42306 11566 42308 11618
rect 42252 11554 42308 11566
rect 41916 11394 42084 11396
rect 41916 11342 42030 11394
rect 42082 11342 42084 11394
rect 41916 11340 42084 11342
rect 41804 10836 41860 10846
rect 41916 10836 41972 11340
rect 42028 11330 42084 11340
rect 41804 10834 41972 10836
rect 41804 10782 41806 10834
rect 41858 10782 41972 10834
rect 41804 10780 41972 10782
rect 42588 10948 42644 10958
rect 41804 10770 41860 10780
rect 42588 9938 42644 10892
rect 43036 10498 43092 12684
rect 43260 12180 43316 13470
rect 43260 12114 43316 12124
rect 43596 13522 43652 13534
rect 43596 13470 43598 13522
rect 43650 13470 43652 13522
rect 43596 12178 43652 13470
rect 43596 12126 43598 12178
rect 43650 12126 43652 12178
rect 43596 12114 43652 12126
rect 43708 12962 43764 12974
rect 43708 12910 43710 12962
rect 43762 12910 43764 12962
rect 43708 12852 43764 12910
rect 43708 12068 43764 12796
rect 44268 12850 44324 13582
rect 44604 13076 44660 13694
rect 45276 13636 45332 13646
rect 44604 13020 45108 13076
rect 44268 12798 44270 12850
rect 44322 12798 44324 12850
rect 44044 12628 44100 12638
rect 44044 12178 44100 12572
rect 44044 12126 44046 12178
rect 44098 12126 44100 12178
rect 44044 12114 44100 12126
rect 44268 12180 44324 12798
rect 44828 12852 44884 12862
rect 44828 12758 44884 12796
rect 44940 12738 44996 12750
rect 44940 12686 44942 12738
rect 44994 12686 44996 12738
rect 44268 12114 44324 12124
rect 44604 12180 44660 12190
rect 44940 12180 44996 12686
rect 44604 12178 44996 12180
rect 44604 12126 44606 12178
rect 44658 12126 44996 12178
rect 44604 12124 44996 12126
rect 45052 12404 45108 13020
rect 45164 12964 45220 12974
rect 45164 12870 45220 12908
rect 44604 12114 44660 12124
rect 43708 12002 43764 12012
rect 45052 12066 45108 12348
rect 45164 12180 45220 12190
rect 45164 12086 45220 12124
rect 45052 12014 45054 12066
rect 45106 12014 45108 12066
rect 45052 12002 45108 12014
rect 45276 11954 45332 13580
rect 45276 11902 45278 11954
rect 45330 11902 45332 11954
rect 45276 11890 45332 11902
rect 43260 11282 43316 11294
rect 43596 11284 43652 11294
rect 43260 11230 43262 11282
rect 43314 11230 43316 11282
rect 43036 10446 43038 10498
rect 43090 10446 43092 10498
rect 43036 10434 43092 10446
rect 43148 11172 43204 11182
rect 42588 9886 42590 9938
rect 42642 9886 42644 9938
rect 42588 9874 42644 9886
rect 43036 9938 43092 9950
rect 43036 9886 43038 9938
rect 43090 9886 43092 9938
rect 41692 9662 41694 9714
rect 41746 9662 41748 9714
rect 41692 9650 41748 9662
rect 40908 9550 40910 9602
rect 40962 9550 40964 9602
rect 40908 9538 40964 9550
rect 41356 9604 41412 9614
rect 41356 9510 41412 9548
rect 40460 9214 40462 9266
rect 40514 9214 40516 9266
rect 40124 9102 40126 9154
rect 40178 9102 40180 9154
rect 40124 9090 40180 9102
rect 39788 8990 39790 9042
rect 39842 8990 39844 9042
rect 39788 8978 39844 8990
rect 40460 8428 40516 9214
rect 39004 8372 39284 8428
rect 40348 8372 40516 8428
rect 41692 9492 41748 9502
rect 38780 8260 38836 8270
rect 38780 8166 38836 8204
rect 38892 8148 38948 8158
rect 39004 8148 39060 8316
rect 39116 8260 39172 8270
rect 39900 8260 39956 8270
rect 39116 8258 39956 8260
rect 39116 8206 39118 8258
rect 39170 8206 39902 8258
rect 39954 8206 39956 8258
rect 39116 8204 39956 8206
rect 39116 8194 39172 8204
rect 39900 8194 39956 8204
rect 40348 8258 40404 8372
rect 40348 8206 40350 8258
rect 40402 8206 40404 8258
rect 40348 8194 40404 8206
rect 38892 8146 39060 8148
rect 38892 8094 38894 8146
rect 38946 8094 39060 8146
rect 38892 8092 39060 8094
rect 40796 8148 40852 8158
rect 40796 8146 40964 8148
rect 40796 8094 40798 8146
rect 40850 8094 40964 8146
rect 40796 8092 40964 8094
rect 38892 8082 38948 8092
rect 40796 8082 40852 8092
rect 39452 8034 39508 8046
rect 39452 7982 39454 8034
rect 39506 7982 39508 8034
rect 38668 7298 38724 7308
rect 38892 7586 38948 7598
rect 38892 7534 38894 7586
rect 38946 7534 38948 7586
rect 38444 6514 38500 6524
rect 38444 6356 38500 6366
rect 38444 5682 38500 6300
rect 38892 6020 38948 7534
rect 39116 7476 39172 7486
rect 39116 6690 39172 7420
rect 39228 7476 39284 7486
rect 39452 7476 39508 7982
rect 39228 7474 39508 7476
rect 39228 7422 39230 7474
rect 39282 7422 39508 7474
rect 39228 7420 39508 7422
rect 39900 7812 39956 7822
rect 39900 7474 39956 7756
rect 40124 7588 40180 7598
rect 40124 7494 40180 7532
rect 39900 7422 39902 7474
rect 39954 7422 39956 7474
rect 39228 6804 39284 7420
rect 39900 7410 39956 7422
rect 40796 7476 40852 7486
rect 40796 7382 40852 7420
rect 40908 7140 40964 8092
rect 41244 8036 41300 8046
rect 41244 8034 41524 8036
rect 41244 7982 41246 8034
rect 41298 7982 41524 8034
rect 41244 7980 41524 7982
rect 41244 7970 41300 7980
rect 41020 7812 41076 7822
rect 41020 7698 41076 7756
rect 41020 7646 41022 7698
rect 41074 7646 41076 7698
rect 41020 7634 41076 7646
rect 41132 7474 41188 7486
rect 41132 7422 41134 7474
rect 41186 7422 41188 7474
rect 41132 7364 41188 7422
rect 41132 7298 41188 7308
rect 41356 7474 41412 7486
rect 41356 7422 41358 7474
rect 41410 7422 41412 7474
rect 40908 7074 40964 7084
rect 41356 6916 41412 7422
rect 39228 6738 39284 6748
rect 40908 6860 41412 6916
rect 40908 6802 40964 6860
rect 40908 6750 40910 6802
rect 40962 6750 40964 6802
rect 39900 6692 39956 6702
rect 40908 6692 40964 6750
rect 39116 6638 39118 6690
rect 39170 6638 39172 6690
rect 39116 6626 39172 6638
rect 39788 6690 39956 6692
rect 39788 6638 39902 6690
rect 39954 6638 39956 6690
rect 39788 6636 39956 6638
rect 39116 6468 39172 6478
rect 39116 6374 39172 6412
rect 39676 6466 39732 6478
rect 39676 6414 39678 6466
rect 39730 6414 39732 6466
rect 39676 6356 39732 6414
rect 39676 6290 39732 6300
rect 38892 5954 38948 5964
rect 39228 6244 39284 6254
rect 38892 5796 38948 5806
rect 38444 5630 38446 5682
rect 38498 5630 38500 5682
rect 38444 5236 38500 5630
rect 38444 5170 38500 5180
rect 38668 5682 38724 5694
rect 38668 5630 38670 5682
rect 38722 5630 38724 5682
rect 38668 5348 38724 5630
rect 38668 5122 38724 5292
rect 38892 5234 38948 5740
rect 38892 5182 38894 5234
rect 38946 5182 38948 5234
rect 38892 5170 38948 5182
rect 38668 5070 38670 5122
rect 38722 5070 38724 5122
rect 38668 5058 38724 5070
rect 39228 4340 39284 6188
rect 39564 6132 39620 6142
rect 39340 5684 39396 5694
rect 39340 5590 39396 5628
rect 39340 5236 39396 5246
rect 39340 5142 39396 5180
rect 39564 5124 39620 6076
rect 39788 5906 39844 6636
rect 39900 6626 39956 6636
rect 40460 6636 40964 6692
rect 41020 6690 41076 6702
rect 41020 6638 41022 6690
rect 41074 6638 41076 6690
rect 40236 6468 40292 6478
rect 40460 6468 40516 6636
rect 40124 6466 40292 6468
rect 40124 6414 40238 6466
rect 40290 6414 40292 6466
rect 40124 6412 40292 6414
rect 39788 5854 39790 5906
rect 39842 5854 39844 5906
rect 39788 5684 39844 5854
rect 40012 6130 40068 6142
rect 40012 6078 40014 6130
rect 40066 6078 40068 6130
rect 40012 5908 40068 6078
rect 40012 5842 40068 5852
rect 40124 5906 40180 6412
rect 40236 6402 40292 6412
rect 40348 6466 40516 6468
rect 40348 6414 40462 6466
rect 40514 6414 40516 6466
rect 40348 6412 40516 6414
rect 40348 6018 40404 6412
rect 40460 6402 40516 6412
rect 40572 6468 40628 6478
rect 41020 6468 41076 6638
rect 40572 6466 40964 6468
rect 40572 6414 40574 6466
rect 40626 6414 40964 6466
rect 40572 6412 40964 6414
rect 40572 6402 40628 6412
rect 40348 5966 40350 6018
rect 40402 5966 40404 6018
rect 40348 5954 40404 5966
rect 40124 5854 40126 5906
rect 40178 5854 40180 5906
rect 39788 5618 39844 5628
rect 39676 5348 39732 5358
rect 40124 5348 40180 5854
rect 40908 5906 40964 6412
rect 41020 6018 41076 6412
rect 41020 5966 41022 6018
rect 41074 5966 41076 6018
rect 41020 5954 41076 5966
rect 41244 6692 41300 6702
rect 40908 5854 40910 5906
rect 40962 5854 40964 5906
rect 40908 5842 40964 5854
rect 40908 5684 40964 5694
rect 39676 5346 40740 5348
rect 39676 5294 39678 5346
rect 39730 5294 40740 5346
rect 39676 5292 40740 5294
rect 39676 5282 39732 5292
rect 40684 5234 40740 5292
rect 40908 5346 40964 5628
rect 40908 5294 40910 5346
rect 40962 5294 40964 5346
rect 40908 5282 40964 5294
rect 41244 5346 41300 6636
rect 41356 6020 41412 6030
rect 41468 6020 41524 7980
rect 41580 7588 41636 7598
rect 41580 7494 41636 7532
rect 41692 7586 41748 9436
rect 42924 9492 42980 9502
rect 42924 9154 42980 9436
rect 43036 9380 43092 9886
rect 43148 9826 43204 11116
rect 43260 10500 43316 11230
rect 43484 11282 43652 11284
rect 43484 11230 43598 11282
rect 43650 11230 43652 11282
rect 43484 11228 43652 11230
rect 43260 10434 43316 10444
rect 43372 11170 43428 11182
rect 43372 11118 43374 11170
rect 43426 11118 43428 11170
rect 43372 10164 43428 11118
rect 43484 11172 43540 11228
rect 43596 11218 43652 11228
rect 45612 11284 45668 11294
rect 45612 11190 45668 11228
rect 43484 11106 43540 11116
rect 44492 11172 44548 11182
rect 44492 10722 44548 11116
rect 45388 11170 45444 11182
rect 45388 11118 45390 11170
rect 45442 11118 45444 11170
rect 44492 10670 44494 10722
rect 44546 10670 44548 10722
rect 44492 10658 44548 10670
rect 45276 11060 45332 11070
rect 43596 10610 43652 10622
rect 43596 10558 43598 10610
rect 43650 10558 43652 10610
rect 43372 10098 43428 10108
rect 43484 10498 43540 10510
rect 43484 10446 43486 10498
rect 43538 10446 43540 10498
rect 43148 9774 43150 9826
rect 43202 9774 43204 9826
rect 43148 9762 43204 9774
rect 43036 9324 43204 9380
rect 42924 9102 42926 9154
rect 42978 9102 42980 9154
rect 42924 9090 42980 9102
rect 43036 9156 43092 9166
rect 43036 9062 43092 9100
rect 43148 9044 43204 9324
rect 43484 9044 43540 10446
rect 43596 10052 43652 10558
rect 44380 10388 44436 10398
rect 44268 10386 44436 10388
rect 44268 10334 44382 10386
rect 44434 10334 44436 10386
rect 44268 10332 44436 10334
rect 43596 9996 44100 10052
rect 44044 9938 44100 9996
rect 44044 9886 44046 9938
rect 44098 9886 44100 9938
rect 44044 9874 44100 9886
rect 44268 9826 44324 10332
rect 44380 10322 44436 10332
rect 45276 9940 45332 11004
rect 45388 10276 45444 11118
rect 45724 10498 45780 15148
rect 46060 14644 46116 14654
rect 46060 14550 46116 14588
rect 46172 14418 46228 15262
rect 46396 15316 46452 15374
rect 46396 15250 46452 15260
rect 46508 15314 46564 15326
rect 46508 15262 46510 15314
rect 46562 15262 46564 15314
rect 46508 15204 46564 15262
rect 46508 15138 46564 15148
rect 46956 14644 47012 15484
rect 47068 15316 47124 15326
rect 47068 15222 47124 15260
rect 46956 14578 47012 14588
rect 46172 14366 46174 14418
rect 46226 14366 46228 14418
rect 46172 14354 46228 14366
rect 46956 13860 47012 13870
rect 47180 13860 47236 15484
rect 47404 15314 47460 15326
rect 47404 15262 47406 15314
rect 47458 15262 47460 15314
rect 47404 14532 47460 15262
rect 47516 15316 47572 15326
rect 47572 15260 47684 15316
rect 47516 15250 47572 15260
rect 47628 15202 47684 15260
rect 47964 15314 48020 15484
rect 48188 15428 48244 19852
rect 48748 18562 48804 18574
rect 48748 18510 48750 18562
rect 48802 18510 48804 18562
rect 48748 17780 48804 18510
rect 48748 17714 48804 17724
rect 48860 18116 48916 19966
rect 48972 18564 49028 20078
rect 49644 19794 49700 20860
rect 49756 20850 49812 20860
rect 50556 20412 50820 20422
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50556 20346 50820 20356
rect 49980 20020 50036 20030
rect 49980 19926 50036 19964
rect 49644 19742 49646 19794
rect 49698 19742 49700 19794
rect 49644 19236 49700 19742
rect 49644 19170 49700 19180
rect 52108 19684 52164 19694
rect 50556 18844 50820 18854
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50556 18778 50820 18788
rect 48972 18498 49028 18508
rect 49084 18452 49140 18462
rect 49084 18450 50036 18452
rect 49084 18398 49086 18450
rect 49138 18398 50036 18450
rect 49084 18396 50036 18398
rect 49084 18386 49140 18396
rect 48860 16882 48916 18060
rect 49084 17444 49140 17454
rect 49084 16994 49140 17388
rect 49980 17106 50036 18396
rect 51660 18450 51716 18462
rect 51660 18398 51662 18450
rect 51714 18398 51716 18450
rect 51212 18340 51268 18350
rect 51100 18004 51156 18014
rect 50764 17892 50820 17902
rect 50764 17798 50820 17836
rect 51100 17890 51156 17948
rect 51100 17838 51102 17890
rect 51154 17838 51156 17890
rect 51100 17826 51156 17838
rect 51212 17890 51268 18284
rect 51548 18228 51604 18238
rect 51548 18134 51604 18172
rect 51212 17838 51214 17890
rect 51266 17838 51268 17890
rect 51212 17826 51268 17838
rect 49980 17054 49982 17106
rect 50034 17054 50036 17106
rect 49980 17042 50036 17054
rect 50204 17778 50260 17790
rect 50204 17726 50206 17778
rect 50258 17726 50260 17778
rect 49084 16942 49086 16994
rect 49138 16942 49140 16994
rect 49084 16930 49140 16942
rect 48860 16830 48862 16882
rect 48914 16830 48916 16882
rect 48860 16818 48916 16830
rect 49644 16658 49700 16670
rect 49644 16606 49646 16658
rect 49698 16606 49700 16658
rect 48188 15362 48244 15372
rect 48636 16210 48692 16222
rect 48636 16158 48638 16210
rect 48690 16158 48692 16210
rect 47964 15262 47966 15314
rect 48018 15262 48020 15314
rect 47964 15250 48020 15262
rect 47628 15150 47630 15202
rect 47682 15150 47684 15202
rect 47628 14756 47684 15150
rect 47964 15092 48020 15102
rect 47964 15090 48580 15092
rect 47964 15038 47966 15090
rect 48018 15038 48580 15090
rect 47964 15036 48580 15038
rect 47964 15026 48020 15036
rect 47628 14700 47908 14756
rect 47740 14532 47796 14542
rect 47404 14530 47796 14532
rect 47404 14478 47742 14530
rect 47794 14478 47796 14530
rect 47404 14476 47796 14478
rect 47740 14466 47796 14476
rect 47852 14196 47908 14700
rect 48412 14644 48468 14654
rect 48412 14550 48468 14588
rect 48524 14530 48580 15036
rect 48524 14478 48526 14530
rect 48578 14478 48580 14530
rect 48524 14466 48580 14478
rect 48636 14196 48692 16158
rect 48748 16100 48804 16110
rect 48748 15426 48804 16044
rect 49644 16100 49700 16606
rect 49644 16034 49700 16044
rect 50204 16100 50260 17726
rect 51660 17778 51716 18398
rect 52108 18450 52164 19628
rect 53228 19684 53284 19694
rect 53228 19346 53284 19628
rect 53228 19294 53230 19346
rect 53282 19294 53284 19346
rect 53228 19282 53284 19294
rect 52780 19122 52836 19134
rect 52780 19070 52782 19122
rect 52834 19070 52836 19122
rect 52668 19012 52724 19022
rect 52108 18398 52110 18450
rect 52162 18398 52164 18450
rect 51996 18340 52052 18350
rect 51996 18246 52052 18284
rect 51660 17726 51662 17778
rect 51714 17726 51716 17778
rect 51660 17714 51716 17726
rect 51772 18004 51828 18014
rect 50876 17666 50932 17678
rect 50876 17614 50878 17666
rect 50930 17614 50932 17666
rect 50876 17444 50932 17614
rect 51548 17554 51604 17566
rect 51548 17502 51550 17554
rect 51602 17502 51604 17554
rect 51548 17444 51604 17502
rect 51772 17444 51828 17948
rect 52108 17444 52164 18398
rect 52220 19010 52724 19012
rect 52220 18958 52670 19010
rect 52722 18958 52724 19010
rect 52220 18956 52724 18958
rect 52220 17892 52276 18956
rect 52668 18946 52724 18956
rect 52220 17666 52276 17836
rect 52220 17614 52222 17666
rect 52274 17614 52276 17666
rect 52220 17602 52276 17614
rect 52668 17668 52724 17678
rect 52668 17574 52724 17612
rect 50876 17388 51716 17444
rect 50556 17276 50820 17286
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50556 17210 50820 17220
rect 50652 16996 50708 17006
rect 50652 16902 50708 16940
rect 51324 16884 51380 16894
rect 51324 16790 51380 16828
rect 50204 16034 50260 16044
rect 51660 15988 51716 17388
rect 51772 17442 51940 17444
rect 51772 17390 51774 17442
rect 51826 17390 51940 17442
rect 51772 17388 51940 17390
rect 52108 17388 52276 17444
rect 51772 17378 51828 17388
rect 51660 15986 51828 15988
rect 51660 15934 51662 15986
rect 51714 15934 51828 15986
rect 51660 15932 51828 15934
rect 51660 15922 51716 15932
rect 50556 15708 50820 15718
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50556 15642 50820 15652
rect 48748 15374 48750 15426
rect 48802 15374 48804 15426
rect 48748 15362 48804 15374
rect 49196 15314 49252 15326
rect 49196 15262 49198 15314
rect 49250 15262 49252 15314
rect 49196 14532 49252 15262
rect 50876 15314 50932 15326
rect 50876 15262 50878 15314
rect 50930 15262 50932 15314
rect 49196 14418 49252 14476
rect 50540 14532 50596 14542
rect 50540 14438 50596 14476
rect 49196 14366 49198 14418
rect 49250 14366 49252 14418
rect 49196 14354 49252 14366
rect 50428 14418 50484 14430
rect 50428 14366 50430 14418
rect 50482 14366 50484 14418
rect 47852 14140 48692 14196
rect 47404 13860 47460 13870
rect 47180 13858 47460 13860
rect 47180 13806 47406 13858
rect 47458 13806 47460 13858
rect 47180 13804 47460 13806
rect 46956 13748 47012 13804
rect 47404 13794 47460 13804
rect 47852 13860 47908 13870
rect 47852 13766 47908 13804
rect 46732 13746 47012 13748
rect 46732 13694 46958 13746
rect 47010 13694 47012 13746
rect 46732 13692 47012 13694
rect 46508 13636 46564 13646
rect 46508 13542 46564 13580
rect 46732 13186 46788 13692
rect 46956 13682 47012 13692
rect 47516 13748 47572 13758
rect 46732 13134 46734 13186
rect 46786 13134 46788 13186
rect 46732 13122 46788 13134
rect 46284 12964 46340 12974
rect 46284 12870 46340 12908
rect 47068 12964 47124 12974
rect 47068 12870 47124 12908
rect 46172 12850 46228 12862
rect 47292 12852 47348 12862
rect 46172 12798 46174 12850
rect 46226 12798 46228 12850
rect 46172 12404 46228 12798
rect 46172 12338 46228 12348
rect 47180 12796 47292 12852
rect 47068 12066 47124 12078
rect 47068 12014 47070 12066
rect 47122 12014 47124 12066
rect 47068 11788 47124 12014
rect 47180 11956 47236 12796
rect 47292 12758 47348 12796
rect 47292 12404 47348 12414
rect 47292 12310 47348 12348
rect 47516 12404 47572 13692
rect 47740 13746 47796 13758
rect 47740 13694 47742 13746
rect 47794 13694 47796 13746
rect 47740 13636 47796 13694
rect 48076 13748 48132 13758
rect 48076 13654 48132 13692
rect 47740 13570 47796 13580
rect 47852 12850 47908 12862
rect 47852 12798 47854 12850
rect 47906 12798 47908 12850
rect 47852 12404 47908 12798
rect 48300 12852 48356 12862
rect 48300 12758 48356 12796
rect 48412 12738 48468 12750
rect 48412 12686 48414 12738
rect 48466 12686 48468 12738
rect 47964 12404 48020 12414
rect 47516 12402 47796 12404
rect 47516 12350 47518 12402
rect 47570 12350 47796 12402
rect 47516 12348 47796 12350
rect 47852 12402 48020 12404
rect 47852 12350 47966 12402
rect 48018 12350 48020 12402
rect 47852 12348 48020 12350
rect 47180 11890 47236 11900
rect 47516 11788 47572 12348
rect 47068 11732 47572 11788
rect 47516 11508 47572 11732
rect 47628 12178 47684 12190
rect 47628 12126 47630 12178
rect 47682 12126 47684 12178
rect 47628 11732 47684 12126
rect 47740 12180 47796 12348
rect 47964 12338 48020 12348
rect 48412 12404 48468 12686
rect 48412 12338 48468 12348
rect 48076 12180 48132 12190
rect 47740 12178 48132 12180
rect 47740 12126 48078 12178
rect 48130 12126 48132 12178
rect 47740 12124 48132 12126
rect 48076 12114 48132 12124
rect 47628 11666 47684 11676
rect 47740 11956 47796 11966
rect 47628 11508 47684 11518
rect 47516 11506 47684 11508
rect 47516 11454 47630 11506
rect 47682 11454 47684 11506
rect 47516 11452 47684 11454
rect 47628 11442 47684 11452
rect 45724 10446 45726 10498
rect 45778 10446 45780 10498
rect 45724 10434 45780 10446
rect 45836 11394 45892 11406
rect 45836 11342 45838 11394
rect 45890 11342 45892 11394
rect 45836 10276 45892 11342
rect 47068 11284 47124 11294
rect 45388 10220 45892 10276
rect 45276 9938 45780 9940
rect 45276 9886 45278 9938
rect 45330 9886 45780 9938
rect 45276 9884 45780 9886
rect 45276 9874 45332 9884
rect 44268 9774 44270 9826
rect 44322 9774 44324 9826
rect 43932 9714 43988 9726
rect 43932 9662 43934 9714
rect 43986 9662 43988 9714
rect 43596 9044 43652 9054
rect 43820 9044 43876 9054
rect 43932 9044 43988 9662
rect 43484 9042 43764 9044
rect 43484 8990 43598 9042
rect 43650 8990 43764 9042
rect 43484 8988 43764 8990
rect 42476 8930 42532 8942
rect 42476 8878 42478 8930
rect 42530 8878 42532 8930
rect 42476 8428 42532 8878
rect 42588 8932 42644 8942
rect 42588 8838 42644 8876
rect 43036 8818 43092 8830
rect 43036 8766 43038 8818
rect 43090 8766 43092 8818
rect 43036 8428 43092 8766
rect 42140 8372 42196 8382
rect 42476 8372 43092 8428
rect 41692 7534 41694 7586
rect 41746 7534 41748 7586
rect 41692 7522 41748 7534
rect 42028 8370 42196 8372
rect 42028 8318 42142 8370
rect 42194 8318 42196 8370
rect 42028 8316 42196 8318
rect 42028 7476 42084 8316
rect 42140 8306 42196 8316
rect 42588 8146 42644 8372
rect 42588 8094 42590 8146
rect 42642 8094 42644 8146
rect 42588 8082 42644 8094
rect 42028 6804 42084 7420
rect 42588 7588 42644 7598
rect 42252 7364 42308 7374
rect 41916 6748 42084 6804
rect 42140 7308 42252 7364
rect 41916 6130 41972 6748
rect 41916 6078 41918 6130
rect 41970 6078 41972 6130
rect 41916 6066 41972 6078
rect 41412 5964 41524 6020
rect 41356 5954 41412 5964
rect 41804 5908 41860 5918
rect 41804 5814 41860 5852
rect 41244 5294 41246 5346
rect 41298 5294 41300 5346
rect 41244 5282 41300 5294
rect 40684 5182 40686 5234
rect 40738 5182 40740 5234
rect 40684 5170 40740 5182
rect 41132 5236 41188 5246
rect 39788 5124 39844 5134
rect 39564 5068 39788 5124
rect 39788 5030 39844 5068
rect 40684 4788 40740 4798
rect 39340 4340 39396 4350
rect 40012 4340 40068 4350
rect 39228 4338 39844 4340
rect 39228 4286 39342 4338
rect 39394 4286 39844 4338
rect 39228 4284 39844 4286
rect 39340 4274 39396 4284
rect 39116 4228 39172 4238
rect 39004 4226 39172 4228
rect 39004 4174 39118 4226
rect 39170 4174 39172 4226
rect 39004 4172 39172 4174
rect 38892 3668 38948 3678
rect 38892 3442 38948 3612
rect 38892 3390 38894 3442
rect 38946 3390 38948 3442
rect 38892 3378 38948 3390
rect 39004 3220 39060 4172
rect 39116 4162 39172 4172
rect 39676 3668 39732 3678
rect 39116 3554 39172 3566
rect 39116 3502 39118 3554
rect 39170 3502 39172 3554
rect 39116 3444 39172 3502
rect 39116 3378 39172 3388
rect 39004 3154 39060 3164
rect 39676 800 39732 3612
rect 39788 3666 39844 4284
rect 40012 4246 40068 4284
rect 40348 3892 40404 3902
rect 40348 3778 40404 3836
rect 40348 3726 40350 3778
rect 40402 3726 40404 3778
rect 40348 3714 40404 3726
rect 39788 3614 39790 3666
rect 39842 3614 39844 3666
rect 39788 3602 39844 3614
rect 40012 3554 40068 3566
rect 40012 3502 40014 3554
rect 40066 3502 40068 3554
rect 40012 3220 40068 3502
rect 40684 3442 40740 4732
rect 40908 4564 40964 4574
rect 40908 4470 40964 4508
rect 40908 4004 40964 4014
rect 40908 3554 40964 3948
rect 40908 3502 40910 3554
rect 40962 3502 40964 3554
rect 40908 3490 40964 3502
rect 40684 3390 40686 3442
rect 40738 3390 40740 3442
rect 40684 3378 40740 3390
rect 41132 3444 41188 5180
rect 41356 5124 41412 5134
rect 41356 4226 41412 5068
rect 42028 4898 42084 4910
rect 42028 4846 42030 4898
rect 42082 4846 42084 4898
rect 42028 4340 42084 4846
rect 42140 4450 42196 7308
rect 42252 7298 42308 7308
rect 42252 6916 42308 6926
rect 42252 5908 42308 6860
rect 42588 6804 42644 7532
rect 42364 6692 42420 6702
rect 42364 6598 42420 6636
rect 42364 5908 42420 5918
rect 42252 5906 42420 5908
rect 42252 5854 42366 5906
rect 42418 5854 42420 5906
rect 42252 5852 42420 5854
rect 42364 5842 42420 5852
rect 42588 5906 42644 6748
rect 43148 6802 43204 8988
rect 43596 8950 43652 8988
rect 43708 8428 43764 8988
rect 43876 8988 43988 9044
rect 44268 9042 44324 9774
rect 45612 9714 45668 9726
rect 45612 9662 45614 9714
rect 45666 9662 45668 9714
rect 45612 9604 45668 9662
rect 45724 9714 45780 9884
rect 45724 9662 45726 9714
rect 45778 9662 45780 9714
rect 45724 9650 45780 9662
rect 44268 8990 44270 9042
rect 44322 8990 44324 9042
rect 43820 8950 43876 8988
rect 44268 8978 44324 8990
rect 44492 9156 44548 9166
rect 44044 8484 44100 8494
rect 43708 8372 43988 8428
rect 43596 8258 43652 8270
rect 43596 8206 43598 8258
rect 43650 8206 43652 8258
rect 43148 6750 43150 6802
rect 43202 6750 43204 6802
rect 43148 6738 43204 6750
rect 43484 7812 43540 7822
rect 42588 5854 42590 5906
rect 42642 5854 42644 5906
rect 42588 5842 42644 5854
rect 43372 5794 43428 5806
rect 43372 5742 43374 5794
rect 43426 5742 43428 5794
rect 42924 5684 42980 5694
rect 42924 5590 42980 5628
rect 43148 5348 43204 5358
rect 43036 5124 43092 5134
rect 42252 4900 42308 4910
rect 42252 4806 42308 4844
rect 42364 4898 42420 4910
rect 42364 4846 42366 4898
rect 42418 4846 42420 4898
rect 42364 4564 42420 4846
rect 42476 4900 42532 4910
rect 42812 4900 42868 4910
rect 42476 4898 42756 4900
rect 42476 4846 42478 4898
rect 42530 4846 42756 4898
rect 42476 4844 42756 4846
rect 42476 4834 42532 4844
rect 42364 4498 42420 4508
rect 42140 4398 42142 4450
rect 42194 4398 42196 4450
rect 42140 4386 42196 4398
rect 42028 4274 42084 4284
rect 42364 4340 42420 4350
rect 42420 4284 42644 4340
rect 42364 4246 42420 4284
rect 41356 4174 41358 4226
rect 41410 4174 41412 4226
rect 41356 4162 41412 4174
rect 42140 4228 42196 4238
rect 42140 3666 42196 4172
rect 42364 3780 42420 3790
rect 42364 3686 42420 3724
rect 42588 3778 42644 4284
rect 42588 3726 42590 3778
rect 42642 3726 42644 3778
rect 42588 3714 42644 3726
rect 42700 3780 42756 4844
rect 42812 4806 42868 4844
rect 42700 3714 42756 3724
rect 43036 3778 43092 5068
rect 43148 5010 43204 5292
rect 43148 4958 43150 5010
rect 43202 4958 43204 5010
rect 43148 4340 43204 4958
rect 43148 4274 43204 4284
rect 43372 4004 43428 5742
rect 43372 3938 43428 3948
rect 43036 3726 43038 3778
rect 43090 3726 43092 3778
rect 43036 3714 43092 3726
rect 42140 3614 42142 3666
rect 42194 3614 42196 3666
rect 42140 3602 42196 3614
rect 41580 3556 41636 3566
rect 41580 3462 41636 3500
rect 41356 3444 41412 3454
rect 41132 3442 41412 3444
rect 41132 3390 41358 3442
rect 41410 3390 41412 3442
rect 41132 3388 41412 3390
rect 41356 3378 41412 3388
rect 43148 3444 43204 3454
rect 43484 3444 43540 7756
rect 43596 7364 43652 8206
rect 43932 8034 43988 8372
rect 43932 7982 43934 8034
rect 43986 7982 43988 8034
rect 43932 7970 43988 7982
rect 43708 7364 43764 7374
rect 43596 7308 43708 7364
rect 43708 7270 43764 7308
rect 44044 6692 44100 8428
rect 44044 6626 44100 6636
rect 44156 7476 44212 7486
rect 44156 5908 44212 7420
rect 44156 5842 44212 5852
rect 44380 5906 44436 5918
rect 44380 5854 44382 5906
rect 44434 5854 44436 5906
rect 43820 5794 43876 5806
rect 43820 5742 43822 5794
rect 43874 5742 43876 5794
rect 43708 5124 43764 5134
rect 43708 5030 43764 5068
rect 43820 3668 43876 5742
rect 44268 5684 44324 5694
rect 44044 5348 44100 5358
rect 44044 5122 44100 5292
rect 44044 5070 44046 5122
rect 44098 5070 44100 5122
rect 44044 5058 44100 5070
rect 44268 5012 44324 5628
rect 44380 5346 44436 5854
rect 44380 5294 44382 5346
rect 44434 5294 44436 5346
rect 44380 5282 44436 5294
rect 44156 5010 44324 5012
rect 44156 4958 44270 5010
rect 44322 4958 44324 5010
rect 44156 4956 44324 4958
rect 44156 4676 44212 4956
rect 44268 4946 44324 4956
rect 44044 4620 44212 4676
rect 44044 4338 44100 4620
rect 44044 4286 44046 4338
rect 44098 4286 44100 4338
rect 44044 4274 44100 4286
rect 44156 4228 44212 4238
rect 44156 4134 44212 4172
rect 43820 3554 43876 3612
rect 43820 3502 43822 3554
rect 43874 3502 43876 3554
rect 43820 3490 43876 3502
rect 43596 3444 43652 3454
rect 43484 3442 43652 3444
rect 43484 3390 43598 3442
rect 43650 3390 43652 3442
rect 43484 3388 43652 3390
rect 40012 3154 40068 3164
rect 43148 1764 43204 3388
rect 43596 3378 43652 3388
rect 44268 3444 44324 3454
rect 44492 3444 44548 9100
rect 45612 9156 45668 9548
rect 45612 9090 45668 9100
rect 45164 9042 45220 9054
rect 45164 8990 45166 9042
rect 45218 8990 45220 9042
rect 45164 8428 45220 8990
rect 45388 8932 45444 8942
rect 45388 8838 45444 8876
rect 45276 8820 45332 8830
rect 45276 8726 45332 8764
rect 44604 8372 45220 8428
rect 44604 7586 44660 8372
rect 44604 7534 44606 7586
rect 44658 7534 44660 7586
rect 44604 7522 44660 7534
rect 45500 6580 45556 6590
rect 45276 6468 45332 6478
rect 45276 6018 45332 6412
rect 45500 6466 45556 6524
rect 45500 6414 45502 6466
rect 45554 6414 45556 6466
rect 45500 6356 45556 6414
rect 45836 6356 45892 10220
rect 46060 10610 46116 10622
rect 46060 10558 46062 10610
rect 46114 10558 46116 10610
rect 45948 9602 46004 9614
rect 45948 9550 45950 9602
rect 46002 9550 46004 9602
rect 45948 9156 46004 9550
rect 45948 8146 46004 9100
rect 46060 8820 46116 10558
rect 46396 10498 46452 10510
rect 46396 10446 46398 10498
rect 46450 10446 46452 10498
rect 46284 10164 46340 10174
rect 46172 9604 46228 9614
rect 46284 9604 46340 10108
rect 46396 9828 46452 10446
rect 46396 9772 46676 9828
rect 46620 9716 46676 9772
rect 46844 9716 46900 9726
rect 46620 9714 46900 9716
rect 46620 9662 46846 9714
rect 46898 9662 46900 9714
rect 46620 9660 46900 9662
rect 46508 9604 46564 9614
rect 46284 9602 46564 9604
rect 46284 9550 46510 9602
rect 46562 9550 46564 9602
rect 46284 9548 46564 9550
rect 46172 9510 46228 9548
rect 46508 8932 46564 9548
rect 46508 8866 46564 8876
rect 46060 8754 46116 8764
rect 46844 8428 46900 9660
rect 46956 9602 47012 9614
rect 46956 9550 46958 9602
rect 47010 9550 47012 9602
rect 46956 8820 47012 9550
rect 47068 8932 47124 11228
rect 47740 10722 47796 11900
rect 47964 11284 48020 11294
rect 47740 10670 47742 10722
rect 47794 10670 47796 10722
rect 47740 10658 47796 10670
rect 47852 11282 48020 11284
rect 47852 11230 47966 11282
rect 48018 11230 48020 11282
rect 47852 11228 48020 11230
rect 47516 10610 47572 10622
rect 47516 10558 47518 10610
rect 47570 10558 47572 10610
rect 47516 10500 47572 10558
rect 47852 10500 47908 11228
rect 47964 11218 48020 11228
rect 48076 11170 48132 11182
rect 48076 11118 48078 11170
rect 48130 11118 48132 11170
rect 47964 10612 48020 10622
rect 48076 10612 48132 11118
rect 48300 11172 48356 11182
rect 48300 11078 48356 11116
rect 48524 10724 48580 14140
rect 48860 13972 48916 13982
rect 48636 13970 48916 13972
rect 48636 13918 48862 13970
rect 48914 13918 48916 13970
rect 48636 13916 48916 13918
rect 48636 12962 48692 13916
rect 48860 13906 48916 13916
rect 50316 13972 50372 13982
rect 50428 13972 50484 14366
rect 50556 14140 50820 14150
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50556 14074 50820 14084
rect 50316 13970 50484 13972
rect 50316 13918 50318 13970
rect 50370 13918 50484 13970
rect 50316 13916 50484 13918
rect 50316 13906 50372 13916
rect 49084 13860 49140 13870
rect 49084 13766 49140 13804
rect 49756 13860 49812 13870
rect 49756 13766 49812 13804
rect 50652 13860 50708 13870
rect 48748 13748 48804 13758
rect 48748 13654 48804 13692
rect 49980 13748 50036 13758
rect 49980 13654 50036 13692
rect 50652 13748 50708 13804
rect 50876 13748 50932 15262
rect 50652 13746 50932 13748
rect 50652 13694 50654 13746
rect 50706 13694 50932 13746
rect 50652 13692 50932 13694
rect 50988 15202 51044 15214
rect 50988 15150 50990 15202
rect 51042 15150 51044 15202
rect 50652 13682 50708 13692
rect 50652 13524 50708 13534
rect 50876 13524 50932 13534
rect 50988 13524 51044 15150
rect 51324 14530 51380 14542
rect 51324 14478 51326 14530
rect 51378 14478 51380 14530
rect 51212 14308 51268 14318
rect 51212 14214 51268 14252
rect 51212 13972 51268 13982
rect 51324 13972 51380 14478
rect 51772 14532 51828 15932
rect 51772 14418 51828 14476
rect 51772 14366 51774 14418
rect 51826 14366 51828 14418
rect 51772 14354 51828 14366
rect 51884 15874 51940 17388
rect 52220 16996 52276 17388
rect 52220 16994 52388 16996
rect 52220 16942 52222 16994
rect 52274 16942 52388 16994
rect 52220 16940 52388 16942
rect 52220 16930 52276 16940
rect 51996 16882 52052 16894
rect 51996 16830 51998 16882
rect 52050 16830 52052 16882
rect 51996 16322 52052 16830
rect 52108 16884 52164 16894
rect 52108 16660 52164 16828
rect 52108 16604 52276 16660
rect 51996 16270 51998 16322
rect 52050 16270 52052 16322
rect 51996 16258 52052 16270
rect 51884 15822 51886 15874
rect 51938 15822 51940 15874
rect 51212 13970 51380 13972
rect 51212 13918 51214 13970
rect 51266 13918 51380 13970
rect 51212 13916 51380 13918
rect 51884 13972 51940 15822
rect 51996 15540 52052 15550
rect 51996 15446 52052 15484
rect 52220 15148 52276 16604
rect 52332 15540 52388 16940
rect 52780 16884 52836 19070
rect 53452 18452 53508 18462
rect 53452 18358 53508 18396
rect 52780 16818 52836 16828
rect 53564 16882 53620 22428
rect 55020 22482 55076 22494
rect 55020 22430 55022 22482
rect 55074 22430 55076 22482
rect 55020 21588 55076 22430
rect 55580 22372 55636 22382
rect 55580 22278 55636 22316
rect 57932 22260 57988 22270
rect 55020 21522 55076 21532
rect 55468 21700 55524 21710
rect 55356 21362 55412 21374
rect 55356 21310 55358 21362
rect 55410 21310 55412 21362
rect 53676 20916 53732 20926
rect 53676 20018 53732 20860
rect 55356 20916 55412 21310
rect 55356 20850 55412 20860
rect 55356 20692 55412 20702
rect 55468 20692 55524 21644
rect 57932 21026 57988 22204
rect 57932 20974 57934 21026
rect 57986 20974 57988 21026
rect 57932 20962 57988 20974
rect 55580 20802 55636 20814
rect 55580 20750 55582 20802
rect 55634 20750 55636 20802
rect 55580 20692 55636 20750
rect 55356 20690 55636 20692
rect 55356 20638 55358 20690
rect 55410 20638 55636 20690
rect 55356 20636 55636 20638
rect 55356 20626 55412 20636
rect 53676 19966 53678 20018
rect 53730 19966 53732 20018
rect 53676 19954 53732 19966
rect 57932 20132 57988 20142
rect 55356 19796 55412 19806
rect 55356 19702 55412 19740
rect 57932 19458 57988 20076
rect 57932 19406 57934 19458
rect 57986 19406 57988 19458
rect 57932 19394 57988 19406
rect 55580 19236 55636 19246
rect 55580 19142 55636 19180
rect 57932 18900 57988 18910
rect 55356 18228 55412 18238
rect 55356 18134 55412 18172
rect 57932 17890 57988 18844
rect 57932 17838 57934 17890
rect 57986 17838 57988 17890
rect 57932 17826 57988 17838
rect 53564 16830 53566 16882
rect 53618 16830 53620 16882
rect 53564 16818 53620 16830
rect 55020 17778 55076 17790
rect 55020 17726 55022 17778
rect 55074 17726 55076 17778
rect 55020 16884 55076 17726
rect 55580 17668 55636 17678
rect 55580 17574 55636 17612
rect 55356 17556 55412 17566
rect 55020 16818 55076 16828
rect 55244 17500 55356 17556
rect 52780 16660 52836 16670
rect 52780 16322 52836 16604
rect 52780 16270 52782 16322
rect 52834 16270 52836 16322
rect 52780 16258 52836 16270
rect 52332 15474 52388 15484
rect 52892 16098 52948 16110
rect 52892 16046 52894 16098
rect 52946 16046 52948 16098
rect 52108 15092 52276 15148
rect 52668 15202 52724 15214
rect 52668 15150 52670 15202
rect 52722 15150 52724 15202
rect 52444 15092 52500 15102
rect 51996 14644 52052 14654
rect 51996 14530 52052 14588
rect 51996 14478 51998 14530
rect 52050 14478 52052 14530
rect 51996 14466 52052 14478
rect 51212 13906 51268 13916
rect 51884 13906 51940 13916
rect 50708 13522 51044 13524
rect 50708 13470 50878 13522
rect 50930 13470 51044 13522
rect 50708 13468 51044 13470
rect 48636 12910 48638 12962
rect 48690 12910 48692 12962
rect 48636 12898 48692 12910
rect 49756 12962 49812 12974
rect 49756 12910 49758 12962
rect 49810 12910 49812 12962
rect 49532 12290 49588 12302
rect 49532 12238 49534 12290
rect 49586 12238 49588 12290
rect 49308 11956 49364 11966
rect 49308 11862 49364 11900
rect 49196 11172 49252 11182
rect 49532 11172 49588 12238
rect 49644 12068 49700 12078
rect 49756 12068 49812 12910
rect 50428 12962 50484 12974
rect 50428 12910 50430 12962
rect 50482 12910 50484 12962
rect 50092 12740 50148 12750
rect 50092 12402 50148 12684
rect 50092 12350 50094 12402
rect 50146 12350 50148 12402
rect 50092 12338 50148 12350
rect 49644 12066 49812 12068
rect 49644 12014 49646 12066
rect 49698 12014 49812 12066
rect 49644 12012 49812 12014
rect 49868 12180 49924 12190
rect 49644 12002 49700 12012
rect 49868 11394 49924 12124
rect 49980 12178 50036 12190
rect 49980 12126 49982 12178
rect 50034 12126 50036 12178
rect 49980 12068 50036 12126
rect 49980 12002 50036 12012
rect 50204 12178 50260 12190
rect 50204 12126 50206 12178
rect 50258 12126 50260 12178
rect 49868 11342 49870 11394
rect 49922 11342 49924 11394
rect 49868 11330 49924 11342
rect 50204 11172 50260 12126
rect 50428 12180 50484 12910
rect 50652 12962 50708 13468
rect 50876 13458 50932 13468
rect 50652 12910 50654 12962
rect 50706 12910 50708 12962
rect 50652 12898 50708 12910
rect 51884 12964 51940 12974
rect 50556 12572 50820 12582
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50556 12506 50820 12516
rect 50652 12180 50708 12190
rect 50428 12178 50708 12180
rect 50428 12126 50654 12178
rect 50706 12126 50708 12178
rect 50428 12124 50708 12126
rect 50652 11844 50708 12124
rect 50988 12180 51044 12190
rect 50988 12066 51044 12124
rect 50988 12014 50990 12066
rect 51042 12014 51044 12066
rect 50988 12002 51044 12014
rect 51436 12178 51492 12190
rect 51436 12126 51438 12178
rect 51490 12126 51492 12178
rect 50652 11778 50708 11788
rect 51100 11732 51156 11742
rect 50428 11394 50484 11406
rect 50428 11342 50430 11394
rect 50482 11342 50484 11394
rect 50316 11284 50372 11294
rect 50316 11190 50372 11228
rect 49532 11170 50260 11172
rect 49532 11118 50206 11170
rect 50258 11118 50260 11170
rect 49532 11116 50260 11118
rect 48748 10724 48804 10734
rect 48524 10722 48804 10724
rect 48524 10670 48750 10722
rect 48802 10670 48804 10722
rect 48524 10668 48804 10670
rect 48748 10658 48804 10668
rect 47964 10610 48132 10612
rect 47964 10558 47966 10610
rect 48018 10558 48132 10610
rect 47964 10556 48132 10558
rect 47964 10546 48020 10556
rect 47516 10444 47908 10500
rect 47180 9828 47236 9838
rect 47516 9828 47572 10444
rect 47180 9826 47572 9828
rect 47180 9774 47182 9826
rect 47234 9774 47572 9826
rect 47180 9772 47572 9774
rect 47180 9762 47236 9772
rect 47180 9604 47236 9614
rect 47180 9154 47236 9548
rect 47516 9324 48020 9380
rect 47516 9266 47572 9324
rect 47516 9214 47518 9266
rect 47570 9214 47572 9266
rect 47516 9202 47572 9214
rect 47180 9102 47182 9154
rect 47234 9102 47236 9154
rect 47180 9090 47236 9102
rect 47292 9154 47348 9166
rect 47292 9102 47294 9154
rect 47346 9102 47348 9154
rect 47292 8932 47348 9102
rect 47852 9156 47908 9166
rect 47852 9062 47908 9100
rect 47068 8876 47348 8932
rect 47740 9042 47796 9054
rect 47740 8990 47742 9042
rect 47794 8990 47796 9042
rect 46956 8754 47012 8764
rect 46844 8372 47460 8428
rect 45948 8094 45950 8146
rect 46002 8094 46004 8146
rect 45948 8082 46004 8094
rect 46396 8258 46452 8270
rect 46396 8206 46398 8258
rect 46450 8206 46452 8258
rect 46396 7476 46452 8206
rect 47404 8034 47460 8372
rect 47404 7982 47406 8034
rect 47458 7982 47460 8034
rect 47404 7970 47460 7982
rect 47516 8146 47572 8158
rect 47516 8094 47518 8146
rect 47570 8094 47572 8146
rect 46396 7410 46452 7420
rect 47180 7476 47236 7486
rect 45500 6300 45892 6356
rect 45276 5966 45278 6018
rect 45330 5966 45332 6018
rect 45276 5954 45332 5966
rect 44828 5908 44884 5918
rect 44828 5814 44884 5852
rect 44940 5794 44996 5806
rect 44940 5742 44942 5794
rect 44994 5742 44996 5794
rect 44940 5234 44996 5742
rect 45276 5684 45332 5694
rect 44940 5182 44942 5234
rect 44994 5182 44996 5234
rect 44940 5170 44996 5182
rect 45164 5348 45220 5358
rect 44716 5124 44772 5134
rect 45164 5124 45220 5292
rect 44716 5030 44772 5068
rect 45052 5122 45220 5124
rect 45052 5070 45166 5122
rect 45218 5070 45220 5122
rect 45052 5068 45220 5070
rect 45276 5124 45332 5628
rect 45388 5124 45444 5134
rect 45276 5122 45444 5124
rect 45276 5070 45390 5122
rect 45442 5070 45444 5122
rect 45276 5068 45444 5070
rect 44940 4340 44996 4350
rect 44940 4246 44996 4284
rect 44716 4228 44772 4238
rect 44716 4134 44772 4172
rect 44604 4114 44660 4126
rect 44604 4062 44606 4114
rect 44658 4062 44660 4114
rect 44604 3780 44660 4062
rect 44604 3714 44660 3724
rect 44268 3442 44548 3444
rect 44268 3390 44270 3442
rect 44322 3390 44548 3442
rect 44268 3388 44548 3390
rect 44604 3444 44660 3454
rect 44268 3378 44324 3388
rect 44604 3350 44660 3388
rect 44940 3444 44996 3454
rect 45052 3444 45108 5068
rect 45164 5058 45220 5068
rect 45388 5058 45444 5068
rect 45724 5124 45780 5134
rect 45164 4564 45220 4574
rect 45164 3556 45220 4508
rect 45724 4450 45780 5068
rect 45836 5012 45892 6300
rect 46060 6804 46116 6814
rect 45948 5012 46004 5022
rect 45836 5010 46004 5012
rect 45836 4958 45950 5010
rect 46002 4958 46004 5010
rect 45836 4956 46004 4958
rect 45948 4946 46004 4956
rect 46060 5010 46116 6748
rect 46284 6692 46340 6702
rect 46284 6132 46340 6636
rect 47180 6468 47236 7420
rect 47516 7474 47572 8094
rect 47628 7588 47684 7598
rect 47740 7588 47796 8990
rect 47964 9044 48020 9324
rect 48076 9266 48132 10556
rect 48188 10610 48244 10622
rect 48188 10558 48190 10610
rect 48242 10558 48244 10610
rect 48188 10500 48244 10558
rect 49196 10610 49252 11116
rect 50204 11106 50260 11116
rect 49196 10558 49198 10610
rect 49250 10558 49252 10610
rect 49196 10546 49252 10558
rect 48188 10434 48244 10444
rect 49644 10500 49700 10510
rect 49700 10444 49812 10500
rect 49644 10406 49700 10444
rect 48524 9826 48580 9838
rect 48524 9774 48526 9826
rect 48578 9774 48580 9826
rect 48076 9214 48078 9266
rect 48130 9214 48132 9266
rect 48076 9202 48132 9214
rect 48188 9714 48244 9726
rect 48188 9662 48190 9714
rect 48242 9662 48244 9714
rect 48188 9044 48244 9662
rect 47964 8988 48244 9044
rect 48524 9716 48580 9774
rect 48524 8428 48580 9660
rect 49756 9602 49812 10444
rect 50428 9938 50484 11342
rect 50556 11004 50820 11014
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50556 10938 50820 10948
rect 51100 10724 51156 11676
rect 51436 11396 51492 12126
rect 51884 12180 51940 12908
rect 51996 12852 52052 12862
rect 51996 12292 52052 12796
rect 52108 12402 52164 15092
rect 52444 14998 52500 15036
rect 52668 14644 52724 15150
rect 52892 15202 52948 16046
rect 52892 15150 52894 15202
rect 52946 15150 52948 15202
rect 52892 14868 52948 15150
rect 52892 14802 52948 14812
rect 53116 16098 53172 16110
rect 53116 16046 53118 16098
rect 53170 16046 53172 16098
rect 53116 15314 53172 16046
rect 55244 15988 55300 17500
rect 55356 17490 55412 17500
rect 57932 17556 57988 17566
rect 55356 16658 55412 16670
rect 55356 16606 55358 16658
rect 55410 16606 55412 16658
rect 55356 16212 55412 16606
rect 57932 16322 57988 17500
rect 57932 16270 57934 16322
rect 57986 16270 57988 16322
rect 57932 16258 57988 16270
rect 55356 16146 55412 16156
rect 55580 16100 55636 16110
rect 55580 16006 55636 16044
rect 55356 15988 55412 15998
rect 55244 15986 55412 15988
rect 55244 15934 55358 15986
rect 55410 15934 55412 15986
rect 55244 15932 55412 15934
rect 55356 15922 55412 15932
rect 54236 15874 54292 15886
rect 54236 15822 54238 15874
rect 54290 15822 54292 15874
rect 54236 15540 54292 15822
rect 54236 15474 54292 15484
rect 57932 15540 57988 15550
rect 53116 15262 53118 15314
rect 53170 15262 53172 15314
rect 53004 14756 53060 14766
rect 53004 14662 53060 14700
rect 52668 14578 52724 14588
rect 52892 14532 52948 14542
rect 52892 14438 52948 14476
rect 53116 14308 53172 15262
rect 53452 15316 53508 15326
rect 53452 15222 53508 15260
rect 53340 15092 53396 15102
rect 53340 14530 53396 15036
rect 55356 15090 55412 15102
rect 55356 15038 55358 15090
rect 55410 15038 55412 15090
rect 54124 14868 54180 14878
rect 54124 14642 54180 14812
rect 55356 14868 55412 15038
rect 55356 14802 55412 14812
rect 55580 15092 55636 15102
rect 54124 14590 54126 14642
rect 54178 14590 54180 14642
rect 53340 14478 53342 14530
rect 53394 14478 53396 14530
rect 53340 14308 53396 14478
rect 53788 14530 53844 14542
rect 53788 14478 53790 14530
rect 53842 14478 53844 14530
rect 53788 14308 53844 14478
rect 54124 14532 54180 14590
rect 54908 14644 54964 14654
rect 54908 14550 54964 14588
rect 55580 14532 55636 15036
rect 57932 14754 57988 15484
rect 57932 14702 57934 14754
rect 57986 14702 57988 14754
rect 57932 14690 57988 14702
rect 54124 14466 54180 14476
rect 55356 14530 55636 14532
rect 55356 14478 55582 14530
rect 55634 14478 55636 14530
rect 55356 14476 55636 14478
rect 54796 14420 54852 14430
rect 53340 14252 53732 14308
rect 53116 14242 53172 14252
rect 53004 13972 53060 13982
rect 53676 13972 53732 14252
rect 53788 14242 53844 14252
rect 54236 14418 54852 14420
rect 54236 14366 54798 14418
rect 54850 14366 54852 14418
rect 54236 14364 54852 14366
rect 53900 13972 53956 13982
rect 53676 13970 53956 13972
rect 53676 13918 53902 13970
rect 53954 13918 53956 13970
rect 53676 13916 53956 13918
rect 52892 13748 52948 13758
rect 52780 13746 52948 13748
rect 52780 13694 52894 13746
rect 52946 13694 52948 13746
rect 52780 13692 52948 13694
rect 52780 13300 52836 13692
rect 52892 13682 52948 13692
rect 52220 13244 52836 13300
rect 52220 12962 52276 13244
rect 53004 13074 53060 13916
rect 53900 13906 53956 13916
rect 53564 13860 53620 13870
rect 53564 13766 53620 13804
rect 54236 13860 54292 14364
rect 54796 14354 54852 14364
rect 53004 13022 53006 13074
rect 53058 13022 53060 13074
rect 53004 13010 53060 13022
rect 53452 13746 53508 13758
rect 53452 13694 53454 13746
rect 53506 13694 53508 13746
rect 52220 12910 52222 12962
rect 52274 12910 52276 12962
rect 52220 12898 52276 12910
rect 52668 12964 52724 12974
rect 52668 12870 52724 12908
rect 53452 12964 53508 13694
rect 54236 13746 54292 13804
rect 54236 13694 54238 13746
rect 54290 13694 54292 13746
rect 54236 13682 54292 13694
rect 55020 14306 55076 14318
rect 55020 14254 55022 14306
rect 55074 14254 55076 14306
rect 54460 13636 54516 13646
rect 55020 13636 55076 14254
rect 55356 13970 55412 14476
rect 55580 14466 55636 14476
rect 56588 14532 56644 14542
rect 55356 13918 55358 13970
rect 55410 13918 55412 13970
rect 55356 13906 55412 13918
rect 56588 13858 56644 14476
rect 56588 13806 56590 13858
rect 56642 13806 56644 13858
rect 56588 13794 56644 13806
rect 57036 13748 57092 13758
rect 54460 13634 55076 13636
rect 54460 13582 54462 13634
rect 54514 13582 55076 13634
rect 54460 13580 55076 13582
rect 56700 13746 57092 13748
rect 56700 13694 57038 13746
rect 57090 13694 57092 13746
rect 56700 13692 57092 13694
rect 53564 12964 53620 12974
rect 53452 12962 53620 12964
rect 53452 12910 53566 12962
rect 53618 12910 53620 12962
rect 53452 12908 53620 12910
rect 52108 12350 52110 12402
rect 52162 12350 52164 12402
rect 52108 12338 52164 12350
rect 53116 12852 53172 12862
rect 51996 12226 52052 12236
rect 52668 12290 52724 12302
rect 52668 12238 52670 12290
rect 52722 12238 52724 12290
rect 51884 12086 51940 12124
rect 51884 11396 51940 11406
rect 51436 11394 52164 11396
rect 51436 11342 51886 11394
rect 51938 11342 52164 11394
rect 51436 11340 52164 11342
rect 51884 11330 51940 11340
rect 51660 11172 51716 11182
rect 51100 10630 51156 10668
rect 51436 11170 51828 11172
rect 51436 11118 51662 11170
rect 51714 11118 51828 11170
rect 51436 11116 51828 11118
rect 50428 9886 50430 9938
rect 50482 9886 50484 9938
rect 50428 9874 50484 9886
rect 49756 9550 49758 9602
rect 49810 9550 49812 9602
rect 49756 9538 49812 9550
rect 49868 9828 49924 9838
rect 49868 9714 49924 9772
rect 50540 9828 50596 9838
rect 50540 9734 50596 9772
rect 50988 9826 51044 9838
rect 50988 9774 50990 9826
rect 51042 9774 51044 9826
rect 49868 9662 49870 9714
rect 49922 9662 49924 9714
rect 49644 9380 49700 9390
rect 47628 7586 47796 7588
rect 47628 7534 47630 7586
rect 47682 7534 47796 7586
rect 47628 7532 47796 7534
rect 48300 8372 48580 8428
rect 49532 8484 49588 8494
rect 47628 7522 47684 7532
rect 47516 7422 47518 7474
rect 47570 7422 47572 7474
rect 47516 6692 47572 7422
rect 47852 6692 47908 6702
rect 47516 6690 48020 6692
rect 47516 6638 47854 6690
rect 47906 6638 48020 6690
rect 47516 6636 48020 6638
rect 47852 6626 47908 6636
rect 47404 6578 47460 6590
rect 47404 6526 47406 6578
rect 47458 6526 47460 6578
rect 47292 6468 47348 6478
rect 47404 6468 47460 6526
rect 47180 6412 47292 6468
rect 47348 6412 47460 6468
rect 47292 6402 47348 6412
rect 46284 5906 46340 6076
rect 47740 6132 47796 6142
rect 47740 6038 47796 6076
rect 46284 5854 46286 5906
rect 46338 5854 46340 5906
rect 46284 5842 46340 5854
rect 47180 5908 47236 5918
rect 47180 5906 47460 5908
rect 47180 5854 47182 5906
rect 47234 5854 47460 5906
rect 47180 5852 47460 5854
rect 47180 5842 47236 5852
rect 46060 4958 46062 5010
rect 46114 4958 46116 5010
rect 46060 4946 46116 4958
rect 46508 5794 46564 5806
rect 46508 5742 46510 5794
rect 46562 5742 46564 5794
rect 46508 5684 46564 5742
rect 45724 4398 45726 4450
rect 45778 4398 45780 4450
rect 45724 4386 45780 4398
rect 45948 4338 46004 4350
rect 45948 4286 45950 4338
rect 46002 4286 46004 4338
rect 45724 3892 45780 3902
rect 45612 3556 45668 3566
rect 45164 3554 45668 3556
rect 45164 3502 45166 3554
rect 45218 3502 45614 3554
rect 45666 3502 45668 3554
rect 45164 3500 45668 3502
rect 45164 3490 45220 3500
rect 45612 3490 45668 3500
rect 44940 3442 45108 3444
rect 44940 3390 44942 3442
rect 44994 3390 45108 3442
rect 44940 3388 45108 3390
rect 45724 3442 45780 3836
rect 45948 3554 46004 4286
rect 45948 3502 45950 3554
rect 46002 3502 46004 3554
rect 45948 3490 46004 3502
rect 46284 3556 46340 3566
rect 46284 3462 46340 3500
rect 45724 3390 45726 3442
rect 45778 3390 45780 3442
rect 44940 3378 44996 3388
rect 45724 3378 45780 3390
rect 46508 3332 46564 5628
rect 46956 5348 47012 5358
rect 46956 5122 47012 5292
rect 47068 5236 47124 5246
rect 47068 5142 47124 5180
rect 47404 5124 47460 5852
rect 47852 5796 47908 5806
rect 47852 5702 47908 5740
rect 47516 5684 47572 5694
rect 47516 5590 47572 5628
rect 47516 5124 47572 5134
rect 46956 5070 46958 5122
rect 47010 5070 47012 5122
rect 46620 5010 46676 5022
rect 46620 4958 46622 5010
rect 46674 4958 46676 5010
rect 46620 3892 46676 4958
rect 46956 5012 47012 5070
rect 47180 5122 47796 5124
rect 47180 5070 47518 5122
rect 47570 5070 47796 5122
rect 47180 5068 47796 5070
rect 46956 4956 47124 5012
rect 47068 4116 47124 4956
rect 47180 4338 47236 5068
rect 47516 5058 47572 5068
rect 47180 4286 47182 4338
rect 47234 4286 47236 4338
rect 47180 4274 47236 4286
rect 47068 4060 47684 4116
rect 46620 3826 46676 3836
rect 47404 3892 47460 3902
rect 47404 3554 47460 3836
rect 47404 3502 47406 3554
rect 47458 3502 47460 3554
rect 47404 3490 47460 3502
rect 47628 3554 47684 4060
rect 47628 3502 47630 3554
rect 47682 3502 47684 3554
rect 47628 3490 47684 3502
rect 47740 3554 47796 5068
rect 47964 4450 48020 6636
rect 48188 6690 48244 6702
rect 48188 6638 48190 6690
rect 48242 6638 48244 6690
rect 48076 5348 48132 5358
rect 48188 5348 48244 6638
rect 48300 6466 48356 8372
rect 49308 8148 49364 8158
rect 48748 7924 48804 7934
rect 48748 7588 48804 7868
rect 49308 7698 49364 8092
rect 49308 7646 49310 7698
rect 49362 7646 49364 7698
rect 49308 7634 49364 7646
rect 48748 7586 49140 7588
rect 48748 7534 48750 7586
rect 48802 7534 49140 7586
rect 48748 7532 49140 7534
rect 48748 7522 48804 7532
rect 48972 7252 49028 7262
rect 48972 6802 49028 7196
rect 48972 6750 48974 6802
rect 49026 6750 49028 6802
rect 48972 6738 49028 6750
rect 49084 6690 49140 7532
rect 49532 7028 49588 8428
rect 49644 8372 49700 9324
rect 49868 8596 49924 9662
rect 50988 9716 51044 9774
rect 50556 9436 50820 9446
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50556 9370 50820 9380
rect 50988 8820 51044 9660
rect 51436 9268 51492 11116
rect 51660 11106 51716 11116
rect 51772 11060 51828 11116
rect 51996 11170 52052 11182
rect 51996 11118 51998 11170
rect 52050 11118 52052 11170
rect 51996 11060 52052 11118
rect 51772 11004 52052 11060
rect 52108 10948 52164 11340
rect 52220 11284 52276 11294
rect 52220 11190 52276 11228
rect 51996 10892 52164 10948
rect 51548 10610 51604 10622
rect 51548 10558 51550 10610
rect 51602 10558 51604 10610
rect 51548 10388 51604 10558
rect 51604 10332 51940 10388
rect 51548 10322 51604 10332
rect 51772 10052 51828 10062
rect 51772 9826 51828 9996
rect 51772 9774 51774 9826
rect 51826 9774 51828 9826
rect 51772 9762 51828 9774
rect 51884 9714 51940 10332
rect 51884 9662 51886 9714
rect 51938 9662 51940 9714
rect 51884 9650 51940 9662
rect 51772 9268 51828 9278
rect 51436 9202 51492 9212
rect 51548 9266 51828 9268
rect 51548 9214 51774 9266
rect 51826 9214 51828 9266
rect 51548 9212 51828 9214
rect 51324 8932 51380 8942
rect 50988 8754 51044 8764
rect 51212 8930 51380 8932
rect 51212 8878 51326 8930
rect 51378 8878 51380 8930
rect 51212 8876 51380 8878
rect 49868 8530 49924 8540
rect 49644 8278 49700 8316
rect 51212 8372 51268 8876
rect 51324 8820 51380 8876
rect 51548 8820 51604 9212
rect 51772 9202 51828 9212
rect 51660 9044 51716 9082
rect 51996 9044 52052 10892
rect 52332 10724 52388 10734
rect 52668 10724 52724 12238
rect 53116 10948 53172 12796
rect 53452 12516 53508 12908
rect 53564 12898 53620 12908
rect 54460 12628 54516 13580
rect 56700 13300 56756 13692
rect 57036 13682 57092 13692
rect 57372 13636 57428 13646
rect 55580 13244 56756 13300
rect 57260 13634 57428 13636
rect 57260 13582 57374 13634
rect 57426 13582 57428 13634
rect 57260 13580 57428 13582
rect 55580 12962 55636 13244
rect 55580 12910 55582 12962
rect 55634 12910 55636 12962
rect 55580 12898 55636 12910
rect 55692 13132 56196 13188
rect 55244 12850 55300 12862
rect 55244 12798 55246 12850
rect 55298 12798 55300 12850
rect 55244 12740 55300 12798
rect 55468 12852 55524 12862
rect 55244 12674 55300 12684
rect 55356 12740 55412 12750
rect 55468 12740 55524 12796
rect 55356 12738 55524 12740
rect 55356 12686 55358 12738
rect 55410 12686 55524 12738
rect 55356 12684 55524 12686
rect 55356 12674 55412 12684
rect 54460 12562 54516 12572
rect 53452 12460 53620 12516
rect 53452 12292 53508 12302
rect 53340 11396 53396 11406
rect 53452 11396 53508 12236
rect 53564 11618 53620 12460
rect 55132 12292 55188 12302
rect 55132 12198 55188 12236
rect 53564 11566 53566 11618
rect 53618 11566 53620 11618
rect 53564 11554 53620 11566
rect 53788 12178 53844 12190
rect 53788 12126 53790 12178
rect 53842 12126 53844 12178
rect 53116 10882 53172 10892
rect 53228 11394 53508 11396
rect 53228 11342 53342 11394
rect 53394 11342 53508 11394
rect 53228 11340 53508 11342
rect 53564 11396 53620 11406
rect 53228 10834 53284 11340
rect 53340 11330 53396 11340
rect 53564 11302 53620 11340
rect 53788 11172 53844 12126
rect 55356 11844 55412 11854
rect 55132 11284 55188 11294
rect 55020 11282 55188 11284
rect 55020 11230 55134 11282
rect 55186 11230 55188 11282
rect 55020 11228 55188 11230
rect 53228 10782 53230 10834
rect 53282 10782 53284 10834
rect 53228 10770 53284 10782
rect 53340 11116 53844 11172
rect 54572 11170 54628 11182
rect 54572 11118 54574 11170
rect 54626 11118 54628 11170
rect 52388 10668 52836 10724
rect 52332 10630 52388 10668
rect 52220 10612 52276 10622
rect 52220 10518 52276 10556
rect 52668 10052 52724 10062
rect 52108 9828 52164 9838
rect 52668 9828 52724 9996
rect 52108 9734 52164 9772
rect 52332 9826 52724 9828
rect 52332 9774 52670 9826
rect 52722 9774 52724 9826
rect 52332 9772 52724 9774
rect 52332 9268 52388 9772
rect 52668 9762 52724 9772
rect 52780 9714 52836 10668
rect 52780 9662 52782 9714
rect 52834 9662 52836 9714
rect 52780 9650 52836 9662
rect 52892 10612 52948 10622
rect 52892 9492 52948 10556
rect 53340 10610 53396 11116
rect 53340 10558 53342 10610
rect 53394 10558 53396 10610
rect 53340 9938 53396 10558
rect 53676 10948 53732 10958
rect 53676 10610 53732 10892
rect 53676 10558 53678 10610
rect 53730 10558 53732 10610
rect 53676 10546 53732 10558
rect 53900 10612 53956 10622
rect 53900 10518 53956 10556
rect 54572 10610 54628 11118
rect 54572 10558 54574 10610
rect 54626 10558 54628 10610
rect 54572 10546 54628 10558
rect 54684 11170 54740 11182
rect 54684 11118 54686 11170
rect 54738 11118 54740 11170
rect 54236 10500 54292 10510
rect 54236 10406 54292 10444
rect 54684 10500 54740 11118
rect 54684 10434 54740 10444
rect 54908 11170 54964 11182
rect 54908 11118 54910 11170
rect 54962 11118 54964 11170
rect 54908 10724 54964 11118
rect 53340 9886 53342 9938
rect 53394 9886 53396 9938
rect 53340 9874 53396 9886
rect 53452 9940 53508 9950
rect 51716 8988 52052 9044
rect 52108 9266 52388 9268
rect 52108 9214 52334 9266
rect 52386 9214 52388 9266
rect 52108 9212 52388 9214
rect 51660 8978 51716 8988
rect 51324 8764 51604 8820
rect 51660 8820 51716 8830
rect 51212 8278 51268 8316
rect 50204 8260 50260 8270
rect 50204 8146 50260 8204
rect 50988 8260 51044 8270
rect 50988 8166 51044 8204
rect 50204 8094 50206 8146
rect 50258 8094 50260 8146
rect 50204 8082 50260 8094
rect 49868 8034 49924 8046
rect 49868 7982 49870 8034
rect 49922 7982 49924 8034
rect 49532 6972 49700 7028
rect 49084 6638 49086 6690
rect 49138 6638 49140 6690
rect 49084 6626 49140 6638
rect 48300 6414 48302 6466
rect 48354 6414 48356 6466
rect 48300 6402 48356 6414
rect 49196 6018 49252 6030
rect 49196 5966 49198 6018
rect 49250 5966 49252 6018
rect 49196 5796 49252 5966
rect 49644 6018 49700 6972
rect 49868 6804 49924 7982
rect 50652 8036 50708 8046
rect 50652 8034 50932 8036
rect 50652 7982 50654 8034
rect 50706 7982 50932 8034
rect 50652 7980 50932 7982
rect 50652 7970 50708 7980
rect 50556 7868 50820 7878
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50556 7802 50820 7812
rect 50652 7700 50708 7710
rect 50876 7700 50932 7980
rect 50652 7698 51044 7700
rect 50652 7646 50654 7698
rect 50706 7646 51044 7698
rect 50652 7644 51044 7646
rect 50652 7634 50708 7644
rect 49868 6738 49924 6748
rect 50204 7474 50260 7486
rect 50204 7422 50206 7474
rect 50258 7422 50260 7474
rect 50204 6692 50260 7422
rect 50428 7474 50484 7486
rect 50428 7422 50430 7474
rect 50482 7422 50484 7474
rect 50428 6804 50484 7422
rect 50876 7474 50932 7486
rect 50876 7422 50878 7474
rect 50930 7422 50932 7474
rect 50764 7364 50820 7374
rect 50876 7364 50932 7422
rect 50764 7362 50932 7364
rect 50764 7310 50766 7362
rect 50818 7310 50932 7362
rect 50764 7308 50932 7310
rect 50764 7298 50820 7308
rect 50428 6738 50484 6748
rect 50204 6626 50260 6636
rect 50876 6692 50932 6702
rect 49756 6580 49812 6590
rect 49756 6486 49812 6524
rect 50428 6580 50484 6590
rect 50092 6466 50148 6478
rect 50092 6414 50094 6466
rect 50146 6414 50148 6466
rect 50092 6020 50148 6414
rect 50204 6468 50260 6478
rect 50204 6374 50260 6412
rect 50316 6466 50372 6478
rect 50316 6414 50318 6466
rect 50370 6414 50372 6466
rect 50316 6020 50372 6414
rect 49644 5966 49646 6018
rect 49698 5966 49700 6018
rect 49644 5954 49700 5966
rect 49756 5964 50148 6020
rect 50204 5964 50372 6020
rect 50428 6468 50484 6524
rect 50540 6468 50596 6478
rect 50428 6466 50596 6468
rect 50428 6414 50542 6466
rect 50594 6414 50596 6466
rect 50428 6412 50596 6414
rect 49196 5730 49252 5740
rect 49308 5908 49364 5918
rect 49308 5794 49364 5852
rect 49308 5742 49310 5794
rect 49362 5742 49364 5794
rect 49308 5730 49364 5742
rect 48076 5346 48244 5348
rect 48076 5294 48078 5346
rect 48130 5294 48244 5346
rect 48076 5292 48244 5294
rect 48972 5682 49028 5694
rect 48972 5630 48974 5682
rect 49026 5630 49028 5682
rect 48076 5282 48132 5292
rect 48412 5236 48468 5246
rect 48412 5142 48468 5180
rect 48972 5236 49028 5630
rect 48972 5170 49028 5180
rect 49756 5236 49812 5964
rect 49756 5170 49812 5180
rect 49868 5796 49924 5806
rect 50204 5796 50260 5964
rect 50428 5908 50484 6412
rect 50540 6402 50596 6412
rect 50556 6300 50820 6310
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50556 6234 50820 6244
rect 49924 5740 50260 5796
rect 50316 5906 50484 5908
rect 50316 5854 50430 5906
rect 50482 5854 50484 5906
rect 50316 5852 50484 5854
rect 49868 5234 49924 5740
rect 50316 5346 50372 5852
rect 50428 5814 50484 5852
rect 50316 5294 50318 5346
rect 50370 5294 50372 5346
rect 50316 5282 50372 5294
rect 50764 5348 50820 5358
rect 50876 5348 50932 6636
rect 50988 6580 51044 7644
rect 51660 7474 51716 8764
rect 51772 8818 51828 8830
rect 51772 8766 51774 8818
rect 51826 8766 51828 8818
rect 51772 8708 51828 8766
rect 51772 8642 51828 8652
rect 51772 8484 51828 8494
rect 51772 8034 51828 8428
rect 52108 8370 52164 9212
rect 52332 9202 52388 9212
rect 52780 9436 52948 9492
rect 52108 8318 52110 8370
rect 52162 8318 52164 8370
rect 52108 8306 52164 8318
rect 52780 9042 52836 9436
rect 52780 8990 52782 9042
rect 52834 8990 52836 9042
rect 52780 8260 52836 8990
rect 52892 9268 52948 9278
rect 52892 9154 52948 9212
rect 53452 9266 53508 9884
rect 54124 9940 54180 9950
rect 53676 9826 53732 9838
rect 53676 9774 53678 9826
rect 53730 9774 53732 9826
rect 53676 9716 53732 9774
rect 53452 9214 53454 9266
rect 53506 9214 53508 9266
rect 53452 9202 53508 9214
rect 53564 9660 53676 9716
rect 53564 9266 53620 9660
rect 53676 9650 53732 9660
rect 53564 9214 53566 9266
rect 53618 9214 53620 9266
rect 53564 9202 53620 9214
rect 54124 9268 54180 9884
rect 54348 9826 54404 9838
rect 54348 9774 54350 9826
rect 54402 9774 54404 9826
rect 54236 9268 54292 9278
rect 54124 9266 54292 9268
rect 54124 9214 54238 9266
rect 54290 9214 54292 9266
rect 54124 9212 54292 9214
rect 54236 9202 54292 9212
rect 52892 9102 52894 9154
rect 52946 9102 52948 9154
rect 52892 8484 52948 9102
rect 53116 9044 53172 9054
rect 53116 9042 53284 9044
rect 53116 8990 53118 9042
rect 53170 8990 53284 9042
rect 53116 8988 53284 8990
rect 53116 8978 53172 8988
rect 52892 8418 52948 8428
rect 53228 8372 53284 8988
rect 54012 9042 54068 9054
rect 54012 8990 54014 9042
rect 54066 8990 54068 9042
rect 53676 8820 53732 8830
rect 54012 8820 54068 8990
rect 54124 9044 54180 9054
rect 54124 8950 54180 8988
rect 53676 8818 54068 8820
rect 53676 8766 53678 8818
rect 53730 8766 54068 8818
rect 53676 8764 54068 8766
rect 53676 8754 53732 8764
rect 54012 8708 54068 8764
rect 54348 8708 54404 9774
rect 54572 9828 54628 9838
rect 54572 9042 54628 9772
rect 54572 8990 54574 9042
rect 54626 8990 54628 9042
rect 54572 8978 54628 8990
rect 54684 9044 54740 9054
rect 54908 9044 54964 10668
rect 55020 10612 55076 11228
rect 55132 11218 55188 11228
rect 55020 10050 55076 10556
rect 55020 9998 55022 10050
rect 55074 9998 55076 10050
rect 55020 9986 55076 9998
rect 54740 8988 54964 9044
rect 54684 8978 54740 8988
rect 54012 8652 54404 8708
rect 53228 8316 53508 8372
rect 52780 8194 52836 8204
rect 52892 8258 52948 8270
rect 52892 8206 52894 8258
rect 52946 8206 52948 8258
rect 51772 7982 51774 8034
rect 51826 7982 51828 8034
rect 51772 7700 51828 7982
rect 52892 8148 52948 8206
rect 53452 8260 53508 8316
rect 51772 7634 51828 7644
rect 51996 7700 52052 7710
rect 51996 7586 52052 7644
rect 51996 7534 51998 7586
rect 52050 7534 52052 7586
rect 51996 7522 52052 7534
rect 51660 7422 51662 7474
rect 51714 7422 51716 7474
rect 51660 7410 51716 7422
rect 51548 7362 51604 7374
rect 51548 7310 51550 7362
rect 51602 7310 51604 7362
rect 51548 7028 51604 7310
rect 51100 6972 51604 7028
rect 51100 6802 51156 6972
rect 52556 6804 52612 6814
rect 51100 6750 51102 6802
rect 51154 6750 51156 6802
rect 51100 6738 51156 6750
rect 51212 6748 51492 6804
rect 51212 6580 51268 6748
rect 51436 6690 51492 6748
rect 51436 6638 51438 6690
rect 51490 6638 51492 6690
rect 50988 6524 51268 6580
rect 51324 6580 51380 6590
rect 51324 6486 51380 6524
rect 51100 5908 51156 5918
rect 51100 5814 51156 5852
rect 51436 5906 51492 6638
rect 52556 6130 52612 6748
rect 52556 6078 52558 6130
rect 52610 6078 52612 6130
rect 52556 6066 52612 6078
rect 52780 6468 52836 6478
rect 52892 6468 52948 8092
rect 53116 8146 53172 8158
rect 53116 8094 53118 8146
rect 53170 8094 53172 8146
rect 53004 6804 53060 6814
rect 53116 6804 53172 8094
rect 53228 8146 53284 8158
rect 53228 8094 53230 8146
rect 53282 8094 53284 8146
rect 53228 7028 53284 8094
rect 53452 7586 53508 8204
rect 53676 8260 53732 8270
rect 54012 8260 54068 8270
rect 53676 8258 54068 8260
rect 53676 8206 53678 8258
rect 53730 8206 54014 8258
rect 54066 8206 54068 8258
rect 53676 8204 54068 8206
rect 53676 8194 53732 8204
rect 54012 8194 54068 8204
rect 54124 8036 54180 8652
rect 54236 8258 54292 8270
rect 54236 8206 54238 8258
rect 54290 8206 54292 8258
rect 54236 8036 54292 8206
rect 54460 8260 54516 8270
rect 55356 8260 55412 11788
rect 55468 9268 55524 12684
rect 55692 12516 55748 13132
rect 56140 12962 56196 13132
rect 56812 13076 56868 13086
rect 56588 13074 56868 13076
rect 56588 13022 56814 13074
rect 56866 13022 56868 13074
rect 56588 13020 56868 13022
rect 56140 12910 56142 12962
rect 56194 12910 56196 12962
rect 56140 12898 56196 12910
rect 56364 12964 56420 12974
rect 56588 12964 56644 13020
rect 56812 13010 56868 13020
rect 56364 12962 56644 12964
rect 56364 12910 56366 12962
rect 56418 12910 56644 12962
rect 56364 12908 56644 12910
rect 56924 12962 56980 12974
rect 56924 12910 56926 12962
rect 56978 12910 56980 12962
rect 56364 12898 56420 12908
rect 55804 12850 55860 12862
rect 55804 12798 55806 12850
rect 55858 12798 55860 12850
rect 55804 12628 55860 12798
rect 56700 12850 56756 12862
rect 56700 12798 56702 12850
rect 56754 12798 56756 12850
rect 56028 12738 56084 12750
rect 56028 12686 56030 12738
rect 56082 12686 56084 12738
rect 56028 12628 56084 12686
rect 56588 12740 56644 12750
rect 56700 12740 56756 12798
rect 56924 12852 56980 12910
rect 56924 12786 56980 12796
rect 57260 12962 57316 13580
rect 57372 13570 57428 13580
rect 57260 12910 57262 12962
rect 57314 12910 57316 12962
rect 56644 12684 56756 12740
rect 56588 12674 56644 12684
rect 55804 12572 55972 12628
rect 55692 12460 55860 12516
rect 55580 12180 55636 12190
rect 55580 11506 55636 12124
rect 55580 11454 55582 11506
rect 55634 11454 55636 11506
rect 55580 10610 55636 11454
rect 55692 12178 55748 12190
rect 55692 12126 55694 12178
rect 55746 12126 55748 12178
rect 55692 11396 55748 12126
rect 55692 10722 55748 11340
rect 55804 11284 55860 12460
rect 55916 12292 55972 12572
rect 56028 12562 56084 12572
rect 56588 12292 56644 12302
rect 55916 12290 56644 12292
rect 55916 12238 56590 12290
rect 56642 12238 56644 12290
rect 55916 12236 56644 12238
rect 56588 12226 56644 12236
rect 57036 12180 57092 12190
rect 57036 12086 57092 12124
rect 55804 11190 55860 11228
rect 57260 11172 57316 12910
rect 57372 12066 57428 12078
rect 57372 12014 57374 12066
rect 57426 12014 57428 12066
rect 57372 11396 57428 12014
rect 57372 11340 57540 11396
rect 57484 11282 57540 11340
rect 57484 11230 57486 11282
rect 57538 11230 57540 11282
rect 57372 11172 57428 11182
rect 57260 11170 57428 11172
rect 57260 11118 57374 11170
rect 57426 11118 57428 11170
rect 57260 11116 57428 11118
rect 57372 11106 57428 11116
rect 56700 10836 56756 10846
rect 55692 10670 55694 10722
rect 55746 10670 55748 10722
rect 55692 10658 55748 10670
rect 55916 10834 56756 10836
rect 55916 10782 56702 10834
rect 56754 10782 56756 10834
rect 55916 10780 56756 10782
rect 55580 10558 55582 10610
rect 55634 10558 55636 10610
rect 55580 10388 55636 10558
rect 55916 10610 55972 10780
rect 56700 10770 56756 10780
rect 56812 10724 56868 10734
rect 55916 10558 55918 10610
rect 55970 10558 55972 10610
rect 55916 10546 55972 10558
rect 56476 10612 56532 10622
rect 56476 10518 56532 10556
rect 56812 10610 56868 10668
rect 56812 10558 56814 10610
rect 56866 10558 56868 10610
rect 56812 10546 56868 10558
rect 57036 10610 57092 10622
rect 57036 10558 57038 10610
rect 57090 10558 57092 10610
rect 56028 10500 56084 10510
rect 55580 10332 55860 10388
rect 55580 9938 55636 9950
rect 55580 9886 55582 9938
rect 55634 9886 55636 9938
rect 55580 9828 55636 9886
rect 55580 9762 55636 9772
rect 55692 9268 55748 9278
rect 55468 9266 55748 9268
rect 55468 9214 55694 9266
rect 55746 9214 55748 9266
rect 55468 9212 55748 9214
rect 55692 9202 55748 9212
rect 55804 8484 55860 10332
rect 56028 9826 56084 10444
rect 57036 10500 57092 10558
rect 57036 10434 57092 10444
rect 57484 10050 57540 11230
rect 57484 9998 57486 10050
rect 57538 9998 57540 10050
rect 57484 9986 57540 9998
rect 56028 9774 56030 9826
rect 56082 9774 56084 9826
rect 56028 9762 56084 9774
rect 57148 9826 57204 9838
rect 57148 9774 57150 9826
rect 57202 9774 57204 9826
rect 57148 9716 57204 9774
rect 57148 9650 57204 9660
rect 55916 9154 55972 9166
rect 55916 9102 55918 9154
rect 55970 9102 55972 9154
rect 55916 8708 55972 9102
rect 56028 9044 56084 9054
rect 56588 9044 56644 9054
rect 56028 9042 56644 9044
rect 56028 8990 56030 9042
rect 56082 8990 56590 9042
rect 56642 8990 56644 9042
rect 56028 8988 56644 8990
rect 56028 8978 56084 8988
rect 56588 8978 56644 8988
rect 56700 9042 56756 9054
rect 56700 8990 56702 9042
rect 56754 8990 56756 9042
rect 55916 8642 55972 8652
rect 55804 8428 56196 8484
rect 55916 8260 55972 8270
rect 55356 8258 55972 8260
rect 55356 8206 55918 8258
rect 55970 8206 55972 8258
rect 55356 8204 55972 8206
rect 54460 8166 54516 8204
rect 55916 8194 55972 8204
rect 53452 7534 53454 7586
rect 53506 7534 53508 7586
rect 53452 7522 53508 7534
rect 54012 7980 54292 8036
rect 54572 8146 54628 8158
rect 54572 8094 54574 8146
rect 54626 8094 54628 8146
rect 53340 7364 53396 7374
rect 53340 7362 53620 7364
rect 53340 7310 53342 7362
rect 53394 7310 53620 7362
rect 53340 7308 53620 7310
rect 53340 7298 53396 7308
rect 53228 6962 53284 6972
rect 53060 6748 53172 6804
rect 53004 6690 53060 6748
rect 53004 6638 53006 6690
rect 53058 6638 53060 6690
rect 53004 6626 53060 6638
rect 53116 6578 53172 6590
rect 53116 6526 53118 6578
rect 53170 6526 53172 6578
rect 53116 6468 53172 6526
rect 52892 6412 53396 6468
rect 51436 5854 51438 5906
rect 51490 5854 51492 5906
rect 51436 5842 51492 5854
rect 52780 6020 52836 6412
rect 53340 6130 53396 6412
rect 53340 6078 53342 6130
rect 53394 6078 53396 6130
rect 53340 6066 53396 6078
rect 53564 6130 53620 7308
rect 53900 7028 53956 7038
rect 53900 6690 53956 6972
rect 53900 6638 53902 6690
rect 53954 6638 53956 6690
rect 53900 6626 53956 6638
rect 54012 6466 54068 7980
rect 54572 7476 54628 8094
rect 56140 7700 56196 8428
rect 56588 8260 56644 8270
rect 56700 8260 56756 8990
rect 57036 9042 57092 9054
rect 57036 8990 57038 9042
rect 57090 8990 57092 9042
rect 57036 8372 57092 8990
rect 57484 8708 57540 8718
rect 57036 8316 57316 8372
rect 56588 8258 57204 8260
rect 56588 8206 56590 8258
rect 56642 8206 57204 8258
rect 56588 8204 57204 8206
rect 56588 8194 56644 8204
rect 56700 7700 56756 7710
rect 56140 7698 56756 7700
rect 56140 7646 56702 7698
rect 56754 7646 56756 7698
rect 56140 7644 56756 7646
rect 56700 7634 56756 7644
rect 55916 7588 55972 7598
rect 55916 7494 55972 7532
rect 57148 7588 57204 8204
rect 54572 7410 54628 7420
rect 54684 7474 54740 7486
rect 54684 7422 54686 7474
rect 54738 7422 54740 7474
rect 54684 7028 54740 7422
rect 56588 7476 56644 7486
rect 56588 7382 56644 7420
rect 57148 7474 57204 7532
rect 57260 8258 57316 8316
rect 57260 8206 57262 8258
rect 57314 8206 57316 8258
rect 57260 7700 57316 8206
rect 57484 8146 57540 8652
rect 57484 8094 57486 8146
rect 57538 8094 57540 8146
rect 57484 8082 57540 8094
rect 57260 7586 57316 7644
rect 57260 7534 57262 7586
rect 57314 7534 57316 7586
rect 57260 7522 57316 7534
rect 57148 7422 57150 7474
rect 57202 7422 57204 7474
rect 57148 7410 57204 7422
rect 54684 6962 54740 6972
rect 54012 6414 54014 6466
rect 54066 6414 54068 6466
rect 54012 6402 54068 6414
rect 53564 6078 53566 6130
rect 53618 6078 53620 6130
rect 53564 6066 53620 6078
rect 53228 6020 53284 6030
rect 52780 6018 53284 6020
rect 52780 5966 53230 6018
rect 53282 5966 53284 6018
rect 52780 5964 53284 5966
rect 52780 5906 52836 5964
rect 53228 5954 53284 5964
rect 52780 5854 52782 5906
rect 52834 5854 52836 5906
rect 52780 5842 52836 5854
rect 50764 5346 50932 5348
rect 50764 5294 50766 5346
rect 50818 5294 50932 5346
rect 50764 5292 50932 5294
rect 50764 5282 50820 5292
rect 49868 5182 49870 5234
rect 49922 5182 49924 5234
rect 49868 5170 49924 5182
rect 50092 5236 50148 5246
rect 50092 5142 50148 5180
rect 48188 5124 48244 5134
rect 48188 5030 48244 5068
rect 48524 5122 48580 5134
rect 48524 5070 48526 5122
rect 48578 5070 48580 5122
rect 47964 4398 47966 4450
rect 48018 4398 48020 4450
rect 47964 4386 48020 4398
rect 48524 3892 48580 5070
rect 50556 4732 50820 4742
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50556 4666 50820 4676
rect 48188 3836 48580 3892
rect 48188 3778 48244 3836
rect 48188 3726 48190 3778
rect 48242 3726 48244 3778
rect 48188 3714 48244 3726
rect 47740 3502 47742 3554
rect 47794 3502 47796 3554
rect 47740 3490 47796 3502
rect 46732 3444 46788 3454
rect 46732 3350 46788 3388
rect 46508 3266 46564 3276
rect 50556 3164 50820 3174
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50556 3098 50820 3108
rect 43036 1708 43204 1764
rect 43036 800 43092 1708
rect 37884 700 38388 756
rect 39648 0 39760 800
rect 43008 0 43120 800
<< via2 >>
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 8204 45778 8260 45780
rect 8204 45726 8206 45778
rect 8206 45726 8258 45778
rect 8258 45726 8260 45778
rect 8204 45724 8260 45726
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 7980 44380 8036 44436
rect 2044 44098 2100 44100
rect 2044 44046 2046 44098
rect 2046 44046 2098 44098
rect 2098 44046 2100 44098
rect 2044 44044 2100 44046
rect 1708 43708 1764 43764
rect 2492 43708 2548 43764
rect 7084 44044 7140 44100
rect 7644 44098 7700 44100
rect 7644 44046 7646 44098
rect 7646 44046 7698 44098
rect 7698 44046 7700 44098
rect 7644 44044 7700 44046
rect 8316 44044 8372 44100
rect 7196 43538 7252 43540
rect 7196 43486 7198 43538
rect 7198 43486 7250 43538
rect 7250 43486 7252 43538
rect 7196 43484 7252 43486
rect 1708 41970 1764 41972
rect 1708 41918 1710 41970
rect 1710 41918 1762 41970
rect 1762 41918 1764 41970
rect 1708 41916 1764 41918
rect 7084 43314 7140 43316
rect 7084 43262 7086 43314
rect 7086 43262 7138 43314
rect 7138 43262 7140 43314
rect 7084 43260 7140 43262
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 9660 46002 9716 46004
rect 9660 45950 9662 46002
rect 9662 45950 9714 46002
rect 9714 45950 9716 46002
rect 9660 45948 9716 45950
rect 11900 45948 11956 46004
rect 10780 45890 10836 45892
rect 10780 45838 10782 45890
rect 10782 45838 10834 45890
rect 10834 45838 10836 45890
rect 10780 45836 10836 45838
rect 11564 45836 11620 45892
rect 12348 45948 12404 46004
rect 14476 46002 14532 46004
rect 14476 45950 14478 46002
rect 14478 45950 14530 46002
rect 14530 45950 14532 46002
rect 14476 45948 14532 45950
rect 16044 46002 16100 46004
rect 16044 45950 16046 46002
rect 16046 45950 16098 46002
rect 16098 45950 16100 46002
rect 16044 45948 16100 45950
rect 16828 45948 16884 46004
rect 13132 45890 13188 45892
rect 13132 45838 13134 45890
rect 13134 45838 13186 45890
rect 13186 45838 13188 45890
rect 13132 45836 13188 45838
rect 10108 45612 10164 45668
rect 9884 45218 9940 45220
rect 9884 45166 9886 45218
rect 9886 45166 9938 45218
rect 9938 45166 9940 45218
rect 9884 45164 9940 45166
rect 8428 43484 8484 43540
rect 8652 44380 8708 44436
rect 7868 43260 7924 43316
rect 8540 43426 8596 43428
rect 8540 43374 8542 43426
rect 8542 43374 8594 43426
rect 8594 43374 8596 43426
rect 8540 43372 8596 43374
rect 7308 42642 7364 42644
rect 7308 42590 7310 42642
rect 7310 42590 7362 42642
rect 7362 42590 7364 42642
rect 7308 42588 7364 42590
rect 9660 44380 9716 44436
rect 9772 44210 9828 44212
rect 9772 44158 9774 44210
rect 9774 44158 9826 44210
rect 9826 44158 9828 44210
rect 9772 44156 9828 44158
rect 8764 44098 8820 44100
rect 8764 44046 8766 44098
rect 8766 44046 8818 44098
rect 8818 44046 8820 44098
rect 8764 44044 8820 44046
rect 8204 42588 8260 42644
rect 8876 43484 8932 43540
rect 2716 42530 2772 42532
rect 2716 42478 2718 42530
rect 2718 42478 2770 42530
rect 2770 42478 2772 42530
rect 2716 42476 2772 42478
rect 2380 42364 2436 42420
rect 2044 42252 2100 42308
rect 1708 41692 1764 41748
rect 2044 41580 2100 41636
rect 2380 41804 2436 41860
rect 2268 41186 2324 41188
rect 2268 41134 2270 41186
rect 2270 41134 2322 41186
rect 2322 41134 2324 41186
rect 2268 41132 2324 41134
rect 2380 41020 2436 41076
rect 1708 40348 1764 40404
rect 7532 42530 7588 42532
rect 7532 42478 7534 42530
rect 7534 42478 7586 42530
rect 7586 42478 7588 42530
rect 7532 42476 7588 42478
rect 4396 42252 4452 42308
rect 3612 41970 3668 41972
rect 3612 41918 3614 41970
rect 3614 41918 3666 41970
rect 3666 41918 3668 41970
rect 3612 41916 3668 41918
rect 3164 41858 3220 41860
rect 3164 41806 3166 41858
rect 3166 41806 3218 41858
rect 3218 41806 3220 41858
rect 3164 41804 3220 41806
rect 2940 41692 2996 41748
rect 3388 41692 3444 41748
rect 4396 41746 4452 41748
rect 4396 41694 4398 41746
rect 4398 41694 4450 41746
rect 4450 41694 4452 41746
rect 4396 41692 4452 41694
rect 4284 41580 4340 41636
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 10556 45666 10612 45668
rect 10556 45614 10558 45666
rect 10558 45614 10610 45666
rect 10610 45614 10612 45666
rect 10556 45612 10612 45614
rect 10444 45330 10500 45332
rect 10444 45278 10446 45330
rect 10446 45278 10498 45330
rect 10498 45278 10500 45330
rect 10444 45276 10500 45278
rect 12572 45778 12628 45780
rect 12572 45726 12574 45778
rect 12574 45726 12626 45778
rect 12626 45726 12628 45778
rect 12572 45724 12628 45726
rect 13244 45778 13300 45780
rect 13244 45726 13246 45778
rect 13246 45726 13298 45778
rect 13298 45726 13300 45778
rect 13244 45724 13300 45726
rect 11116 45164 11172 45220
rect 10220 44380 10276 44436
rect 10556 44434 10612 44436
rect 10556 44382 10558 44434
rect 10558 44382 10610 44434
rect 10610 44382 10612 44434
rect 10556 44380 10612 44382
rect 12124 45276 12180 45332
rect 12236 45218 12292 45220
rect 12236 45166 12238 45218
rect 12238 45166 12290 45218
rect 12290 45166 12292 45218
rect 12236 45164 12292 45166
rect 16492 45890 16548 45892
rect 16492 45838 16494 45890
rect 16494 45838 16546 45890
rect 16546 45838 16548 45890
rect 16492 45836 16548 45838
rect 26236 46060 26292 46116
rect 17500 45836 17556 45892
rect 13804 45276 13860 45332
rect 13916 45724 13972 45780
rect 13468 45164 13524 45220
rect 11564 44994 11620 44996
rect 11564 44942 11566 44994
rect 11566 44942 11618 44994
rect 11618 44942 11620 44994
rect 11564 44940 11620 44942
rect 12460 44940 12516 44996
rect 11340 44156 11396 44212
rect 10108 44044 10164 44100
rect 9996 43708 10052 43764
rect 10332 43148 10388 43204
rect 9100 42700 9156 42756
rect 9436 42700 9492 42756
rect 5964 41692 6020 41748
rect 5292 41356 5348 41412
rect 2716 41020 2772 41076
rect 1708 39676 1764 39732
rect 1708 39004 1764 39060
rect 2044 39058 2100 39060
rect 2044 39006 2046 39058
rect 2046 39006 2098 39058
rect 2098 39006 2100 39058
rect 2044 39004 2100 39006
rect 2604 40236 2660 40292
rect 3276 40236 3332 40292
rect 2940 39788 2996 39844
rect 2268 39618 2324 39620
rect 2268 39566 2270 39618
rect 2270 39566 2322 39618
rect 2322 39566 2324 39618
rect 2268 39564 2324 39566
rect 2156 38108 2212 38164
rect 4060 39788 4116 39844
rect 3724 39564 3780 39620
rect 3052 39228 3108 39284
rect 2716 39116 2772 39172
rect 2380 37826 2436 37828
rect 2380 37774 2382 37826
rect 2382 37774 2434 37826
rect 2434 37774 2436 37826
rect 2380 37772 2436 37774
rect 2268 37660 2324 37716
rect 3724 39058 3780 39060
rect 3724 39006 3726 39058
rect 3726 39006 3778 39058
rect 3778 39006 3780 39058
rect 3724 39004 3780 39006
rect 5068 41244 5124 41300
rect 5292 40626 5348 40628
rect 5292 40574 5294 40626
rect 5294 40574 5346 40626
rect 5346 40574 5348 40626
rect 5292 40572 5348 40574
rect 6412 41244 6468 41300
rect 6972 41186 7028 41188
rect 6972 41134 6974 41186
rect 6974 41134 7026 41186
rect 7026 41134 7028 41186
rect 6972 41132 7028 41134
rect 7644 41692 7700 41748
rect 8540 42252 8596 42308
rect 9212 42530 9268 42532
rect 9212 42478 9214 42530
rect 9214 42478 9266 42530
rect 9266 42478 9268 42530
rect 9212 42476 9268 42478
rect 8988 41916 9044 41972
rect 7196 41074 7252 41076
rect 7196 41022 7198 41074
rect 7198 41022 7250 41074
rect 7250 41022 7252 41074
rect 7196 41020 7252 41022
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 4396 39788 4452 39844
rect 4732 39676 4788 39732
rect 4844 39506 4900 39508
rect 4844 39454 4846 39506
rect 4846 39454 4898 39506
rect 4898 39454 4900 39506
rect 4844 39452 4900 39454
rect 4060 38780 4116 38836
rect 3500 38668 3556 38724
rect 4284 38834 4340 38836
rect 4284 38782 4286 38834
rect 4286 38782 4338 38834
rect 4338 38782 4340 38834
rect 4284 38780 4340 38782
rect 3164 38556 3220 38612
rect 2828 38108 2884 38164
rect 2716 37660 2772 37716
rect 2044 35980 2100 36036
rect 1708 35644 1764 35700
rect 2044 34354 2100 34356
rect 2044 34302 2046 34354
rect 2046 34302 2098 34354
rect 2098 34302 2100 34354
rect 2044 34300 2100 34302
rect 1708 33628 1764 33684
rect 2940 37772 2996 37828
rect 4956 39004 5012 39060
rect 5068 40124 5124 40180
rect 5852 40626 5908 40628
rect 5852 40574 5854 40626
rect 5854 40574 5906 40626
rect 5906 40574 5908 40626
rect 5852 40572 5908 40574
rect 5628 40124 5684 40180
rect 5740 39730 5796 39732
rect 5740 39678 5742 39730
rect 5742 39678 5794 39730
rect 5794 39678 5796 39730
rect 5740 39676 5796 39678
rect 4844 38668 4900 38724
rect 5852 39452 5908 39508
rect 6524 39730 6580 39732
rect 6524 39678 6526 39730
rect 6526 39678 6578 39730
rect 6578 39678 6580 39730
rect 6524 39676 6580 39678
rect 6412 39452 6468 39508
rect 5068 38668 5124 38724
rect 2492 35810 2548 35812
rect 2492 35758 2494 35810
rect 2494 35758 2546 35810
rect 2546 35758 2548 35810
rect 2492 35756 2548 35758
rect 4732 38610 4788 38612
rect 4732 38558 4734 38610
rect 4734 38558 4786 38610
rect 4786 38558 4788 38610
rect 4732 38556 4788 38558
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 5740 38668 5796 38724
rect 5852 38780 5908 38836
rect 5068 37938 5124 37940
rect 5068 37886 5070 37938
rect 5070 37886 5122 37938
rect 5122 37886 5124 37938
rect 5068 37884 5124 37886
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 3948 35868 4004 35924
rect 3164 35644 3220 35700
rect 2492 33628 2548 33684
rect 2716 33068 2772 33124
rect 3276 33068 3332 33124
rect 4396 35698 4452 35700
rect 4396 35646 4398 35698
rect 4398 35646 4450 35698
rect 4450 35646 4452 35698
rect 4396 35644 4452 35646
rect 4172 35308 4228 35364
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4956 35810 5012 35812
rect 4956 35758 4958 35810
rect 4958 35758 5010 35810
rect 5010 35758 5012 35810
rect 4956 35756 5012 35758
rect 3724 33404 3780 33460
rect 5068 34914 5124 34916
rect 5068 34862 5070 34914
rect 5070 34862 5122 34914
rect 5122 34862 5124 34914
rect 5068 34860 5124 34862
rect 6076 35810 6132 35812
rect 6076 35758 6078 35810
rect 6078 35758 6130 35810
rect 6130 35758 6132 35810
rect 6076 35756 6132 35758
rect 6188 34300 6244 34356
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 2716 31500 2772 31556
rect 3164 31500 3220 31556
rect 2828 31106 2884 31108
rect 2828 31054 2830 31106
rect 2830 31054 2882 31106
rect 2882 31054 2884 31106
rect 2828 31052 2884 31054
rect 2380 30268 2436 30324
rect 3724 31500 3780 31556
rect 4508 31836 4564 31892
rect 4172 31612 4228 31668
rect 3276 31052 3332 31108
rect 3500 30994 3556 30996
rect 3500 30942 3502 30994
rect 3502 30942 3554 30994
rect 3554 30942 3556 30994
rect 3500 30940 3556 30942
rect 4284 31164 4340 31220
rect 4172 31052 4228 31108
rect 4844 31724 4900 31780
rect 5068 33628 5124 33684
rect 5964 33458 6020 33460
rect 5964 33406 5966 33458
rect 5966 33406 6018 33458
rect 6018 33406 6020 33458
rect 5964 33404 6020 33406
rect 5964 32956 6020 33012
rect 8876 41244 8932 41300
rect 10108 42754 10164 42756
rect 10108 42702 10110 42754
rect 10110 42702 10162 42754
rect 10162 42702 10164 42754
rect 10108 42700 10164 42702
rect 11340 43596 11396 43652
rect 12124 44434 12180 44436
rect 12124 44382 12126 44434
rect 12126 44382 12178 44434
rect 12178 44382 12180 44434
rect 12124 44380 12180 44382
rect 12124 44210 12180 44212
rect 12124 44158 12126 44210
rect 12126 44158 12178 44210
rect 12178 44158 12180 44210
rect 12124 44156 12180 44158
rect 13804 44604 13860 44660
rect 12684 44044 12740 44100
rect 12124 43596 12180 43652
rect 10668 43148 10724 43204
rect 10444 42588 10500 42644
rect 10332 42476 10388 42532
rect 9996 41970 10052 41972
rect 9996 41918 9998 41970
rect 9998 41918 10050 41970
rect 10050 41918 10052 41970
rect 9996 41916 10052 41918
rect 9548 41244 9604 41300
rect 10668 41298 10724 41300
rect 10668 41246 10670 41298
rect 10670 41246 10722 41298
rect 10722 41246 10724 41298
rect 10668 41244 10724 41246
rect 7980 40962 8036 40964
rect 7980 40910 7982 40962
rect 7982 40910 8034 40962
rect 8034 40910 8036 40962
rect 7980 40908 8036 40910
rect 7196 40460 7252 40516
rect 7868 40514 7924 40516
rect 7868 40462 7870 40514
rect 7870 40462 7922 40514
rect 7922 40462 7924 40514
rect 7868 40460 7924 40462
rect 6524 37660 6580 37716
rect 6412 36316 6468 36372
rect 6860 39452 6916 39508
rect 7084 39452 7140 39508
rect 7308 39228 7364 39284
rect 6748 38668 6804 38724
rect 7644 39676 7700 39732
rect 6636 35980 6692 36036
rect 6188 33068 6244 33124
rect 5068 31836 5124 31892
rect 5964 32508 6020 32564
rect 4620 31106 4676 31108
rect 4620 31054 4622 31106
rect 4622 31054 4674 31106
rect 4674 31054 4676 31106
rect 4620 31052 4676 31054
rect 4172 30716 4228 30772
rect 3836 30380 3892 30436
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4508 30434 4564 30436
rect 4508 30382 4510 30434
rect 4510 30382 4562 30434
rect 4562 30382 4564 30434
rect 4508 30380 4564 30382
rect 6412 33346 6468 33348
rect 6412 33294 6414 33346
rect 6414 33294 6466 33346
rect 6466 33294 6468 33346
rect 6412 33292 6468 33294
rect 6412 32956 6468 33012
rect 7084 37660 7140 37716
rect 7420 36482 7476 36484
rect 7420 36430 7422 36482
rect 7422 36430 7474 36482
rect 7474 36430 7476 36482
rect 7420 36428 7476 36430
rect 6860 35532 6916 35588
rect 6972 35980 7028 36036
rect 7308 35980 7364 36036
rect 7084 35756 7140 35812
rect 7420 35868 7476 35924
rect 7308 35698 7364 35700
rect 7308 35646 7310 35698
rect 7310 35646 7362 35698
rect 7362 35646 7364 35698
rect 7308 35644 7364 35646
rect 7196 35532 7252 35588
rect 6860 34802 6916 34804
rect 6860 34750 6862 34802
rect 6862 34750 6914 34802
rect 6914 34750 6916 34802
rect 6860 34748 6916 34750
rect 7420 35586 7476 35588
rect 7420 35534 7422 35586
rect 7422 35534 7474 35586
rect 7474 35534 7476 35586
rect 7420 35532 7476 35534
rect 7420 34636 7476 34692
rect 6860 33292 6916 33348
rect 7196 33628 7252 33684
rect 9772 40572 9828 40628
rect 8316 39394 8372 39396
rect 8316 39342 8318 39394
rect 8318 39342 8370 39394
rect 8370 39342 8372 39394
rect 8316 39340 8372 39342
rect 8652 39618 8708 39620
rect 8652 39566 8654 39618
rect 8654 39566 8706 39618
rect 8706 39566 8708 39618
rect 8652 39564 8708 39566
rect 9660 39618 9716 39620
rect 9660 39566 9662 39618
rect 9662 39566 9714 39618
rect 9714 39566 9716 39618
rect 9660 39564 9716 39566
rect 8988 39340 9044 39396
rect 8764 39228 8820 39284
rect 7980 36428 8036 36484
rect 8204 35810 8260 35812
rect 8204 35758 8206 35810
rect 8206 35758 8258 35810
rect 8258 35758 8260 35810
rect 8204 35756 8260 35758
rect 8652 35756 8708 35812
rect 8540 35532 8596 35588
rect 8876 35420 8932 35476
rect 9660 38050 9716 38052
rect 9660 37998 9662 38050
rect 9662 37998 9714 38050
rect 9714 37998 9716 38050
rect 9660 37996 9716 37998
rect 11452 42866 11508 42868
rect 11452 42814 11454 42866
rect 11454 42814 11506 42866
rect 11506 42814 11508 42866
rect 11452 42812 11508 42814
rect 11676 42700 11732 42756
rect 13244 44380 13300 44436
rect 14140 45218 14196 45220
rect 14140 45166 14142 45218
rect 14142 45166 14194 45218
rect 14194 45166 14196 45218
rect 14140 45164 14196 45166
rect 14364 45276 14420 45332
rect 14812 45330 14868 45332
rect 14812 45278 14814 45330
rect 14814 45278 14866 45330
rect 14866 45278 14868 45330
rect 14812 45276 14868 45278
rect 14252 44828 14308 44884
rect 16828 45388 16884 45444
rect 16268 45276 16324 45332
rect 15596 45106 15652 45108
rect 15596 45054 15598 45106
rect 15598 45054 15650 45106
rect 15650 45054 15652 45106
rect 15596 45052 15652 45054
rect 15708 44994 15764 44996
rect 15708 44942 15710 44994
rect 15710 44942 15762 44994
rect 15762 44942 15764 44994
rect 15708 44940 15764 44942
rect 15372 44380 15428 44436
rect 15596 44716 15652 44772
rect 14924 44268 14980 44324
rect 16604 45218 16660 45220
rect 16604 45166 16606 45218
rect 16606 45166 16658 45218
rect 16658 45166 16660 45218
rect 16604 45164 16660 45166
rect 16492 44882 16548 44884
rect 16492 44830 16494 44882
rect 16494 44830 16546 44882
rect 16546 44830 16548 44882
rect 16492 44828 16548 44830
rect 16828 44492 16884 44548
rect 15484 44268 15540 44324
rect 13356 44156 13412 44212
rect 13468 44098 13524 44100
rect 13468 44046 13470 44098
rect 13470 44046 13522 44098
rect 13522 44046 13524 44098
rect 13468 44044 13524 44046
rect 13468 43708 13524 43764
rect 12684 43596 12740 43652
rect 12796 43372 12852 43428
rect 10892 42642 10948 42644
rect 10892 42590 10894 42642
rect 10894 42590 10946 42642
rect 10946 42590 10948 42642
rect 10892 42588 10948 42590
rect 10108 40460 10164 40516
rect 10332 40348 10388 40404
rect 9660 37378 9716 37380
rect 9660 37326 9662 37378
rect 9662 37326 9714 37378
rect 9714 37326 9716 37378
rect 9884 39116 9940 39172
rect 10556 39340 10612 39396
rect 9660 37324 9716 37326
rect 9772 37100 9828 37156
rect 9660 37042 9716 37044
rect 9660 36990 9662 37042
rect 9662 36990 9714 37042
rect 9714 36990 9716 37042
rect 9660 36988 9716 36990
rect 9100 35196 9156 35252
rect 9772 36204 9828 36260
rect 9212 35084 9268 35140
rect 9100 34748 9156 34804
rect 8988 34300 9044 34356
rect 8652 33964 8708 34020
rect 7308 33122 7364 33124
rect 7308 33070 7310 33122
rect 7310 33070 7362 33122
rect 7362 33070 7364 33122
rect 7308 33068 7364 33070
rect 7532 33122 7588 33124
rect 7532 33070 7534 33122
rect 7534 33070 7586 33122
rect 7586 33070 7588 33122
rect 7532 33068 7588 33070
rect 6860 32732 6916 32788
rect 7980 33346 8036 33348
rect 7980 33294 7982 33346
rect 7982 33294 8034 33346
rect 8034 33294 8036 33346
rect 7980 33292 8036 33294
rect 7980 32786 8036 32788
rect 7980 32734 7982 32786
rect 7982 32734 8034 32786
rect 8034 32734 8036 32786
rect 7980 32732 8036 32734
rect 7084 32562 7140 32564
rect 7084 32510 7086 32562
rect 7086 32510 7138 32562
rect 7138 32510 7140 32562
rect 7084 32508 7140 32510
rect 6412 31554 6468 31556
rect 6412 31502 6414 31554
rect 6414 31502 6466 31554
rect 6466 31502 6468 31554
rect 6412 31500 6468 31502
rect 4956 31388 5012 31444
rect 7308 31948 7364 32004
rect 7196 31890 7252 31892
rect 7196 31838 7198 31890
rect 7198 31838 7250 31890
rect 7250 31838 7252 31890
rect 7196 31836 7252 31838
rect 5404 30994 5460 30996
rect 5404 30942 5406 30994
rect 5406 30942 5458 30994
rect 5458 30942 5460 30994
rect 5404 30940 5460 30942
rect 6188 30882 6244 30884
rect 6188 30830 6190 30882
rect 6190 30830 6242 30882
rect 6242 30830 6244 30882
rect 6188 30828 6244 30830
rect 6076 30380 6132 30436
rect 4732 30268 4788 30324
rect 6972 30716 7028 30772
rect 6636 30210 6692 30212
rect 6636 30158 6638 30210
rect 6638 30158 6690 30210
rect 6690 30158 6692 30210
rect 6636 30156 6692 30158
rect 7196 30828 7252 30884
rect 8652 33234 8708 33236
rect 8652 33182 8654 33234
rect 8654 33182 8706 33234
rect 8706 33182 8708 33234
rect 8652 33180 8708 33182
rect 8988 33346 9044 33348
rect 8988 33294 8990 33346
rect 8990 33294 9042 33346
rect 9042 33294 9044 33346
rect 8988 33292 9044 33294
rect 8204 31948 8260 32004
rect 7868 31666 7924 31668
rect 7868 31614 7870 31666
rect 7870 31614 7922 31666
rect 7922 31614 7924 31666
rect 7868 31612 7924 31614
rect 8428 31612 8484 31668
rect 8764 31724 8820 31780
rect 7756 30716 7812 30772
rect 8540 31554 8596 31556
rect 8540 31502 8542 31554
rect 8542 31502 8594 31554
rect 8594 31502 8596 31554
rect 8540 31500 8596 31502
rect 7756 30156 7812 30212
rect 6524 29372 6580 29428
rect 4732 29314 4788 29316
rect 4732 29262 4734 29314
rect 4734 29262 4786 29314
rect 4786 29262 4788 29314
rect 4732 29260 4788 29262
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4956 28812 5012 28868
rect 7308 29426 7364 29428
rect 7308 29374 7310 29426
rect 7310 29374 7362 29426
rect 7362 29374 7364 29426
rect 7308 29372 7364 29374
rect 7756 29426 7812 29428
rect 7756 29374 7758 29426
rect 7758 29374 7810 29426
rect 7810 29374 7812 29426
rect 7756 29372 7812 29374
rect 7084 28700 7140 28756
rect 6972 28642 7028 28644
rect 6972 28590 6974 28642
rect 6974 28590 7026 28642
rect 7026 28590 7028 28642
rect 6972 28588 7028 28590
rect 9660 35196 9716 35252
rect 9996 38556 10052 38612
rect 11004 42028 11060 42084
rect 11004 40572 11060 40628
rect 11676 42476 11732 42532
rect 11452 41916 11508 41972
rect 15036 43708 15092 43764
rect 14140 43426 14196 43428
rect 14140 43374 14142 43426
rect 14142 43374 14194 43426
rect 14194 43374 14196 43426
rect 14140 43372 14196 43374
rect 16380 44322 16436 44324
rect 16380 44270 16382 44322
rect 16382 44270 16434 44322
rect 16434 44270 16436 44322
rect 16380 44268 16436 44270
rect 17724 45218 17780 45220
rect 17724 45166 17726 45218
rect 17726 45166 17778 45218
rect 17778 45166 17780 45218
rect 17724 45164 17780 45166
rect 17612 44604 17668 44660
rect 17052 44322 17108 44324
rect 17052 44270 17054 44322
rect 17054 44270 17106 44322
rect 17106 44270 17108 44322
rect 17052 44268 17108 44270
rect 18172 45276 18228 45332
rect 18060 44604 18116 44660
rect 16268 44098 16324 44100
rect 16268 44046 16270 44098
rect 16270 44046 16322 44098
rect 16322 44046 16324 44098
rect 16268 44044 16324 44046
rect 15260 43372 15316 43428
rect 16268 43426 16324 43428
rect 16268 43374 16270 43426
rect 16270 43374 16322 43426
rect 16322 43374 16324 43426
rect 16268 43372 16324 43374
rect 17836 44210 17892 44212
rect 17836 44158 17838 44210
rect 17838 44158 17890 44210
rect 17890 44158 17892 44210
rect 17836 44156 17892 44158
rect 11900 42028 11956 42084
rect 12908 42028 12964 42084
rect 12796 41468 12852 41524
rect 13244 42028 13300 42084
rect 13132 41804 13188 41860
rect 12572 41074 12628 41076
rect 12572 41022 12574 41074
rect 12574 41022 12626 41074
rect 12626 41022 12628 41074
rect 12572 41020 12628 41022
rect 12796 40962 12852 40964
rect 12796 40910 12798 40962
rect 12798 40910 12850 40962
rect 12850 40910 12852 40962
rect 12796 40908 12852 40910
rect 11900 40572 11956 40628
rect 11116 39788 11172 39844
rect 10780 39452 10836 39508
rect 11452 40348 11508 40404
rect 13020 40460 13076 40516
rect 10892 38722 10948 38724
rect 10892 38670 10894 38722
rect 10894 38670 10946 38722
rect 10946 38670 10948 38722
rect 10892 38668 10948 38670
rect 11900 40402 11956 40404
rect 11900 40350 11902 40402
rect 11902 40350 11954 40402
rect 11954 40350 11956 40402
rect 11900 40348 11956 40350
rect 12236 40348 12292 40404
rect 12012 39506 12068 39508
rect 12012 39454 12014 39506
rect 12014 39454 12066 39506
rect 12066 39454 12068 39506
rect 12012 39452 12068 39454
rect 12012 38834 12068 38836
rect 12012 38782 12014 38834
rect 12014 38782 12066 38834
rect 12066 38782 12068 38834
rect 12012 38780 12068 38782
rect 11900 38722 11956 38724
rect 11900 38670 11902 38722
rect 11902 38670 11954 38722
rect 11954 38670 11956 38722
rect 11900 38668 11956 38670
rect 10108 38108 10164 38164
rect 9996 37884 10052 37940
rect 9772 34860 9828 34916
rect 9660 34748 9716 34804
rect 9884 34802 9940 34804
rect 9884 34750 9886 34802
rect 9886 34750 9938 34802
rect 9938 34750 9940 34802
rect 9884 34748 9940 34750
rect 9884 34412 9940 34468
rect 9436 34300 9492 34356
rect 9772 34354 9828 34356
rect 9772 34302 9774 34354
rect 9774 34302 9826 34354
rect 9826 34302 9828 34354
rect 9772 34300 9828 34302
rect 9548 34130 9604 34132
rect 9548 34078 9550 34130
rect 9550 34078 9602 34130
rect 9602 34078 9604 34130
rect 9548 34076 9604 34078
rect 9660 33122 9716 33124
rect 9660 33070 9662 33122
rect 9662 33070 9714 33122
rect 9714 33070 9716 33122
rect 9660 33068 9716 33070
rect 9436 32732 9492 32788
rect 9996 33122 10052 33124
rect 9996 33070 9998 33122
rect 9998 33070 10050 33122
rect 10050 33070 10052 33122
rect 9996 33068 10052 33070
rect 11116 38162 11172 38164
rect 11116 38110 11118 38162
rect 11118 38110 11170 38162
rect 11170 38110 11172 38162
rect 11116 38108 11172 38110
rect 11116 37772 11172 37828
rect 10220 36988 10276 37044
rect 10220 36482 10276 36484
rect 10220 36430 10222 36482
rect 10222 36430 10274 36482
rect 10274 36430 10276 36482
rect 10220 36428 10276 36430
rect 10332 36370 10388 36372
rect 10332 36318 10334 36370
rect 10334 36318 10386 36370
rect 10386 36318 10388 36370
rect 10332 36316 10388 36318
rect 10780 36316 10836 36372
rect 10668 34914 10724 34916
rect 10668 34862 10670 34914
rect 10670 34862 10722 34914
rect 10722 34862 10724 34914
rect 10668 34860 10724 34862
rect 10556 34748 10612 34804
rect 10668 34242 10724 34244
rect 10668 34190 10670 34242
rect 10670 34190 10722 34242
rect 10722 34190 10724 34242
rect 10668 34188 10724 34190
rect 10556 33068 10612 33124
rect 10332 32956 10388 33012
rect 10892 36258 10948 36260
rect 10892 36206 10894 36258
rect 10894 36206 10946 36258
rect 10946 36206 10948 36258
rect 10892 36204 10948 36206
rect 11452 37100 11508 37156
rect 11004 34748 11060 34804
rect 11564 36428 11620 36484
rect 13468 42252 13524 42308
rect 13692 42530 13748 42532
rect 13692 42478 13694 42530
rect 13694 42478 13746 42530
rect 13746 42478 13748 42530
rect 13692 42476 13748 42478
rect 14588 42252 14644 42308
rect 13580 42140 13636 42196
rect 13468 41804 13524 41860
rect 13244 41468 13300 41524
rect 13580 41298 13636 41300
rect 13580 41246 13582 41298
rect 13582 41246 13634 41298
rect 13634 41246 13636 41298
rect 13580 41244 13636 41246
rect 14028 41244 14084 41300
rect 13804 41074 13860 41076
rect 13804 41022 13806 41074
rect 13806 41022 13858 41074
rect 13858 41022 13860 41074
rect 13804 41020 13860 41022
rect 14252 40908 14308 40964
rect 13020 39564 13076 39620
rect 13692 39004 13748 39060
rect 12796 38834 12852 38836
rect 12796 38782 12798 38834
rect 12798 38782 12850 38834
rect 12850 38782 12852 38834
rect 12796 38780 12852 38782
rect 11900 36204 11956 36260
rect 12236 37548 12292 37604
rect 13804 38668 13860 38724
rect 13916 38780 13972 38836
rect 14476 42082 14532 42084
rect 14476 42030 14478 42082
rect 14478 42030 14530 42082
rect 14530 42030 14532 42082
rect 14476 42028 14532 42030
rect 15372 42082 15428 42084
rect 15372 42030 15374 42082
rect 15374 42030 15426 42082
rect 15426 42030 15428 42082
rect 15372 42028 15428 42030
rect 16268 42028 16324 42084
rect 15596 41970 15652 41972
rect 15596 41918 15598 41970
rect 15598 41918 15650 41970
rect 15650 41918 15652 41970
rect 15596 41916 15652 41918
rect 14588 41020 14644 41076
rect 16492 41916 16548 41972
rect 16604 42140 16660 42196
rect 16380 41244 16436 41300
rect 16604 41356 16660 41412
rect 16380 41074 16436 41076
rect 16380 41022 16382 41074
rect 16382 41022 16434 41074
rect 16434 41022 16436 41074
rect 16380 41020 16436 41022
rect 16156 40908 16212 40964
rect 16716 40962 16772 40964
rect 16716 40910 16718 40962
rect 16718 40910 16770 40962
rect 16770 40910 16772 40962
rect 16716 40908 16772 40910
rect 18060 41298 18116 41300
rect 18060 41246 18062 41298
rect 18062 41246 18114 41298
rect 18114 41246 18116 41298
rect 18060 41244 18116 41246
rect 17500 41132 17556 41188
rect 17948 41020 18004 41076
rect 16604 40572 16660 40628
rect 14700 40402 14756 40404
rect 14700 40350 14702 40402
rect 14702 40350 14754 40402
rect 14754 40350 14756 40402
rect 14700 40348 14756 40350
rect 14588 39564 14644 39620
rect 14364 39004 14420 39060
rect 13468 37490 13524 37492
rect 13468 37438 13470 37490
rect 13470 37438 13522 37490
rect 13522 37438 13524 37490
rect 13468 37436 13524 37438
rect 14700 39340 14756 39396
rect 15372 39340 15428 39396
rect 14588 38780 14644 38836
rect 17388 40402 17444 40404
rect 17388 40350 17390 40402
rect 17390 40350 17442 40402
rect 17442 40350 17444 40402
rect 17388 40348 17444 40350
rect 19628 45612 19684 45668
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 21084 45666 21140 45668
rect 21084 45614 21086 45666
rect 21086 45614 21138 45666
rect 21138 45614 21140 45666
rect 21084 45612 21140 45614
rect 20748 45276 20804 45332
rect 26796 46002 26852 46004
rect 26796 45950 26798 46002
rect 26798 45950 26850 46002
rect 26850 45950 26852 46002
rect 26796 45948 26852 45950
rect 27132 45890 27188 45892
rect 27132 45838 27134 45890
rect 27134 45838 27186 45890
rect 27186 45838 27188 45890
rect 27132 45836 27188 45838
rect 18956 45106 19012 45108
rect 18956 45054 18958 45106
rect 18958 45054 19010 45106
rect 19010 45054 19012 45106
rect 18956 45052 19012 45054
rect 19292 45052 19348 45108
rect 18956 44828 19012 44884
rect 19628 44268 19684 44324
rect 20188 45106 20244 45108
rect 20188 45054 20190 45106
rect 20190 45054 20242 45106
rect 20242 45054 20244 45106
rect 20188 45052 20244 45054
rect 20748 45052 20804 45108
rect 20636 44994 20692 44996
rect 20636 44942 20638 44994
rect 20638 44942 20690 44994
rect 20690 44942 20692 44994
rect 20636 44940 20692 44942
rect 20412 44882 20468 44884
rect 20412 44830 20414 44882
rect 20414 44830 20466 44882
rect 20466 44830 20468 44882
rect 20412 44828 20468 44830
rect 19964 44492 20020 44548
rect 20524 44492 20580 44548
rect 20412 44322 20468 44324
rect 20412 44270 20414 44322
rect 20414 44270 20466 44322
rect 20466 44270 20468 44322
rect 20412 44268 20468 44270
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 20748 44044 20804 44100
rect 21308 44994 21364 44996
rect 21308 44942 21310 44994
rect 21310 44942 21362 44994
rect 21362 44942 21364 44994
rect 21308 44940 21364 44942
rect 21532 44828 21588 44884
rect 21308 44492 21364 44548
rect 21980 45106 22036 45108
rect 21980 45054 21982 45106
rect 21982 45054 22034 45106
rect 22034 45054 22036 45106
rect 21980 45052 22036 45054
rect 21644 43708 21700 43764
rect 21868 44268 21924 44324
rect 19516 43372 19572 43428
rect 22092 44156 22148 44212
rect 22204 44098 22260 44100
rect 22204 44046 22206 44098
rect 22206 44046 22258 44098
rect 22258 44046 22260 44098
rect 22204 44044 22260 44046
rect 26796 45052 26852 45108
rect 22540 43708 22596 43764
rect 21420 43314 21476 43316
rect 21420 43262 21422 43314
rect 21422 43262 21474 43314
rect 21474 43262 21476 43314
rect 21420 43260 21476 43262
rect 20972 42812 21028 42868
rect 22764 43260 22820 43316
rect 19516 42252 19572 42308
rect 23436 44156 23492 44212
rect 24332 43708 24388 43764
rect 23436 43260 23492 43316
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 18732 41132 18788 41188
rect 18284 40796 18340 40852
rect 17724 39676 17780 39732
rect 16828 39452 16884 39508
rect 16044 38722 16100 38724
rect 16044 38670 16046 38722
rect 16046 38670 16098 38722
rect 16098 38670 16100 38722
rect 16044 38668 16100 38670
rect 18396 40572 18452 40628
rect 18172 39228 18228 39284
rect 17948 39116 18004 39172
rect 19292 41132 19348 41188
rect 18732 39788 18788 39844
rect 19516 41186 19572 41188
rect 19516 41134 19518 41186
rect 19518 41134 19570 41186
rect 19570 41134 19572 41186
rect 19516 41132 19572 41134
rect 19964 42140 20020 42196
rect 20636 41970 20692 41972
rect 20636 41918 20638 41970
rect 20638 41918 20690 41970
rect 20690 41918 20692 41970
rect 20636 41916 20692 41918
rect 22204 41970 22260 41972
rect 22204 41918 22206 41970
rect 22206 41918 22258 41970
rect 22258 41918 22260 41970
rect 22204 41916 22260 41918
rect 21196 41804 21252 41860
rect 19964 41356 20020 41412
rect 19852 40962 19908 40964
rect 19852 40910 19854 40962
rect 19854 40910 19906 40962
rect 19906 40910 19908 40962
rect 19852 40908 19908 40910
rect 19068 40796 19124 40852
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 19068 40402 19124 40404
rect 19068 40350 19070 40402
rect 19070 40350 19122 40402
rect 19122 40350 19124 40402
rect 19068 40348 19124 40350
rect 20972 40572 21028 40628
rect 19628 40514 19684 40516
rect 19628 40462 19630 40514
rect 19630 40462 19682 40514
rect 19682 40462 19684 40514
rect 19628 40460 19684 40462
rect 19852 40514 19908 40516
rect 19852 40462 19854 40514
rect 19854 40462 19906 40514
rect 19906 40462 19908 40514
rect 19852 40460 19908 40462
rect 19404 40348 19460 40404
rect 20188 40402 20244 40404
rect 20188 40350 20190 40402
rect 20190 40350 20242 40402
rect 20242 40350 20244 40402
rect 20188 40348 20244 40350
rect 18844 39676 18900 39732
rect 19180 39788 19236 39844
rect 18620 39506 18676 39508
rect 18620 39454 18622 39506
rect 18622 39454 18674 39506
rect 18674 39454 18676 39506
rect 18620 39452 18676 39454
rect 18844 39394 18900 39396
rect 18844 39342 18846 39394
rect 18846 39342 18898 39394
rect 18898 39342 18900 39394
rect 18844 39340 18900 39342
rect 18620 39116 18676 39172
rect 16268 38444 16324 38500
rect 14476 37548 14532 37604
rect 12460 37378 12516 37380
rect 12460 37326 12462 37378
rect 12462 37326 12514 37378
rect 12514 37326 12516 37378
rect 12460 37324 12516 37326
rect 11452 34412 11508 34468
rect 11228 34354 11284 34356
rect 11228 34302 11230 34354
rect 11230 34302 11282 34354
rect 11282 34302 11284 34354
rect 11228 34300 11284 34302
rect 11788 34242 11844 34244
rect 11788 34190 11790 34242
rect 11790 34190 11842 34242
rect 11842 34190 11844 34242
rect 11788 34188 11844 34190
rect 11116 34130 11172 34132
rect 11116 34078 11118 34130
rect 11118 34078 11170 34130
rect 11170 34078 11172 34130
rect 11116 34076 11172 34078
rect 11228 33964 11284 34020
rect 11228 32732 11284 32788
rect 12348 37212 12404 37268
rect 13244 37212 13300 37268
rect 12460 36482 12516 36484
rect 12460 36430 12462 36482
rect 12462 36430 12514 36482
rect 12514 36430 12516 36482
rect 12460 36428 12516 36430
rect 12908 36258 12964 36260
rect 12908 36206 12910 36258
rect 12910 36206 12962 36258
rect 12962 36206 12964 36258
rect 12908 36204 12964 36206
rect 14028 37266 14084 37268
rect 14028 37214 14030 37266
rect 14030 37214 14082 37266
rect 14082 37214 14084 37266
rect 14028 37212 14084 37214
rect 14140 36428 14196 36484
rect 13916 35922 13972 35924
rect 13916 35870 13918 35922
rect 13918 35870 13970 35922
rect 13970 35870 13972 35922
rect 13916 35868 13972 35870
rect 14588 37436 14644 37492
rect 15820 37324 15876 37380
rect 15820 37100 15876 37156
rect 15036 36988 15092 37044
rect 15148 36482 15204 36484
rect 15148 36430 15150 36482
rect 15150 36430 15202 36482
rect 15202 36430 15204 36482
rect 15148 36428 15204 36430
rect 14364 35644 14420 35700
rect 14028 35420 14084 35476
rect 14476 36204 14532 36260
rect 14700 35868 14756 35924
rect 14252 34690 14308 34692
rect 14252 34638 14254 34690
rect 14254 34638 14306 34690
rect 14306 34638 14308 34690
rect 14252 34636 14308 34638
rect 13132 34300 13188 34356
rect 11788 32732 11844 32788
rect 10556 31836 10612 31892
rect 9660 31724 9716 31780
rect 9884 31612 9940 31668
rect 9100 31388 9156 31444
rect 9548 31388 9604 31444
rect 9660 30994 9716 30996
rect 9660 30942 9662 30994
rect 9662 30942 9714 30994
rect 9714 30942 9716 30994
rect 9660 30940 9716 30942
rect 11004 31836 11060 31892
rect 11564 31666 11620 31668
rect 11564 31614 11566 31666
rect 11566 31614 11618 31666
rect 11618 31614 11620 31666
rect 11564 31612 11620 31614
rect 10892 31500 10948 31556
rect 11228 31276 11284 31332
rect 9884 30716 9940 30772
rect 14364 34300 14420 34356
rect 13580 34130 13636 34132
rect 13580 34078 13582 34130
rect 13582 34078 13634 34130
rect 13634 34078 13636 34130
rect 13580 34076 13636 34078
rect 12684 33404 12740 33460
rect 13132 33404 13188 33460
rect 13580 33458 13636 33460
rect 13580 33406 13582 33458
rect 13582 33406 13634 33458
rect 13634 33406 13636 33458
rect 13580 33404 13636 33406
rect 14812 35420 14868 35476
rect 15036 34860 15092 34916
rect 14700 34130 14756 34132
rect 14700 34078 14702 34130
rect 14702 34078 14754 34130
rect 14754 34078 14756 34130
rect 14700 34076 14756 34078
rect 15260 34076 15316 34132
rect 13916 33404 13972 33460
rect 14028 33346 14084 33348
rect 14028 33294 14030 33346
rect 14030 33294 14082 33346
rect 14082 33294 14084 33346
rect 14028 33292 14084 33294
rect 14924 32674 14980 32676
rect 14924 32622 14926 32674
rect 14926 32622 14978 32674
rect 14978 32622 14980 32674
rect 14924 32620 14980 32622
rect 15148 32956 15204 33012
rect 14924 31836 14980 31892
rect 12124 31778 12180 31780
rect 12124 31726 12126 31778
rect 12126 31726 12178 31778
rect 12178 31726 12180 31778
rect 12124 31724 12180 31726
rect 12572 31778 12628 31780
rect 12572 31726 12574 31778
rect 12574 31726 12626 31778
rect 12626 31726 12628 31778
rect 12572 31724 12628 31726
rect 14140 31666 14196 31668
rect 14140 31614 14142 31666
rect 14142 31614 14194 31666
rect 14194 31614 14196 31666
rect 14140 31612 14196 31614
rect 14476 31612 14532 31668
rect 12012 31554 12068 31556
rect 12012 31502 12014 31554
rect 12014 31502 12066 31554
rect 12066 31502 12068 31554
rect 12012 31500 12068 31502
rect 12460 31106 12516 31108
rect 12460 31054 12462 31106
rect 12462 31054 12514 31106
rect 12514 31054 12516 31106
rect 12460 31052 12516 31054
rect 12348 30940 12404 30996
rect 11676 30716 11732 30772
rect 13468 30940 13524 30996
rect 12684 30716 12740 30772
rect 8988 30434 9044 30436
rect 8988 30382 8990 30434
rect 8990 30382 9042 30434
rect 9042 30382 9044 30434
rect 8988 30380 9044 30382
rect 9884 30380 9940 30436
rect 7868 28700 7924 28756
rect 8092 29260 8148 29316
rect 8316 29202 8372 29204
rect 8316 29150 8318 29202
rect 8318 29150 8370 29202
rect 8370 29150 8372 29202
rect 8316 29148 8372 29150
rect 8540 29314 8596 29316
rect 8540 29262 8542 29314
rect 8542 29262 8594 29314
rect 8594 29262 8596 29314
rect 8540 29260 8596 29262
rect 9212 30210 9268 30212
rect 9212 30158 9214 30210
rect 9214 30158 9266 30210
rect 9266 30158 9268 30210
rect 9212 30156 9268 30158
rect 8764 29372 8820 29428
rect 10444 30380 10500 30436
rect 13804 30828 13860 30884
rect 10556 29148 10612 29204
rect 12796 29986 12852 29988
rect 12796 29934 12798 29986
rect 12798 29934 12850 29986
rect 12850 29934 12852 29986
rect 12796 29932 12852 29934
rect 13580 29986 13636 29988
rect 13580 29934 13582 29986
rect 13582 29934 13634 29986
rect 13634 29934 13636 29986
rect 13580 29932 13636 29934
rect 11452 29820 11508 29876
rect 8652 28588 8708 28644
rect 8988 27858 9044 27860
rect 8988 27806 8990 27858
rect 8990 27806 9042 27858
rect 9042 27806 9044 27858
rect 8988 27804 9044 27806
rect 11228 28642 11284 28644
rect 11228 28590 11230 28642
rect 11230 28590 11282 28642
rect 11282 28590 11284 28642
rect 11228 28588 11284 28590
rect 12124 28588 12180 28644
rect 12572 28642 12628 28644
rect 12572 28590 12574 28642
rect 12574 28590 12626 28642
rect 12626 28590 12628 28642
rect 12572 28588 12628 28590
rect 12348 28530 12404 28532
rect 12348 28478 12350 28530
rect 12350 28478 12402 28530
rect 12402 28478 12404 28530
rect 12348 28476 12404 28478
rect 12012 28364 12068 28420
rect 12796 28642 12852 28644
rect 12796 28590 12798 28642
rect 12798 28590 12850 28642
rect 12850 28590 12852 28642
rect 12796 28588 12852 28590
rect 14364 30882 14420 30884
rect 14364 30830 14366 30882
rect 14366 30830 14418 30882
rect 14418 30830 14420 30882
rect 14364 30828 14420 30830
rect 15036 31666 15092 31668
rect 15036 31614 15038 31666
rect 15038 31614 15090 31666
rect 15090 31614 15092 31666
rect 15036 31612 15092 31614
rect 14588 30098 14644 30100
rect 14588 30046 14590 30098
rect 14590 30046 14642 30098
rect 14642 30046 14644 30098
rect 14588 30044 14644 30046
rect 15708 33570 15764 33572
rect 15708 33518 15710 33570
rect 15710 33518 15762 33570
rect 15762 33518 15764 33570
rect 15708 33516 15764 33518
rect 15708 32562 15764 32564
rect 15708 32510 15710 32562
rect 15710 32510 15762 32562
rect 15762 32510 15764 32562
rect 15708 32508 15764 32510
rect 16492 37548 16548 37604
rect 16716 37324 16772 37380
rect 16268 37266 16324 37268
rect 16268 37214 16270 37266
rect 16270 37214 16322 37266
rect 16322 37214 16324 37266
rect 16268 37212 16324 37214
rect 16380 37154 16436 37156
rect 16380 37102 16382 37154
rect 16382 37102 16434 37154
rect 16434 37102 16436 37154
rect 16380 37100 16436 37102
rect 16156 36988 16212 37044
rect 16268 35698 16324 35700
rect 16268 35646 16270 35698
rect 16270 35646 16322 35698
rect 16322 35646 16324 35698
rect 16268 35644 16324 35646
rect 16604 35810 16660 35812
rect 16604 35758 16606 35810
rect 16606 35758 16658 35810
rect 16658 35758 16660 35810
rect 16604 35756 16660 35758
rect 16492 35420 16548 35476
rect 16492 33458 16548 33460
rect 16492 33406 16494 33458
rect 16494 33406 16546 33458
rect 16546 33406 16548 33458
rect 16492 33404 16548 33406
rect 16716 33740 16772 33796
rect 16828 33346 16884 33348
rect 16828 33294 16830 33346
rect 16830 33294 16882 33346
rect 16882 33294 16884 33346
rect 16828 33292 16884 33294
rect 16380 33180 16436 33236
rect 16492 32844 16548 32900
rect 16380 32674 16436 32676
rect 16380 32622 16382 32674
rect 16382 32622 16434 32674
rect 16434 32622 16436 32674
rect 16380 32620 16436 32622
rect 16716 32508 16772 32564
rect 16268 31836 16324 31892
rect 15596 31724 15652 31780
rect 15484 31666 15540 31668
rect 15484 31614 15486 31666
rect 15486 31614 15538 31666
rect 15538 31614 15540 31666
rect 15484 31612 15540 31614
rect 15932 31218 15988 31220
rect 15932 31166 15934 31218
rect 15934 31166 15986 31218
rect 15986 31166 15988 31218
rect 15932 31164 15988 31166
rect 15596 31106 15652 31108
rect 15596 31054 15598 31106
rect 15598 31054 15650 31106
rect 15650 31054 15652 31106
rect 15596 31052 15652 31054
rect 17388 37826 17444 37828
rect 17388 37774 17390 37826
rect 17390 37774 17442 37826
rect 17442 37774 17444 37826
rect 17388 37772 17444 37774
rect 17500 37660 17556 37716
rect 17388 36988 17444 37044
rect 17612 37212 17668 37268
rect 18060 37548 18116 37604
rect 17948 37154 18004 37156
rect 17948 37102 17950 37154
rect 17950 37102 18002 37154
rect 18002 37102 18004 37154
rect 17948 37100 18004 37102
rect 17948 35756 18004 35812
rect 18060 35644 18116 35700
rect 18172 37212 18228 37268
rect 17836 35196 17892 35252
rect 17948 35420 18004 35476
rect 17388 34914 17444 34916
rect 17388 34862 17390 34914
rect 17390 34862 17442 34914
rect 17442 34862 17444 34914
rect 17388 34860 17444 34862
rect 17276 33346 17332 33348
rect 17276 33294 17278 33346
rect 17278 33294 17330 33346
rect 17330 33294 17332 33346
rect 17276 33292 17332 33294
rect 17500 33516 17556 33572
rect 17948 33964 18004 34020
rect 17948 33516 18004 33572
rect 17836 33180 17892 33236
rect 17724 33068 17780 33124
rect 17164 31724 17220 31780
rect 17836 32562 17892 32564
rect 17836 32510 17838 32562
rect 17838 32510 17890 32562
rect 17890 32510 17892 32562
rect 17836 32508 17892 32510
rect 18508 38668 18564 38724
rect 19180 39228 19236 39284
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 19852 38668 19908 38724
rect 20412 38668 20468 38724
rect 19292 38444 19348 38500
rect 20076 38444 20132 38500
rect 19068 37266 19124 37268
rect 19068 37214 19070 37266
rect 19070 37214 19122 37266
rect 19122 37214 19124 37266
rect 19068 37212 19124 37214
rect 19628 37660 19684 37716
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 20300 37266 20356 37268
rect 20300 37214 20302 37266
rect 20302 37214 20354 37266
rect 20354 37214 20356 37266
rect 20300 37212 20356 37214
rect 19180 36652 19236 36708
rect 18620 36594 18676 36596
rect 18620 36542 18622 36594
rect 18622 36542 18674 36594
rect 18674 36542 18676 36594
rect 18620 36540 18676 36542
rect 18284 36370 18340 36372
rect 18284 36318 18286 36370
rect 18286 36318 18338 36370
rect 18338 36318 18340 36370
rect 18284 36316 18340 36318
rect 19516 36540 19572 36596
rect 18956 36370 19012 36372
rect 18956 36318 18958 36370
rect 18958 36318 19010 36370
rect 19010 36318 19012 36370
rect 18956 36316 19012 36318
rect 18508 35756 18564 35812
rect 18396 34748 18452 34804
rect 18620 35698 18676 35700
rect 18620 35646 18622 35698
rect 18622 35646 18674 35698
rect 18674 35646 18676 35698
rect 18620 35644 18676 35646
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19292 35420 19348 35476
rect 20188 35698 20244 35700
rect 20188 35646 20190 35698
rect 20190 35646 20242 35698
rect 20242 35646 20244 35698
rect 20188 35644 20244 35646
rect 20076 35420 20132 35476
rect 18844 35196 18900 35252
rect 18956 34690 19012 34692
rect 18956 34638 18958 34690
rect 18958 34638 19010 34690
rect 19010 34638 19012 34690
rect 18956 34636 19012 34638
rect 19516 34802 19572 34804
rect 19516 34750 19518 34802
rect 19518 34750 19570 34802
rect 19570 34750 19572 34802
rect 19516 34748 19572 34750
rect 20076 34802 20132 34804
rect 20076 34750 20078 34802
rect 20078 34750 20130 34802
rect 20130 34750 20132 34802
rect 20076 34748 20132 34750
rect 18844 34018 18900 34020
rect 18844 33966 18846 34018
rect 18846 33966 18898 34018
rect 18898 33966 18900 34018
rect 18844 33964 18900 33966
rect 18508 33740 18564 33796
rect 18844 33740 18900 33796
rect 19068 33122 19124 33124
rect 19068 33070 19070 33122
rect 19070 33070 19122 33122
rect 19122 33070 19124 33122
rect 19068 33068 19124 33070
rect 18620 32844 18676 32900
rect 18396 32786 18452 32788
rect 18396 32734 18398 32786
rect 18398 32734 18450 32786
rect 18450 32734 18452 32786
rect 18396 32732 18452 32734
rect 18284 32674 18340 32676
rect 18284 32622 18286 32674
rect 18286 32622 18338 32674
rect 18338 32622 18340 32674
rect 18284 32620 18340 32622
rect 18172 31778 18228 31780
rect 18172 31726 18174 31778
rect 18174 31726 18226 31778
rect 18226 31726 18228 31778
rect 18172 31724 18228 31726
rect 19404 33346 19460 33348
rect 19404 33294 19406 33346
rect 19406 33294 19458 33346
rect 19458 33294 19460 33346
rect 19404 33292 19460 33294
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 20300 34130 20356 34132
rect 20300 34078 20302 34130
rect 20302 34078 20354 34130
rect 20354 34078 20356 34130
rect 20300 34076 20356 34078
rect 20860 38108 20916 38164
rect 20748 36594 20804 36596
rect 20748 36542 20750 36594
rect 20750 36542 20802 36594
rect 20802 36542 20804 36594
rect 20748 36540 20804 36542
rect 20636 36316 20692 36372
rect 20524 35698 20580 35700
rect 20524 35646 20526 35698
rect 20526 35646 20578 35698
rect 20578 35646 20580 35698
rect 20524 35644 20580 35646
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 19180 32620 19236 32676
rect 19964 32562 20020 32564
rect 19964 32510 19966 32562
rect 19966 32510 20018 32562
rect 20018 32510 20020 32562
rect 19964 32508 20020 32510
rect 19292 31666 19348 31668
rect 19292 31614 19294 31666
rect 19294 31614 19346 31666
rect 19346 31614 19348 31666
rect 19292 31612 19348 31614
rect 16268 31052 16324 31108
rect 16828 31276 16884 31332
rect 16492 30940 16548 30996
rect 15260 30156 15316 30212
rect 16044 30268 16100 30324
rect 14028 29260 14084 29316
rect 14140 29148 14196 29204
rect 13580 28530 13636 28532
rect 13580 28478 13582 28530
rect 13582 28478 13634 28530
rect 13634 28478 13636 28530
rect 13580 28476 13636 28478
rect 12908 28364 12964 28420
rect 13804 28364 13860 28420
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 1932 27186 1988 27188
rect 1932 27134 1934 27186
rect 1934 27134 1986 27186
rect 1986 27134 1988 27186
rect 1932 27132 1988 27134
rect 14364 28642 14420 28644
rect 14364 28590 14366 28642
rect 14366 28590 14418 28642
rect 14418 28590 14420 28642
rect 14364 28588 14420 28590
rect 14140 27244 14196 27300
rect 12348 26962 12404 26964
rect 12348 26910 12350 26962
rect 12350 26910 12402 26962
rect 12402 26910 12404 26962
rect 12348 26908 12404 26910
rect 15932 29650 15988 29652
rect 15932 29598 15934 29650
rect 15934 29598 15986 29650
rect 15986 29598 15988 29650
rect 15932 29596 15988 29598
rect 16604 31164 16660 31220
rect 16268 29932 16324 29988
rect 16604 30210 16660 30212
rect 16604 30158 16606 30210
rect 16606 30158 16658 30210
rect 16658 30158 16660 30210
rect 16604 30156 16660 30158
rect 16940 30380 16996 30436
rect 16380 29484 16436 29540
rect 15708 29426 15764 29428
rect 15708 29374 15710 29426
rect 15710 29374 15762 29426
rect 15762 29374 15764 29426
rect 15708 29372 15764 29374
rect 17164 31164 17220 31220
rect 17612 31218 17668 31220
rect 17612 31166 17614 31218
rect 17614 31166 17666 31218
rect 17666 31166 17668 31218
rect 17612 31164 17668 31166
rect 17388 31106 17444 31108
rect 17388 31054 17390 31106
rect 17390 31054 17442 31106
rect 17442 31054 17444 31106
rect 17388 31052 17444 31054
rect 17836 30994 17892 30996
rect 17836 30942 17838 30994
rect 17838 30942 17890 30994
rect 17890 30942 17892 30994
rect 17836 30940 17892 30942
rect 17612 30322 17668 30324
rect 17612 30270 17614 30322
rect 17614 30270 17666 30322
rect 17666 30270 17668 30322
rect 17612 30268 17668 30270
rect 17388 30210 17444 30212
rect 17388 30158 17390 30210
rect 17390 30158 17442 30210
rect 17442 30158 17444 30210
rect 17388 30156 17444 30158
rect 19292 30940 19348 30996
rect 20412 33068 20468 33124
rect 20524 35308 20580 35364
rect 20076 31554 20132 31556
rect 20076 31502 20078 31554
rect 20078 31502 20130 31554
rect 20130 31502 20132 31554
rect 20076 31500 20132 31502
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 17948 30380 18004 30436
rect 16716 29484 16772 29540
rect 14924 27858 14980 27860
rect 14924 27806 14926 27858
rect 14926 27806 14978 27858
rect 14978 27806 14980 27858
rect 14924 27804 14980 27806
rect 14700 27468 14756 27524
rect 15260 28252 15316 28308
rect 4284 26460 4340 26516
rect 8652 26460 8708 26516
rect 1932 26178 1988 26180
rect 1932 26126 1934 26178
rect 1934 26126 1986 26178
rect 1986 26126 1988 26178
rect 1932 26124 1988 26126
rect 4284 26124 4340 26180
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 1932 25618 1988 25620
rect 1932 25566 1934 25618
rect 1934 25566 1986 25618
rect 1986 25566 1988 25618
rect 1932 25564 1988 25566
rect 12236 26850 12292 26852
rect 12236 26798 12238 26850
rect 12238 26798 12290 26850
rect 12290 26798 12292 26850
rect 12236 26796 12292 26798
rect 13580 26796 13636 26852
rect 12908 26348 12964 26404
rect 11564 26236 11620 26292
rect 4284 25506 4340 25508
rect 4284 25454 4286 25506
rect 4286 25454 4338 25506
rect 4338 25454 4340 25506
rect 4284 25452 4340 25454
rect 9548 25452 9604 25508
rect 12460 26290 12516 26292
rect 12460 26238 12462 26290
rect 12462 26238 12514 26290
rect 12514 26238 12516 26290
rect 12460 26236 12516 26238
rect 12908 26178 12964 26180
rect 12908 26126 12910 26178
rect 12910 26126 12962 26178
rect 12962 26126 12964 26178
rect 12908 26124 12964 26126
rect 10780 25394 10836 25396
rect 10780 25342 10782 25394
rect 10782 25342 10834 25394
rect 10834 25342 10836 25394
rect 10780 25340 10836 25342
rect 8652 25228 8708 25284
rect 12124 25282 12180 25284
rect 12124 25230 12126 25282
rect 12126 25230 12178 25282
rect 12178 25230 12180 25282
rect 12124 25228 12180 25230
rect 12460 25394 12516 25396
rect 12460 25342 12462 25394
rect 12462 25342 12514 25394
rect 12514 25342 12516 25394
rect 12460 25340 12516 25342
rect 14252 25788 14308 25844
rect 14140 25676 14196 25732
rect 13468 25564 13524 25620
rect 12796 25506 12852 25508
rect 12796 25454 12798 25506
rect 12798 25454 12850 25506
rect 12850 25454 12852 25506
rect 12796 25452 12852 25454
rect 12348 25228 12404 25284
rect 13132 25228 13188 25284
rect 1932 24892 1988 24948
rect 4284 24892 4340 24948
rect 4732 24946 4788 24948
rect 4732 24894 4734 24946
rect 4734 24894 4786 24946
rect 4786 24894 4788 24946
rect 4732 24892 4788 24894
rect 13692 25228 13748 25284
rect 17388 29426 17444 29428
rect 17388 29374 17390 29426
rect 17390 29374 17442 29426
rect 17442 29374 17444 29426
rect 17388 29372 17444 29374
rect 16380 28754 16436 28756
rect 16380 28702 16382 28754
rect 16382 28702 16434 28754
rect 16434 28702 16436 28754
rect 16380 28700 16436 28702
rect 16716 28476 16772 28532
rect 17052 29260 17108 29316
rect 16940 28418 16996 28420
rect 16940 28366 16942 28418
rect 16942 28366 16994 28418
rect 16994 28366 16996 28418
rect 16940 28364 16996 28366
rect 15820 27970 15876 27972
rect 15820 27918 15822 27970
rect 15822 27918 15874 27970
rect 15874 27918 15876 27970
rect 15820 27916 15876 27918
rect 16268 27298 16324 27300
rect 16268 27246 16270 27298
rect 16270 27246 16322 27298
rect 16322 27246 16324 27298
rect 16268 27244 16324 27246
rect 15260 26012 15316 26068
rect 15484 27132 15540 27188
rect 16268 26402 16324 26404
rect 16268 26350 16270 26402
rect 16270 26350 16322 26402
rect 16322 26350 16324 26402
rect 16268 26348 16324 26350
rect 16492 26348 16548 26404
rect 15708 26290 15764 26292
rect 15708 26238 15710 26290
rect 15710 26238 15762 26290
rect 15762 26238 15764 26290
rect 15708 26236 15764 26238
rect 17500 29314 17556 29316
rect 17500 29262 17502 29314
rect 17502 29262 17554 29314
rect 17554 29262 17556 29314
rect 17500 29260 17556 29262
rect 20188 30380 20244 30436
rect 19740 30210 19796 30212
rect 19740 30158 19742 30210
rect 19742 30158 19794 30210
rect 19794 30158 19796 30210
rect 19740 30156 19796 30158
rect 18732 29596 18788 29652
rect 18396 29426 18452 29428
rect 18396 29374 18398 29426
rect 18398 29374 18450 29426
rect 18450 29374 18452 29426
rect 18396 29372 18452 29374
rect 18060 28924 18116 28980
rect 18620 29148 18676 29204
rect 18060 28530 18116 28532
rect 18060 28478 18062 28530
rect 18062 28478 18114 28530
rect 18114 28478 18116 28530
rect 18060 28476 18116 28478
rect 17276 28418 17332 28420
rect 17276 28366 17278 28418
rect 17278 28366 17330 28418
rect 17330 28366 17332 28418
rect 17276 28364 17332 28366
rect 17500 28082 17556 28084
rect 17500 28030 17502 28082
rect 17502 28030 17554 28082
rect 17554 28030 17556 28082
rect 17500 28028 17556 28030
rect 17164 26572 17220 26628
rect 16828 26402 16884 26404
rect 16828 26350 16830 26402
rect 16830 26350 16882 26402
rect 16882 26350 16884 26402
rect 16828 26348 16884 26350
rect 16604 25452 16660 25508
rect 16716 25676 16772 25732
rect 18172 28418 18228 28420
rect 18172 28366 18174 28418
rect 18174 28366 18226 28418
rect 18226 28366 18228 28418
rect 18172 28364 18228 28366
rect 19628 29820 19684 29876
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19964 29484 20020 29540
rect 19292 29426 19348 29428
rect 19292 29374 19294 29426
rect 19294 29374 19346 29426
rect 19346 29374 19348 29426
rect 19292 29372 19348 29374
rect 19516 29148 19572 29204
rect 20860 34188 20916 34244
rect 20972 33292 21028 33348
rect 20972 30994 21028 30996
rect 20972 30942 20974 30994
rect 20974 30942 21026 30994
rect 21026 30942 21028 30994
rect 20972 30940 21028 30942
rect 21980 41858 22036 41860
rect 21980 41806 21982 41858
rect 21982 41806 22034 41858
rect 22034 41806 22036 41858
rect 21980 41804 22036 41806
rect 22652 41804 22708 41860
rect 21420 41020 21476 41076
rect 23324 41970 23380 41972
rect 23324 41918 23326 41970
rect 23326 41918 23378 41970
rect 23378 41918 23380 41970
rect 23324 41916 23380 41918
rect 23660 41970 23716 41972
rect 23660 41918 23662 41970
rect 23662 41918 23714 41970
rect 23714 41918 23716 41970
rect 23660 41916 23716 41918
rect 23100 41186 23156 41188
rect 23100 41134 23102 41186
rect 23102 41134 23154 41186
rect 23154 41134 23156 41186
rect 23100 41132 23156 41134
rect 22316 41074 22372 41076
rect 22316 41022 22318 41074
rect 22318 41022 22370 41074
rect 22370 41022 22372 41074
rect 22316 41020 22372 41022
rect 21644 40572 21700 40628
rect 22428 40908 22484 40964
rect 21532 40514 21588 40516
rect 21532 40462 21534 40514
rect 21534 40462 21586 40514
rect 21586 40462 21588 40514
rect 21532 40460 21588 40462
rect 22652 40348 22708 40404
rect 21980 39564 22036 39620
rect 21868 39506 21924 39508
rect 21868 39454 21870 39506
rect 21870 39454 21922 39506
rect 21922 39454 21924 39506
rect 21868 39452 21924 39454
rect 22540 39452 22596 39508
rect 21308 36652 21364 36708
rect 21532 36482 21588 36484
rect 21532 36430 21534 36482
rect 21534 36430 21586 36482
rect 21586 36430 21588 36482
rect 21532 36428 21588 36430
rect 21756 36540 21812 36596
rect 21980 38162 22036 38164
rect 21980 38110 21982 38162
rect 21982 38110 22034 38162
rect 22034 38110 22036 38162
rect 21980 38108 22036 38110
rect 22316 39340 22372 39396
rect 23660 41020 23716 41076
rect 23548 40514 23604 40516
rect 23548 40462 23550 40514
rect 23550 40462 23602 40514
rect 23602 40462 23604 40514
rect 23548 40460 23604 40462
rect 23436 40348 23492 40404
rect 23324 39564 23380 39620
rect 23100 39340 23156 39396
rect 23660 39452 23716 39508
rect 23548 38722 23604 38724
rect 23548 38670 23550 38722
rect 23550 38670 23602 38722
rect 23602 38670 23604 38722
rect 23548 38668 23604 38670
rect 23212 37436 23268 37492
rect 22092 36652 22148 36708
rect 21980 36428 22036 36484
rect 23548 37436 23604 37492
rect 23324 37266 23380 37268
rect 23324 37214 23326 37266
rect 23326 37214 23378 37266
rect 23378 37214 23380 37266
rect 23324 37212 23380 37214
rect 21868 35308 21924 35364
rect 24108 38050 24164 38052
rect 24108 37998 24110 38050
rect 24110 37998 24162 38050
rect 24162 37998 24164 38050
rect 24108 37996 24164 37998
rect 23884 37772 23940 37828
rect 23996 37042 24052 37044
rect 23996 36990 23998 37042
rect 23998 36990 24050 37042
rect 24050 36990 24052 37042
rect 23996 36988 24052 36990
rect 24332 38892 24388 38948
rect 25452 38946 25508 38948
rect 25452 38894 25454 38946
rect 25454 38894 25506 38946
rect 25506 38894 25508 38946
rect 25452 38892 25508 38894
rect 25004 38050 25060 38052
rect 25004 37998 25006 38050
rect 25006 37998 25058 38050
rect 25058 37998 25060 38050
rect 25004 37996 25060 37998
rect 25228 37772 25284 37828
rect 24444 37212 24500 37268
rect 25228 37266 25284 37268
rect 25228 37214 25230 37266
rect 25230 37214 25282 37266
rect 25282 37214 25284 37266
rect 25228 37212 25284 37214
rect 24556 36988 24612 37044
rect 25340 36988 25396 37044
rect 25788 36988 25844 37044
rect 22316 34972 22372 35028
rect 21644 34748 21700 34804
rect 21532 34242 21588 34244
rect 21532 34190 21534 34242
rect 21534 34190 21586 34242
rect 21586 34190 21588 34242
rect 21532 34188 21588 34190
rect 21420 33292 21476 33348
rect 21420 31052 21476 31108
rect 22316 34242 22372 34244
rect 22316 34190 22318 34242
rect 22318 34190 22370 34242
rect 22370 34190 22372 34242
rect 22316 34188 22372 34190
rect 22764 34860 22820 34916
rect 22988 34972 23044 35028
rect 22652 34802 22708 34804
rect 22652 34750 22654 34802
rect 22654 34750 22706 34802
rect 22706 34750 22708 34802
rect 22652 34748 22708 34750
rect 24444 35084 24500 35140
rect 23548 34972 23604 35028
rect 23772 34914 23828 34916
rect 23772 34862 23774 34914
rect 23774 34862 23826 34914
rect 23826 34862 23828 34914
rect 23772 34860 23828 34862
rect 23324 34748 23380 34804
rect 22540 33346 22596 33348
rect 22540 33294 22542 33346
rect 22542 33294 22594 33346
rect 22594 33294 22596 33346
rect 22540 33292 22596 33294
rect 21868 31052 21924 31108
rect 21644 30882 21700 30884
rect 21644 30830 21646 30882
rect 21646 30830 21698 30882
rect 21698 30830 21700 30882
rect 21644 30828 21700 30830
rect 21420 30434 21476 30436
rect 21420 30382 21422 30434
rect 21422 30382 21474 30434
rect 21474 30382 21476 30434
rect 21420 30380 21476 30382
rect 21532 30156 21588 30212
rect 18732 28588 18788 28644
rect 21420 29260 21476 29316
rect 18060 27970 18116 27972
rect 18060 27918 18062 27970
rect 18062 27918 18114 27970
rect 18114 27918 18116 27970
rect 18060 27916 18116 27918
rect 17948 27858 18004 27860
rect 17948 27806 17950 27858
rect 17950 27806 18002 27858
rect 18002 27806 18004 27858
rect 17948 27804 18004 27806
rect 17948 27186 18004 27188
rect 17948 27134 17950 27186
rect 17950 27134 18002 27186
rect 18002 27134 18004 27186
rect 17948 27132 18004 27134
rect 18956 27970 19012 27972
rect 18956 27918 18958 27970
rect 18958 27918 19010 27970
rect 19010 27918 19012 27970
rect 18956 27916 19012 27918
rect 17836 26236 17892 26292
rect 17388 25618 17444 25620
rect 17388 25566 17390 25618
rect 17390 25566 17442 25618
rect 17442 25566 17444 25618
rect 17388 25564 17444 25566
rect 18844 27858 18900 27860
rect 18844 27806 18846 27858
rect 18846 27806 18898 27858
rect 18898 27806 18900 27858
rect 18844 27804 18900 27806
rect 20188 28812 20244 28868
rect 20412 28642 20468 28644
rect 20412 28590 20414 28642
rect 20414 28590 20466 28642
rect 20466 28590 20468 28642
rect 20412 28588 20468 28590
rect 20076 28476 20132 28532
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 22204 30044 22260 30100
rect 22092 29372 22148 29428
rect 22428 30156 22484 30212
rect 22652 30940 22708 30996
rect 22988 32060 23044 32116
rect 21980 29260 22036 29316
rect 22652 29426 22708 29428
rect 22652 29374 22654 29426
rect 22654 29374 22706 29426
rect 22706 29374 22708 29426
rect 22652 29372 22708 29374
rect 22428 29148 22484 29204
rect 23212 32732 23268 32788
rect 24556 34860 24612 34916
rect 24332 34748 24388 34804
rect 24332 34130 24388 34132
rect 24332 34078 24334 34130
rect 24334 34078 24386 34130
rect 24386 34078 24388 34130
rect 24332 34076 24388 34078
rect 24780 35698 24836 35700
rect 24780 35646 24782 35698
rect 24782 35646 24834 35698
rect 24834 35646 24836 35698
rect 24780 35644 24836 35646
rect 25340 35698 25396 35700
rect 25340 35646 25342 35698
rect 25342 35646 25394 35698
rect 25394 35646 25396 35698
rect 25340 35644 25396 35646
rect 26236 36370 26292 36372
rect 26236 36318 26238 36370
rect 26238 36318 26290 36370
rect 26290 36318 26292 36370
rect 26236 36316 26292 36318
rect 25116 35084 25172 35140
rect 24892 34972 24948 35028
rect 25340 34914 25396 34916
rect 25340 34862 25342 34914
rect 25342 34862 25394 34914
rect 25394 34862 25396 34914
rect 25340 34860 25396 34862
rect 25564 34748 25620 34804
rect 26124 34860 26180 34916
rect 25900 34412 25956 34468
rect 24892 34076 24948 34132
rect 25228 34130 25284 34132
rect 25228 34078 25230 34130
rect 25230 34078 25282 34130
rect 25282 34078 25284 34130
rect 25228 34076 25284 34078
rect 23324 32450 23380 32452
rect 23324 32398 23326 32450
rect 23326 32398 23378 32450
rect 23378 32398 23380 32450
rect 23324 32396 23380 32398
rect 23548 31106 23604 31108
rect 23548 31054 23550 31106
rect 23550 31054 23602 31106
rect 23602 31054 23604 31106
rect 23548 31052 23604 31054
rect 23324 30994 23380 30996
rect 23324 30942 23326 30994
rect 23326 30942 23378 30994
rect 23378 30942 23380 30994
rect 23324 30940 23380 30942
rect 23548 30322 23604 30324
rect 23548 30270 23550 30322
rect 23550 30270 23602 30322
rect 23602 30270 23604 30322
rect 23548 30268 23604 30270
rect 23212 30156 23268 30212
rect 23324 30044 23380 30100
rect 21644 28364 21700 28420
rect 18732 27692 18788 27748
rect 20636 27746 20692 27748
rect 20636 27694 20638 27746
rect 20638 27694 20690 27746
rect 20690 27694 20692 27746
rect 20636 27692 20692 27694
rect 21532 27746 21588 27748
rect 21532 27694 21534 27746
rect 21534 27694 21586 27746
rect 21586 27694 21588 27746
rect 21532 27692 21588 27694
rect 19180 27020 19236 27076
rect 17836 25564 17892 25620
rect 17276 25506 17332 25508
rect 17276 25454 17278 25506
rect 17278 25454 17330 25506
rect 17330 25454 17332 25506
rect 17276 25452 17332 25454
rect 14252 24892 14308 24948
rect 4476 24330 4532 24332
rect 1932 24220 1988 24276
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 5292 24332 5348 24388
rect 4284 23996 4340 24052
rect 3052 23772 3108 23828
rect 1932 23548 1988 23604
rect 4620 23826 4676 23828
rect 4620 23774 4622 23826
rect 4622 23774 4674 23826
rect 4674 23774 4676 23826
rect 4620 23772 4676 23774
rect 4284 23660 4340 23716
rect 2268 22370 2324 22372
rect 2268 22318 2270 22370
rect 2270 22318 2322 22370
rect 2322 22318 2324 22370
rect 2268 22316 2324 22318
rect 2828 22370 2884 22372
rect 2828 22318 2830 22370
rect 2830 22318 2882 22370
rect 2882 22318 2884 22370
rect 2828 22316 2884 22318
rect 2492 22258 2548 22260
rect 2492 22206 2494 22258
rect 2494 22206 2546 22258
rect 2546 22206 2548 22258
rect 2492 22204 2548 22206
rect 2268 21698 2324 21700
rect 2268 21646 2270 21698
rect 2270 21646 2322 21698
rect 2322 21646 2324 21698
rect 2268 21644 2324 21646
rect 3388 22988 3444 23044
rect 3052 21644 3108 21700
rect 3164 21756 3220 21812
rect 2716 21586 2772 21588
rect 2716 21534 2718 21586
rect 2718 21534 2770 21586
rect 2770 21534 2772 21586
rect 2716 21532 2772 21534
rect 4844 23714 4900 23716
rect 4844 23662 4846 23714
rect 4846 23662 4898 23714
rect 4898 23662 4900 23714
rect 4844 23660 4900 23662
rect 4284 23154 4340 23156
rect 4284 23102 4286 23154
rect 4286 23102 4338 23154
rect 4338 23102 4340 23154
rect 4284 23100 4340 23102
rect 4732 23042 4788 23044
rect 4732 22990 4734 23042
rect 4734 22990 4786 23042
rect 4786 22990 4788 23042
rect 4732 22988 4788 22990
rect 4844 22876 4900 22932
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4732 22540 4788 22596
rect 4508 22482 4564 22484
rect 4508 22430 4510 22482
rect 4510 22430 4562 22482
rect 4562 22430 4564 22482
rect 4508 22428 4564 22430
rect 4172 22204 4228 22260
rect 3612 21644 3668 21700
rect 2940 21474 2996 21476
rect 2940 21422 2942 21474
rect 2942 21422 2994 21474
rect 2994 21422 2996 21474
rect 2940 21420 2996 21422
rect 2044 19010 2100 19012
rect 2044 18958 2046 19010
rect 2046 18958 2098 19010
rect 2098 18958 2100 19010
rect 2044 18956 2100 18958
rect 1708 18844 1764 18900
rect 2828 19068 2884 19124
rect 3276 21532 3332 21588
rect 5068 22428 5124 22484
rect 4620 21586 4676 21588
rect 4620 21534 4622 21586
rect 4622 21534 4674 21586
rect 4674 21534 4676 21586
rect 4620 21532 4676 21534
rect 4844 21586 4900 21588
rect 4844 21534 4846 21586
rect 4846 21534 4898 21586
rect 4898 21534 4900 21586
rect 4844 21532 4900 21534
rect 4284 21308 4340 21364
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 3052 20188 3108 20244
rect 3500 20188 3556 20244
rect 2716 18732 2772 18788
rect 3052 18732 3108 18788
rect 2044 18508 2100 18564
rect 1708 17500 1764 17556
rect 2604 16716 2660 16772
rect 1708 16156 1764 16212
rect 3388 19122 3444 19124
rect 3388 19070 3390 19122
rect 3390 19070 3442 19122
rect 3442 19070 3444 19122
rect 3388 19068 3444 19070
rect 2940 18562 2996 18564
rect 2940 18510 2942 18562
rect 2942 18510 2994 18562
rect 2994 18510 2996 18562
rect 2940 18508 2996 18510
rect 3388 17836 3444 17892
rect 5068 21810 5124 21812
rect 5068 21758 5070 21810
rect 5070 21758 5122 21810
rect 5122 21758 5124 21810
rect 5068 21756 5124 21758
rect 5292 23100 5348 23156
rect 5628 22540 5684 22596
rect 6972 23884 7028 23940
rect 5180 21308 5236 21364
rect 4620 20524 4676 20580
rect 6636 23660 6692 23716
rect 6188 22428 6244 22484
rect 6524 22258 6580 22260
rect 6524 22206 6526 22258
rect 6526 22206 6578 22258
rect 6578 22206 6580 22258
rect 6524 22204 6580 22206
rect 6636 21980 6692 22036
rect 5740 20524 5796 20580
rect 6188 21308 6244 21364
rect 5516 20188 5572 20244
rect 4732 20018 4788 20020
rect 4732 19966 4734 20018
rect 4734 19966 4786 20018
rect 4786 19966 4788 20018
rect 4732 19964 4788 19966
rect 5516 20018 5572 20020
rect 5516 19966 5518 20018
rect 5518 19966 5570 20018
rect 5570 19966 5572 20018
rect 5516 19964 5572 19966
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 4508 19234 4564 19236
rect 4508 19182 4510 19234
rect 4510 19182 4562 19234
rect 4562 19182 4564 19234
rect 4508 19180 4564 19182
rect 4396 19122 4452 19124
rect 4396 19070 4398 19122
rect 4398 19070 4450 19122
rect 4450 19070 4452 19122
rect 4396 19068 4452 19070
rect 3724 18732 3780 18788
rect 8540 23826 8596 23828
rect 8540 23774 8542 23826
rect 8542 23774 8594 23826
rect 8594 23774 8596 23826
rect 8540 23772 8596 23774
rect 10108 23884 10164 23940
rect 11116 23714 11172 23716
rect 11116 23662 11118 23714
rect 11118 23662 11170 23714
rect 11170 23662 11172 23714
rect 11116 23660 11172 23662
rect 7868 22876 7924 22932
rect 7196 22540 7252 22596
rect 8428 22540 8484 22596
rect 6412 20188 6468 20244
rect 8316 22204 8372 22260
rect 8092 21420 8148 21476
rect 7084 20524 7140 20580
rect 8204 20412 8260 20468
rect 6636 19964 6692 20020
rect 6524 19852 6580 19908
rect 7756 19852 7812 19908
rect 5068 19180 5124 19236
rect 5628 19122 5684 19124
rect 5628 19070 5630 19122
rect 5630 19070 5682 19122
rect 5682 19070 5684 19122
rect 5628 19068 5684 19070
rect 4956 18844 5012 18900
rect 3052 17052 3108 17108
rect 2940 16716 2996 16772
rect 3388 16716 3444 16772
rect 3500 17612 3556 17668
rect 3388 16098 3444 16100
rect 3388 16046 3390 16098
rect 3390 16046 3442 16098
rect 3442 16046 3444 16098
rect 3388 16044 3444 16046
rect 2044 15986 2100 15988
rect 2044 15934 2046 15986
rect 2046 15934 2098 15986
rect 2098 15934 2100 15986
rect 2044 15932 2100 15934
rect 2156 15820 2212 15876
rect 2716 15874 2772 15876
rect 2716 15822 2718 15874
rect 2718 15822 2770 15874
rect 2770 15822 2772 15874
rect 2716 15820 2772 15822
rect 2604 15314 2660 15316
rect 2604 15262 2606 15314
rect 2606 15262 2658 15314
rect 2658 15262 2660 15314
rect 2604 15260 2660 15262
rect 1820 14812 1876 14868
rect 3388 15484 3444 15540
rect 4172 17836 4228 17892
rect 4284 18396 4340 18452
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 4396 17836 4452 17892
rect 3948 17106 4004 17108
rect 3948 17054 3950 17106
rect 3950 17054 4002 17106
rect 4002 17054 4004 17106
rect 3948 17052 4004 17054
rect 3836 15874 3892 15876
rect 3836 15822 3838 15874
rect 3838 15822 3890 15874
rect 3890 15822 3892 15874
rect 3836 15820 3892 15822
rect 3612 15708 3668 15764
rect 5180 18732 5236 18788
rect 5964 19010 6020 19012
rect 5964 18958 5966 19010
rect 5966 18958 6018 19010
rect 6018 18958 6020 19010
rect 5964 18956 6020 18958
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 4620 16098 4676 16100
rect 4620 16046 4622 16098
rect 4622 16046 4674 16098
rect 4674 16046 4676 16098
rect 4620 16044 4676 16046
rect 2044 14252 2100 14308
rect 3724 14306 3780 14308
rect 3724 14254 3726 14306
rect 3726 14254 3778 14306
rect 3778 14254 3780 14306
rect 3724 14252 3780 14254
rect 2380 14140 2436 14196
rect 3164 14140 3220 14196
rect 2716 14028 2772 14084
rect 4956 16882 5012 16884
rect 4956 16830 4958 16882
rect 4958 16830 5010 16882
rect 5010 16830 5012 16882
rect 4956 16828 5012 16830
rect 4956 15538 5012 15540
rect 4956 15486 4958 15538
rect 4958 15486 5010 15538
rect 5010 15486 5012 15538
rect 4956 15484 5012 15486
rect 4284 15036 4340 15092
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 4956 14476 5012 14532
rect 4284 14252 4340 14308
rect 1932 13692 1988 13748
rect 1708 13468 1764 13524
rect 2044 13468 2100 13524
rect 1708 12684 1764 12740
rect 1708 12124 1764 12180
rect 1708 10780 1764 10836
rect 2380 12850 2436 12852
rect 2380 12798 2382 12850
rect 2382 12798 2434 12850
rect 2434 12798 2436 12850
rect 2380 12796 2436 12798
rect 3724 13692 3780 13748
rect 4732 13970 4788 13972
rect 4732 13918 4734 13970
rect 4734 13918 4786 13970
rect 4786 13918 4788 13970
rect 4732 13916 4788 13918
rect 5180 13916 5236 13972
rect 3948 13468 4004 13524
rect 3388 12572 3444 12628
rect 2044 12290 2100 12292
rect 2044 12238 2046 12290
rect 2046 12238 2098 12290
rect 2098 12238 2100 12290
rect 2044 12236 2100 12238
rect 2380 12012 2436 12068
rect 2380 11452 2436 11508
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 4508 12850 4564 12852
rect 4508 12798 4510 12850
rect 4510 12798 4562 12850
rect 4562 12798 4564 12850
rect 4508 12796 4564 12798
rect 4956 12738 5012 12740
rect 4956 12686 4958 12738
rect 4958 12686 5010 12738
rect 5010 12686 5012 12738
rect 4956 12684 5012 12686
rect 4284 12572 4340 12628
rect 4620 12402 4676 12404
rect 4620 12350 4622 12402
rect 4622 12350 4674 12402
rect 4674 12350 4676 12402
rect 4620 12348 4676 12350
rect 3612 11900 3668 11956
rect 2716 11116 2772 11172
rect 2044 10780 2100 10836
rect 3388 11282 3444 11284
rect 3388 11230 3390 11282
rect 3390 11230 3442 11282
rect 3442 11230 3444 11282
rect 3388 11228 3444 11230
rect 2828 10780 2884 10836
rect 2492 10722 2548 10724
rect 2492 10670 2494 10722
rect 2494 10670 2546 10722
rect 2546 10670 2548 10722
rect 2492 10668 2548 10670
rect 1820 10332 1876 10388
rect 1708 10108 1764 10164
rect 2492 10108 2548 10164
rect 1708 9436 1764 9492
rect 2044 9154 2100 9156
rect 2044 9102 2046 9154
rect 2046 9102 2098 9154
rect 2098 9102 2100 9154
rect 2044 9100 2100 9102
rect 2380 8764 2436 8820
rect 1708 8146 1764 8148
rect 1708 8094 1710 8146
rect 1710 8094 1762 8146
rect 1762 8094 1764 8146
rect 1708 8092 1764 8094
rect 3612 11452 3668 11508
rect 3052 10108 3108 10164
rect 3164 10332 3220 10388
rect 2716 9714 2772 9716
rect 2716 9662 2718 9714
rect 2718 9662 2770 9714
rect 2770 9662 2772 9714
rect 2716 9660 2772 9662
rect 3276 9324 3332 9380
rect 3500 10834 3556 10836
rect 3500 10782 3502 10834
rect 3502 10782 3554 10834
rect 3554 10782 3556 10834
rect 3500 10780 3556 10782
rect 5180 12066 5236 12068
rect 5180 12014 5182 12066
rect 5182 12014 5234 12066
rect 5234 12014 5236 12066
rect 5180 12012 5236 12014
rect 5628 18562 5684 18564
rect 5628 18510 5630 18562
rect 5630 18510 5682 18562
rect 5682 18510 5684 18562
rect 5628 18508 5684 18510
rect 6636 18060 6692 18116
rect 5628 17612 5684 17668
rect 5628 16828 5684 16884
rect 6076 16268 6132 16324
rect 5628 15932 5684 15988
rect 5628 15484 5684 15540
rect 6300 15986 6356 15988
rect 6300 15934 6302 15986
rect 6302 15934 6354 15986
rect 6354 15934 6356 15986
rect 6300 15932 6356 15934
rect 6524 16268 6580 16324
rect 7196 19068 7252 19124
rect 7532 19010 7588 19012
rect 7532 18958 7534 19010
rect 7534 18958 7586 19010
rect 7586 18958 7588 19010
rect 7532 18956 7588 18958
rect 8540 21644 8596 21700
rect 8876 22204 8932 22260
rect 8652 21420 8708 21476
rect 7868 19010 7924 19012
rect 7868 18958 7870 19010
rect 7870 18958 7922 19010
rect 7922 18958 7924 19010
rect 7868 18956 7924 18958
rect 7532 18562 7588 18564
rect 7532 18510 7534 18562
rect 7534 18510 7586 18562
rect 7586 18510 7588 18562
rect 7532 18508 7588 18510
rect 6972 18060 7028 18116
rect 6860 17836 6916 17892
rect 7308 17666 7364 17668
rect 7308 17614 7310 17666
rect 7310 17614 7362 17666
rect 7362 17614 7364 17666
rect 7308 17612 7364 17614
rect 6972 17164 7028 17220
rect 6748 16716 6804 16772
rect 7308 16098 7364 16100
rect 7308 16046 7310 16098
rect 7310 16046 7362 16098
rect 7362 16046 7364 16098
rect 7308 16044 7364 16046
rect 6300 14530 6356 14532
rect 6300 14478 6302 14530
rect 6302 14478 6354 14530
rect 6354 14478 6356 14530
rect 6300 14476 6356 14478
rect 6748 15036 6804 15092
rect 7420 15932 7476 15988
rect 7532 15708 7588 15764
rect 8316 18508 8372 18564
rect 8092 18060 8148 18116
rect 7980 17836 8036 17892
rect 8316 16994 8372 16996
rect 8316 16942 8318 16994
rect 8318 16942 8370 16994
rect 8370 16942 8372 16994
rect 8316 16940 8372 16942
rect 7868 16604 7924 16660
rect 7868 15820 7924 15876
rect 8092 15708 8148 15764
rect 9436 19852 9492 19908
rect 8764 16828 8820 16884
rect 9100 16882 9156 16884
rect 9100 16830 9102 16882
rect 9102 16830 9154 16882
rect 9154 16830 9156 16882
rect 9100 16828 9156 16830
rect 9212 16098 9268 16100
rect 9212 16046 9214 16098
rect 9214 16046 9266 16098
rect 9266 16046 9268 16098
rect 9212 16044 9268 16046
rect 8652 15372 8708 15428
rect 7868 15314 7924 15316
rect 7868 15262 7870 15314
rect 7870 15262 7922 15314
rect 7922 15262 7924 15314
rect 7868 15260 7924 15262
rect 7644 14252 7700 14308
rect 7308 14028 7364 14084
rect 10220 22092 10276 22148
rect 10108 21420 10164 21476
rect 10220 20524 10276 20580
rect 9996 18844 10052 18900
rect 9884 18732 9940 18788
rect 11228 23100 11284 23156
rect 11788 23660 11844 23716
rect 12572 24610 12628 24612
rect 12572 24558 12574 24610
rect 12574 24558 12626 24610
rect 12626 24558 12628 24610
rect 12572 24556 12628 24558
rect 14028 23938 14084 23940
rect 14028 23886 14030 23938
rect 14030 23886 14082 23938
rect 14082 23886 14084 23938
rect 14028 23884 14084 23886
rect 14252 23826 14308 23828
rect 14252 23774 14254 23826
rect 14254 23774 14306 23826
rect 14306 23774 14308 23826
rect 14252 23772 14308 23774
rect 13804 23378 13860 23380
rect 13804 23326 13806 23378
rect 13806 23326 13858 23378
rect 13858 23326 13860 23378
rect 13804 23324 13860 23326
rect 11116 22930 11172 22932
rect 11116 22878 11118 22930
rect 11118 22878 11170 22930
rect 11170 22878 11172 22930
rect 11116 22876 11172 22878
rect 13468 23154 13524 23156
rect 13468 23102 13470 23154
rect 13470 23102 13522 23154
rect 13522 23102 13524 23154
rect 13468 23100 13524 23102
rect 12124 22876 12180 22932
rect 12124 22482 12180 22484
rect 12124 22430 12126 22482
rect 12126 22430 12178 22482
rect 12178 22430 12180 22482
rect 12124 22428 12180 22430
rect 13580 22482 13636 22484
rect 13580 22430 13582 22482
rect 13582 22430 13634 22482
rect 13634 22430 13636 22482
rect 13580 22428 13636 22430
rect 12572 22370 12628 22372
rect 12572 22318 12574 22370
rect 12574 22318 12626 22370
rect 12626 22318 12628 22370
rect 12572 22316 12628 22318
rect 14028 22370 14084 22372
rect 14028 22318 14030 22370
rect 14030 22318 14082 22370
rect 14082 22318 14084 22370
rect 14028 22316 14084 22318
rect 11004 21980 11060 22036
rect 12124 22092 12180 22148
rect 10332 18620 10388 18676
rect 9996 18562 10052 18564
rect 9996 18510 9998 18562
rect 9998 18510 10050 18562
rect 10050 18510 10052 18562
rect 9996 18508 10052 18510
rect 11004 20524 11060 20580
rect 11564 20524 11620 20580
rect 11116 19404 11172 19460
rect 11116 18620 11172 18676
rect 10220 18284 10276 18340
rect 9772 16994 9828 16996
rect 9772 16942 9774 16994
rect 9774 16942 9826 16994
rect 9826 16942 9828 16994
rect 9772 16940 9828 16942
rect 9884 17554 9940 17556
rect 9884 17502 9886 17554
rect 9886 17502 9938 17554
rect 9938 17502 9940 17554
rect 9884 17500 9940 17502
rect 10108 17612 10164 17668
rect 10332 17500 10388 17556
rect 9996 17388 10052 17444
rect 10220 17276 10276 17332
rect 10668 17442 10724 17444
rect 10668 17390 10670 17442
rect 10670 17390 10722 17442
rect 10722 17390 10724 17442
rect 10668 17388 10724 17390
rect 11340 19234 11396 19236
rect 11340 19182 11342 19234
rect 11342 19182 11394 19234
rect 11394 19182 11396 19234
rect 11340 19180 11396 19182
rect 12348 21644 12404 21700
rect 13580 21698 13636 21700
rect 13580 21646 13582 21698
rect 13582 21646 13634 21698
rect 13634 21646 13636 21698
rect 13580 21644 13636 21646
rect 12348 21026 12404 21028
rect 12348 20974 12350 21026
rect 12350 20974 12402 21026
rect 12402 20974 12404 21026
rect 12348 20972 12404 20974
rect 14588 23772 14644 23828
rect 15148 23324 15204 23380
rect 15484 23324 15540 23380
rect 16156 23266 16212 23268
rect 16156 23214 16158 23266
rect 16158 23214 16210 23266
rect 16210 23214 16212 23266
rect 16156 23212 16212 23214
rect 16828 23938 16884 23940
rect 16828 23886 16830 23938
rect 16830 23886 16882 23938
rect 16882 23886 16884 23938
rect 16828 23884 16884 23886
rect 18732 26908 18788 26964
rect 18396 25452 18452 25508
rect 19852 27074 19908 27076
rect 19852 27022 19854 27074
rect 19854 27022 19906 27074
rect 19906 27022 19908 27074
rect 19852 27020 19908 27022
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 20748 27074 20804 27076
rect 20748 27022 20750 27074
rect 20750 27022 20802 27074
rect 20802 27022 20804 27074
rect 20748 27020 20804 27022
rect 21868 27804 21924 27860
rect 18732 24892 18788 24948
rect 19068 25116 19124 25172
rect 18844 24834 18900 24836
rect 18844 24782 18846 24834
rect 18846 24782 18898 24834
rect 18898 24782 18900 24834
rect 18844 24780 18900 24782
rect 19740 25506 19796 25508
rect 19740 25454 19742 25506
rect 19742 25454 19794 25506
rect 19794 25454 19796 25506
rect 19740 25452 19796 25454
rect 19292 25340 19348 25396
rect 20076 25452 20132 25508
rect 20300 25788 20356 25844
rect 21868 25618 21924 25620
rect 21868 25566 21870 25618
rect 21870 25566 21922 25618
rect 21922 25566 21924 25618
rect 21868 25564 21924 25566
rect 22764 28700 22820 28756
rect 22540 28530 22596 28532
rect 22540 28478 22542 28530
rect 22542 28478 22594 28530
rect 22594 28478 22596 28530
rect 22540 28476 22596 28478
rect 22316 28418 22372 28420
rect 22316 28366 22318 28418
rect 22318 28366 22370 28418
rect 22370 28366 22372 28418
rect 22316 28364 22372 28366
rect 22316 27746 22372 27748
rect 22316 27694 22318 27746
rect 22318 27694 22370 27746
rect 22370 27694 22372 27746
rect 22316 27692 22372 27694
rect 22540 27858 22596 27860
rect 22540 27806 22542 27858
rect 22542 27806 22594 27858
rect 22594 27806 22596 27858
rect 22540 27804 22596 27806
rect 22428 27468 22484 27524
rect 22876 28642 22932 28644
rect 22876 28590 22878 28642
rect 22878 28590 22930 28642
rect 22930 28590 22932 28642
rect 22876 28588 22932 28590
rect 23772 32450 23828 32452
rect 23772 32398 23774 32450
rect 23774 32398 23826 32450
rect 23826 32398 23828 32450
rect 23772 32396 23828 32398
rect 24444 31666 24500 31668
rect 24444 31614 24446 31666
rect 24446 31614 24498 31666
rect 24498 31614 24500 31666
rect 24444 31612 24500 31614
rect 24220 31554 24276 31556
rect 24220 31502 24222 31554
rect 24222 31502 24274 31554
rect 24274 31502 24276 31554
rect 24220 31500 24276 31502
rect 24668 31500 24724 31556
rect 24332 30882 24388 30884
rect 24332 30830 24334 30882
rect 24334 30830 24386 30882
rect 24386 30830 24388 30882
rect 24332 30828 24388 30830
rect 24668 30882 24724 30884
rect 24668 30830 24670 30882
rect 24670 30830 24722 30882
rect 24722 30830 24724 30882
rect 24668 30828 24724 30830
rect 26684 34914 26740 34916
rect 26684 34862 26686 34914
rect 26686 34862 26738 34914
rect 26738 34862 26740 34914
rect 26684 34860 26740 34862
rect 26348 34412 26404 34468
rect 25900 34130 25956 34132
rect 25900 34078 25902 34130
rect 25902 34078 25954 34130
rect 25954 34078 25956 34130
rect 25900 34076 25956 34078
rect 24332 30268 24388 30324
rect 24108 30210 24164 30212
rect 24108 30158 24110 30210
rect 24110 30158 24162 30210
rect 24162 30158 24164 30210
rect 24108 30156 24164 30158
rect 25340 31612 25396 31668
rect 25228 30716 25284 30772
rect 25340 30156 25396 30212
rect 24892 30044 24948 30100
rect 23660 28476 23716 28532
rect 22988 27634 23044 27636
rect 22988 27582 22990 27634
rect 22990 27582 23042 27634
rect 23042 27582 23044 27634
rect 22988 27580 23044 27582
rect 22764 26684 22820 26740
rect 23100 26962 23156 26964
rect 23100 26910 23102 26962
rect 23102 26910 23154 26962
rect 23154 26910 23156 26962
rect 23100 26908 23156 26910
rect 22428 26178 22484 26180
rect 22428 26126 22430 26178
rect 22430 26126 22482 26178
rect 22482 26126 22484 26178
rect 22428 26124 22484 26126
rect 23324 27020 23380 27076
rect 22876 25788 22932 25844
rect 23772 26962 23828 26964
rect 23772 26910 23774 26962
rect 23774 26910 23826 26962
rect 23826 26910 23828 26962
rect 23772 26908 23828 26910
rect 24668 28028 24724 28084
rect 25340 28082 25396 28084
rect 25340 28030 25342 28082
rect 25342 28030 25394 28082
rect 25394 28030 25396 28082
rect 25340 28028 25396 28030
rect 25900 31500 25956 31556
rect 26684 33180 26740 33236
rect 25676 30882 25732 30884
rect 25676 30830 25678 30882
rect 25678 30830 25730 30882
rect 25730 30830 25732 30882
rect 25676 30828 25732 30830
rect 26236 30828 26292 30884
rect 26572 31778 26628 31780
rect 26572 31726 26574 31778
rect 26574 31726 26626 31778
rect 26626 31726 26628 31778
rect 26572 31724 26628 31726
rect 26572 30882 26628 30884
rect 26572 30830 26574 30882
rect 26574 30830 26626 30882
rect 26626 30830 26628 30882
rect 26572 30828 26628 30830
rect 25676 28588 25732 28644
rect 24220 27074 24276 27076
rect 24220 27022 24222 27074
rect 24222 27022 24274 27074
rect 24274 27022 24276 27074
rect 24220 27020 24276 27022
rect 24332 26908 24388 26964
rect 23436 26572 23492 26628
rect 24108 26572 24164 26628
rect 23100 25564 23156 25620
rect 23212 25900 23268 25956
rect 22204 25452 22260 25508
rect 22652 25340 22708 25396
rect 19516 25116 19572 25172
rect 19516 24892 19572 24948
rect 19068 23884 19124 23940
rect 16716 23100 16772 23156
rect 16492 22988 16548 23044
rect 14252 22316 14308 22372
rect 14140 21196 14196 21252
rect 14476 22370 14532 22372
rect 14476 22318 14478 22370
rect 14478 22318 14530 22370
rect 14530 22318 14532 22370
rect 14476 22316 14532 22318
rect 14924 22428 14980 22484
rect 14700 21756 14756 21812
rect 15708 22482 15764 22484
rect 15708 22430 15710 22482
rect 15710 22430 15762 22482
rect 15762 22430 15764 22482
rect 15708 22428 15764 22430
rect 15148 21756 15204 21812
rect 15932 21756 15988 21812
rect 16604 22482 16660 22484
rect 16604 22430 16606 22482
rect 16606 22430 16658 22482
rect 16658 22430 16660 22482
rect 16604 22428 16660 22430
rect 17500 22204 17556 22260
rect 17612 22146 17668 22148
rect 17612 22094 17614 22146
rect 17614 22094 17666 22146
rect 17666 22094 17668 22146
rect 17612 22092 17668 22094
rect 17724 21868 17780 21924
rect 13916 20690 13972 20692
rect 13916 20638 13918 20690
rect 13918 20638 13970 20690
rect 13970 20638 13972 20690
rect 13916 20636 13972 20638
rect 13244 19906 13300 19908
rect 13244 19854 13246 19906
rect 13246 19854 13298 19906
rect 13298 19854 13300 19906
rect 13244 19852 13300 19854
rect 14252 20130 14308 20132
rect 14252 20078 14254 20130
rect 14254 20078 14306 20130
rect 14306 20078 14308 20130
rect 14252 20076 14308 20078
rect 11676 19122 11732 19124
rect 11676 19070 11678 19122
rect 11678 19070 11730 19122
rect 11730 19070 11732 19122
rect 11676 19068 11732 19070
rect 11452 18844 11508 18900
rect 11452 18172 11508 18228
rect 11788 18396 11844 18452
rect 10892 17442 10948 17444
rect 10892 17390 10894 17442
rect 10894 17390 10946 17442
rect 10946 17390 10948 17442
rect 10892 17388 10948 17390
rect 9996 16770 10052 16772
rect 9996 16718 9998 16770
rect 9998 16718 10050 16770
rect 10050 16718 10052 16770
rect 9996 16716 10052 16718
rect 9548 15820 9604 15876
rect 9884 15820 9940 15876
rect 9660 15708 9716 15764
rect 10220 15820 10276 15876
rect 8204 14028 8260 14084
rect 8316 14252 8372 14308
rect 5964 13916 6020 13972
rect 6972 13970 7028 13972
rect 6972 13918 6974 13970
rect 6974 13918 7026 13970
rect 7026 13918 7028 13970
rect 6972 13916 7028 13918
rect 5516 12290 5572 12292
rect 5516 12238 5518 12290
rect 5518 12238 5570 12290
rect 5570 12238 5572 12290
rect 5516 12236 5572 12238
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4844 11788 4900 11844
rect 3948 11170 4004 11172
rect 3948 11118 3950 11170
rect 3950 11118 4002 11170
rect 4002 11118 4004 11170
rect 3948 11116 4004 11118
rect 4956 11506 5012 11508
rect 4956 11454 4958 11506
rect 4958 11454 5010 11506
rect 5010 11454 5012 11506
rect 4956 11452 5012 11454
rect 4060 10556 4116 10612
rect 3836 9996 3892 10052
rect 3500 9212 3556 9268
rect 3836 8988 3892 9044
rect 4172 9660 4228 9716
rect 4508 10444 4564 10500
rect 5068 10722 5124 10724
rect 5068 10670 5070 10722
rect 5070 10670 5122 10722
rect 5122 10670 5124 10722
rect 5068 10668 5124 10670
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 5068 10444 5124 10500
rect 4956 9938 5012 9940
rect 4956 9886 4958 9938
rect 4958 9886 5010 9938
rect 5010 9886 5012 9938
rect 4956 9884 5012 9886
rect 4284 9154 4340 9156
rect 4284 9102 4286 9154
rect 4286 9102 4338 9154
rect 4338 9102 4340 9154
rect 4284 9100 4340 9102
rect 3612 8764 3668 8820
rect 4620 9042 4676 9044
rect 4620 8990 4622 9042
rect 4622 8990 4674 9042
rect 4674 8990 4676 9042
rect 4620 8988 4676 8990
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 4956 9548 5012 9604
rect 6300 12460 6356 12516
rect 6972 13522 7028 13524
rect 6972 13470 6974 13522
rect 6974 13470 7026 13522
rect 7026 13470 7028 13522
rect 6972 13468 7028 13470
rect 6412 12236 6468 12292
rect 6300 12178 6356 12180
rect 6300 12126 6302 12178
rect 6302 12126 6354 12178
rect 6354 12126 6356 12178
rect 6300 12124 6356 12126
rect 5740 12012 5796 12068
rect 6300 11788 6356 11844
rect 5740 11564 5796 11620
rect 5740 11282 5796 11284
rect 5740 11230 5742 11282
rect 5742 11230 5794 11282
rect 5794 11230 5796 11282
rect 5740 11228 5796 11230
rect 5852 10610 5908 10612
rect 5852 10558 5854 10610
rect 5854 10558 5906 10610
rect 5906 10558 5908 10610
rect 5852 10556 5908 10558
rect 5180 9324 5236 9380
rect 5292 10108 5348 10164
rect 6412 11394 6468 11396
rect 6412 11342 6414 11394
rect 6414 11342 6466 11394
rect 6466 11342 6468 11394
rect 6412 11340 6468 11342
rect 7868 13020 7924 13076
rect 6636 12124 6692 12180
rect 6748 12012 6804 12068
rect 7084 12850 7140 12852
rect 7084 12798 7086 12850
rect 7086 12798 7138 12850
rect 7138 12798 7140 12850
rect 7084 12796 7140 12798
rect 7420 12460 7476 12516
rect 7532 12908 7588 12964
rect 7644 11788 7700 11844
rect 6972 11340 7028 11396
rect 6524 11228 6580 11284
rect 6412 10108 6468 10164
rect 5404 9266 5460 9268
rect 5404 9214 5406 9266
rect 5406 9214 5458 9266
rect 5458 9214 5460 9266
rect 5404 9212 5460 9214
rect 5292 9154 5348 9156
rect 5292 9102 5294 9154
rect 5294 9102 5346 9154
rect 5346 9102 5348 9154
rect 5292 9100 5348 9102
rect 5068 9042 5124 9044
rect 5068 8990 5070 9042
rect 5070 8990 5122 9042
rect 5122 8990 5124 9042
rect 5068 8988 5124 8990
rect 2940 8146 2996 8148
rect 2940 8094 2942 8146
rect 2942 8094 2994 8146
rect 2994 8094 2996 8146
rect 2940 8092 2996 8094
rect 6972 9884 7028 9940
rect 6748 9714 6804 9716
rect 6748 9662 6750 9714
rect 6750 9662 6802 9714
rect 6802 9662 6804 9714
rect 6748 9660 6804 9662
rect 7084 9548 7140 9604
rect 6636 9266 6692 9268
rect 6636 9214 6638 9266
rect 6638 9214 6690 9266
rect 6690 9214 6692 9266
rect 6636 9212 6692 9214
rect 6412 9042 6468 9044
rect 6412 8990 6414 9042
rect 6414 8990 6466 9042
rect 6466 8990 6468 9042
rect 6412 8988 6468 8990
rect 8204 12236 8260 12292
rect 7980 12066 8036 12068
rect 7980 12014 7982 12066
rect 7982 12014 8034 12066
rect 8034 12014 8036 12066
rect 7980 12012 8036 12014
rect 8204 12012 8260 12068
rect 9212 13356 9268 13412
rect 8540 13244 8596 13300
rect 8652 12962 8708 12964
rect 8652 12910 8654 12962
rect 8654 12910 8706 12962
rect 8706 12910 8708 12962
rect 8652 12908 8708 12910
rect 8876 12962 8932 12964
rect 8876 12910 8878 12962
rect 8878 12910 8930 12962
rect 8930 12910 8932 12962
rect 8876 12908 8932 12910
rect 8876 12572 8932 12628
rect 8540 12460 8596 12516
rect 9212 12796 9268 12852
rect 8764 12178 8820 12180
rect 8764 12126 8766 12178
rect 8766 12126 8818 12178
rect 8818 12126 8820 12178
rect 8764 12124 8820 12126
rect 9548 12850 9604 12852
rect 9548 12798 9550 12850
rect 9550 12798 9602 12850
rect 9602 12798 9604 12850
rect 9548 12796 9604 12798
rect 9548 12572 9604 12628
rect 8316 11788 8372 11844
rect 9212 11900 9268 11956
rect 8988 10498 9044 10500
rect 8988 10446 8990 10498
rect 8990 10446 9042 10498
rect 9042 10446 9044 10498
rect 8988 10444 9044 10446
rect 7756 9660 7812 9716
rect 7196 8988 7252 9044
rect 4732 8258 4788 8260
rect 4732 8206 4734 8258
rect 4734 8206 4786 8258
rect 4786 8206 4788 8258
rect 4732 8204 4788 8206
rect 5404 8204 5460 8260
rect 2044 7420 2100 7476
rect 5964 8258 6020 8260
rect 5964 8206 5966 8258
rect 5966 8206 6018 8258
rect 6018 8206 6020 8258
rect 5964 8204 6020 8206
rect 6636 8258 6692 8260
rect 6636 8206 6638 8258
rect 6638 8206 6690 8258
rect 6690 8206 6692 8258
rect 6636 8204 6692 8206
rect 7084 8204 7140 8260
rect 8204 9884 8260 9940
rect 9996 13356 10052 13412
rect 10444 16268 10500 16324
rect 10892 14306 10948 14308
rect 10892 14254 10894 14306
rect 10894 14254 10946 14306
rect 10946 14254 10948 14306
rect 10892 14252 10948 14254
rect 10556 14140 10612 14196
rect 9884 12290 9940 12292
rect 9884 12238 9886 12290
rect 9886 12238 9938 12290
rect 9938 12238 9940 12290
rect 9884 12236 9940 12238
rect 9772 12124 9828 12180
rect 9660 11900 9716 11956
rect 9660 10722 9716 10724
rect 9660 10670 9662 10722
rect 9662 10670 9714 10722
rect 9714 10670 9716 10722
rect 9660 10668 9716 10670
rect 8092 9212 8148 9268
rect 10556 12850 10612 12852
rect 10556 12798 10558 12850
rect 10558 12798 10610 12850
rect 10610 12798 10612 12850
rect 10556 12796 10612 12798
rect 11900 18172 11956 18228
rect 12124 19458 12180 19460
rect 12124 19406 12126 19458
rect 12126 19406 12178 19458
rect 12178 19406 12180 19458
rect 12124 19404 12180 19406
rect 12572 19234 12628 19236
rect 12572 19182 12574 19234
rect 12574 19182 12626 19234
rect 12626 19182 12628 19234
rect 12572 19180 12628 19182
rect 12124 19010 12180 19012
rect 12124 18958 12126 19010
rect 12126 18958 12178 19010
rect 12178 18958 12180 19010
rect 12124 18956 12180 18958
rect 12236 18732 12292 18788
rect 12684 18620 12740 18676
rect 13468 18844 13524 18900
rect 13356 18562 13412 18564
rect 13356 18510 13358 18562
rect 13358 18510 13410 18562
rect 13410 18510 13412 18562
rect 13356 18508 13412 18510
rect 12460 18060 12516 18116
rect 11788 17388 11844 17444
rect 11340 17276 11396 17332
rect 11900 17052 11956 17108
rect 11788 15820 11844 15876
rect 11228 15036 11284 15092
rect 10332 12290 10388 12292
rect 10332 12238 10334 12290
rect 10334 12238 10386 12290
rect 10386 12238 10388 12290
rect 10332 12236 10388 12238
rect 10108 11228 10164 11284
rect 10668 12124 10724 12180
rect 9884 10444 9940 10500
rect 10332 9996 10388 10052
rect 9772 9660 9828 9716
rect 10444 9714 10500 9716
rect 10444 9662 10446 9714
rect 10446 9662 10498 9714
rect 10498 9662 10500 9714
rect 10444 9660 10500 9662
rect 10780 11170 10836 11172
rect 10780 11118 10782 11170
rect 10782 11118 10834 11170
rect 10834 11118 10836 11170
rect 10780 11116 10836 11118
rect 11004 10668 11060 10724
rect 11452 11788 11508 11844
rect 11340 11282 11396 11284
rect 11340 11230 11342 11282
rect 11342 11230 11394 11282
rect 11394 11230 11396 11282
rect 11340 11228 11396 11230
rect 9884 9266 9940 9268
rect 9884 9214 9886 9266
rect 9886 9214 9938 9266
rect 9938 9214 9940 9266
rect 9884 9212 9940 9214
rect 7420 8316 7476 8372
rect 7420 8034 7476 8036
rect 7420 7982 7422 8034
rect 7422 7982 7474 8034
rect 7474 7982 7476 8034
rect 7420 7980 7476 7982
rect 5964 7250 6020 7252
rect 5964 7198 5966 7250
rect 5966 7198 6018 7250
rect 6018 7198 6020 7250
rect 5964 7196 6020 7198
rect 9548 8316 9604 8372
rect 8316 8092 8372 8148
rect 8428 8204 8484 8260
rect 9436 8258 9492 8260
rect 9436 8206 9438 8258
rect 9438 8206 9490 8258
rect 9490 8206 9492 8258
rect 9436 8204 9492 8206
rect 8876 7698 8932 7700
rect 8876 7646 8878 7698
rect 8878 7646 8930 7698
rect 8930 7646 8932 7698
rect 8876 7644 8932 7646
rect 10220 8370 10276 8372
rect 10220 8318 10222 8370
rect 10222 8318 10274 8370
rect 10274 8318 10276 8370
rect 10220 8316 10276 8318
rect 10108 8092 10164 8148
rect 9772 7474 9828 7476
rect 9772 7422 9774 7474
rect 9774 7422 9826 7474
rect 9826 7422 9828 7474
rect 9772 7420 9828 7422
rect 12012 16380 12068 16436
rect 12236 17052 12292 17108
rect 12124 15932 12180 15988
rect 12236 16882 12292 16884
rect 12236 16830 12238 16882
rect 12238 16830 12290 16882
rect 12290 16830 12292 16882
rect 12236 16828 12292 16830
rect 13468 18396 13524 18452
rect 14588 20412 14644 20468
rect 14812 20748 14868 20804
rect 13916 18284 13972 18340
rect 14476 20188 14532 20244
rect 13468 18226 13524 18228
rect 13468 18174 13470 18226
rect 13470 18174 13522 18226
rect 13522 18174 13524 18226
rect 13468 18172 13524 18174
rect 12796 17164 12852 17220
rect 12348 16380 12404 16436
rect 12796 16156 12852 16212
rect 12684 16098 12740 16100
rect 12684 16046 12686 16098
rect 12686 16046 12738 16098
rect 12738 16046 12740 16098
rect 12684 16044 12740 16046
rect 12796 15874 12852 15876
rect 12796 15822 12798 15874
rect 12798 15822 12850 15874
rect 12850 15822 12852 15874
rect 12796 15820 12852 15822
rect 13692 17666 13748 17668
rect 13692 17614 13694 17666
rect 13694 17614 13746 17666
rect 13746 17614 13748 17666
rect 13692 17612 13748 17614
rect 13356 17388 13412 17444
rect 12684 15036 12740 15092
rect 12796 15260 12852 15316
rect 12684 14140 12740 14196
rect 14028 16882 14084 16884
rect 14028 16830 14030 16882
rect 14030 16830 14082 16882
rect 14082 16830 14084 16882
rect 14028 16828 14084 16830
rect 13692 15314 13748 15316
rect 13692 15262 13694 15314
rect 13694 15262 13746 15314
rect 13746 15262 13748 15314
rect 13692 15260 13748 15262
rect 13356 14140 13412 14196
rect 12684 13746 12740 13748
rect 12684 13694 12686 13746
rect 12686 13694 12738 13746
rect 12738 13694 12740 13746
rect 12684 13692 12740 13694
rect 12908 13468 12964 13524
rect 12124 13244 12180 13300
rect 12012 12348 12068 12404
rect 12012 12012 12068 12068
rect 12124 12684 12180 12740
rect 12124 11788 12180 11844
rect 13916 13468 13972 13524
rect 14700 20018 14756 20020
rect 14700 19966 14702 20018
rect 14702 19966 14754 20018
rect 14754 19966 14756 20018
rect 14700 19964 14756 19966
rect 14364 16268 14420 16324
rect 14476 16716 14532 16772
rect 16156 21026 16212 21028
rect 16156 20974 16158 21026
rect 16158 20974 16210 21026
rect 16210 20974 16212 21026
rect 16156 20972 16212 20974
rect 15596 20802 15652 20804
rect 15596 20750 15598 20802
rect 15598 20750 15650 20802
rect 15650 20750 15652 20802
rect 15596 20748 15652 20750
rect 15820 20412 15876 20468
rect 15260 20130 15316 20132
rect 15260 20078 15262 20130
rect 15262 20078 15314 20130
rect 15314 20078 15316 20130
rect 15260 20076 15316 20078
rect 15484 19852 15540 19908
rect 17388 20802 17444 20804
rect 17388 20750 17390 20802
rect 17390 20750 17442 20802
rect 17442 20750 17444 20802
rect 17388 20748 17444 20750
rect 16268 20076 16324 20132
rect 15932 19740 15988 19796
rect 15148 18450 15204 18452
rect 15148 18398 15150 18450
rect 15150 18398 15202 18450
rect 15202 18398 15204 18450
rect 15148 18396 15204 18398
rect 15820 18620 15876 18676
rect 15036 18172 15092 18228
rect 14924 17388 14980 17444
rect 14700 17106 14756 17108
rect 14700 17054 14702 17106
rect 14702 17054 14754 17106
rect 14754 17054 14756 17106
rect 14700 17052 14756 17054
rect 14924 16828 14980 16884
rect 15148 16268 15204 16324
rect 14812 16210 14868 16212
rect 14812 16158 14814 16210
rect 14814 16158 14866 16210
rect 14866 16158 14868 16210
rect 14812 16156 14868 16158
rect 14588 16098 14644 16100
rect 14588 16046 14590 16098
rect 14590 16046 14642 16098
rect 14642 16046 14644 16098
rect 14588 16044 14644 16046
rect 14476 15986 14532 15988
rect 14476 15934 14478 15986
rect 14478 15934 14530 15986
rect 14530 15934 14532 15986
rect 14476 15932 14532 15934
rect 15932 18284 15988 18340
rect 16268 18396 16324 18452
rect 15932 17164 15988 17220
rect 16268 17612 16324 17668
rect 16268 17052 16324 17108
rect 16940 20076 16996 20132
rect 17948 22092 18004 22148
rect 17948 20748 18004 20804
rect 17276 19964 17332 20020
rect 17612 20018 17668 20020
rect 17612 19966 17614 20018
rect 17614 19966 17666 20018
rect 17666 19966 17668 20018
rect 17612 19964 17668 19966
rect 17612 18844 17668 18900
rect 16828 18508 16884 18564
rect 17500 18508 17556 18564
rect 16716 18284 16772 18340
rect 16268 16658 16324 16660
rect 16268 16606 16270 16658
rect 16270 16606 16322 16658
rect 16322 16606 16324 16658
rect 16268 16604 16324 16606
rect 16044 16268 16100 16324
rect 16716 16604 16772 16660
rect 16492 16492 16548 16548
rect 15148 15314 15204 15316
rect 15148 15262 15150 15314
rect 15150 15262 15202 15314
rect 15202 15262 15204 15314
rect 15148 15260 15204 15262
rect 14140 13746 14196 13748
rect 14140 13694 14142 13746
rect 14142 13694 14194 13746
rect 14194 13694 14196 13746
rect 14140 13692 14196 13694
rect 14700 14530 14756 14532
rect 14700 14478 14702 14530
rect 14702 14478 14754 14530
rect 14754 14478 14756 14530
rect 14700 14476 14756 14478
rect 14476 14418 14532 14420
rect 14476 14366 14478 14418
rect 14478 14366 14530 14418
rect 14530 14366 14532 14418
rect 14476 14364 14532 14366
rect 14476 13522 14532 13524
rect 14476 13470 14478 13522
rect 14478 13470 14530 13522
rect 14530 13470 14532 13522
rect 14476 13468 14532 13470
rect 12572 11394 12628 11396
rect 12572 11342 12574 11394
rect 12574 11342 12626 11394
rect 12626 11342 12628 11394
rect 12572 11340 12628 11342
rect 13580 11564 13636 11620
rect 12460 11116 12516 11172
rect 13804 12402 13860 12404
rect 13804 12350 13806 12402
rect 13806 12350 13858 12402
rect 13858 12350 13860 12402
rect 13804 12348 13860 12350
rect 13916 12178 13972 12180
rect 13916 12126 13918 12178
rect 13918 12126 13970 12178
rect 13970 12126 13972 12178
rect 13916 12124 13972 12126
rect 12796 10892 12852 10948
rect 14588 12908 14644 12964
rect 14700 12738 14756 12740
rect 14700 12686 14702 12738
rect 14702 12686 14754 12738
rect 14754 12686 14756 12738
rect 14700 12684 14756 12686
rect 15596 15426 15652 15428
rect 15596 15374 15598 15426
rect 15598 15374 15650 15426
rect 15650 15374 15652 15426
rect 15596 15372 15652 15374
rect 15372 14364 15428 14420
rect 15484 14588 15540 14644
rect 15372 14140 15428 14196
rect 15932 15372 15988 15428
rect 16156 15538 16212 15540
rect 16156 15486 16158 15538
rect 16158 15486 16210 15538
rect 16210 15486 16212 15538
rect 16156 15484 16212 15486
rect 16044 14588 16100 14644
rect 15596 13804 15652 13860
rect 14812 12348 14868 12404
rect 15708 14140 15764 14196
rect 16716 16156 16772 16212
rect 16940 16658 16996 16660
rect 16940 16606 16942 16658
rect 16942 16606 16994 16658
rect 16994 16606 16996 16658
rect 16940 16604 16996 16606
rect 16380 13580 16436 13636
rect 17388 14530 17444 14532
rect 17388 14478 17390 14530
rect 17390 14478 17442 14530
rect 17442 14478 17444 14530
rect 17388 14476 17444 14478
rect 16940 13746 16996 13748
rect 16940 13694 16942 13746
rect 16942 13694 16994 13746
rect 16994 13694 16996 13746
rect 16940 13692 16996 13694
rect 15708 13468 15764 13524
rect 15596 12908 15652 12964
rect 15372 12402 15428 12404
rect 15372 12350 15374 12402
rect 15374 12350 15426 12402
rect 15426 12350 15428 12402
rect 15372 12348 15428 12350
rect 14588 12124 14644 12180
rect 13916 11340 13972 11396
rect 11452 9212 11508 9268
rect 12236 10332 12292 10388
rect 12124 10050 12180 10052
rect 12124 9998 12126 10050
rect 12126 9998 12178 10050
rect 12178 9998 12180 10050
rect 12124 9996 12180 9998
rect 13692 10892 13748 10948
rect 14476 11116 14532 11172
rect 16268 12348 16324 12404
rect 15820 11900 15876 11956
rect 15932 11506 15988 11508
rect 15932 11454 15934 11506
rect 15934 11454 15986 11506
rect 15986 11454 15988 11506
rect 15932 11452 15988 11454
rect 15484 11394 15540 11396
rect 15484 11342 15486 11394
rect 15486 11342 15538 11394
rect 15538 11342 15540 11394
rect 15484 11340 15540 11342
rect 14476 10386 14532 10388
rect 14476 10334 14478 10386
rect 14478 10334 14530 10386
rect 14530 10334 14532 10386
rect 14476 10332 14532 10334
rect 14924 10332 14980 10388
rect 13580 9324 13636 9380
rect 14588 9996 14644 10052
rect 16380 11618 16436 11620
rect 16380 11566 16382 11618
rect 16382 11566 16434 11618
rect 16434 11566 16436 11618
rect 16380 11564 16436 11566
rect 16492 11340 16548 11396
rect 16828 11900 16884 11956
rect 18508 23042 18564 23044
rect 18508 22990 18510 23042
rect 18510 22990 18562 23042
rect 18562 22990 18564 23042
rect 18508 22988 18564 22990
rect 18620 22930 18676 22932
rect 18620 22878 18622 22930
rect 18622 22878 18674 22930
rect 18674 22878 18676 22930
rect 18620 22876 18676 22878
rect 18172 22204 18228 22260
rect 18732 21868 18788 21924
rect 18060 20076 18116 20132
rect 18508 18956 18564 19012
rect 19292 22930 19348 22932
rect 19292 22878 19294 22930
rect 19294 22878 19346 22930
rect 19346 22878 19348 22930
rect 19292 22876 19348 22878
rect 18732 20578 18788 20580
rect 18732 20526 18734 20578
rect 18734 20526 18786 20578
rect 18786 20526 18788 20578
rect 18732 20524 18788 20526
rect 19180 20578 19236 20580
rect 19180 20526 19182 20578
rect 19182 20526 19234 20578
rect 19234 20526 19236 20578
rect 19180 20524 19236 20526
rect 19068 19964 19124 20020
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 20300 24834 20356 24836
rect 20300 24782 20302 24834
rect 20302 24782 20354 24834
rect 20354 24782 20356 24834
rect 20300 24780 20356 24782
rect 19852 24722 19908 24724
rect 19852 24670 19854 24722
rect 19854 24670 19906 24722
rect 19906 24670 19908 24722
rect 19852 24668 19908 24670
rect 19740 23884 19796 23940
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 20636 24834 20692 24836
rect 20636 24782 20638 24834
rect 20638 24782 20690 24834
rect 20690 24782 20692 24834
rect 20636 24780 20692 24782
rect 21084 24834 21140 24836
rect 21084 24782 21086 24834
rect 21086 24782 21138 24834
rect 21138 24782 21140 24834
rect 21084 24780 21140 24782
rect 21532 24722 21588 24724
rect 21532 24670 21534 24722
rect 21534 24670 21586 24722
rect 21586 24670 21588 24722
rect 21532 24668 21588 24670
rect 21308 24332 21364 24388
rect 20636 24050 20692 24052
rect 20636 23998 20638 24050
rect 20638 23998 20690 24050
rect 20690 23998 20692 24050
rect 20636 23996 20692 23998
rect 21308 23772 21364 23828
rect 22764 24108 22820 24164
rect 21532 23548 21588 23604
rect 20412 23212 20468 23268
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 20748 21698 20804 21700
rect 20748 21646 20750 21698
rect 20750 21646 20802 21698
rect 20802 21646 20804 21698
rect 20748 21644 20804 21646
rect 21644 21644 21700 21700
rect 21420 20860 21476 20916
rect 19740 20636 19796 20692
rect 18732 19180 18788 19236
rect 19404 19234 19460 19236
rect 19404 19182 19406 19234
rect 19406 19182 19458 19234
rect 19458 19182 19460 19234
rect 19404 19180 19460 19182
rect 19180 19068 19236 19124
rect 18620 18674 18676 18676
rect 18620 18622 18622 18674
rect 18622 18622 18674 18674
rect 18674 18622 18676 18674
rect 18620 18620 18676 18622
rect 19404 18956 19460 19012
rect 19180 18674 19236 18676
rect 19180 18622 19182 18674
rect 19182 18622 19234 18674
rect 19234 18622 19236 18674
rect 19180 18620 19236 18622
rect 21196 20690 21252 20692
rect 21196 20638 21198 20690
rect 21198 20638 21250 20690
rect 21250 20638 21252 20690
rect 21196 20636 21252 20638
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 19740 19068 19796 19124
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 17948 17612 18004 17668
rect 17836 17388 17892 17444
rect 17612 16940 17668 16996
rect 18060 17052 18116 17108
rect 17724 16828 17780 16884
rect 17724 16492 17780 16548
rect 17836 16604 17892 16660
rect 17724 15148 17780 15204
rect 18284 16604 18340 16660
rect 18396 16044 18452 16100
rect 18060 13804 18116 13860
rect 18284 15260 18340 15316
rect 19068 16994 19124 16996
rect 19068 16942 19070 16994
rect 19070 16942 19122 16994
rect 19122 16942 19124 16994
rect 19068 16940 19124 16942
rect 22092 20748 22148 20804
rect 22428 23154 22484 23156
rect 22428 23102 22430 23154
rect 22430 23102 22482 23154
rect 22482 23102 22484 23154
rect 22428 23100 22484 23102
rect 22540 22988 22596 23044
rect 22764 22540 22820 22596
rect 23660 26178 23716 26180
rect 23660 26126 23662 26178
rect 23662 26126 23714 26178
rect 23714 26126 23716 26178
rect 23660 26124 23716 26126
rect 23548 25116 23604 25172
rect 23772 24892 23828 24948
rect 24220 24946 24276 24948
rect 24220 24894 24222 24946
rect 24222 24894 24274 24946
rect 24274 24894 24276 24946
rect 24220 24892 24276 24894
rect 24444 25116 24500 25172
rect 27580 45948 27636 46004
rect 28364 45890 28420 45892
rect 28364 45838 28366 45890
rect 28366 45838 28418 45890
rect 28418 45838 28420 45890
rect 28364 45836 28420 45838
rect 27020 36316 27076 36372
rect 26908 34972 26964 35028
rect 26908 32674 26964 32676
rect 26908 32622 26910 32674
rect 26910 32622 26962 32674
rect 26962 32622 26964 32674
rect 26908 32620 26964 32622
rect 26908 31052 26964 31108
rect 27132 31500 27188 31556
rect 26796 29148 26852 29204
rect 26908 29036 26964 29092
rect 29372 46114 29428 46116
rect 29372 46062 29374 46114
rect 29374 46062 29426 46114
rect 29426 46062 29428 46114
rect 29372 46060 29428 46062
rect 29260 45106 29316 45108
rect 29260 45054 29262 45106
rect 29262 45054 29314 45106
rect 29314 45054 29316 45106
rect 29260 45052 29316 45054
rect 28700 42364 28756 42420
rect 28364 40796 28420 40852
rect 28028 40236 28084 40292
rect 28812 40236 28868 40292
rect 28700 40124 28756 40180
rect 28700 39618 28756 39620
rect 28700 39566 28702 39618
rect 28702 39566 28754 39618
rect 28754 39566 28756 39618
rect 28700 39564 28756 39566
rect 28700 39058 28756 39060
rect 28700 39006 28702 39058
rect 28702 39006 28754 39058
rect 28754 39006 28756 39058
rect 28700 39004 28756 39006
rect 28812 38892 28868 38948
rect 28588 37826 28644 37828
rect 28588 37774 28590 37826
rect 28590 37774 28642 37826
rect 28642 37774 28644 37826
rect 28588 37772 28644 37774
rect 28476 37378 28532 37380
rect 28476 37326 28478 37378
rect 28478 37326 28530 37378
rect 28530 37326 28532 37378
rect 28476 37324 28532 37326
rect 28252 36540 28308 36596
rect 27916 35196 27972 35252
rect 27804 34972 27860 35028
rect 27692 34242 27748 34244
rect 27692 34190 27694 34242
rect 27694 34190 27746 34242
rect 27746 34190 27748 34242
rect 27692 34188 27748 34190
rect 27356 31164 27412 31220
rect 27468 34130 27524 34132
rect 27468 34078 27470 34130
rect 27470 34078 27522 34130
rect 27522 34078 27524 34130
rect 27468 34076 27524 34078
rect 30044 42364 30100 42420
rect 30156 42642 30212 42644
rect 30156 42590 30158 42642
rect 30158 42590 30210 42642
rect 30210 42590 30212 42642
rect 30156 42588 30212 42590
rect 30380 44940 30436 44996
rect 30492 42588 30548 42644
rect 30380 42530 30436 42532
rect 30380 42478 30382 42530
rect 30382 42478 30434 42530
rect 30434 42478 30436 42530
rect 30380 42476 30436 42478
rect 29708 41132 29764 41188
rect 29708 40796 29764 40852
rect 29820 41356 29876 41412
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 35084 46002 35140 46004
rect 35084 45950 35086 46002
rect 35086 45950 35138 46002
rect 35138 45950 35140 46002
rect 35084 45948 35140 45950
rect 36988 45948 37044 46004
rect 36540 45890 36596 45892
rect 36540 45838 36542 45890
rect 36542 45838 36594 45890
rect 36594 45838 36596 45890
rect 36540 45836 36596 45838
rect 38108 45890 38164 45892
rect 38108 45838 38110 45890
rect 38110 45838 38162 45890
rect 38162 45838 38164 45890
rect 38108 45836 38164 45838
rect 35532 45778 35588 45780
rect 35532 45726 35534 45778
rect 35534 45726 35586 45778
rect 35586 45726 35588 45778
rect 35532 45724 35588 45726
rect 36316 45052 36372 45108
rect 36204 44940 36260 44996
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 32172 43036 32228 43092
rect 37212 45612 37268 45668
rect 36316 44210 36372 44212
rect 36316 44158 36318 44210
rect 36318 44158 36370 44210
rect 36370 44158 36372 44210
rect 36316 44156 36372 44158
rect 33516 43372 33572 43428
rect 33628 42924 33684 42980
rect 31276 42588 31332 42644
rect 31724 42642 31780 42644
rect 31724 42590 31726 42642
rect 31726 42590 31778 42642
rect 31778 42590 31780 42642
rect 31724 42588 31780 42590
rect 31948 42476 32004 42532
rect 33292 42588 33348 42644
rect 30716 42364 30772 42420
rect 32508 41916 32564 41972
rect 31052 41244 31108 41300
rect 33404 42476 33460 42532
rect 33628 42364 33684 42420
rect 32508 41356 32564 41412
rect 32172 41186 32228 41188
rect 32172 41134 32174 41186
rect 32174 41134 32226 41186
rect 32226 41134 32228 41186
rect 32172 41132 32228 41134
rect 31164 40684 31220 40740
rect 29484 39564 29540 39620
rect 29932 39116 29988 39172
rect 29372 39004 29428 39060
rect 29820 38946 29876 38948
rect 29820 38894 29822 38946
rect 29822 38894 29874 38946
rect 29874 38894 29876 38946
rect 29820 38892 29876 38894
rect 29372 37436 29428 37492
rect 29260 37378 29316 37380
rect 29260 37326 29262 37378
rect 29262 37326 29314 37378
rect 29314 37326 29316 37378
rect 29260 37324 29316 37326
rect 29708 37772 29764 37828
rect 29484 36594 29540 36596
rect 29484 36542 29486 36594
rect 29486 36542 29538 36594
rect 29538 36542 29540 36594
rect 29484 36540 29540 36542
rect 29932 37436 29988 37492
rect 28588 35698 28644 35700
rect 28588 35646 28590 35698
rect 28590 35646 28642 35698
rect 28642 35646 28644 35698
rect 28588 35644 28644 35646
rect 28364 35196 28420 35252
rect 28476 34636 28532 34692
rect 27580 33180 27636 33236
rect 27692 31948 27748 32004
rect 28924 34524 28980 34580
rect 28812 34300 28868 34356
rect 28924 34242 28980 34244
rect 28924 34190 28926 34242
rect 28926 34190 28978 34242
rect 28978 34190 28980 34242
rect 28924 34188 28980 34190
rect 28588 34130 28644 34132
rect 28588 34078 28590 34130
rect 28590 34078 28642 34130
rect 28642 34078 28644 34130
rect 28588 34076 28644 34078
rect 27020 28642 27076 28644
rect 27020 28590 27022 28642
rect 27022 28590 27074 28642
rect 27074 28590 27076 28642
rect 27020 28588 27076 28590
rect 27244 28530 27300 28532
rect 27244 28478 27246 28530
rect 27246 28478 27298 28530
rect 27298 28478 27300 28530
rect 27244 28476 27300 28478
rect 27356 28028 27412 28084
rect 27916 31218 27972 31220
rect 27916 31166 27918 31218
rect 27918 31166 27970 31218
rect 27970 31166 27972 31218
rect 27916 31164 27972 31166
rect 27132 27186 27188 27188
rect 27132 27134 27134 27186
rect 27134 27134 27186 27186
rect 27186 27134 27188 27186
rect 27132 27132 27188 27134
rect 27580 29372 27636 29428
rect 26460 26908 26516 26964
rect 25004 25676 25060 25732
rect 25676 25340 25732 25396
rect 25900 25676 25956 25732
rect 25564 24892 25620 24948
rect 24332 24780 24388 24836
rect 25452 24668 25508 24724
rect 24668 24556 24724 24612
rect 24780 24332 24836 24388
rect 24444 24108 24500 24164
rect 22876 22428 22932 22484
rect 25004 24108 25060 24164
rect 24332 23772 24388 23828
rect 24220 23436 24276 23492
rect 22988 20748 23044 20804
rect 22540 20636 22596 20692
rect 20524 19292 20580 19348
rect 21420 19292 21476 19348
rect 20412 19180 20468 19236
rect 21756 19234 21812 19236
rect 21756 19182 21758 19234
rect 21758 19182 21810 19234
rect 21810 19182 21812 19234
rect 21756 19180 21812 19182
rect 20412 18620 20468 18676
rect 20300 18508 20356 18564
rect 19628 17500 19684 17556
rect 20636 17554 20692 17556
rect 20636 17502 20638 17554
rect 20638 17502 20690 17554
rect 20690 17502 20692 17554
rect 20636 17500 20692 17502
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19516 16828 19572 16884
rect 18844 16380 18900 16436
rect 20636 16322 20692 16324
rect 20636 16270 20638 16322
rect 20638 16270 20690 16322
rect 20690 16270 20692 16322
rect 20636 16268 20692 16270
rect 19180 16098 19236 16100
rect 19180 16046 19182 16098
rect 19182 16046 19234 16098
rect 19234 16046 19236 16098
rect 19180 16044 19236 16046
rect 18844 15820 18900 15876
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 20524 15484 20580 15540
rect 21308 17388 21364 17444
rect 20972 17052 21028 17108
rect 21980 17500 22036 17556
rect 21868 16044 21924 16100
rect 20636 15596 20692 15652
rect 21532 15820 21588 15876
rect 21196 15372 21252 15428
rect 19292 15202 19348 15204
rect 19292 15150 19294 15202
rect 19294 15150 19346 15202
rect 19346 15150 19348 15202
rect 19292 15148 19348 15150
rect 21308 15314 21364 15316
rect 21308 15262 21310 15314
rect 21310 15262 21362 15314
rect 21362 15262 21364 15314
rect 21308 15260 21364 15262
rect 22204 15314 22260 15316
rect 22204 15262 22206 15314
rect 22206 15262 22258 15314
rect 22258 15262 22260 15314
rect 22204 15260 22260 15262
rect 23100 20636 23156 20692
rect 24108 22540 24164 22596
rect 23884 22316 23940 22372
rect 24668 23826 24724 23828
rect 24668 23774 24670 23826
rect 24670 23774 24722 23826
rect 24722 23774 24724 23826
rect 24668 23772 24724 23774
rect 24780 23548 24836 23604
rect 24444 23266 24500 23268
rect 24444 23214 24446 23266
rect 24446 23214 24498 23266
rect 24498 23214 24500 23266
rect 24444 23212 24500 23214
rect 23660 21644 23716 21700
rect 25340 24610 25396 24612
rect 25340 24558 25342 24610
rect 25342 24558 25394 24610
rect 25394 24558 25396 24610
rect 25340 24556 25396 24558
rect 25340 23996 25396 24052
rect 25228 23436 25284 23492
rect 25676 23826 25732 23828
rect 25676 23774 25678 23826
rect 25678 23774 25730 23826
rect 25730 23774 25732 23826
rect 25676 23772 25732 23774
rect 26124 22988 26180 23044
rect 26348 25340 26404 25396
rect 25900 22316 25956 22372
rect 26348 24780 26404 24836
rect 26684 24892 26740 24948
rect 27804 29148 27860 29204
rect 27804 28700 27860 28756
rect 28140 31948 28196 32004
rect 27804 28530 27860 28532
rect 27804 28478 27806 28530
rect 27806 28478 27858 28530
rect 27858 28478 27860 28530
rect 27804 28476 27860 28478
rect 27804 28028 27860 28084
rect 27356 26962 27412 26964
rect 27356 26910 27358 26962
rect 27358 26910 27410 26962
rect 27410 26910 27412 26962
rect 27356 26908 27412 26910
rect 27244 24892 27300 24948
rect 27356 25116 27412 25172
rect 26796 23436 26852 23492
rect 26796 23154 26852 23156
rect 26796 23102 26798 23154
rect 26798 23102 26850 23154
rect 26850 23102 26852 23154
rect 26796 23100 26852 23102
rect 26460 22428 26516 22484
rect 25564 21868 25620 21924
rect 25340 21644 25396 21700
rect 24668 21196 24724 21252
rect 23996 20802 24052 20804
rect 23996 20750 23998 20802
rect 23998 20750 24050 20802
rect 24050 20750 24052 20802
rect 23996 20748 24052 20750
rect 23884 20188 23940 20244
rect 23212 20076 23268 20132
rect 23212 19292 23268 19348
rect 22764 18508 22820 18564
rect 22876 17836 22932 17892
rect 23548 18508 23604 18564
rect 23436 17836 23492 17892
rect 22540 17612 22596 17668
rect 23212 17666 23268 17668
rect 23212 17614 23214 17666
rect 23214 17614 23266 17666
rect 23266 17614 23268 17666
rect 23212 17612 23268 17614
rect 23212 16994 23268 16996
rect 23212 16942 23214 16994
rect 23214 16942 23266 16994
rect 23266 16942 23268 16994
rect 23212 16940 23268 16942
rect 23772 16268 23828 16324
rect 22428 16098 22484 16100
rect 22428 16046 22430 16098
rect 22430 16046 22482 16098
rect 22482 16046 22484 16098
rect 22428 16044 22484 16046
rect 22540 15708 22596 15764
rect 18396 14642 18452 14644
rect 18396 14590 18398 14642
rect 18398 14590 18450 14642
rect 18450 14590 18452 14642
rect 18396 14588 18452 14590
rect 19068 14642 19124 14644
rect 19068 14590 19070 14642
rect 19070 14590 19122 14642
rect 19122 14590 19124 14642
rect 19068 14588 19124 14590
rect 19068 13804 19124 13860
rect 18732 13746 18788 13748
rect 18732 13694 18734 13746
rect 18734 13694 18786 13746
rect 18786 13694 18788 13746
rect 18732 13692 18788 13694
rect 16940 11452 16996 11508
rect 17164 11564 17220 11620
rect 16940 10556 16996 10612
rect 16492 10498 16548 10500
rect 16492 10446 16494 10498
rect 16494 10446 16546 10498
rect 16546 10446 16548 10498
rect 16492 10444 16548 10446
rect 14812 9714 14868 9716
rect 14812 9662 14814 9714
rect 14814 9662 14866 9714
rect 14866 9662 14868 9714
rect 14812 9660 14868 9662
rect 13244 8316 13300 8372
rect 13580 8370 13636 8372
rect 13580 8318 13582 8370
rect 13582 8318 13634 8370
rect 13634 8318 13636 8370
rect 13580 8316 13636 8318
rect 12572 8204 12628 8260
rect 13804 8258 13860 8260
rect 13804 8206 13806 8258
rect 13806 8206 13858 8258
rect 13858 8206 13860 8258
rect 13804 8204 13860 8206
rect 11228 7868 11284 7924
rect 11116 7644 11172 7700
rect 11676 8146 11732 8148
rect 11676 8094 11678 8146
rect 11678 8094 11730 8146
rect 11730 8094 11732 8146
rect 11676 8092 11732 8094
rect 11452 7532 11508 7588
rect 11004 7420 11060 7476
rect 13580 7532 13636 7588
rect 12572 7474 12628 7476
rect 12572 7422 12574 7474
rect 12574 7422 12626 7474
rect 12626 7422 12628 7474
rect 12572 7420 12628 7422
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 13916 7980 13972 8036
rect 14028 7250 14084 7252
rect 14028 7198 14030 7250
rect 14030 7198 14082 7250
rect 14082 7198 14084 7250
rect 14028 7196 14084 7198
rect 13916 6748 13972 6804
rect 14588 9154 14644 9156
rect 14588 9102 14590 9154
rect 14590 9102 14642 9154
rect 14642 9102 14644 9154
rect 14588 9100 14644 9102
rect 14812 9100 14868 9156
rect 14924 8092 14980 8148
rect 14812 7868 14868 7924
rect 14588 7644 14644 7700
rect 14700 7586 14756 7588
rect 14700 7534 14702 7586
rect 14702 7534 14754 7586
rect 14754 7534 14756 7586
rect 14700 7532 14756 7534
rect 15148 7532 15204 7588
rect 14476 7308 14532 7364
rect 14700 6748 14756 6804
rect 15260 7362 15316 7364
rect 15260 7310 15262 7362
rect 15262 7310 15314 7362
rect 15314 7310 15316 7362
rect 15260 7308 15316 7310
rect 17724 11564 17780 11620
rect 17612 11340 17668 11396
rect 18732 13468 18788 13524
rect 19292 13468 19348 13524
rect 19628 14252 19684 14308
rect 18396 12348 18452 12404
rect 17948 11900 18004 11956
rect 18284 11788 18340 11844
rect 17724 10498 17780 10500
rect 17724 10446 17726 10498
rect 17726 10446 17778 10498
rect 17778 10446 17780 10498
rect 17724 10444 17780 10446
rect 17612 9826 17668 9828
rect 17612 9774 17614 9826
rect 17614 9774 17666 9826
rect 17666 9774 17668 9826
rect 17612 9772 17668 9774
rect 20412 14306 20468 14308
rect 20412 14254 20414 14306
rect 20414 14254 20466 14306
rect 20466 14254 20468 14306
rect 20412 14252 20468 14254
rect 20636 14306 20692 14308
rect 20636 14254 20638 14306
rect 20638 14254 20690 14306
rect 20690 14254 20692 14306
rect 20636 14252 20692 14254
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 20860 13916 20916 13972
rect 19740 13804 19796 13860
rect 20412 13804 20468 13860
rect 20076 13468 20132 13524
rect 20748 13580 20804 13636
rect 20748 12962 20804 12964
rect 20748 12910 20750 12962
rect 20750 12910 20802 12962
rect 20802 12910 20804 12962
rect 20748 12908 20804 12910
rect 20748 12684 20804 12740
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19964 12348 20020 12404
rect 19516 12290 19572 12292
rect 19516 12238 19518 12290
rect 19518 12238 19570 12290
rect 19570 12238 19572 12290
rect 19516 12236 19572 12238
rect 20076 12290 20132 12292
rect 20076 12238 20078 12290
rect 20078 12238 20130 12290
rect 20130 12238 20132 12290
rect 20076 12236 20132 12238
rect 22428 15484 22484 15540
rect 21756 14418 21812 14420
rect 21756 14366 21758 14418
rect 21758 14366 21810 14418
rect 21810 14366 21812 14418
rect 21756 14364 21812 14366
rect 21420 12684 21476 12740
rect 20748 12290 20804 12292
rect 20748 12238 20750 12290
rect 20750 12238 20802 12290
rect 20802 12238 20804 12290
rect 20748 12236 20804 12238
rect 19180 11788 19236 11844
rect 20300 11564 20356 11620
rect 20188 11452 20244 11508
rect 19180 11394 19236 11396
rect 19180 11342 19182 11394
rect 19182 11342 19234 11394
rect 19234 11342 19236 11394
rect 19180 11340 19236 11342
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 21420 11452 21476 11508
rect 21532 11564 21588 11620
rect 22764 15986 22820 15988
rect 22764 15934 22766 15986
rect 22766 15934 22818 15986
rect 22818 15934 22820 15986
rect 22764 15932 22820 15934
rect 23100 15874 23156 15876
rect 23100 15822 23102 15874
rect 23102 15822 23154 15874
rect 23154 15822 23156 15874
rect 23100 15820 23156 15822
rect 23660 15820 23716 15876
rect 22652 15372 22708 15428
rect 25452 20690 25508 20692
rect 25452 20638 25454 20690
rect 25454 20638 25506 20690
rect 25506 20638 25508 20690
rect 25452 20636 25508 20638
rect 24556 20130 24612 20132
rect 24556 20078 24558 20130
rect 24558 20078 24610 20130
rect 24610 20078 24612 20130
rect 24556 20076 24612 20078
rect 24108 19794 24164 19796
rect 24108 19742 24110 19794
rect 24110 19742 24162 19794
rect 24162 19742 24164 19794
rect 24108 19740 24164 19742
rect 26460 21868 26516 21924
rect 25676 21756 25732 21812
rect 25676 20524 25732 20580
rect 25900 20300 25956 20356
rect 26796 21196 26852 21252
rect 27020 23826 27076 23828
rect 27020 23774 27022 23826
rect 27022 23774 27074 23826
rect 27074 23774 27076 23826
rect 27020 23772 27076 23774
rect 27580 27132 27636 27188
rect 27692 26572 27748 26628
rect 28700 32060 28756 32116
rect 28588 31948 28644 32004
rect 28364 31612 28420 31668
rect 28252 31500 28308 31556
rect 28364 31164 28420 31220
rect 28252 30994 28308 30996
rect 28252 30942 28254 30994
rect 28254 30942 28306 30994
rect 28306 30942 28308 30994
rect 28252 30940 28308 30942
rect 28924 31218 28980 31220
rect 28924 31166 28926 31218
rect 28926 31166 28978 31218
rect 28978 31166 28980 31218
rect 28924 31164 28980 31166
rect 29260 35420 29316 35476
rect 29148 35196 29204 35252
rect 30044 36652 30100 36708
rect 29820 35810 29876 35812
rect 29820 35758 29822 35810
rect 29822 35758 29874 35810
rect 29874 35758 29876 35810
rect 29820 35756 29876 35758
rect 29372 35196 29428 35252
rect 29820 35196 29876 35252
rect 29484 34690 29540 34692
rect 29484 34638 29486 34690
rect 29486 34638 29538 34690
rect 29538 34638 29540 34690
rect 29484 34636 29540 34638
rect 29596 34524 29652 34580
rect 29596 34354 29652 34356
rect 29596 34302 29598 34354
rect 29598 34302 29650 34354
rect 29650 34302 29652 34354
rect 29596 34300 29652 34302
rect 29372 34076 29428 34132
rect 29820 34130 29876 34132
rect 29820 34078 29822 34130
rect 29822 34078 29874 34130
rect 29874 34078 29876 34130
rect 29820 34076 29876 34078
rect 29372 32620 29428 32676
rect 29148 31666 29204 31668
rect 29148 31614 29150 31666
rect 29150 31614 29202 31666
rect 29202 31614 29204 31666
rect 29148 31612 29204 31614
rect 28924 30994 28980 30996
rect 28924 30942 28926 30994
rect 28926 30942 28978 30994
rect 28978 30942 28980 30994
rect 28924 30940 28980 30942
rect 28476 30828 28532 30884
rect 28364 30380 28420 30436
rect 29036 30268 29092 30324
rect 28140 29650 28196 29652
rect 28140 29598 28142 29650
rect 28142 29598 28194 29650
rect 28194 29598 28196 29650
rect 28140 29596 28196 29598
rect 28028 28812 28084 28868
rect 28140 27916 28196 27972
rect 27468 24780 27524 24836
rect 27916 25618 27972 25620
rect 27916 25566 27918 25618
rect 27918 25566 27970 25618
rect 27970 25566 27972 25618
rect 27916 25564 27972 25566
rect 27356 24722 27412 24724
rect 27356 24670 27358 24722
rect 27358 24670 27410 24722
rect 27410 24670 27412 24722
rect 27356 24668 27412 24670
rect 27244 24498 27300 24500
rect 27244 24446 27246 24498
rect 27246 24446 27298 24498
rect 27298 24446 27300 24498
rect 27244 24444 27300 24446
rect 29820 32562 29876 32564
rect 29820 32510 29822 32562
rect 29822 32510 29874 32562
rect 29874 32510 29876 32562
rect 29820 32508 29876 32510
rect 29708 31724 29764 31780
rect 29708 30940 29764 30996
rect 29820 31164 29876 31220
rect 29596 30828 29652 30884
rect 29260 30770 29316 30772
rect 29260 30718 29262 30770
rect 29262 30718 29314 30770
rect 29314 30718 29316 30770
rect 29260 30716 29316 30718
rect 29036 29986 29092 29988
rect 29036 29934 29038 29986
rect 29038 29934 29090 29986
rect 29090 29934 29092 29986
rect 29036 29932 29092 29934
rect 29372 29708 29428 29764
rect 28476 29596 28532 29652
rect 28812 29596 28868 29652
rect 28588 29484 28644 29540
rect 28476 28700 28532 28756
rect 29148 29426 29204 29428
rect 29148 29374 29150 29426
rect 29150 29374 29202 29426
rect 29202 29374 29204 29426
rect 29148 29372 29204 29374
rect 28812 29314 28868 29316
rect 28812 29262 28814 29314
rect 28814 29262 28866 29314
rect 28866 29262 28868 29314
rect 28812 29260 28868 29262
rect 28364 27916 28420 27972
rect 28588 27074 28644 27076
rect 28588 27022 28590 27074
rect 28590 27022 28642 27074
rect 28642 27022 28644 27074
rect 28588 27020 28644 27022
rect 29708 30322 29764 30324
rect 29708 30270 29710 30322
rect 29710 30270 29762 30322
rect 29762 30270 29764 30322
rect 29708 30268 29764 30270
rect 29596 29260 29652 29316
rect 29708 29036 29764 29092
rect 29484 28924 29540 28980
rect 30044 35532 30100 35588
rect 31052 40460 31108 40516
rect 30380 40402 30436 40404
rect 30380 40350 30382 40402
rect 30382 40350 30434 40402
rect 30434 40350 30436 40402
rect 30380 40348 30436 40350
rect 30380 40124 30436 40180
rect 30380 39116 30436 39172
rect 31836 40684 31892 40740
rect 31500 40402 31556 40404
rect 31500 40350 31502 40402
rect 31502 40350 31554 40402
rect 31554 40350 31556 40402
rect 31500 40348 31556 40350
rect 31948 39618 32004 39620
rect 31948 39566 31950 39618
rect 31950 39566 32002 39618
rect 32002 39566 32004 39618
rect 31948 39564 32004 39566
rect 30940 37996 30996 38052
rect 30492 37490 30548 37492
rect 30492 37438 30494 37490
rect 30494 37438 30546 37490
rect 30546 37438 30548 37490
rect 30492 37436 30548 37438
rect 30940 37490 30996 37492
rect 30940 37438 30942 37490
rect 30942 37438 30994 37490
rect 30994 37438 30996 37490
rect 30940 37436 30996 37438
rect 30268 36652 30324 36708
rect 30828 37324 30884 37380
rect 30156 34860 30212 34916
rect 31052 36258 31108 36260
rect 31052 36206 31054 36258
rect 31054 36206 31106 36258
rect 31106 36206 31108 36258
rect 31052 36204 31108 36206
rect 30492 35532 30548 35588
rect 30380 35420 30436 35476
rect 30828 34130 30884 34132
rect 30828 34078 30830 34130
rect 30830 34078 30882 34130
rect 30882 34078 30884 34130
rect 30828 34076 30884 34078
rect 30380 33964 30436 34020
rect 30380 32508 30436 32564
rect 31500 34914 31556 34916
rect 31500 34862 31502 34914
rect 31502 34862 31554 34914
rect 31554 34862 31556 34914
rect 31500 34860 31556 34862
rect 31276 34636 31332 34692
rect 32620 39618 32676 39620
rect 32620 39566 32622 39618
rect 32622 39566 32674 39618
rect 32674 39566 32676 39618
rect 32620 39564 32676 39566
rect 31948 37660 32004 37716
rect 32060 37490 32116 37492
rect 32060 37438 32062 37490
rect 32062 37438 32114 37490
rect 32114 37438 32116 37490
rect 32060 37436 32116 37438
rect 31948 36204 32004 36260
rect 31836 35420 31892 35476
rect 31948 35196 32004 35252
rect 31948 34748 32004 34804
rect 31612 34130 31668 34132
rect 31612 34078 31614 34130
rect 31614 34078 31666 34130
rect 31666 34078 31668 34130
rect 31612 34076 31668 34078
rect 31388 33964 31444 34020
rect 31052 33740 31108 33796
rect 31052 33516 31108 33572
rect 32396 37378 32452 37380
rect 32396 37326 32398 37378
rect 32398 37326 32450 37378
rect 32450 37326 32452 37378
rect 32396 37324 32452 37326
rect 32508 37436 32564 37492
rect 33404 39228 33460 39284
rect 34300 43426 34356 43428
rect 34300 43374 34302 43426
rect 34302 43374 34354 43426
rect 34354 43374 34356 43426
rect 34300 43372 34356 43374
rect 34636 43314 34692 43316
rect 34636 43262 34638 43314
rect 34638 43262 34690 43314
rect 34690 43262 34692 43314
rect 34636 43260 34692 43262
rect 34412 42978 34468 42980
rect 34412 42926 34414 42978
rect 34414 42926 34466 42978
rect 34466 42926 34468 42978
rect 34412 42924 34468 42926
rect 34748 43036 34804 43092
rect 34188 42364 34244 42420
rect 33964 40402 34020 40404
rect 33964 40350 33966 40402
rect 33966 40350 34018 40402
rect 34018 40350 34020 40402
rect 33964 40348 34020 40350
rect 33516 38220 33572 38276
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 35308 42642 35364 42644
rect 35308 42590 35310 42642
rect 35310 42590 35362 42642
rect 35362 42590 35364 42642
rect 35308 42588 35364 42590
rect 35196 42530 35252 42532
rect 35196 42478 35198 42530
rect 35198 42478 35250 42530
rect 35250 42478 35252 42530
rect 35196 42476 35252 42478
rect 35084 41916 35140 41972
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 35084 40514 35140 40516
rect 35084 40462 35086 40514
rect 35086 40462 35138 40514
rect 35138 40462 35140 40514
rect 35084 40460 35140 40462
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 35196 39340 35252 39396
rect 33404 37996 33460 38052
rect 33292 37938 33348 37940
rect 33292 37886 33294 37938
rect 33294 37886 33346 37938
rect 33346 37886 33348 37938
rect 33292 37884 33348 37886
rect 33292 37324 33348 37380
rect 32732 36988 32788 37044
rect 32396 35420 32452 35476
rect 32172 35084 32228 35140
rect 32396 34914 32452 34916
rect 32396 34862 32398 34914
rect 32398 34862 32450 34914
rect 32450 34862 32452 34914
rect 32396 34860 32452 34862
rect 32284 34802 32340 34804
rect 32284 34750 32286 34802
rect 32286 34750 32338 34802
rect 32338 34750 32340 34802
rect 32284 34748 32340 34750
rect 32172 34690 32228 34692
rect 32172 34638 32174 34690
rect 32174 34638 32226 34690
rect 32226 34638 32228 34690
rect 32172 34636 32228 34638
rect 32060 33516 32116 33572
rect 31836 33458 31892 33460
rect 31836 33406 31838 33458
rect 31838 33406 31890 33458
rect 31890 33406 31892 33458
rect 31836 33404 31892 33406
rect 33404 37266 33460 37268
rect 33404 37214 33406 37266
rect 33406 37214 33458 37266
rect 33458 37214 33460 37266
rect 33404 37212 33460 37214
rect 33740 38108 33796 38164
rect 33628 37378 33684 37380
rect 33628 37326 33630 37378
rect 33630 37326 33682 37378
rect 33682 37326 33684 37378
rect 33628 37324 33684 37326
rect 33964 37884 34020 37940
rect 33852 37826 33908 37828
rect 33852 37774 33854 37826
rect 33854 37774 33906 37826
rect 33906 37774 33908 37826
rect 33852 37772 33908 37774
rect 34300 37324 34356 37380
rect 35868 43538 35924 43540
rect 35868 43486 35870 43538
rect 35870 43486 35922 43538
rect 35922 43486 35924 43538
rect 35868 43484 35924 43486
rect 37212 42924 37268 42980
rect 37324 43484 37380 43540
rect 37212 42754 37268 42756
rect 37212 42702 37214 42754
rect 37214 42702 37266 42754
rect 37266 42702 37268 42754
rect 37212 42700 37268 42702
rect 36540 41804 36596 41860
rect 36540 41244 36596 41300
rect 36204 41186 36260 41188
rect 36204 41134 36206 41186
rect 36206 41134 36258 41186
rect 36258 41134 36260 41186
rect 36204 41132 36260 41134
rect 36428 40962 36484 40964
rect 36428 40910 36430 40962
rect 36430 40910 36482 40962
rect 36482 40910 36484 40962
rect 36428 40908 36484 40910
rect 36764 40908 36820 40964
rect 37548 44940 37604 44996
rect 39004 45724 39060 45780
rect 40012 45724 40068 45780
rect 38668 45612 38724 45668
rect 38108 44940 38164 44996
rect 37548 44210 37604 44212
rect 37548 44158 37550 44210
rect 37550 44158 37602 44210
rect 37602 44158 37604 44210
rect 37548 44156 37604 44158
rect 37660 43484 37716 43540
rect 37436 43260 37492 43316
rect 37772 42700 37828 42756
rect 37548 42364 37604 42420
rect 37884 41580 37940 41636
rect 37772 41244 37828 41300
rect 37324 41186 37380 41188
rect 37324 41134 37326 41186
rect 37326 41134 37378 41186
rect 37378 41134 37380 41186
rect 37324 41132 37380 41134
rect 37548 41074 37604 41076
rect 37548 41022 37550 41074
rect 37550 41022 37602 41074
rect 37602 41022 37604 41074
rect 37548 41020 37604 41022
rect 37884 40962 37940 40964
rect 37884 40910 37886 40962
rect 37886 40910 37938 40962
rect 37938 40910 37940 40962
rect 37884 40908 37940 40910
rect 38220 44156 38276 44212
rect 38332 41186 38388 41188
rect 38332 41134 38334 41186
rect 38334 41134 38386 41186
rect 38386 41134 38388 41186
rect 38332 41132 38388 41134
rect 39564 45106 39620 45108
rect 39564 45054 39566 45106
rect 39566 45054 39618 45106
rect 39618 45054 39620 45106
rect 39564 45052 39620 45054
rect 39116 44156 39172 44212
rect 39116 43260 39172 43316
rect 39004 42924 39060 42980
rect 39676 44322 39732 44324
rect 39676 44270 39678 44322
rect 39678 44270 39730 44322
rect 39730 44270 39732 44322
rect 39676 44268 39732 44270
rect 40236 45052 40292 45108
rect 40348 44940 40404 44996
rect 40236 44882 40292 44884
rect 40236 44830 40238 44882
rect 40238 44830 40290 44882
rect 40290 44830 40292 44882
rect 40236 44828 40292 44830
rect 40348 44716 40404 44772
rect 40236 44156 40292 44212
rect 38556 41074 38612 41076
rect 38556 41022 38558 41074
rect 38558 41022 38610 41074
rect 38610 41022 38612 41074
rect 38556 41020 38612 41022
rect 39004 40908 39060 40964
rect 36540 40012 36596 40068
rect 35868 39506 35924 39508
rect 35868 39454 35870 39506
rect 35870 39454 35922 39506
rect 35922 39454 35924 39506
rect 35868 39452 35924 39454
rect 36540 39452 36596 39508
rect 36652 39676 36708 39732
rect 37100 40236 37156 40292
rect 37100 39788 37156 39844
rect 37660 40348 37716 40404
rect 36988 39564 37044 39620
rect 39340 42642 39396 42644
rect 39340 42590 39342 42642
rect 39342 42590 39394 42642
rect 39394 42590 39396 42642
rect 39340 42588 39396 42590
rect 39788 43372 39844 43428
rect 40124 43650 40180 43652
rect 40124 43598 40126 43650
rect 40126 43598 40178 43650
rect 40178 43598 40180 43650
rect 40124 43596 40180 43598
rect 40012 43260 40068 43316
rect 40348 43596 40404 43652
rect 39676 42364 39732 42420
rect 39900 42252 39956 42308
rect 39788 41580 39844 41636
rect 39452 41244 39508 41300
rect 39788 40572 39844 40628
rect 36652 38892 36708 38948
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 34524 37266 34580 37268
rect 34524 37214 34526 37266
rect 34526 37214 34578 37266
rect 34578 37214 34580 37266
rect 34524 37212 34580 37214
rect 34076 37042 34132 37044
rect 34076 36990 34078 37042
rect 34078 36990 34130 37042
rect 34130 36990 34132 37042
rect 34076 36988 34132 36990
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 34972 35980 35028 36036
rect 35644 36764 35700 36820
rect 33404 35138 33460 35140
rect 33404 35086 33406 35138
rect 33406 35086 33458 35138
rect 33458 35086 33460 35138
rect 33404 35084 33460 35086
rect 33628 35532 33684 35588
rect 33964 35084 34020 35140
rect 34412 35586 34468 35588
rect 34412 35534 34414 35586
rect 34414 35534 34466 35586
rect 34466 35534 34468 35586
rect 34412 35532 34468 35534
rect 35420 35532 35476 35588
rect 33628 35026 33684 35028
rect 33628 34974 33630 35026
rect 33630 34974 33682 35026
rect 33682 34974 33684 35026
rect 33628 34972 33684 34974
rect 33740 34242 33796 34244
rect 33740 34190 33742 34242
rect 33742 34190 33794 34242
rect 33794 34190 33796 34242
rect 33740 34188 33796 34190
rect 33628 33740 33684 33796
rect 32732 33516 32788 33572
rect 33516 33516 33572 33572
rect 32844 33404 32900 33460
rect 30604 31948 30660 32004
rect 30044 31836 30100 31892
rect 30044 31500 30100 31556
rect 30940 32396 30996 32452
rect 31724 32450 31780 32452
rect 31724 32398 31726 32450
rect 31726 32398 31778 32450
rect 31778 32398 31780 32450
rect 31724 32396 31780 32398
rect 31836 32508 31892 32564
rect 29932 30716 29988 30772
rect 29932 30044 29988 30100
rect 29932 29596 29988 29652
rect 30044 30940 30100 30996
rect 30492 30434 30548 30436
rect 30492 30382 30494 30434
rect 30494 30382 30546 30434
rect 30546 30382 30548 30434
rect 30492 30380 30548 30382
rect 30268 30098 30324 30100
rect 30268 30046 30270 30098
rect 30270 30046 30322 30098
rect 30322 30046 30324 30098
rect 30268 30044 30324 30046
rect 31388 30940 31444 30996
rect 32060 32450 32116 32452
rect 32060 32398 32062 32450
rect 32062 32398 32114 32450
rect 32114 32398 32116 32450
rect 32060 32396 32116 32398
rect 33628 32284 33684 32340
rect 32284 30994 32340 30996
rect 32284 30942 32286 30994
rect 32286 30942 32338 30994
rect 32338 30942 32340 30994
rect 32284 30940 32340 30942
rect 30828 29484 30884 29540
rect 32284 30380 32340 30436
rect 33292 31948 33348 32004
rect 32508 31106 32564 31108
rect 32508 31054 32510 31106
rect 32510 31054 32562 31106
rect 32562 31054 32564 31106
rect 32508 31052 32564 31054
rect 31612 30322 31668 30324
rect 31612 30270 31614 30322
rect 31614 30270 31666 30322
rect 31666 30270 31668 30322
rect 31612 30268 31668 30270
rect 32060 30156 32116 30212
rect 30716 28924 30772 28980
rect 30380 28642 30436 28644
rect 30380 28590 30382 28642
rect 30382 28590 30434 28642
rect 30434 28590 30436 28642
rect 30380 28588 30436 28590
rect 30156 28418 30212 28420
rect 30156 28366 30158 28418
rect 30158 28366 30210 28418
rect 30210 28366 30212 28418
rect 30156 28364 30212 28366
rect 29484 28252 29540 28308
rect 31052 29036 31108 29092
rect 30828 28642 30884 28644
rect 30828 28590 30830 28642
rect 30830 28590 30882 28642
rect 30882 28590 30884 28642
rect 30828 28588 30884 28590
rect 29484 27132 29540 27188
rect 27244 23938 27300 23940
rect 27244 23886 27246 23938
rect 27246 23886 27298 23938
rect 27298 23886 27300 23938
rect 27244 23884 27300 23886
rect 27244 22876 27300 22932
rect 27804 24892 27860 24948
rect 28028 24892 28084 24948
rect 27916 24722 27972 24724
rect 27916 24670 27918 24722
rect 27918 24670 27970 24722
rect 27970 24670 27972 24722
rect 27916 24668 27972 24670
rect 27804 24556 27860 24612
rect 28028 24108 28084 24164
rect 27692 23772 27748 23828
rect 27020 21756 27076 21812
rect 28252 25900 28308 25956
rect 28252 25394 28308 25396
rect 28252 25342 28254 25394
rect 28254 25342 28306 25394
rect 28306 25342 28308 25394
rect 28252 25340 28308 25342
rect 28364 25228 28420 25284
rect 28924 26796 28980 26852
rect 28588 26402 28644 26404
rect 28588 26350 28590 26402
rect 28590 26350 28642 26402
rect 28642 26350 28644 26402
rect 28588 26348 28644 26350
rect 29148 26514 29204 26516
rect 29148 26462 29150 26514
rect 29150 26462 29202 26514
rect 29202 26462 29204 26514
rect 29148 26460 29204 26462
rect 29260 26402 29316 26404
rect 29260 26350 29262 26402
rect 29262 26350 29314 26402
rect 29314 26350 29316 26402
rect 29260 26348 29316 26350
rect 28924 25564 28980 25620
rect 29036 26012 29092 26068
rect 28588 25282 28644 25284
rect 28588 25230 28590 25282
rect 28590 25230 28642 25282
rect 28642 25230 28644 25282
rect 28588 25228 28644 25230
rect 28588 25004 28644 25060
rect 28812 24834 28868 24836
rect 28812 24782 28814 24834
rect 28814 24782 28866 24834
rect 28866 24782 28868 24834
rect 28812 24780 28868 24782
rect 28588 23996 28644 24052
rect 28364 23548 28420 23604
rect 29596 27074 29652 27076
rect 29596 27022 29598 27074
rect 29598 27022 29650 27074
rect 29650 27022 29652 27074
rect 29596 27020 29652 27022
rect 30940 28082 30996 28084
rect 30940 28030 30942 28082
rect 30942 28030 30994 28082
rect 30994 28030 30996 28082
rect 30940 28028 30996 28030
rect 30380 27580 30436 27636
rect 30156 27186 30212 27188
rect 30156 27134 30158 27186
rect 30158 27134 30210 27186
rect 30210 27134 30212 27186
rect 30156 27132 30212 27134
rect 29932 27020 29988 27076
rect 29820 26908 29876 26964
rect 29484 25452 29540 25508
rect 29596 26012 29652 26068
rect 29148 25282 29204 25284
rect 29148 25230 29150 25282
rect 29150 25230 29202 25282
rect 29202 25230 29204 25282
rect 29148 25228 29204 25230
rect 29484 24556 29540 24612
rect 29148 24444 29204 24500
rect 29708 25676 29764 25732
rect 29596 24332 29652 24388
rect 29708 24668 29764 24724
rect 29372 23714 29428 23716
rect 29372 23662 29374 23714
rect 29374 23662 29426 23714
rect 29426 23662 29428 23714
rect 29372 23660 29428 23662
rect 28588 22652 28644 22708
rect 27020 21026 27076 21028
rect 27020 20974 27022 21026
rect 27022 20974 27074 21026
rect 27074 20974 27076 21026
rect 27020 20972 27076 20974
rect 26124 20524 26180 20580
rect 26908 20578 26964 20580
rect 26908 20526 26910 20578
rect 26910 20526 26962 20578
rect 26962 20526 26964 20578
rect 26908 20524 26964 20526
rect 26012 20188 26068 20244
rect 26236 20412 26292 20468
rect 26124 20076 26180 20132
rect 26012 20018 26068 20020
rect 26012 19966 26014 20018
rect 26014 19966 26066 20018
rect 26066 19966 26068 20018
rect 26012 19964 26068 19966
rect 25788 19740 25844 19796
rect 27020 20076 27076 20132
rect 28140 21196 28196 21252
rect 28140 21026 28196 21028
rect 28140 20974 28142 21026
rect 28142 20974 28194 21026
rect 28194 20974 28196 21026
rect 28140 20972 28196 20974
rect 27580 20690 27636 20692
rect 27580 20638 27582 20690
rect 27582 20638 27634 20690
rect 27634 20638 27636 20690
rect 27580 20636 27636 20638
rect 27804 20690 27860 20692
rect 27804 20638 27806 20690
rect 27806 20638 27858 20690
rect 27858 20638 27860 20690
rect 27804 20636 27860 20638
rect 28252 20578 28308 20580
rect 28252 20526 28254 20578
rect 28254 20526 28306 20578
rect 28306 20526 28308 20578
rect 28252 20524 28308 20526
rect 27692 20130 27748 20132
rect 27692 20078 27694 20130
rect 27694 20078 27746 20130
rect 27746 20078 27748 20130
rect 27692 20076 27748 20078
rect 28924 22988 28980 23044
rect 28700 22146 28756 22148
rect 28700 22094 28702 22146
rect 28702 22094 28754 22146
rect 28754 22094 28756 22146
rect 28700 22092 28756 22094
rect 28812 21644 28868 21700
rect 29596 22988 29652 23044
rect 30044 26460 30100 26516
rect 30492 27074 30548 27076
rect 30492 27022 30494 27074
rect 30494 27022 30546 27074
rect 30546 27022 30548 27074
rect 30492 27020 30548 27022
rect 30716 26348 30772 26404
rect 30044 24332 30100 24388
rect 30492 25452 30548 25508
rect 30716 25340 30772 25396
rect 29820 21644 29876 21700
rect 29932 23772 29988 23828
rect 29260 21196 29316 21252
rect 29036 20690 29092 20692
rect 29036 20638 29038 20690
rect 29038 20638 29090 20690
rect 29090 20638 29092 20690
rect 29036 20636 29092 20638
rect 28924 20524 28980 20580
rect 29148 20524 29204 20580
rect 29036 20018 29092 20020
rect 29036 19966 29038 20018
rect 29038 19966 29090 20018
rect 29090 19966 29092 20018
rect 29036 19964 29092 19966
rect 25228 19122 25284 19124
rect 25228 19070 25230 19122
rect 25230 19070 25282 19122
rect 25282 19070 25284 19122
rect 25228 19068 25284 19070
rect 25900 19122 25956 19124
rect 25900 19070 25902 19122
rect 25902 19070 25954 19122
rect 25954 19070 25956 19122
rect 25900 19068 25956 19070
rect 23996 16940 24052 16996
rect 23996 15986 24052 15988
rect 23996 15934 23998 15986
rect 23998 15934 24050 15986
rect 24050 15934 24052 15986
rect 23996 15932 24052 15934
rect 26572 18508 26628 18564
rect 27132 19292 27188 19348
rect 27356 19068 27412 19124
rect 27244 18396 27300 18452
rect 24668 17500 24724 17556
rect 24780 16940 24836 16996
rect 26796 17612 26852 17668
rect 25564 17442 25620 17444
rect 25564 17390 25566 17442
rect 25566 17390 25618 17442
rect 25618 17390 25620 17442
rect 25564 17388 25620 17390
rect 26460 17388 26516 17444
rect 26572 17500 26628 17556
rect 25004 16268 25060 16324
rect 23884 15538 23940 15540
rect 23884 15486 23886 15538
rect 23886 15486 23938 15538
rect 23938 15486 23940 15538
rect 23884 15484 23940 15486
rect 23996 15426 24052 15428
rect 23996 15374 23998 15426
rect 23998 15374 24050 15426
rect 24050 15374 24052 15426
rect 23996 15372 24052 15374
rect 23548 15260 23604 15316
rect 22428 14418 22484 14420
rect 22428 14366 22430 14418
rect 22430 14366 22482 14418
rect 22482 14366 22484 14418
rect 22428 14364 22484 14366
rect 25676 15986 25732 15988
rect 25676 15934 25678 15986
rect 25678 15934 25730 15986
rect 25730 15934 25732 15986
rect 25676 15932 25732 15934
rect 26236 15932 26292 15988
rect 25900 15538 25956 15540
rect 25900 15486 25902 15538
rect 25902 15486 25954 15538
rect 25954 15486 25956 15538
rect 25900 15484 25956 15486
rect 27020 17666 27076 17668
rect 27020 17614 27022 17666
rect 27022 17614 27074 17666
rect 27074 17614 27076 17666
rect 27020 17612 27076 17614
rect 27244 17666 27300 17668
rect 27244 17614 27246 17666
rect 27246 17614 27298 17666
rect 27298 17614 27300 17666
rect 27244 17612 27300 17614
rect 26348 15148 26404 15204
rect 27692 19292 27748 19348
rect 28140 19234 28196 19236
rect 28140 19182 28142 19234
rect 28142 19182 28194 19234
rect 28194 19182 28196 19234
rect 28140 19180 28196 19182
rect 28476 19292 28532 19348
rect 28588 19122 28644 19124
rect 28588 19070 28590 19122
rect 28590 19070 28642 19122
rect 28642 19070 28644 19122
rect 28588 19068 28644 19070
rect 29372 20690 29428 20692
rect 29372 20638 29374 20690
rect 29374 20638 29426 20690
rect 29426 20638 29428 20690
rect 29372 20636 29428 20638
rect 29036 19180 29092 19236
rect 29820 20300 29876 20356
rect 30044 23660 30100 23716
rect 30380 25004 30436 25060
rect 30828 24780 30884 24836
rect 30940 25282 30996 25284
rect 30940 25230 30942 25282
rect 30942 25230 30994 25282
rect 30994 25230 30996 25282
rect 30940 25228 30996 25230
rect 30604 23884 30660 23940
rect 30828 23884 30884 23940
rect 30940 23660 30996 23716
rect 31164 26684 31220 26740
rect 31500 30098 31556 30100
rect 31500 30046 31502 30098
rect 31502 30046 31554 30098
rect 31554 30046 31556 30098
rect 31500 30044 31556 30046
rect 31948 30098 32004 30100
rect 31948 30046 31950 30098
rect 31950 30046 32002 30098
rect 32002 30046 32004 30098
rect 31948 30044 32004 30046
rect 32508 30210 32564 30212
rect 32508 30158 32510 30210
rect 32510 30158 32562 30210
rect 32562 30158 32564 30210
rect 32508 30156 32564 30158
rect 33068 30156 33124 30212
rect 32172 30098 32228 30100
rect 32172 30046 32174 30098
rect 32174 30046 32226 30098
rect 32226 30046 32228 30098
rect 32172 30044 32228 30046
rect 31388 29260 31444 29316
rect 32284 29372 32340 29428
rect 31724 28700 31780 28756
rect 31836 29260 31892 29316
rect 31612 26908 31668 26964
rect 32060 29148 32116 29204
rect 31836 26572 31892 26628
rect 31948 28364 32004 28420
rect 31276 26460 31332 26516
rect 31612 26236 31668 26292
rect 33180 29148 33236 29204
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 34748 34860 34804 34916
rect 34524 34802 34580 34804
rect 34524 34750 34526 34802
rect 34526 34750 34578 34802
rect 34578 34750 34580 34802
rect 34524 34748 34580 34750
rect 34748 34188 34804 34244
rect 33964 34130 34020 34132
rect 33964 34078 33966 34130
rect 33966 34078 34018 34130
rect 34018 34078 34020 34130
rect 33964 34076 34020 34078
rect 34636 34130 34692 34132
rect 34636 34078 34638 34130
rect 34638 34078 34690 34130
rect 34690 34078 34692 34130
rect 34636 34076 34692 34078
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 34748 33404 34804 33460
rect 34300 33346 34356 33348
rect 34300 33294 34302 33346
rect 34302 33294 34354 33346
rect 34354 33294 34356 33346
rect 34300 33292 34356 33294
rect 34524 31890 34580 31892
rect 34524 31838 34526 31890
rect 34526 31838 34578 31890
rect 34578 31838 34580 31890
rect 34524 31836 34580 31838
rect 34748 31612 34804 31668
rect 35532 33404 35588 33460
rect 34972 33180 35028 33236
rect 35644 33346 35700 33348
rect 35644 33294 35646 33346
rect 35646 33294 35698 33346
rect 35698 33294 35700 33346
rect 35644 33292 35700 33294
rect 35756 33180 35812 33236
rect 35084 32284 35140 32340
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35196 31836 35252 31892
rect 34972 31500 35028 31556
rect 34188 30940 34244 30996
rect 33740 29708 33796 29764
rect 32396 28812 32452 28868
rect 32732 28700 32788 28756
rect 32396 28028 32452 28084
rect 32732 28028 32788 28084
rect 32060 26290 32116 26292
rect 32060 26238 32062 26290
rect 32062 26238 32114 26290
rect 32114 26238 32116 26290
rect 32060 26236 32116 26238
rect 32396 26348 32452 26404
rect 31612 25340 31668 25396
rect 31276 23996 31332 24052
rect 32060 25004 32116 25060
rect 32284 25228 32340 25284
rect 31836 24892 31892 24948
rect 31612 23660 31668 23716
rect 31164 23436 31220 23492
rect 31836 23660 31892 23716
rect 32060 23996 32116 24052
rect 31724 23436 31780 23492
rect 31948 22988 32004 23044
rect 32172 23938 32228 23940
rect 32172 23886 32174 23938
rect 32174 23886 32226 23938
rect 32226 23886 32228 23938
rect 32172 23884 32228 23886
rect 32732 24892 32788 24948
rect 33180 28082 33236 28084
rect 33180 28030 33182 28082
rect 33182 28030 33234 28082
rect 33234 28030 33236 28082
rect 33180 28028 33236 28030
rect 33628 29426 33684 29428
rect 33628 29374 33630 29426
rect 33630 29374 33682 29426
rect 33682 29374 33684 29426
rect 33628 29372 33684 29374
rect 33852 29426 33908 29428
rect 33852 29374 33854 29426
rect 33854 29374 33906 29426
rect 33906 29374 33908 29426
rect 33852 29372 33908 29374
rect 34076 29148 34132 29204
rect 33516 28476 33572 28532
rect 33628 28252 33684 28308
rect 33404 26572 33460 26628
rect 36316 37266 36372 37268
rect 36316 37214 36318 37266
rect 36318 37214 36370 37266
rect 36370 37214 36372 37266
rect 36316 37212 36372 37214
rect 39116 39394 39172 39396
rect 39116 39342 39118 39394
rect 39118 39342 39170 39394
rect 39170 39342 39172 39394
rect 39116 39340 39172 39342
rect 36540 38722 36596 38724
rect 36540 38670 36542 38722
rect 36542 38670 36594 38722
rect 36594 38670 36596 38722
rect 36540 38668 36596 38670
rect 37100 38108 37156 38164
rect 37100 37212 37156 37268
rect 37212 37772 37268 37828
rect 36092 35756 36148 35812
rect 36540 35810 36596 35812
rect 36540 35758 36542 35810
rect 36542 35758 36594 35810
rect 36594 35758 36596 35810
rect 36540 35756 36596 35758
rect 36876 35698 36932 35700
rect 36876 35646 36878 35698
rect 36878 35646 36930 35698
rect 36930 35646 36932 35698
rect 36876 35644 36932 35646
rect 36316 35532 36372 35588
rect 36092 34914 36148 34916
rect 36092 34862 36094 34914
rect 36094 34862 36146 34914
rect 36146 34862 36148 34914
rect 36092 34860 36148 34862
rect 35980 34802 36036 34804
rect 35980 34750 35982 34802
rect 35982 34750 36034 34802
rect 36034 34750 36036 34802
rect 35980 34748 36036 34750
rect 37100 35532 37156 35588
rect 36652 35474 36708 35476
rect 36652 35422 36654 35474
rect 36654 35422 36706 35474
rect 36706 35422 36708 35474
rect 36652 35420 36708 35422
rect 36316 35084 36372 35140
rect 37772 38668 37828 38724
rect 39676 39618 39732 39620
rect 39676 39566 39678 39618
rect 39678 39566 39730 39618
rect 39730 39566 39732 39618
rect 39676 39564 39732 39566
rect 39788 39340 39844 39396
rect 38444 38108 38500 38164
rect 39340 38220 39396 38276
rect 37772 36876 37828 36932
rect 38332 37324 38388 37380
rect 40348 42588 40404 42644
rect 40124 42364 40180 42420
rect 40236 42140 40292 42196
rect 41020 45836 41076 45892
rect 41356 46060 41412 46116
rect 40572 44268 40628 44324
rect 40684 45164 40740 45220
rect 40684 43708 40740 43764
rect 40124 40962 40180 40964
rect 40124 40910 40126 40962
rect 40126 40910 40178 40962
rect 40178 40910 40180 40962
rect 40124 40908 40180 40910
rect 40012 38780 40068 38836
rect 40124 39788 40180 39844
rect 39900 38220 39956 38276
rect 39788 37490 39844 37492
rect 39788 37438 39790 37490
rect 39790 37438 39842 37490
rect 39842 37438 39844 37490
rect 39788 37436 39844 37438
rect 41020 45276 41076 45332
rect 41020 44716 41076 44772
rect 41356 44994 41412 44996
rect 41356 44942 41358 44994
rect 41358 44942 41410 44994
rect 41410 44942 41412 44994
rect 41356 44940 41412 44942
rect 41356 44044 41412 44100
rect 40908 43708 40964 43764
rect 41244 43596 41300 43652
rect 41132 42978 41188 42980
rect 41132 42926 41134 42978
rect 41134 42926 41186 42978
rect 41186 42926 41188 42978
rect 41132 42924 41188 42926
rect 41020 42028 41076 42084
rect 41132 42588 41188 42644
rect 41356 43538 41412 43540
rect 41356 43486 41358 43538
rect 41358 43486 41410 43538
rect 41410 43486 41412 43538
rect 41356 43484 41412 43486
rect 41580 45052 41636 45108
rect 42252 46172 42308 46228
rect 44380 46844 44436 46900
rect 42588 46060 42644 46116
rect 42364 45778 42420 45780
rect 42364 45726 42366 45778
rect 42366 45726 42418 45778
rect 42418 45726 42420 45778
rect 42364 45724 42420 45726
rect 42252 45218 42308 45220
rect 42252 45166 42254 45218
rect 42254 45166 42306 45218
rect 42306 45166 42308 45218
rect 42252 45164 42308 45166
rect 41804 45052 41860 45108
rect 41692 44604 41748 44660
rect 41916 44044 41972 44100
rect 42028 43932 42084 43988
rect 42588 45052 42644 45108
rect 41244 42140 41300 42196
rect 41580 43484 41636 43540
rect 41804 43538 41860 43540
rect 41804 43486 41806 43538
rect 41806 43486 41858 43538
rect 41858 43486 41860 43538
rect 41804 43484 41860 43486
rect 41804 42754 41860 42756
rect 41804 42702 41806 42754
rect 41806 42702 41858 42754
rect 41858 42702 41860 42754
rect 41804 42700 41860 42702
rect 43036 45724 43092 45780
rect 43596 45724 43652 45780
rect 43148 45666 43204 45668
rect 43148 45614 43150 45666
rect 43150 45614 43202 45666
rect 43202 45614 43204 45666
rect 43148 45612 43204 45614
rect 42924 45106 42980 45108
rect 42924 45054 42926 45106
rect 42926 45054 42978 45106
rect 42978 45054 42980 45106
rect 42924 45052 42980 45054
rect 42812 44210 42868 44212
rect 42812 44158 42814 44210
rect 42814 44158 42866 44210
rect 42866 44158 42868 44210
rect 42812 44156 42868 44158
rect 42700 43652 42756 43708
rect 42924 44044 42980 44100
rect 43372 44994 43428 44996
rect 43372 44942 43374 44994
rect 43374 44942 43426 44994
rect 43426 44942 43428 44994
rect 43372 44940 43428 44942
rect 43036 43708 43092 43764
rect 43708 44492 43764 44548
rect 44268 45164 44324 45220
rect 44156 45106 44212 45108
rect 44156 45054 44158 45106
rect 44158 45054 44210 45106
rect 44210 45054 44212 45106
rect 44156 45052 44212 45054
rect 44604 46060 44660 46116
rect 44380 44828 44436 44884
rect 44940 45164 44996 45220
rect 44156 44156 44212 44212
rect 44156 43652 44212 43708
rect 42140 43036 42196 43092
rect 42812 42700 42868 42756
rect 42028 42588 42084 42644
rect 41692 42476 41748 42532
rect 42700 42642 42756 42644
rect 42700 42590 42702 42642
rect 42702 42590 42754 42642
rect 42754 42590 42756 42642
rect 42700 42588 42756 42590
rect 41804 42028 41860 42084
rect 40348 40684 40404 40740
rect 40348 40236 40404 40292
rect 40460 40572 40516 40628
rect 41356 40962 41412 40964
rect 41356 40910 41358 40962
rect 41358 40910 41410 40962
rect 41410 40910 41412 40962
rect 41356 40908 41412 40910
rect 41580 40796 41636 40852
rect 41692 40684 41748 40740
rect 41132 40124 41188 40180
rect 40684 39730 40740 39732
rect 40684 39678 40686 39730
rect 40686 39678 40738 39730
rect 40738 39678 40740 39730
rect 40684 39676 40740 39678
rect 42700 42364 42756 42420
rect 42476 42028 42532 42084
rect 42812 42028 42868 42084
rect 42364 41804 42420 41860
rect 42476 41746 42532 41748
rect 42476 41694 42478 41746
rect 42478 41694 42530 41746
rect 42530 41694 42532 41746
rect 42476 41692 42532 41694
rect 43820 42476 43876 42532
rect 44268 43484 44324 43540
rect 45276 44380 45332 44436
rect 44604 43708 44660 43764
rect 44380 42924 44436 42980
rect 43372 42082 43428 42084
rect 43372 42030 43374 42082
rect 43374 42030 43426 42082
rect 43426 42030 43428 42082
rect 43372 42028 43428 42030
rect 43148 41970 43204 41972
rect 43148 41918 43150 41970
rect 43150 41918 43202 41970
rect 43202 41918 43204 41970
rect 43148 41916 43204 41918
rect 42364 41356 42420 41412
rect 42140 40124 42196 40180
rect 42588 40962 42644 40964
rect 42588 40910 42590 40962
rect 42590 40910 42642 40962
rect 42642 40910 42644 40962
rect 42588 40908 42644 40910
rect 43036 40684 43092 40740
rect 43372 40684 43428 40740
rect 42364 40348 42420 40404
rect 40908 38834 40964 38836
rect 40908 38782 40910 38834
rect 40910 38782 40962 38834
rect 40962 38782 40964 38834
rect 40908 38780 40964 38782
rect 40236 38332 40292 38388
rect 40012 37996 40068 38052
rect 39452 37324 39508 37380
rect 41244 39676 41300 39732
rect 40348 38108 40404 38164
rect 40236 37884 40292 37940
rect 40460 37884 40516 37940
rect 37660 35980 37716 36036
rect 37324 35810 37380 35812
rect 37324 35758 37326 35810
rect 37326 35758 37378 35810
rect 37378 35758 37380 35810
rect 37324 35756 37380 35758
rect 37436 35698 37492 35700
rect 37436 35646 37438 35698
rect 37438 35646 37490 35698
rect 37490 35646 37492 35698
rect 37436 35644 37492 35646
rect 37436 35420 37492 35476
rect 38108 35756 38164 35812
rect 37996 35644 38052 35700
rect 38444 35420 38500 35476
rect 38556 35532 38612 35588
rect 38332 34860 38388 34916
rect 36316 33852 36372 33908
rect 36876 34130 36932 34132
rect 36876 34078 36878 34130
rect 36878 34078 36930 34130
rect 36930 34078 36932 34130
rect 36876 34076 36932 34078
rect 36540 33404 36596 33460
rect 38780 35698 38836 35700
rect 38780 35646 38782 35698
rect 38782 35646 38834 35698
rect 38834 35646 38836 35698
rect 38780 35644 38836 35646
rect 39228 35698 39284 35700
rect 39228 35646 39230 35698
rect 39230 35646 39282 35698
rect 39282 35646 39284 35698
rect 39228 35644 39284 35646
rect 42252 39452 42308 39508
rect 41468 39394 41524 39396
rect 41468 39342 41470 39394
rect 41470 39342 41522 39394
rect 41522 39342 41524 39394
rect 41468 39340 41524 39342
rect 42252 39116 42308 39172
rect 43260 40402 43316 40404
rect 43260 40350 43262 40402
rect 43262 40350 43314 40402
rect 43314 40350 43316 40402
rect 43260 40348 43316 40350
rect 42700 40124 42756 40180
rect 43820 41970 43876 41972
rect 43820 41918 43822 41970
rect 43822 41918 43874 41970
rect 43874 41918 43876 41970
rect 43820 41916 43876 41918
rect 43708 41804 43764 41860
rect 43596 41692 43652 41748
rect 44828 42194 44884 42196
rect 44828 42142 44830 42194
rect 44830 42142 44882 42194
rect 44882 42142 44884 42194
rect 44828 42140 44884 42142
rect 44156 41410 44212 41412
rect 44156 41358 44158 41410
rect 44158 41358 44210 41410
rect 44210 41358 44212 41410
rect 44156 41356 44212 41358
rect 43596 40572 43652 40628
rect 44268 40796 44324 40852
rect 44156 40626 44212 40628
rect 44156 40574 44158 40626
rect 44158 40574 44210 40626
rect 44210 40574 44212 40626
rect 44156 40572 44212 40574
rect 43148 39506 43204 39508
rect 43148 39454 43150 39506
rect 43150 39454 43202 39506
rect 43202 39454 43204 39506
rect 43148 39452 43204 39454
rect 44044 40290 44100 40292
rect 44044 40238 44046 40290
rect 44046 40238 44098 40290
rect 44098 40238 44100 40290
rect 44044 40236 44100 40238
rect 41916 38834 41972 38836
rect 41916 38782 41918 38834
rect 41918 38782 41970 38834
rect 41970 38782 41972 38834
rect 41916 38780 41972 38782
rect 41580 38668 41636 38724
rect 42924 39058 42980 39060
rect 42924 39006 42926 39058
rect 42926 39006 42978 39058
rect 42978 39006 42980 39058
rect 42924 39004 42980 39006
rect 42252 38668 42308 38724
rect 41580 38050 41636 38052
rect 41580 37998 41582 38050
rect 41582 37998 41634 38050
rect 41634 37998 41636 38050
rect 41580 37996 41636 37998
rect 41804 37996 41860 38052
rect 41132 36652 41188 36708
rect 40012 35756 40068 35812
rect 41468 36594 41524 36596
rect 41468 36542 41470 36594
rect 41470 36542 41522 36594
rect 41522 36542 41524 36594
rect 41468 36540 41524 36542
rect 41580 36876 41636 36932
rect 41356 36092 41412 36148
rect 42700 37996 42756 38052
rect 42476 37938 42532 37940
rect 42476 37886 42478 37938
rect 42478 37886 42530 37938
rect 42530 37886 42532 37938
rect 42476 37884 42532 37886
rect 42028 36540 42084 36596
rect 44716 41580 44772 41636
rect 45052 43708 45108 43764
rect 45388 42978 45444 42980
rect 45388 42926 45390 42978
rect 45390 42926 45442 42978
rect 45442 42926 45444 42978
rect 45388 42924 45444 42926
rect 45164 42476 45220 42532
rect 45052 41858 45108 41860
rect 45052 41806 45054 41858
rect 45054 41806 45106 41858
rect 45106 41806 45108 41858
rect 45052 41804 45108 41806
rect 44716 40684 44772 40740
rect 44604 40402 44660 40404
rect 44604 40350 44606 40402
rect 44606 40350 44658 40402
rect 44658 40350 44660 40402
rect 44604 40348 44660 40350
rect 44940 40236 44996 40292
rect 44828 39058 44884 39060
rect 44828 39006 44830 39058
rect 44830 39006 44882 39058
rect 44882 39006 44884 39058
rect 44828 39004 44884 39006
rect 45276 41916 45332 41972
rect 51436 46844 51492 46900
rect 46396 45836 46452 45892
rect 47404 46172 47460 46228
rect 45724 45164 45780 45220
rect 45612 43538 45668 43540
rect 45612 43486 45614 43538
rect 45614 43486 45666 43538
rect 45666 43486 45668 43538
rect 45612 43484 45668 43486
rect 45836 43596 45892 43652
rect 46732 45778 46788 45780
rect 46732 45726 46734 45778
rect 46734 45726 46786 45778
rect 46786 45726 46788 45778
rect 46732 45724 46788 45726
rect 46284 45612 46340 45668
rect 46396 45276 46452 45332
rect 47628 44940 47684 44996
rect 46060 43484 46116 43540
rect 45948 43372 46004 43428
rect 45836 42530 45892 42532
rect 45836 42478 45838 42530
rect 45838 42478 45890 42530
rect 45890 42478 45892 42530
rect 45836 42476 45892 42478
rect 45724 42140 45780 42196
rect 46956 43596 47012 43652
rect 46284 43148 46340 43204
rect 46508 43372 46564 43428
rect 45948 41916 46004 41972
rect 45724 41410 45780 41412
rect 45724 41358 45726 41410
rect 45726 41358 45778 41410
rect 45778 41358 45780 41410
rect 45724 41356 45780 41358
rect 45836 41244 45892 41300
rect 45948 40626 46004 40628
rect 45948 40574 45950 40626
rect 45950 40574 46002 40626
rect 46002 40574 46004 40626
rect 45948 40572 46004 40574
rect 45724 39340 45780 39396
rect 43596 38332 43652 38388
rect 43372 37548 43428 37604
rect 43484 37996 43540 38052
rect 43820 37826 43876 37828
rect 43820 37774 43822 37826
rect 43822 37774 43874 37826
rect 43874 37774 43876 37826
rect 43820 37772 43876 37774
rect 44044 37826 44100 37828
rect 44044 37774 44046 37826
rect 44046 37774 44098 37826
rect 44098 37774 44100 37826
rect 44044 37772 44100 37774
rect 44156 37548 44212 37604
rect 43708 37100 43764 37156
rect 43260 36652 43316 36708
rect 41244 35810 41300 35812
rect 41244 35758 41246 35810
rect 41246 35758 41298 35810
rect 41298 35758 41300 35810
rect 41244 35756 41300 35758
rect 40124 35698 40180 35700
rect 40124 35646 40126 35698
rect 40126 35646 40178 35698
rect 40178 35646 40180 35698
rect 40124 35644 40180 35646
rect 39900 34860 39956 34916
rect 40908 35698 40964 35700
rect 40908 35646 40910 35698
rect 40910 35646 40962 35698
rect 40962 35646 40964 35698
rect 40908 35644 40964 35646
rect 43596 36370 43652 36372
rect 43596 36318 43598 36370
rect 43598 36318 43650 36370
rect 43650 36318 43652 36370
rect 43596 36316 43652 36318
rect 39900 34636 39956 34692
rect 37100 33964 37156 34020
rect 37100 33458 37156 33460
rect 37100 33406 37102 33458
rect 37102 33406 37154 33458
rect 37154 33406 37156 33458
rect 37100 33404 37156 33406
rect 37660 34018 37716 34020
rect 37660 33966 37662 34018
rect 37662 33966 37714 34018
rect 37714 33966 37716 34018
rect 37660 33964 37716 33966
rect 38780 33964 38836 34020
rect 39004 34076 39060 34132
rect 38220 33628 38276 33684
rect 37660 32562 37716 32564
rect 37660 32510 37662 32562
rect 37662 32510 37714 32562
rect 37714 32510 37716 32562
rect 37660 32508 37716 32510
rect 38668 33628 38724 33684
rect 41132 34690 41188 34692
rect 41132 34638 41134 34690
rect 41134 34638 41186 34690
rect 41186 34638 41188 34690
rect 41132 34636 41188 34638
rect 44940 37826 44996 37828
rect 44940 37774 44942 37826
rect 44942 37774 44994 37826
rect 44994 37774 44996 37826
rect 44940 37772 44996 37774
rect 45948 39394 46004 39396
rect 45948 39342 45950 39394
rect 45950 39342 46002 39394
rect 46002 39342 46004 39394
rect 45948 39340 46004 39342
rect 46060 39004 46116 39060
rect 45836 38834 45892 38836
rect 45836 38782 45838 38834
rect 45838 38782 45890 38834
rect 45890 38782 45892 38834
rect 45836 38780 45892 38782
rect 47740 44604 47796 44660
rect 48188 44604 48244 44660
rect 47964 43538 48020 43540
rect 47964 43486 47966 43538
rect 47966 43486 48018 43538
rect 48018 43486 48020 43538
rect 47964 43484 48020 43486
rect 47180 42700 47236 42756
rect 46508 41916 46564 41972
rect 46620 41356 46676 41412
rect 47964 42476 48020 42532
rect 48076 42082 48132 42084
rect 48076 42030 48078 42082
rect 48078 42030 48130 42082
rect 48130 42030 48132 42082
rect 48076 42028 48132 42030
rect 48748 45666 48804 45668
rect 48748 45614 48750 45666
rect 48750 45614 48802 45666
rect 48802 45614 48804 45666
rect 48748 45612 48804 45614
rect 48412 44828 48468 44884
rect 49084 45276 49140 45332
rect 48860 44380 48916 44436
rect 49532 44380 49588 44436
rect 49084 44044 49140 44100
rect 48300 41970 48356 41972
rect 48300 41918 48302 41970
rect 48302 41918 48354 41970
rect 48354 41918 48356 41970
rect 48300 41916 48356 41918
rect 48748 43372 48804 43428
rect 48748 43148 48804 43204
rect 48860 42476 48916 42532
rect 49308 43538 49364 43540
rect 49308 43486 49310 43538
rect 49310 43486 49362 43538
rect 49362 43486 49364 43538
rect 49308 43484 49364 43486
rect 49532 43708 49588 43764
rect 49756 44268 49812 44324
rect 48972 42364 49028 42420
rect 49532 42754 49588 42756
rect 49532 42702 49534 42754
rect 49534 42702 49586 42754
rect 49586 42702 49588 42754
rect 49532 42700 49588 42702
rect 49980 44716 50036 44772
rect 50092 44492 50148 44548
rect 51436 45948 51492 46004
rect 53788 46002 53844 46004
rect 53788 45950 53790 46002
rect 53790 45950 53842 46002
rect 53842 45950 53844 46002
rect 53788 45948 53844 45950
rect 50556 45498 50612 45500
rect 50556 45446 50558 45498
rect 50558 45446 50610 45498
rect 50610 45446 50612 45498
rect 50556 45444 50612 45446
rect 50660 45498 50716 45500
rect 50660 45446 50662 45498
rect 50662 45446 50714 45498
rect 50714 45446 50716 45498
rect 50660 45444 50716 45446
rect 50764 45498 50820 45500
rect 50764 45446 50766 45498
rect 50766 45446 50818 45498
rect 50818 45446 50820 45498
rect 50764 45444 50820 45446
rect 50204 44322 50260 44324
rect 50204 44270 50206 44322
rect 50206 44270 50258 44322
rect 50258 44270 50260 44322
rect 50204 44268 50260 44270
rect 49980 43596 50036 43652
rect 50092 43708 50148 43764
rect 48412 41580 48468 41636
rect 46284 40514 46340 40516
rect 46284 40462 46286 40514
rect 46286 40462 46338 40514
rect 46338 40462 46340 40514
rect 46284 40460 46340 40462
rect 46284 39618 46340 39620
rect 46284 39566 46286 39618
rect 46286 39566 46338 39618
rect 46338 39566 46340 39618
rect 46284 39564 46340 39566
rect 49644 41804 49700 41860
rect 49308 41020 49364 41076
rect 47404 40572 47460 40628
rect 46956 39900 47012 39956
rect 46732 39228 46788 39284
rect 46508 38892 46564 38948
rect 45724 38220 45780 38276
rect 46396 38444 46452 38500
rect 45500 37772 45556 37828
rect 46732 39004 46788 39060
rect 46732 38780 46788 38836
rect 49084 40962 49140 40964
rect 49084 40910 49086 40962
rect 49086 40910 49138 40962
rect 49138 40910 49140 40962
rect 49084 40908 49140 40910
rect 49308 40572 49364 40628
rect 49308 40290 49364 40292
rect 49308 40238 49310 40290
rect 49310 40238 49362 40290
rect 49362 40238 49364 40290
rect 49308 40236 49364 40238
rect 48860 39564 48916 39620
rect 47292 39228 47348 39284
rect 47068 38946 47124 38948
rect 47068 38894 47070 38946
rect 47070 38894 47122 38946
rect 47122 38894 47124 38946
rect 47068 38892 47124 38894
rect 49532 40796 49588 40852
rect 49420 38892 49476 38948
rect 47740 38668 47796 38724
rect 46620 38332 46676 38388
rect 44828 37548 44884 37604
rect 44716 37154 44772 37156
rect 44716 37102 44718 37154
rect 44718 37102 44770 37154
rect 44770 37102 44772 37154
rect 44716 37100 44772 37102
rect 44156 36652 44212 36708
rect 43932 36316 43988 36372
rect 44380 36482 44436 36484
rect 44380 36430 44382 36482
rect 44382 36430 44434 36482
rect 44434 36430 44436 36482
rect 44380 36428 44436 36430
rect 41244 34076 41300 34132
rect 41580 34300 41636 34356
rect 42252 34130 42308 34132
rect 42252 34078 42254 34130
rect 42254 34078 42306 34130
rect 42306 34078 42308 34130
rect 42252 34076 42308 34078
rect 40124 33740 40180 33796
rect 41020 33740 41076 33796
rect 39676 33458 39732 33460
rect 39676 33406 39678 33458
rect 39678 33406 39730 33458
rect 39730 33406 39732 33458
rect 39676 33404 39732 33406
rect 38892 32844 38948 32900
rect 37884 32396 37940 32452
rect 36092 31890 36148 31892
rect 36092 31838 36094 31890
rect 36094 31838 36146 31890
rect 36146 31838 36148 31890
rect 36092 31836 36148 31838
rect 36204 31724 36260 31780
rect 36428 31666 36484 31668
rect 36428 31614 36430 31666
rect 36430 31614 36482 31666
rect 36482 31614 36484 31666
rect 36428 31612 36484 31614
rect 35868 30940 35924 30996
rect 36092 31052 36148 31108
rect 37100 31724 37156 31780
rect 37212 31612 37268 31668
rect 37324 31500 37380 31556
rect 37212 31218 37268 31220
rect 37212 31166 37214 31218
rect 37214 31166 37266 31218
rect 37266 31166 37268 31218
rect 37212 31164 37268 31166
rect 35196 30770 35252 30772
rect 35196 30718 35198 30770
rect 35198 30718 35250 30770
rect 35250 30718 35252 30770
rect 35196 30716 35252 30718
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35308 30098 35364 30100
rect 35308 30046 35310 30098
rect 35310 30046 35362 30098
rect 35362 30046 35364 30098
rect 35308 30044 35364 30046
rect 34748 28588 34804 28644
rect 34524 28530 34580 28532
rect 34524 28478 34526 28530
rect 34526 28478 34578 28530
rect 34578 28478 34580 28530
rect 34524 28476 34580 28478
rect 34300 28418 34356 28420
rect 34300 28366 34302 28418
rect 34302 28366 34354 28418
rect 34354 28366 34356 28418
rect 34300 28364 34356 28366
rect 34188 27970 34244 27972
rect 34188 27918 34190 27970
rect 34190 27918 34242 27970
rect 34242 27918 34244 27970
rect 34188 27916 34244 27918
rect 35756 29932 35812 29988
rect 35868 30716 35924 30772
rect 35196 29708 35252 29764
rect 36204 30210 36260 30212
rect 36204 30158 36206 30210
rect 36206 30158 36258 30210
rect 36258 30158 36260 30210
rect 36204 30156 36260 30158
rect 36204 29932 36260 29988
rect 35980 29708 36036 29764
rect 36204 29596 36260 29652
rect 36988 30210 37044 30212
rect 36988 30158 36990 30210
rect 36990 30158 37042 30210
rect 37042 30158 37044 30210
rect 36988 30156 37044 30158
rect 39676 32844 39732 32900
rect 40236 32844 40292 32900
rect 38556 31778 38612 31780
rect 38556 31726 38558 31778
rect 38558 31726 38610 31778
rect 38610 31726 38612 31778
rect 38556 31724 38612 31726
rect 42812 34300 42868 34356
rect 45612 36764 45668 36820
rect 45052 36428 45108 36484
rect 45724 36482 45780 36484
rect 45724 36430 45726 36482
rect 45726 36430 45778 36482
rect 45778 36430 45780 36482
rect 45724 36428 45780 36430
rect 46732 37266 46788 37268
rect 46732 37214 46734 37266
rect 46734 37214 46786 37266
rect 46786 37214 46788 37266
rect 46732 37212 46788 37214
rect 46396 37042 46452 37044
rect 46396 36990 46398 37042
rect 46398 36990 46450 37042
rect 46450 36990 46452 37042
rect 46396 36988 46452 36990
rect 46284 36482 46340 36484
rect 46284 36430 46286 36482
rect 46286 36430 46338 36482
rect 46338 36430 46340 36482
rect 46284 36428 46340 36430
rect 47404 37938 47460 37940
rect 47404 37886 47406 37938
rect 47406 37886 47458 37938
rect 47458 37886 47460 37938
rect 47404 37884 47460 37886
rect 47180 37212 47236 37268
rect 47292 37324 47348 37380
rect 45276 36370 45332 36372
rect 45276 36318 45278 36370
rect 45278 36318 45330 36370
rect 45330 36318 45332 36370
rect 45276 36316 45332 36318
rect 44044 35308 44100 35364
rect 42588 34242 42644 34244
rect 42588 34190 42590 34242
rect 42590 34190 42642 34242
rect 42642 34190 42644 34242
rect 42588 34188 42644 34190
rect 43148 34130 43204 34132
rect 43148 34078 43150 34130
rect 43150 34078 43202 34130
rect 43202 34078 43204 34130
rect 43148 34076 43204 34078
rect 45836 36258 45892 36260
rect 45836 36206 45838 36258
rect 45838 36206 45890 36258
rect 45890 36206 45892 36258
rect 45836 36204 45892 36206
rect 45612 35698 45668 35700
rect 45612 35646 45614 35698
rect 45614 35646 45666 35698
rect 45666 35646 45668 35698
rect 45612 35644 45668 35646
rect 44940 34860 44996 34916
rect 45836 35308 45892 35364
rect 45836 34860 45892 34916
rect 43932 33852 43988 33908
rect 43036 33740 43092 33796
rect 44380 33516 44436 33572
rect 44268 33234 44324 33236
rect 44268 33182 44270 33234
rect 44270 33182 44322 33234
rect 44322 33182 44324 33234
rect 44268 33180 44324 33182
rect 45836 34300 45892 34356
rect 45052 34130 45108 34132
rect 45052 34078 45054 34130
rect 45054 34078 45106 34130
rect 45106 34078 45108 34130
rect 45052 34076 45108 34078
rect 45052 33180 45108 33236
rect 41580 32620 41636 32676
rect 41468 32562 41524 32564
rect 41468 32510 41470 32562
rect 41470 32510 41522 32562
rect 41522 32510 41524 32562
rect 41468 32508 41524 32510
rect 45500 34242 45556 34244
rect 45500 34190 45502 34242
rect 45502 34190 45554 34242
rect 45554 34190 45556 34242
rect 45500 34188 45556 34190
rect 45276 33516 45332 33572
rect 45388 34076 45444 34132
rect 45724 33852 45780 33908
rect 46732 33852 46788 33908
rect 45164 32732 45220 32788
rect 43260 32674 43316 32676
rect 43260 32622 43262 32674
rect 43262 32622 43314 32674
rect 43314 32622 43316 32674
rect 43260 32620 43316 32622
rect 43596 32620 43652 32676
rect 42924 32562 42980 32564
rect 42924 32510 42926 32562
rect 42926 32510 42978 32562
rect 42978 32510 42980 32562
rect 42924 32508 42980 32510
rect 43148 32562 43204 32564
rect 43148 32510 43150 32562
rect 43150 32510 43202 32562
rect 43202 32510 43204 32562
rect 43148 32508 43204 32510
rect 39228 31890 39284 31892
rect 39228 31838 39230 31890
rect 39230 31838 39282 31890
rect 39282 31838 39284 31890
rect 39228 31836 39284 31838
rect 38108 31500 38164 31556
rect 39004 31612 39060 31668
rect 39676 31666 39732 31668
rect 39676 31614 39678 31666
rect 39678 31614 39730 31666
rect 39730 31614 39732 31666
rect 39676 31612 39732 31614
rect 41356 31836 41412 31892
rect 38108 31218 38164 31220
rect 38108 31166 38110 31218
rect 38110 31166 38162 31218
rect 38162 31166 38164 31218
rect 38108 31164 38164 31166
rect 38668 31164 38724 31220
rect 39900 31276 39956 31332
rect 39788 31218 39844 31220
rect 39788 31166 39790 31218
rect 39790 31166 39842 31218
rect 39842 31166 39844 31218
rect 39788 31164 39844 31166
rect 37884 30380 37940 30436
rect 38668 30492 38724 30548
rect 37100 30044 37156 30100
rect 36764 29932 36820 29988
rect 37324 30098 37380 30100
rect 37324 30046 37326 30098
rect 37326 30046 37378 30098
rect 37378 30046 37380 30098
rect 37324 30044 37380 30046
rect 36876 29314 36932 29316
rect 36876 29262 36878 29314
rect 36878 29262 36930 29314
rect 36930 29262 36932 29314
rect 36876 29260 36932 29262
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 34748 28418 34804 28420
rect 34748 28366 34750 28418
rect 34750 28366 34802 28418
rect 34802 28366 34804 28418
rect 34748 28364 34804 28366
rect 35308 28812 35364 28868
rect 34412 27916 34468 27972
rect 32956 25228 33012 25284
rect 33740 27132 33796 27188
rect 34748 27132 34804 27188
rect 34524 26796 34580 26852
rect 35532 28588 35588 28644
rect 35532 27970 35588 27972
rect 35532 27918 35534 27970
rect 35534 27918 35586 27970
rect 35586 27918 35588 27970
rect 35532 27916 35588 27918
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 35084 26850 35140 26852
rect 35084 26798 35086 26850
rect 35086 26798 35138 26850
rect 35138 26798 35140 26850
rect 35084 26796 35140 26798
rect 33404 25004 33460 25060
rect 32956 23826 33012 23828
rect 32956 23774 32958 23826
rect 32958 23774 33010 23826
rect 33010 23774 33012 23826
rect 32956 23772 33012 23774
rect 32620 23436 32676 23492
rect 32172 23212 32228 23268
rect 32396 23266 32452 23268
rect 32396 23214 32398 23266
rect 32398 23214 32450 23266
rect 32450 23214 32452 23266
rect 32396 23212 32452 23214
rect 30828 22316 30884 22372
rect 30604 21756 30660 21812
rect 30156 21644 30212 21700
rect 28812 18956 28868 19012
rect 28252 18620 28308 18676
rect 27916 18562 27972 18564
rect 27916 18510 27918 18562
rect 27918 18510 27970 18562
rect 27970 18510 27972 18562
rect 27916 18508 27972 18510
rect 28028 18396 28084 18452
rect 28588 18450 28644 18452
rect 28588 18398 28590 18450
rect 28590 18398 28642 18450
rect 28642 18398 28644 18450
rect 28588 18396 28644 18398
rect 27356 15148 27412 15204
rect 22204 13916 22260 13972
rect 22316 13580 22372 13636
rect 23100 13858 23156 13860
rect 23100 13806 23102 13858
rect 23102 13806 23154 13858
rect 23154 13806 23156 13858
rect 23100 13804 23156 13806
rect 23436 13804 23492 13860
rect 23100 13074 23156 13076
rect 23100 13022 23102 13074
rect 23102 13022 23154 13074
rect 23154 13022 23156 13074
rect 23100 13020 23156 13022
rect 23212 12962 23268 12964
rect 23212 12910 23214 12962
rect 23214 12910 23266 12962
rect 23266 12910 23268 12962
rect 23212 12908 23268 12910
rect 23548 13692 23604 13748
rect 23772 12908 23828 12964
rect 22876 11452 22932 11508
rect 19180 10610 19236 10612
rect 19180 10558 19182 10610
rect 19182 10558 19234 10610
rect 19234 10558 19236 10610
rect 19180 10556 19236 10558
rect 18284 9772 18340 9828
rect 17948 9602 18004 9604
rect 17948 9550 17950 9602
rect 17950 9550 18002 9602
rect 18002 9550 18004 9602
rect 17948 9548 18004 9550
rect 18732 9548 18788 9604
rect 18844 9100 18900 9156
rect 15820 8146 15876 8148
rect 15820 8094 15822 8146
rect 15822 8094 15874 8146
rect 15874 8094 15876 8146
rect 15820 8092 15876 8094
rect 15484 7644 15540 7700
rect 16268 7868 16324 7924
rect 16492 8988 16548 9044
rect 17948 9042 18004 9044
rect 17948 8990 17950 9042
rect 17950 8990 18002 9042
rect 18002 8990 18004 9042
rect 17948 8988 18004 8990
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 18172 8370 18228 8372
rect 18172 8318 18174 8370
rect 18174 8318 18226 8370
rect 18226 8318 18228 8370
rect 18172 8316 18228 8318
rect 16828 7868 16884 7924
rect 19964 9100 20020 9156
rect 19404 8316 19460 8372
rect 15708 7362 15764 7364
rect 15708 7310 15710 7362
rect 15710 7310 15762 7362
rect 15762 7310 15764 7362
rect 15708 7308 15764 7310
rect 21532 9660 21588 9716
rect 22092 9660 22148 9716
rect 20972 9548 21028 9604
rect 21196 9154 21252 9156
rect 21196 9102 21198 9154
rect 21198 9102 21250 9154
rect 21250 9102 21252 9154
rect 21196 9100 21252 9102
rect 24220 14530 24276 14532
rect 24220 14478 24222 14530
rect 24222 14478 24274 14530
rect 24274 14478 24276 14530
rect 24220 14476 24276 14478
rect 24780 14306 24836 14308
rect 24780 14254 24782 14306
rect 24782 14254 24834 14306
rect 24834 14254 24836 14306
rect 24780 14252 24836 14254
rect 25340 14252 25396 14308
rect 24668 13692 24724 13748
rect 25116 13746 25172 13748
rect 25116 13694 25118 13746
rect 25118 13694 25170 13746
rect 25170 13694 25172 13746
rect 25116 13692 25172 13694
rect 25676 14476 25732 14532
rect 26012 14476 26068 14532
rect 25900 12738 25956 12740
rect 25900 12686 25902 12738
rect 25902 12686 25954 12738
rect 25954 12686 25956 12738
rect 25900 12684 25956 12686
rect 26908 12850 26964 12852
rect 26908 12798 26910 12850
rect 26910 12798 26962 12850
rect 26962 12798 26964 12850
rect 26908 12796 26964 12798
rect 27580 14530 27636 14532
rect 27580 14478 27582 14530
rect 27582 14478 27634 14530
rect 27634 14478 27636 14530
rect 27580 14476 27636 14478
rect 27132 12684 27188 12740
rect 26908 12124 26964 12180
rect 25116 11282 25172 11284
rect 25116 11230 25118 11282
rect 25118 11230 25170 11282
rect 25170 11230 25172 11282
rect 25116 11228 25172 11230
rect 26572 10780 26628 10836
rect 25788 10556 25844 10612
rect 25564 9938 25620 9940
rect 25564 9886 25566 9938
rect 25566 9886 25618 9938
rect 25618 9886 25620 9938
rect 25564 9884 25620 9886
rect 22764 9772 22820 9828
rect 23772 9826 23828 9828
rect 23772 9774 23774 9826
rect 23774 9774 23826 9826
rect 23826 9774 23828 9826
rect 23772 9772 23828 9774
rect 26460 10610 26516 10612
rect 26460 10558 26462 10610
rect 26462 10558 26514 10610
rect 26514 10558 26516 10610
rect 26460 10556 26516 10558
rect 26348 10498 26404 10500
rect 26348 10446 26350 10498
rect 26350 10446 26402 10498
rect 26402 10446 26404 10498
rect 26348 10444 26404 10446
rect 23212 9714 23268 9716
rect 23212 9662 23214 9714
rect 23214 9662 23266 9714
rect 23266 9662 23268 9714
rect 23212 9660 23268 9662
rect 21980 9154 22036 9156
rect 21980 9102 21982 9154
rect 21982 9102 22034 9154
rect 22034 9102 22036 9154
rect 21980 9100 22036 9102
rect 22092 8988 22148 9044
rect 20188 8428 20244 8484
rect 23436 8988 23492 9044
rect 22092 8428 22148 8484
rect 24668 8482 24724 8484
rect 24668 8430 24670 8482
rect 24670 8430 24722 8482
rect 24722 8430 24724 8482
rect 24668 8428 24724 8430
rect 25004 8370 25060 8372
rect 25004 8318 25006 8370
rect 25006 8318 25058 8370
rect 25058 8318 25060 8370
rect 25004 8316 25060 8318
rect 22876 7980 22932 8036
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 23212 7474 23268 7476
rect 23212 7422 23214 7474
rect 23214 7422 23266 7474
rect 23266 7422 23268 7474
rect 23212 7420 23268 7422
rect 18844 7196 18900 7252
rect 24668 7980 24724 8036
rect 26460 10332 26516 10388
rect 25788 8428 25844 8484
rect 25900 8316 25956 8372
rect 28140 14364 28196 14420
rect 28476 14476 28532 14532
rect 27356 12124 27412 12180
rect 27132 11900 27188 11956
rect 28812 14252 28868 14308
rect 28364 12348 28420 12404
rect 28252 12178 28308 12180
rect 28252 12126 28254 12178
rect 28254 12126 28306 12178
rect 28306 12126 28308 12178
rect 28252 12124 28308 12126
rect 28476 12124 28532 12180
rect 28252 11900 28308 11956
rect 27804 11394 27860 11396
rect 27804 11342 27806 11394
rect 27806 11342 27858 11394
rect 27858 11342 27860 11394
rect 27804 11340 27860 11342
rect 27356 11116 27412 11172
rect 28028 10834 28084 10836
rect 28028 10782 28030 10834
rect 28030 10782 28082 10834
rect 28082 10782 28084 10834
rect 28028 10780 28084 10782
rect 28588 11676 28644 11732
rect 28476 10834 28532 10836
rect 28476 10782 28478 10834
rect 28478 10782 28530 10834
rect 28530 10782 28532 10834
rect 28476 10780 28532 10782
rect 27468 10610 27524 10612
rect 27468 10558 27470 10610
rect 27470 10558 27522 10610
rect 27522 10558 27524 10610
rect 27468 10556 27524 10558
rect 27692 10498 27748 10500
rect 27692 10446 27694 10498
rect 27694 10446 27746 10498
rect 27746 10446 27748 10498
rect 27692 10444 27748 10446
rect 27020 10332 27076 10388
rect 29484 18732 29540 18788
rect 30380 20802 30436 20804
rect 30380 20750 30382 20802
rect 30382 20750 30434 20802
rect 30434 20750 30436 20802
rect 30380 20748 30436 20750
rect 31164 20690 31220 20692
rect 31164 20638 31166 20690
rect 31166 20638 31218 20690
rect 31218 20638 31220 20690
rect 31164 20636 31220 20638
rect 31052 20188 31108 20244
rect 30380 20018 30436 20020
rect 30380 19966 30382 20018
rect 30382 19966 30434 20018
rect 30434 19966 30436 20018
rect 30380 19964 30436 19966
rect 30492 19906 30548 19908
rect 30492 19854 30494 19906
rect 30494 19854 30546 19906
rect 30546 19854 30548 19906
rect 30492 19852 30548 19854
rect 29708 19122 29764 19124
rect 29708 19070 29710 19122
rect 29710 19070 29762 19122
rect 29762 19070 29764 19122
rect 29708 19068 29764 19070
rect 29932 19010 29988 19012
rect 29932 18958 29934 19010
rect 29934 18958 29986 19010
rect 29986 18958 29988 19010
rect 29932 18956 29988 18958
rect 29596 18620 29652 18676
rect 30268 18620 30324 18676
rect 30716 18956 30772 19012
rect 31052 18620 31108 18676
rect 30604 18396 30660 18452
rect 29708 17836 29764 17892
rect 31388 17500 31444 17556
rect 29372 15874 29428 15876
rect 29372 15822 29374 15874
rect 29374 15822 29426 15874
rect 29426 15822 29428 15874
rect 29372 15820 29428 15822
rect 30380 15820 30436 15876
rect 30044 15372 30100 15428
rect 29148 14418 29204 14420
rect 29148 14366 29150 14418
rect 29150 14366 29202 14418
rect 29202 14366 29204 14418
rect 29148 14364 29204 14366
rect 29484 14252 29540 14308
rect 30604 15596 30660 15652
rect 31388 16268 31444 16324
rect 33516 24946 33572 24948
rect 33516 24894 33518 24946
rect 33518 24894 33570 24946
rect 33570 24894 33572 24946
rect 33516 24892 33572 24894
rect 33516 24220 33572 24276
rect 33292 24108 33348 24164
rect 33180 22428 33236 22484
rect 32060 21698 32116 21700
rect 32060 21646 32062 21698
rect 32062 21646 32114 21698
rect 32114 21646 32116 21698
rect 32060 21644 32116 21646
rect 32508 21698 32564 21700
rect 32508 21646 32510 21698
rect 32510 21646 32562 21698
rect 32562 21646 32564 21698
rect 32508 21644 32564 21646
rect 33068 21644 33124 21700
rect 32060 21196 32116 21252
rect 33516 23884 33572 23940
rect 33516 23212 33572 23268
rect 33292 20802 33348 20804
rect 33292 20750 33294 20802
rect 33294 20750 33346 20802
rect 33346 20750 33348 20802
rect 33292 20748 33348 20750
rect 32060 20188 32116 20244
rect 31948 20076 32004 20132
rect 33740 25004 33796 25060
rect 33740 23996 33796 24052
rect 35196 26290 35252 26292
rect 35196 26238 35198 26290
rect 35198 26238 35250 26290
rect 35250 26238 35252 26290
rect 35196 26236 35252 26238
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 34076 25116 34132 25172
rect 33964 24108 34020 24164
rect 34188 25004 34244 25060
rect 36204 29148 36260 29204
rect 35868 28588 35924 28644
rect 35532 24892 35588 24948
rect 34636 24332 34692 24388
rect 34188 24220 34244 24276
rect 34748 24108 34804 24164
rect 34748 23772 34804 23828
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 34972 23996 35028 24052
rect 35644 24050 35700 24052
rect 35644 23998 35646 24050
rect 35646 23998 35698 24050
rect 35698 23998 35700 24050
rect 35644 23996 35700 23998
rect 34636 23100 34692 23156
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 35420 22540 35476 22596
rect 35196 22316 35252 22372
rect 33964 21196 34020 21252
rect 34076 22092 34132 22148
rect 34188 21980 34244 22036
rect 33964 20860 34020 20916
rect 34412 21756 34468 21812
rect 35756 22146 35812 22148
rect 35756 22094 35758 22146
rect 35758 22094 35810 22146
rect 35810 22094 35812 22146
rect 35756 22092 35812 22094
rect 35420 21980 35476 22036
rect 34972 20972 35028 21028
rect 35196 21868 35252 21924
rect 34860 20860 34916 20916
rect 34636 20578 34692 20580
rect 34636 20526 34638 20578
rect 34638 20526 34690 20578
rect 34690 20526 34692 20578
rect 34636 20524 34692 20526
rect 34972 20578 35028 20580
rect 34972 20526 34974 20578
rect 34974 20526 35026 20578
rect 35026 20526 35028 20578
rect 34972 20524 35028 20526
rect 34748 19740 34804 19796
rect 31948 17778 32004 17780
rect 31948 17726 31950 17778
rect 31950 17726 32002 17778
rect 32002 17726 32004 17778
rect 31948 17724 32004 17726
rect 33516 17106 33572 17108
rect 33516 17054 33518 17106
rect 33518 17054 33570 17106
rect 33570 17054 33572 17106
rect 33516 17052 33572 17054
rect 31500 16156 31556 16212
rect 30828 14530 30884 14532
rect 30828 14478 30830 14530
rect 30830 14478 30882 14530
rect 30882 14478 30884 14530
rect 30828 14476 30884 14478
rect 31276 14476 31332 14532
rect 29820 14418 29876 14420
rect 29820 14366 29822 14418
rect 29822 14366 29874 14418
rect 29874 14366 29876 14418
rect 29820 14364 29876 14366
rect 29596 12236 29652 12292
rect 29036 11282 29092 11284
rect 29036 11230 29038 11282
rect 29038 11230 29090 11282
rect 29090 11230 29092 11282
rect 29036 11228 29092 11230
rect 29372 11282 29428 11284
rect 29372 11230 29374 11282
rect 29374 11230 29426 11282
rect 29426 11230 29428 11282
rect 29372 11228 29428 11230
rect 29820 11900 29876 11956
rect 30604 13634 30660 13636
rect 30604 13582 30606 13634
rect 30606 13582 30658 13634
rect 30658 13582 30660 13634
rect 30604 13580 30660 13582
rect 30156 12402 30212 12404
rect 30156 12350 30158 12402
rect 30158 12350 30210 12402
rect 30210 12350 30212 12402
rect 30156 12348 30212 12350
rect 30380 11676 30436 11732
rect 30716 12684 30772 12740
rect 29596 10834 29652 10836
rect 29596 10782 29598 10834
rect 29598 10782 29650 10834
rect 29650 10782 29652 10834
rect 29596 10780 29652 10782
rect 29708 11228 29764 11284
rect 26796 9884 26852 9940
rect 28588 9772 28644 9828
rect 28476 9660 28532 9716
rect 27580 9100 27636 9156
rect 27468 8988 27524 9044
rect 26908 8764 26964 8820
rect 26236 7980 26292 8036
rect 24444 7420 24500 7476
rect 24220 6636 24276 6692
rect 27244 8204 27300 8260
rect 26460 7084 26516 7140
rect 24668 6636 24724 6692
rect 25340 6636 25396 6692
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 26124 6636 26180 6692
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 25676 5906 25732 5908
rect 25676 5854 25678 5906
rect 25678 5854 25730 5906
rect 25730 5854 25732 5906
rect 25676 5852 25732 5854
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 25116 3554 25172 3556
rect 25116 3502 25118 3554
rect 25118 3502 25170 3554
rect 25170 3502 25172 3554
rect 25116 3500 25172 3502
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 26460 6076 26516 6132
rect 27020 7196 27076 7252
rect 27916 8764 27972 8820
rect 28140 8370 28196 8372
rect 28140 8318 28142 8370
rect 28142 8318 28194 8370
rect 28194 8318 28196 8370
rect 28140 8316 28196 8318
rect 28252 8204 28308 8260
rect 27468 7980 27524 8036
rect 28028 8034 28084 8036
rect 28028 7982 28030 8034
rect 28030 7982 28082 8034
rect 28082 7982 28084 8034
rect 28028 7980 28084 7982
rect 27132 6860 27188 6916
rect 26796 6412 26852 6468
rect 27580 7084 27636 7140
rect 26908 6636 26964 6692
rect 26572 6188 26628 6244
rect 27468 6748 27524 6804
rect 27132 6188 27188 6244
rect 26460 5852 26516 5908
rect 27244 6412 27300 6468
rect 27356 6188 27412 6244
rect 27244 5628 27300 5684
rect 26012 3554 26068 3556
rect 26012 3502 26014 3554
rect 26014 3502 26066 3554
rect 26066 3502 26068 3554
rect 26012 3500 26068 3502
rect 28028 6748 28084 6804
rect 27916 6524 27972 6580
rect 28364 6860 28420 6916
rect 28588 9042 28644 9044
rect 28588 8990 28590 9042
rect 28590 8990 28642 9042
rect 28642 8990 28644 9042
rect 28588 8988 28644 8990
rect 29260 9660 29316 9716
rect 29036 8930 29092 8932
rect 29036 8878 29038 8930
rect 29038 8878 29090 8930
rect 29090 8878 29092 8930
rect 29036 8876 29092 8878
rect 28812 8764 28868 8820
rect 29036 7980 29092 8036
rect 29372 6860 29428 6916
rect 28252 6466 28308 6468
rect 28252 6414 28254 6466
rect 28254 6414 28306 6466
rect 28306 6414 28308 6466
rect 28252 6412 28308 6414
rect 30380 10892 30436 10948
rect 29708 9324 29764 9380
rect 29820 9996 29876 10052
rect 31500 15314 31556 15316
rect 31500 15262 31502 15314
rect 31502 15262 31554 15314
rect 31554 15262 31556 15314
rect 31500 15260 31556 15262
rect 31500 14252 31556 14308
rect 31388 12290 31444 12292
rect 31388 12238 31390 12290
rect 31390 12238 31442 12290
rect 31442 12238 31444 12290
rect 31388 12236 31444 12238
rect 30940 11900 30996 11956
rect 30492 9996 30548 10052
rect 31052 9714 31108 9716
rect 31052 9662 31054 9714
rect 31054 9662 31106 9714
rect 31106 9662 31108 9714
rect 31052 9660 31108 9662
rect 30716 9212 30772 9268
rect 29820 7308 29876 7364
rect 29596 6690 29652 6692
rect 29596 6638 29598 6690
rect 29598 6638 29650 6690
rect 29650 6638 29652 6690
rect 29596 6636 29652 6638
rect 29596 6412 29652 6468
rect 28812 4956 28868 5012
rect 28364 3442 28420 3444
rect 28364 3390 28366 3442
rect 28366 3390 28418 3442
rect 28418 3390 28420 3442
rect 28364 3388 28420 3390
rect 29372 5010 29428 5012
rect 29372 4958 29374 5010
rect 29374 4958 29426 5010
rect 29426 4958 29428 5010
rect 29372 4956 29428 4958
rect 29484 4508 29540 4564
rect 29372 3164 29428 3220
rect 31164 8988 31220 9044
rect 30268 8876 30324 8932
rect 30492 8146 30548 8148
rect 30492 8094 30494 8146
rect 30494 8094 30546 8146
rect 30546 8094 30548 8146
rect 30492 8092 30548 8094
rect 30940 8092 30996 8148
rect 30380 8034 30436 8036
rect 30380 7982 30382 8034
rect 30382 7982 30434 8034
rect 30434 7982 30436 8034
rect 30380 7980 30436 7982
rect 30604 7586 30660 7588
rect 30604 7534 30606 7586
rect 30606 7534 30658 7586
rect 30658 7534 30660 7586
rect 30604 7532 30660 7534
rect 30380 7474 30436 7476
rect 30380 7422 30382 7474
rect 30382 7422 30434 7474
rect 30434 7422 30436 7474
rect 30380 7420 30436 7422
rect 31052 5852 31108 5908
rect 33292 16882 33348 16884
rect 33292 16830 33294 16882
rect 33294 16830 33346 16882
rect 33346 16830 33348 16882
rect 33292 16828 33348 16830
rect 33068 16716 33124 16772
rect 32060 16268 32116 16324
rect 32956 16210 33012 16212
rect 32956 16158 32958 16210
rect 32958 16158 33010 16210
rect 33010 16158 33012 16210
rect 32956 16156 33012 16158
rect 32844 15596 32900 15652
rect 33180 16098 33236 16100
rect 33180 16046 33182 16098
rect 33182 16046 33234 16098
rect 33234 16046 33236 16098
rect 33180 16044 33236 16046
rect 32956 15148 33012 15204
rect 33180 15260 33236 15316
rect 33180 14530 33236 14532
rect 33180 14478 33182 14530
rect 33182 14478 33234 14530
rect 33234 14478 33236 14530
rect 33180 14476 33236 14478
rect 33740 18284 33796 18340
rect 34412 17724 34468 17780
rect 34076 17052 34132 17108
rect 34412 16940 34468 16996
rect 34076 16882 34132 16884
rect 34076 16830 34078 16882
rect 34078 16830 34130 16882
rect 34130 16830 34132 16882
rect 34076 16828 34132 16830
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 36092 28588 36148 28644
rect 37100 29538 37156 29540
rect 37100 29486 37102 29538
rect 37102 29486 37154 29538
rect 37154 29486 37156 29538
rect 37100 29484 37156 29486
rect 38892 30492 38948 30548
rect 38780 30380 38836 30436
rect 37660 29932 37716 29988
rect 37884 29986 37940 29988
rect 37884 29934 37886 29986
rect 37886 29934 37938 29986
rect 37938 29934 37940 29986
rect 37884 29932 37940 29934
rect 37884 29484 37940 29540
rect 37212 29260 37268 29316
rect 38444 29596 38500 29652
rect 39004 30156 39060 30212
rect 38668 29260 38724 29316
rect 37548 28700 37604 28756
rect 36988 27916 37044 27972
rect 36204 24444 36260 24500
rect 35980 22652 36036 22708
rect 36092 22092 36148 22148
rect 37436 27804 37492 27860
rect 37100 27132 37156 27188
rect 37660 28642 37716 28644
rect 37660 28590 37662 28642
rect 37662 28590 37714 28642
rect 37714 28590 37716 28642
rect 37660 28588 37716 28590
rect 38108 28642 38164 28644
rect 38108 28590 38110 28642
rect 38110 28590 38162 28642
rect 38162 28590 38164 28642
rect 38108 28588 38164 28590
rect 38220 28364 38276 28420
rect 38668 28418 38724 28420
rect 38668 28366 38670 28418
rect 38670 28366 38722 28418
rect 38722 28366 38724 28418
rect 38668 28364 38724 28366
rect 38668 27970 38724 27972
rect 38668 27918 38670 27970
rect 38670 27918 38722 27970
rect 38722 27918 38724 27970
rect 38668 27916 38724 27918
rect 42364 31890 42420 31892
rect 42364 31838 42366 31890
rect 42366 31838 42418 31890
rect 42418 31838 42420 31890
rect 42364 31836 42420 31838
rect 41916 31164 41972 31220
rect 40460 30716 40516 30772
rect 40124 30156 40180 30212
rect 39116 29596 39172 29652
rect 39228 30044 39284 30100
rect 39340 29708 39396 29764
rect 39004 28700 39060 28756
rect 37996 27858 38052 27860
rect 37996 27806 37998 27858
rect 37998 27806 38050 27858
rect 38050 27806 38052 27858
rect 37996 27804 38052 27806
rect 37772 26850 37828 26852
rect 37772 26798 37774 26850
rect 37774 26798 37826 26850
rect 37826 26798 37828 26850
rect 37772 26796 37828 26798
rect 36428 25618 36484 25620
rect 36428 25566 36430 25618
rect 36430 25566 36482 25618
rect 36482 25566 36484 25618
rect 36428 25564 36484 25566
rect 36764 25564 36820 25620
rect 36988 26236 37044 26292
rect 37212 25564 37268 25620
rect 36876 25116 36932 25172
rect 37548 24498 37604 24500
rect 37548 24446 37550 24498
rect 37550 24446 37602 24498
rect 37602 24446 37604 24498
rect 37548 24444 37604 24446
rect 37436 24332 37492 24388
rect 37324 22988 37380 23044
rect 36988 22482 37044 22484
rect 36988 22430 36990 22482
rect 36990 22430 37042 22482
rect 37042 22430 37044 22482
rect 36988 22428 37044 22430
rect 36316 21868 36372 21924
rect 37212 22370 37268 22372
rect 37212 22318 37214 22370
rect 37214 22318 37266 22370
rect 37266 22318 37268 22370
rect 37212 22316 37268 22318
rect 35980 20914 36036 20916
rect 35980 20862 35982 20914
rect 35982 20862 36034 20914
rect 36034 20862 36036 20914
rect 35980 20860 36036 20862
rect 35420 20802 35476 20804
rect 35420 20750 35422 20802
rect 35422 20750 35474 20802
rect 35474 20750 35476 20802
rect 35420 20748 35476 20750
rect 35644 20076 35700 20132
rect 35196 19740 35252 19796
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 35084 18396 35140 18452
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 36988 20914 37044 20916
rect 36988 20862 36990 20914
rect 36990 20862 37042 20914
rect 37042 20862 37044 20914
rect 36988 20860 37044 20862
rect 36540 20578 36596 20580
rect 36540 20526 36542 20578
rect 36542 20526 36594 20578
rect 36594 20526 36596 20578
rect 36540 20524 36596 20526
rect 36316 20076 36372 20132
rect 35756 19740 35812 19796
rect 38220 27132 38276 27188
rect 38108 26796 38164 26852
rect 38108 25506 38164 25508
rect 38108 25454 38110 25506
rect 38110 25454 38162 25506
rect 38162 25454 38164 25506
rect 38108 25452 38164 25454
rect 39228 27970 39284 27972
rect 39228 27918 39230 27970
rect 39230 27918 39282 27970
rect 39282 27918 39284 27970
rect 39228 27916 39284 27918
rect 39228 27074 39284 27076
rect 39228 27022 39230 27074
rect 39230 27022 39282 27074
rect 39282 27022 39284 27074
rect 39228 27020 39284 27022
rect 38444 26796 38500 26852
rect 38780 26348 38836 26404
rect 39004 26290 39060 26292
rect 39004 26238 39006 26290
rect 39006 26238 39058 26290
rect 39058 26238 39060 26290
rect 39004 26236 39060 26238
rect 39564 28700 39620 28756
rect 39564 28364 39620 28420
rect 39676 27970 39732 27972
rect 39676 27918 39678 27970
rect 39678 27918 39730 27970
rect 39730 27918 39732 27970
rect 39676 27916 39732 27918
rect 39004 26012 39060 26068
rect 39004 25506 39060 25508
rect 39004 25454 39006 25506
rect 39006 25454 39058 25506
rect 39058 25454 39060 25506
rect 39004 25452 39060 25454
rect 38892 25340 38948 25396
rect 40124 25676 40180 25732
rect 40460 30044 40516 30100
rect 41132 30268 41188 30324
rect 42812 31164 42868 31220
rect 43148 31164 43204 31220
rect 43372 31052 43428 31108
rect 41916 30268 41972 30324
rect 41244 30098 41300 30100
rect 41244 30046 41246 30098
rect 41246 30046 41298 30098
rect 41298 30046 41300 30098
rect 41244 30044 41300 30046
rect 42476 30098 42532 30100
rect 42476 30046 42478 30098
rect 42478 30046 42530 30098
rect 42530 30046 42532 30098
rect 42476 30044 42532 30046
rect 40908 29986 40964 29988
rect 40908 29934 40910 29986
rect 40910 29934 40962 29986
rect 40962 29934 40964 29986
rect 40908 29932 40964 29934
rect 40908 29426 40964 29428
rect 40908 29374 40910 29426
rect 40910 29374 40962 29426
rect 40962 29374 40964 29426
rect 40908 29372 40964 29374
rect 43372 30322 43428 30324
rect 43372 30270 43374 30322
rect 43374 30270 43426 30322
rect 43426 30270 43428 30322
rect 43372 30268 43428 30270
rect 42924 29372 42980 29428
rect 45388 32562 45444 32564
rect 45388 32510 45390 32562
rect 45390 32510 45442 32562
rect 45442 32510 45444 32562
rect 45388 32508 45444 32510
rect 43708 31836 43764 31892
rect 44156 31554 44212 31556
rect 44156 31502 44158 31554
rect 44158 31502 44210 31554
rect 44210 31502 44212 31554
rect 44156 31500 44212 31502
rect 44044 30434 44100 30436
rect 44044 30382 44046 30434
rect 44046 30382 44098 30434
rect 44098 30382 44100 30434
rect 44044 30380 44100 30382
rect 43820 30322 43876 30324
rect 43820 30270 43822 30322
rect 43822 30270 43874 30322
rect 43874 30270 43876 30322
rect 43820 30268 43876 30270
rect 43708 30210 43764 30212
rect 43708 30158 43710 30210
rect 43710 30158 43762 30210
rect 43762 30158 43764 30210
rect 43708 30156 43764 30158
rect 43820 29820 43876 29876
rect 44940 31724 44996 31780
rect 45836 31778 45892 31780
rect 45836 31726 45838 31778
rect 45838 31726 45890 31778
rect 45890 31726 45892 31778
rect 45836 31724 45892 31726
rect 45164 31666 45220 31668
rect 45164 31614 45166 31666
rect 45166 31614 45218 31666
rect 45218 31614 45220 31666
rect 45164 31612 45220 31614
rect 44604 31106 44660 31108
rect 44604 31054 44606 31106
rect 44606 31054 44658 31106
rect 44658 31054 44660 31106
rect 44604 31052 44660 31054
rect 45276 31500 45332 31556
rect 44940 30268 44996 30324
rect 44156 29372 44212 29428
rect 41020 28364 41076 28420
rect 42140 28364 42196 28420
rect 40796 27970 40852 27972
rect 40796 27918 40798 27970
rect 40798 27918 40850 27970
rect 40850 27918 40852 27970
rect 40796 27916 40852 27918
rect 40348 26460 40404 26516
rect 43708 28700 43764 28756
rect 43260 28082 43316 28084
rect 43260 28030 43262 28082
rect 43262 28030 43314 28082
rect 43314 28030 43316 28082
rect 43260 28028 43316 28030
rect 42924 27858 42980 27860
rect 42924 27806 42926 27858
rect 42926 27806 42978 27858
rect 42978 27806 42980 27858
rect 42924 27804 42980 27806
rect 41132 26348 41188 26404
rect 41020 26290 41076 26292
rect 41020 26238 41022 26290
rect 41022 26238 41074 26290
rect 41074 26238 41076 26290
rect 41020 26236 41076 26238
rect 39788 25394 39844 25396
rect 39788 25342 39790 25394
rect 39790 25342 39842 25394
rect 39842 25342 39844 25394
rect 39788 25340 39844 25342
rect 38892 24946 38948 24948
rect 38892 24894 38894 24946
rect 38894 24894 38946 24946
rect 38946 24894 38948 24946
rect 38892 24892 38948 24894
rect 39228 24834 39284 24836
rect 39228 24782 39230 24834
rect 39230 24782 39282 24834
rect 39282 24782 39284 24834
rect 39228 24780 39284 24782
rect 37548 23660 37604 23716
rect 38556 23938 38612 23940
rect 38556 23886 38558 23938
rect 38558 23886 38610 23938
rect 38610 23886 38612 23938
rect 38556 23884 38612 23886
rect 37660 23378 37716 23380
rect 37660 23326 37662 23378
rect 37662 23326 37714 23378
rect 37714 23326 37716 23378
rect 37660 23324 37716 23326
rect 38332 23324 38388 23380
rect 37884 22988 37940 23044
rect 38108 23100 38164 23156
rect 38556 23378 38612 23380
rect 38556 23326 38558 23378
rect 38558 23326 38610 23378
rect 38610 23326 38612 23378
rect 38556 23324 38612 23326
rect 37884 22540 37940 22596
rect 38108 22428 38164 22484
rect 38668 22428 38724 22484
rect 38780 23100 38836 23156
rect 37660 22316 37716 22372
rect 37548 22092 37604 22148
rect 38220 22092 38276 22148
rect 38668 21644 38724 21700
rect 38220 20748 38276 20804
rect 37212 19852 37268 19908
rect 37996 20524 38052 20580
rect 36988 19628 37044 19684
rect 36428 19122 36484 19124
rect 36428 19070 36430 19122
rect 36430 19070 36482 19122
rect 36482 19070 36484 19122
rect 36428 19068 36484 19070
rect 35756 18284 35812 18340
rect 36316 17724 36372 17780
rect 38108 19628 38164 19684
rect 37100 19122 37156 19124
rect 37100 19070 37102 19122
rect 37102 19070 37154 19122
rect 37154 19070 37156 19122
rect 37100 19068 37156 19070
rect 37212 18396 37268 18452
rect 37100 17612 37156 17668
rect 34748 17052 34804 17108
rect 35196 17500 35252 17556
rect 34748 16716 34804 16772
rect 35756 16994 35812 16996
rect 35756 16942 35758 16994
rect 35758 16942 35810 16994
rect 35810 16942 35812 16994
rect 35756 16940 35812 16942
rect 35644 16828 35700 16884
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 35756 16716 35812 16772
rect 32172 14418 32228 14420
rect 32172 14366 32174 14418
rect 32174 14366 32226 14418
rect 32226 14366 32228 14418
rect 32172 14364 32228 14366
rect 32284 14252 32340 14308
rect 32284 13692 32340 13748
rect 31948 12684 32004 12740
rect 33516 13020 33572 13076
rect 33068 11900 33124 11956
rect 32508 11340 32564 11396
rect 33404 12012 33460 12068
rect 33292 11788 33348 11844
rect 33180 11506 33236 11508
rect 33180 11454 33182 11506
rect 33182 11454 33234 11506
rect 33234 11454 33236 11506
rect 33180 11452 33236 11454
rect 33628 11452 33684 11508
rect 33404 11228 33460 11284
rect 33628 10780 33684 10836
rect 31836 9996 31892 10052
rect 31836 9772 31892 9828
rect 32284 10556 32340 10612
rect 31388 9100 31444 9156
rect 31612 8876 31668 8932
rect 31836 8428 31892 8484
rect 31948 9100 32004 9156
rect 33628 10610 33684 10612
rect 33628 10558 33630 10610
rect 33630 10558 33682 10610
rect 33682 10558 33684 10610
rect 33628 10556 33684 10558
rect 33516 8428 33572 8484
rect 33292 8316 33348 8372
rect 31836 8092 31892 8148
rect 31724 7308 31780 7364
rect 31388 6636 31444 6692
rect 32284 7532 32340 7588
rect 32172 6524 32228 6580
rect 32508 7308 32564 7364
rect 33068 7980 33124 8036
rect 33068 7084 33124 7140
rect 31500 6076 31556 6132
rect 32284 6188 32340 6244
rect 30940 5794 30996 5796
rect 30940 5742 30942 5794
rect 30942 5742 30994 5794
rect 30994 5742 30996 5794
rect 30940 5740 30996 5742
rect 31500 5906 31556 5908
rect 31500 5854 31502 5906
rect 31502 5854 31554 5906
rect 31554 5854 31556 5906
rect 31500 5852 31556 5854
rect 30604 5234 30660 5236
rect 30604 5182 30606 5234
rect 30606 5182 30658 5234
rect 30658 5182 30660 5234
rect 30604 5180 30660 5182
rect 30940 5122 30996 5124
rect 30940 5070 30942 5122
rect 30942 5070 30994 5122
rect 30994 5070 30996 5122
rect 30940 5068 30996 5070
rect 31388 5628 31444 5684
rect 31388 4562 31444 4564
rect 31388 4510 31390 4562
rect 31390 4510 31442 4562
rect 31442 4510 31444 4562
rect 31388 4508 31444 4510
rect 30268 3388 30324 3444
rect 31612 5740 31668 5796
rect 31948 5740 32004 5796
rect 31724 5292 31780 5348
rect 33068 6466 33124 6468
rect 33068 6414 33070 6466
rect 33070 6414 33122 6466
rect 33122 6414 33124 6466
rect 33068 6412 33124 6414
rect 32844 6076 32900 6132
rect 32732 5292 32788 5348
rect 32956 5404 33012 5460
rect 32620 5122 32676 5124
rect 32620 5070 32622 5122
rect 32622 5070 32674 5122
rect 32674 5070 32676 5122
rect 32620 5068 32676 5070
rect 33628 8204 33684 8260
rect 33628 7980 33684 8036
rect 33628 7362 33684 7364
rect 33628 7310 33630 7362
rect 33630 7310 33682 7362
rect 33682 7310 33684 7362
rect 33628 7308 33684 7310
rect 34076 15484 34132 15540
rect 35420 16098 35476 16100
rect 35420 16046 35422 16098
rect 35422 16046 35474 16098
rect 35474 16046 35476 16098
rect 35420 16044 35476 16046
rect 34972 15596 35028 15652
rect 34972 15260 35028 15316
rect 35084 15484 35140 15540
rect 34412 15036 34468 15092
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 38108 18508 38164 18564
rect 37436 18396 37492 18452
rect 37324 17836 37380 17892
rect 39004 22988 39060 23044
rect 39004 22540 39060 22596
rect 38668 19964 38724 20020
rect 36204 16882 36260 16884
rect 36204 16830 36206 16882
rect 36206 16830 36258 16882
rect 36258 16830 36260 16882
rect 36204 16828 36260 16830
rect 36540 16882 36596 16884
rect 36540 16830 36542 16882
rect 36542 16830 36594 16882
rect 36594 16830 36596 16882
rect 36540 16828 36596 16830
rect 37548 17276 37604 17332
rect 37436 16882 37492 16884
rect 37436 16830 37438 16882
rect 37438 16830 37490 16882
rect 37490 16830 37492 16882
rect 37436 16828 37492 16830
rect 37100 16044 37156 16100
rect 37324 16716 37380 16772
rect 36988 15372 37044 15428
rect 36092 15260 36148 15316
rect 36204 14530 36260 14532
rect 36204 14478 36206 14530
rect 36206 14478 36258 14530
rect 36258 14478 36260 14530
rect 36204 14476 36260 14478
rect 35308 14306 35364 14308
rect 35308 14254 35310 14306
rect 35310 14254 35362 14306
rect 35362 14254 35364 14306
rect 35308 14252 35364 14254
rect 35644 14418 35700 14420
rect 35644 14366 35646 14418
rect 35646 14366 35698 14418
rect 35698 14366 35700 14418
rect 35644 14364 35700 14366
rect 37436 16380 37492 16436
rect 38780 20076 38836 20132
rect 39340 23996 39396 24052
rect 39228 23548 39284 23604
rect 40236 24780 40292 24836
rect 40684 24556 40740 24612
rect 40908 23996 40964 24052
rect 40236 23938 40292 23940
rect 40236 23886 40238 23938
rect 40238 23886 40290 23938
rect 40290 23886 40292 23938
rect 40236 23884 40292 23886
rect 39452 23212 39508 23268
rect 39676 23042 39732 23044
rect 39676 22990 39678 23042
rect 39678 22990 39730 23042
rect 39730 22990 39732 23042
rect 39676 22988 39732 22990
rect 39564 22764 39620 22820
rect 39564 22370 39620 22372
rect 39564 22318 39566 22370
rect 39566 22318 39618 22370
rect 39618 22318 39620 22370
rect 39564 22316 39620 22318
rect 39004 22146 39060 22148
rect 39004 22094 39006 22146
rect 39006 22094 39058 22146
rect 39058 22094 39060 22146
rect 39004 22092 39060 22094
rect 39228 21644 39284 21700
rect 40012 22764 40068 22820
rect 40012 22540 40068 22596
rect 39900 22316 39956 22372
rect 39676 21698 39732 21700
rect 39676 21646 39678 21698
rect 39678 21646 39730 21698
rect 39730 21646 39732 21698
rect 39676 21644 39732 21646
rect 38892 19628 38948 19684
rect 38444 18396 38500 18452
rect 38556 17836 38612 17892
rect 38220 17500 38276 17556
rect 38332 17724 38388 17780
rect 38668 17442 38724 17444
rect 38668 17390 38670 17442
rect 38670 17390 38722 17442
rect 38722 17390 38724 17442
rect 38668 17388 38724 17390
rect 37996 17052 38052 17108
rect 39228 18508 39284 18564
rect 39004 18172 39060 18228
rect 39452 20130 39508 20132
rect 39452 20078 39454 20130
rect 39454 20078 39506 20130
rect 39506 20078 39508 20130
rect 39452 20076 39508 20078
rect 39452 19292 39508 19348
rect 39900 21868 39956 21924
rect 42588 26236 42644 26292
rect 41356 25788 41412 25844
rect 41132 25676 41188 25732
rect 42700 26012 42756 26068
rect 44268 29932 44324 29988
rect 44380 30156 44436 30212
rect 43820 27916 43876 27972
rect 45724 31276 45780 31332
rect 45388 30434 45444 30436
rect 45388 30382 45390 30434
rect 45390 30382 45442 30434
rect 45442 30382 45444 30434
rect 45388 30380 45444 30382
rect 45948 31666 46004 31668
rect 45948 31614 45950 31666
rect 45950 31614 46002 31666
rect 46002 31614 46004 31666
rect 45948 31612 46004 31614
rect 46060 31276 46116 31332
rect 46508 32562 46564 32564
rect 46508 32510 46510 32562
rect 46510 32510 46562 32562
rect 46562 32510 46564 32562
rect 46508 32508 46564 32510
rect 46396 31724 46452 31780
rect 46732 32786 46788 32788
rect 46732 32734 46734 32786
rect 46734 32734 46786 32786
rect 46786 32734 46788 32786
rect 46732 32732 46788 32734
rect 46732 32060 46788 32116
rect 45388 29820 45444 29876
rect 45500 30044 45556 30100
rect 46060 29986 46116 29988
rect 46060 29934 46062 29986
rect 46062 29934 46114 29986
rect 46114 29934 46116 29986
rect 46060 29932 46116 29934
rect 46284 29932 46340 29988
rect 45948 29820 46004 29876
rect 45612 29596 45668 29652
rect 45388 29202 45444 29204
rect 45388 29150 45390 29202
rect 45390 29150 45442 29202
rect 45442 29150 45444 29202
rect 45388 29148 45444 29150
rect 44604 28812 44660 28868
rect 44940 28754 44996 28756
rect 44940 28702 44942 28754
rect 44942 28702 44994 28754
rect 44994 28702 44996 28754
rect 44940 28700 44996 28702
rect 44716 28028 44772 28084
rect 45052 28028 45108 28084
rect 44828 27970 44884 27972
rect 44828 27918 44830 27970
rect 44830 27918 44882 27970
rect 44882 27918 44884 27970
rect 44828 27916 44884 27918
rect 43932 27580 43988 27636
rect 43820 27468 43876 27524
rect 45948 28476 46004 28532
rect 44380 27746 44436 27748
rect 44380 27694 44382 27746
rect 44382 27694 44434 27746
rect 44434 27694 44436 27746
rect 44380 27692 44436 27694
rect 45500 27692 45556 27748
rect 45612 27580 45668 27636
rect 45052 27468 45108 27524
rect 43372 26348 43428 26404
rect 42588 25900 42644 25956
rect 41356 25116 41412 25172
rect 43036 25394 43092 25396
rect 43036 25342 43038 25394
rect 43038 25342 43090 25394
rect 43090 25342 43092 25394
rect 43036 25340 43092 25342
rect 44156 26348 44212 26404
rect 44940 26572 44996 26628
rect 43820 25900 43876 25956
rect 43932 25340 43988 25396
rect 41132 24722 41188 24724
rect 41132 24670 41134 24722
rect 41134 24670 41186 24722
rect 41186 24670 41188 24722
rect 41132 24668 41188 24670
rect 41468 23884 41524 23940
rect 43932 24834 43988 24836
rect 43932 24782 43934 24834
rect 43934 24782 43986 24834
rect 43986 24782 43988 24834
rect 43932 24780 43988 24782
rect 41244 23154 41300 23156
rect 41244 23102 41246 23154
rect 41246 23102 41298 23154
rect 41298 23102 41300 23154
rect 41244 23100 41300 23102
rect 41916 24556 41972 24612
rect 40236 22370 40292 22372
rect 40236 22318 40238 22370
rect 40238 22318 40290 22370
rect 40290 22318 40292 22370
rect 40236 22316 40292 22318
rect 40348 21756 40404 21812
rect 40236 20076 40292 20132
rect 39900 20018 39956 20020
rect 39900 19966 39902 20018
rect 39902 19966 39954 20018
rect 39954 19966 39956 20018
rect 39900 19964 39956 19966
rect 39788 18060 39844 18116
rect 38780 16380 38836 16436
rect 38556 16268 38612 16324
rect 38556 15538 38612 15540
rect 38556 15486 38558 15538
rect 38558 15486 38610 15538
rect 38610 15486 38612 15538
rect 38556 15484 38612 15486
rect 38780 16044 38836 16100
rect 39340 17442 39396 17444
rect 39340 17390 39342 17442
rect 39342 17390 39394 17442
rect 39394 17390 39396 17442
rect 39340 17388 39396 17390
rect 39788 17666 39844 17668
rect 39788 17614 39790 17666
rect 39790 17614 39842 17666
rect 39842 17614 39844 17666
rect 39788 17612 39844 17614
rect 40908 22428 40964 22484
rect 41244 22428 41300 22484
rect 41244 22258 41300 22260
rect 41244 22206 41246 22258
rect 41246 22206 41298 22258
rect 41298 22206 41300 22258
rect 41244 22204 41300 22206
rect 41132 20860 41188 20916
rect 41804 22258 41860 22260
rect 41804 22206 41806 22258
rect 41806 22206 41858 22258
rect 41858 22206 41860 22258
rect 41804 22204 41860 22206
rect 41468 22092 41524 22148
rect 41692 21308 41748 21364
rect 41692 20914 41748 20916
rect 41692 20862 41694 20914
rect 41694 20862 41746 20914
rect 41746 20862 41748 20914
rect 41692 20860 41748 20862
rect 41356 20412 41412 20468
rect 40908 20130 40964 20132
rect 40908 20078 40910 20130
rect 40910 20078 40962 20130
rect 40962 20078 40964 20130
rect 40908 20076 40964 20078
rect 41132 18562 41188 18564
rect 41132 18510 41134 18562
rect 41134 18510 41186 18562
rect 41186 18510 41188 18562
rect 41132 18508 41188 18510
rect 41244 18396 41300 18452
rect 41804 18284 41860 18340
rect 39452 17276 39508 17332
rect 41020 18060 41076 18116
rect 40460 17388 40516 17444
rect 40684 17442 40740 17444
rect 40684 17390 40686 17442
rect 40686 17390 40738 17442
rect 40738 17390 40740 17442
rect 40684 17388 40740 17390
rect 40460 17164 40516 17220
rect 39340 16044 39396 16100
rect 39788 16770 39844 16772
rect 39788 16718 39790 16770
rect 39790 16718 39842 16770
rect 39842 16718 39844 16770
rect 39788 16716 39844 16718
rect 37772 15372 37828 15428
rect 36316 14418 36372 14420
rect 36316 14366 36318 14418
rect 36318 14366 36370 14418
rect 36370 14366 36372 14418
rect 36316 14364 36372 14366
rect 33852 11788 33908 11844
rect 36876 14252 36932 14308
rect 36316 13468 36372 13524
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 37100 13020 37156 13076
rect 35980 12402 36036 12404
rect 35980 12350 35982 12402
rect 35982 12350 36034 12402
rect 36034 12350 36036 12402
rect 35980 12348 36036 12350
rect 35084 12290 35140 12292
rect 35084 12238 35086 12290
rect 35086 12238 35138 12290
rect 35138 12238 35140 12290
rect 35084 12236 35140 12238
rect 33964 12012 34020 12068
rect 33964 11116 34020 11172
rect 34188 11788 34244 11844
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 34524 11564 34580 11620
rect 33964 10780 34020 10836
rect 34972 11452 35028 11508
rect 34860 10780 34916 10836
rect 34524 10722 34580 10724
rect 34524 10670 34526 10722
rect 34526 10670 34578 10722
rect 34578 10670 34580 10722
rect 34524 10668 34580 10670
rect 33964 9548 34020 9604
rect 34412 9602 34468 9604
rect 34412 9550 34414 9602
rect 34414 9550 34466 9602
rect 34466 9550 34468 9602
rect 34412 9548 34468 9550
rect 33852 8316 33908 8372
rect 33964 8540 34020 8596
rect 33740 7084 33796 7140
rect 33292 6188 33348 6244
rect 33180 5516 33236 5572
rect 32732 5010 32788 5012
rect 32732 4958 32734 5010
rect 32734 4958 32786 5010
rect 32786 4958 32788 5010
rect 32732 4956 32788 4958
rect 32060 4562 32116 4564
rect 32060 4510 32062 4562
rect 32062 4510 32114 4562
rect 32114 4510 32116 4562
rect 32060 4508 32116 4510
rect 33068 4844 33124 4900
rect 33180 4620 33236 4676
rect 33740 5852 33796 5908
rect 33404 5628 33460 5684
rect 33628 5628 33684 5684
rect 33516 5404 33572 5460
rect 33516 5234 33572 5236
rect 33516 5182 33518 5234
rect 33518 5182 33570 5234
rect 33570 5182 33572 5234
rect 33516 5180 33572 5182
rect 33628 4844 33684 4900
rect 33628 4060 33684 4116
rect 33516 3554 33572 3556
rect 33516 3502 33518 3554
rect 33518 3502 33570 3554
rect 33570 3502 33572 3554
rect 33516 3500 33572 3502
rect 33292 3276 33348 3332
rect 34412 8204 34468 8260
rect 34748 9436 34804 9492
rect 34636 8540 34692 8596
rect 34076 8146 34132 8148
rect 34076 8094 34078 8146
rect 34078 8094 34130 8146
rect 34130 8094 34132 8146
rect 34076 8092 34132 8094
rect 34188 7420 34244 7476
rect 34300 7980 34356 8036
rect 35420 11564 35476 11620
rect 35644 11618 35700 11620
rect 35644 11566 35646 11618
rect 35646 11566 35698 11618
rect 35698 11566 35700 11618
rect 35644 11564 35700 11566
rect 36428 11564 36484 11620
rect 35868 11228 35924 11284
rect 35644 10556 35700 10612
rect 35084 10332 35140 10388
rect 34972 9714 35028 9716
rect 34972 9662 34974 9714
rect 34974 9662 35026 9714
rect 35026 9662 35028 9714
rect 34972 9660 35028 9662
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35868 10332 35924 10388
rect 35644 9826 35700 9828
rect 35644 9774 35646 9826
rect 35646 9774 35698 9826
rect 35698 9774 35700 9826
rect 35644 9772 35700 9774
rect 36540 10386 36596 10388
rect 36540 10334 36542 10386
rect 36542 10334 36594 10386
rect 36594 10334 36596 10386
rect 36540 10332 36596 10334
rect 36652 10220 36708 10276
rect 37212 12178 37268 12180
rect 37212 12126 37214 12178
rect 37214 12126 37266 12178
rect 37266 12126 37268 12178
rect 37212 12124 37268 12126
rect 35308 9436 35364 9492
rect 35756 9602 35812 9604
rect 35756 9550 35758 9602
rect 35758 9550 35810 9602
rect 35810 9550 35812 9602
rect 35756 9548 35812 9550
rect 36316 9714 36372 9716
rect 36316 9662 36318 9714
rect 36318 9662 36370 9714
rect 36370 9662 36372 9714
rect 36316 9660 36372 9662
rect 36204 9436 36260 9492
rect 36876 9436 36932 9492
rect 35308 9154 35364 9156
rect 35308 9102 35310 9154
rect 35310 9102 35362 9154
rect 35362 9102 35364 9154
rect 35308 9100 35364 9102
rect 34748 8204 34804 8260
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35084 8092 35140 8148
rect 34636 7756 34692 7812
rect 35308 7698 35364 7700
rect 35308 7646 35310 7698
rect 35310 7646 35362 7698
rect 35362 7646 35364 7698
rect 35308 7644 35364 7646
rect 36428 9212 36484 9268
rect 35980 9154 36036 9156
rect 35980 9102 35982 9154
rect 35982 9102 36034 9154
rect 36034 9102 36036 9154
rect 35980 9100 36036 9102
rect 36316 9100 36372 9156
rect 36092 9042 36148 9044
rect 36092 8990 36094 9042
rect 36094 8990 36146 9042
rect 36146 8990 36148 9042
rect 36092 8988 36148 8990
rect 35420 7532 35476 7588
rect 34300 6860 34356 6916
rect 34412 7308 34468 7364
rect 35980 8146 36036 8148
rect 35980 8094 35982 8146
rect 35982 8094 36034 8146
rect 36034 8094 36036 8146
rect 35980 8092 36036 8094
rect 36204 8034 36260 8036
rect 36204 7982 36206 8034
rect 36206 7982 36258 8034
rect 36258 7982 36260 8034
rect 36204 7980 36260 7982
rect 34636 6412 34692 6468
rect 33964 5516 34020 5572
rect 34524 5906 34580 5908
rect 34524 5854 34526 5906
rect 34526 5854 34578 5906
rect 34578 5854 34580 5906
rect 34524 5852 34580 5854
rect 33964 5292 34020 5348
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35868 7644 35924 7700
rect 35756 6802 35812 6804
rect 35756 6750 35758 6802
rect 35758 6750 35810 6802
rect 35810 6750 35812 6802
rect 35756 6748 35812 6750
rect 35420 6578 35476 6580
rect 35420 6526 35422 6578
rect 35422 6526 35474 6578
rect 35474 6526 35476 6578
rect 35420 6524 35476 6526
rect 35644 6466 35700 6468
rect 35644 6414 35646 6466
rect 35646 6414 35698 6466
rect 35698 6414 35700 6466
rect 35644 6412 35700 6414
rect 35196 6188 35252 6244
rect 35532 6300 35588 6356
rect 36652 8204 36708 8260
rect 36652 7644 36708 7700
rect 36764 7586 36820 7588
rect 36764 7534 36766 7586
rect 36766 7534 36818 7586
rect 36818 7534 36820 7586
rect 36764 7532 36820 7534
rect 36540 6690 36596 6692
rect 36540 6638 36542 6690
rect 36542 6638 36594 6690
rect 36594 6638 36596 6690
rect 36540 6636 36596 6638
rect 36428 6524 36484 6580
rect 36204 6300 36260 6356
rect 35644 5852 35700 5908
rect 35196 5628 35252 5684
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 34748 5292 34804 5348
rect 34972 5292 35028 5348
rect 34636 5122 34692 5124
rect 34636 5070 34638 5122
rect 34638 5070 34690 5122
rect 34690 5070 34692 5122
rect 34636 5068 34692 5070
rect 34300 4956 34356 5012
rect 36316 6076 36372 6132
rect 35868 5122 35924 5124
rect 35868 5070 35870 5122
rect 35870 5070 35922 5122
rect 35922 5070 35924 5122
rect 35868 5068 35924 5070
rect 36092 5852 36148 5908
rect 36428 5516 36484 5572
rect 36316 5068 36372 5124
rect 34636 3500 34692 3556
rect 34748 4620 34804 4676
rect 35644 4956 35700 5012
rect 35420 4898 35476 4900
rect 35420 4846 35422 4898
rect 35422 4846 35474 4898
rect 35474 4846 35476 4898
rect 35420 4844 35476 4846
rect 35196 4284 35252 4340
rect 34860 4114 34916 4116
rect 34860 4062 34862 4114
rect 34862 4062 34914 4114
rect 34914 4062 34916 4114
rect 34860 4060 34916 4062
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 35084 3778 35140 3780
rect 35084 3726 35086 3778
rect 35086 3726 35138 3778
rect 35138 3726 35140 3778
rect 35084 3724 35140 3726
rect 34972 3612 35028 3668
rect 34860 3554 34916 3556
rect 34860 3502 34862 3554
rect 34862 3502 34914 3554
rect 34914 3502 34916 3554
rect 34860 3500 34916 3502
rect 33964 3388 34020 3444
rect 34412 3388 34468 3444
rect 35532 3442 35588 3444
rect 35532 3390 35534 3442
rect 35534 3390 35586 3442
rect 35586 3390 35588 3442
rect 35532 3388 35588 3390
rect 37212 7196 37268 7252
rect 36764 5906 36820 5908
rect 36764 5854 36766 5906
rect 36766 5854 36818 5906
rect 36818 5854 36820 5906
rect 36764 5852 36820 5854
rect 36876 5516 36932 5572
rect 36988 6412 37044 6468
rect 37212 6300 37268 6356
rect 37660 14530 37716 14532
rect 37660 14478 37662 14530
rect 37662 14478 37714 14530
rect 37714 14478 37716 14530
rect 37660 14476 37716 14478
rect 38332 14418 38388 14420
rect 38332 14366 38334 14418
rect 38334 14366 38386 14418
rect 38386 14366 38388 14418
rect 38332 14364 38388 14366
rect 39004 15932 39060 15988
rect 39004 14924 39060 14980
rect 39340 15314 39396 15316
rect 39340 15262 39342 15314
rect 39342 15262 39394 15314
rect 39394 15262 39396 15314
rect 39340 15260 39396 15262
rect 39564 15932 39620 15988
rect 40124 16604 40180 16660
rect 39900 16098 39956 16100
rect 39900 16046 39902 16098
rect 39902 16046 39954 16098
rect 39954 16046 39956 16098
rect 39900 16044 39956 16046
rect 37660 13692 37716 13748
rect 37548 11394 37604 11396
rect 37548 11342 37550 11394
rect 37550 11342 37602 11394
rect 37602 11342 37604 11394
rect 37548 11340 37604 11342
rect 37996 13692 38052 13748
rect 38444 13692 38500 13748
rect 38332 12796 38388 12852
rect 38108 12738 38164 12740
rect 38108 12686 38110 12738
rect 38110 12686 38162 12738
rect 38162 12686 38164 12738
rect 38108 12684 38164 12686
rect 38220 12572 38276 12628
rect 38444 11228 38500 11284
rect 38108 10834 38164 10836
rect 38108 10782 38110 10834
rect 38110 10782 38162 10834
rect 38162 10782 38164 10834
rect 38108 10780 38164 10782
rect 38892 12572 38948 12628
rect 39228 13692 39284 13748
rect 39676 14924 39732 14980
rect 40236 16044 40292 16100
rect 39900 15314 39956 15316
rect 39900 15262 39902 15314
rect 39902 15262 39954 15314
rect 39954 15262 39956 15314
rect 39900 15260 39956 15262
rect 40012 15036 40068 15092
rect 39900 14140 39956 14196
rect 39116 12684 39172 12740
rect 38892 11340 38948 11396
rect 38444 10668 38500 10724
rect 38668 11004 38724 11060
rect 38780 10780 38836 10836
rect 37996 10444 38052 10500
rect 38668 10332 38724 10388
rect 37436 6802 37492 6804
rect 37436 6750 37438 6802
rect 37438 6750 37490 6802
rect 37490 6750 37492 6802
rect 37436 6748 37492 6750
rect 37548 6524 37604 6580
rect 37324 6188 37380 6244
rect 37100 6076 37156 6132
rect 38444 9826 38500 9828
rect 38444 9774 38446 9826
rect 38446 9774 38498 9826
rect 38498 9774 38500 9826
rect 38444 9772 38500 9774
rect 38220 9436 38276 9492
rect 39228 11116 39284 11172
rect 39116 11004 39172 11060
rect 39564 11340 39620 11396
rect 40796 16716 40852 16772
rect 40908 16658 40964 16660
rect 40908 16606 40910 16658
rect 40910 16606 40962 16658
rect 40962 16606 40964 16658
rect 40908 16604 40964 16606
rect 40908 16380 40964 16436
rect 42252 23100 42308 23156
rect 42140 22988 42196 23044
rect 42028 20690 42084 20692
rect 42028 20638 42030 20690
rect 42030 20638 42082 20690
rect 42082 20638 42084 20690
rect 42028 20636 42084 20638
rect 42476 22540 42532 22596
rect 43036 22482 43092 22484
rect 43036 22430 43038 22482
rect 43038 22430 43090 22482
rect 43090 22430 43092 22482
rect 43036 22428 43092 22430
rect 42700 22370 42756 22372
rect 42700 22318 42702 22370
rect 42702 22318 42754 22370
rect 42754 22318 42756 22370
rect 42700 22316 42756 22318
rect 45500 27356 45556 27412
rect 46284 28364 46340 28420
rect 46060 28082 46116 28084
rect 46060 28030 46062 28082
rect 46062 28030 46114 28082
rect 46114 28030 46116 28082
rect 46060 28028 46116 28030
rect 47068 36482 47124 36484
rect 47068 36430 47070 36482
rect 47070 36430 47122 36482
rect 47122 36430 47124 36482
rect 47068 36428 47124 36430
rect 47292 36204 47348 36260
rect 47404 35868 47460 35924
rect 47628 35756 47684 35812
rect 47516 35644 47572 35700
rect 48748 38722 48804 38724
rect 48748 38670 48750 38722
rect 48750 38670 48802 38722
rect 48802 38670 48804 38722
rect 48748 38668 48804 38670
rect 48300 38444 48356 38500
rect 48524 37772 48580 37828
rect 49868 40236 49924 40292
rect 50092 41804 50148 41860
rect 50556 43930 50612 43932
rect 50556 43878 50558 43930
rect 50558 43878 50610 43930
rect 50610 43878 50612 43930
rect 50556 43876 50612 43878
rect 50660 43930 50716 43932
rect 50660 43878 50662 43930
rect 50662 43878 50714 43930
rect 50714 43878 50716 43930
rect 50660 43876 50716 43878
rect 50764 43930 50820 43932
rect 50764 43878 50766 43930
rect 50766 43878 50818 43930
rect 50818 43878 50820 43930
rect 50764 43876 50820 43878
rect 50428 43260 50484 43316
rect 51212 45052 51268 45108
rect 51772 45052 51828 45108
rect 51548 44994 51604 44996
rect 51548 44942 51550 44994
rect 51550 44942 51602 44994
rect 51602 44942 51604 44994
rect 51548 44940 51604 44942
rect 52780 45890 52836 45892
rect 52780 45838 52782 45890
rect 52782 45838 52834 45890
rect 52834 45838 52836 45890
rect 52780 45836 52836 45838
rect 54236 45890 54292 45892
rect 54236 45838 54238 45890
rect 54238 45838 54290 45890
rect 54290 45838 54292 45890
rect 54236 45836 54292 45838
rect 53340 45778 53396 45780
rect 53340 45726 53342 45778
rect 53342 45726 53394 45778
rect 53394 45726 53396 45778
rect 53340 45724 53396 45726
rect 52220 45330 52276 45332
rect 52220 45278 52222 45330
rect 52222 45278 52274 45330
rect 52274 45278 52276 45330
rect 52220 45276 52276 45278
rect 52108 45164 52164 45220
rect 51996 45106 52052 45108
rect 51996 45054 51998 45106
rect 51998 45054 52050 45106
rect 52050 45054 52052 45106
rect 51996 45052 52052 45054
rect 52108 44994 52164 44996
rect 52108 44942 52110 44994
rect 52110 44942 52162 44994
rect 52162 44942 52164 44994
rect 52108 44940 52164 44942
rect 51772 44380 51828 44436
rect 50988 44044 51044 44100
rect 51548 43596 51604 43652
rect 51212 43538 51268 43540
rect 51212 43486 51214 43538
rect 51214 43486 51266 43538
rect 51266 43486 51268 43538
rect 51212 43484 51268 43486
rect 51884 43484 51940 43540
rect 51548 43260 51604 43316
rect 50876 43036 50932 43092
rect 51324 43036 51380 43092
rect 50556 42362 50612 42364
rect 50556 42310 50558 42362
rect 50558 42310 50610 42362
rect 50610 42310 50612 42362
rect 50556 42308 50612 42310
rect 50660 42362 50716 42364
rect 50660 42310 50662 42362
rect 50662 42310 50714 42362
rect 50714 42310 50716 42362
rect 50660 42308 50716 42310
rect 50764 42362 50820 42364
rect 50764 42310 50766 42362
rect 50766 42310 50818 42362
rect 50818 42310 50820 42362
rect 50764 42308 50820 42310
rect 50764 41804 50820 41860
rect 51436 41132 51492 41188
rect 50652 41074 50708 41076
rect 50652 41022 50654 41074
rect 50654 41022 50706 41074
rect 50706 41022 50708 41074
rect 50652 41020 50708 41022
rect 50556 40794 50612 40796
rect 50556 40742 50558 40794
rect 50558 40742 50610 40794
rect 50610 40742 50612 40794
rect 50556 40740 50612 40742
rect 50660 40794 50716 40796
rect 50660 40742 50662 40794
rect 50662 40742 50714 40794
rect 50714 40742 50716 40794
rect 50660 40740 50716 40742
rect 50764 40794 50820 40796
rect 50764 40742 50766 40794
rect 50766 40742 50818 40794
rect 50818 40742 50820 40794
rect 50764 40740 50820 40742
rect 50204 40402 50260 40404
rect 50204 40350 50206 40402
rect 50206 40350 50258 40402
rect 50258 40350 50260 40402
rect 50204 40348 50260 40350
rect 51100 40348 51156 40404
rect 49196 37884 49252 37940
rect 48300 37212 48356 37268
rect 49420 37884 49476 37940
rect 48188 35868 48244 35924
rect 47852 35698 47908 35700
rect 47852 35646 47854 35698
rect 47854 35646 47906 35698
rect 47906 35646 47908 35698
rect 47852 35644 47908 35646
rect 48300 35756 48356 35812
rect 48188 35532 48244 35588
rect 47516 34242 47572 34244
rect 47516 34190 47518 34242
rect 47518 34190 47570 34242
rect 47570 34190 47572 34242
rect 47516 34188 47572 34190
rect 47180 33404 47236 33460
rect 47404 33180 47460 33236
rect 47852 34300 47908 34356
rect 48076 34300 48132 34356
rect 48524 36258 48580 36260
rect 48524 36206 48526 36258
rect 48526 36206 48578 36258
rect 48578 36206 48580 36258
rect 48524 36204 48580 36206
rect 49084 36204 49140 36260
rect 49308 35810 49364 35812
rect 49308 35758 49310 35810
rect 49310 35758 49362 35810
rect 49362 35758 49364 35810
rect 49308 35756 49364 35758
rect 48636 35698 48692 35700
rect 48636 35646 48638 35698
rect 48638 35646 48690 35698
rect 48690 35646 48692 35698
rect 48636 35644 48692 35646
rect 48300 34076 48356 34132
rect 48748 34412 48804 34468
rect 48972 34300 49028 34356
rect 49196 34242 49252 34244
rect 49196 34190 49198 34242
rect 49198 34190 49250 34242
rect 49250 34190 49252 34242
rect 49196 34188 49252 34190
rect 49308 34130 49364 34132
rect 49308 34078 49310 34130
rect 49310 34078 49362 34130
rect 49362 34078 49364 34130
rect 49308 34076 49364 34078
rect 48748 33458 48804 33460
rect 48748 33406 48750 33458
rect 48750 33406 48802 33458
rect 48802 33406 48804 33458
rect 48748 33404 48804 33406
rect 48972 33346 49028 33348
rect 48972 33294 48974 33346
rect 48974 33294 49026 33346
rect 49026 33294 49028 33346
rect 48972 33292 49028 33294
rect 48412 33234 48468 33236
rect 48412 33182 48414 33234
rect 48414 33182 48466 33234
rect 48466 33182 48468 33234
rect 48412 33180 48468 33182
rect 48188 33068 48244 33124
rect 47628 32844 47684 32900
rect 46844 31890 46900 31892
rect 46844 31838 46846 31890
rect 46846 31838 46898 31890
rect 46898 31838 46900 31890
rect 46844 31836 46900 31838
rect 47068 31948 47124 32004
rect 46732 28028 46788 28084
rect 47964 31836 48020 31892
rect 47964 31388 48020 31444
rect 47292 31052 47348 31108
rect 49644 38108 49700 38164
rect 50204 38220 50260 38276
rect 51884 42700 51940 42756
rect 51660 41356 51716 41412
rect 51660 40908 51716 40964
rect 51772 40348 51828 40404
rect 51996 40908 52052 40964
rect 51100 39340 51156 39396
rect 50556 39226 50612 39228
rect 50556 39174 50558 39226
rect 50558 39174 50610 39226
rect 50610 39174 50612 39226
rect 50556 39172 50612 39174
rect 50660 39226 50716 39228
rect 50660 39174 50662 39226
rect 50662 39174 50714 39226
rect 50714 39174 50716 39226
rect 50660 39172 50716 39174
rect 50764 39226 50820 39228
rect 50764 39174 50766 39226
rect 50766 39174 50818 39226
rect 50818 39174 50820 39226
rect 50764 39172 50820 39174
rect 51100 38668 51156 38724
rect 51548 38946 51604 38948
rect 51548 38894 51550 38946
rect 51550 38894 51602 38946
rect 51602 38894 51604 38946
rect 51548 38892 51604 38894
rect 50316 38108 50372 38164
rect 51212 38220 51268 38276
rect 50316 37826 50372 37828
rect 50316 37774 50318 37826
rect 50318 37774 50370 37826
rect 50370 37774 50372 37826
rect 50316 37772 50372 37774
rect 50204 37436 50260 37492
rect 49980 35698 50036 35700
rect 49980 35646 49982 35698
rect 49982 35646 50034 35698
rect 50034 35646 50036 35698
rect 49980 35644 50036 35646
rect 49980 35420 50036 35476
rect 49644 34300 49700 34356
rect 49756 34130 49812 34132
rect 49756 34078 49758 34130
rect 49758 34078 49810 34130
rect 49810 34078 49812 34130
rect 49756 34076 49812 34078
rect 49532 33068 49588 33124
rect 48636 31778 48692 31780
rect 48636 31726 48638 31778
rect 48638 31726 48690 31778
rect 48690 31726 48692 31778
rect 48636 31724 48692 31726
rect 49308 31890 49364 31892
rect 49308 31838 49310 31890
rect 49310 31838 49362 31890
rect 49362 31838 49364 31890
rect 49308 31836 49364 31838
rect 48860 31388 48916 31444
rect 48524 31052 48580 31108
rect 48860 31164 48916 31220
rect 48188 30994 48244 30996
rect 48188 30942 48190 30994
rect 48190 30942 48242 30994
rect 48242 30942 48244 30994
rect 48188 30940 48244 30942
rect 47628 30492 47684 30548
rect 47852 30322 47908 30324
rect 47852 30270 47854 30322
rect 47854 30270 47906 30322
rect 47906 30270 47908 30322
rect 47852 30268 47908 30270
rect 48748 30268 48804 30324
rect 47292 29708 47348 29764
rect 47068 27356 47124 27412
rect 46508 27186 46564 27188
rect 46508 27134 46510 27186
rect 46510 27134 46562 27186
rect 46562 27134 46564 27186
rect 46508 27132 46564 27134
rect 47516 27186 47572 27188
rect 47516 27134 47518 27186
rect 47518 27134 47570 27186
rect 47570 27134 47572 27186
rect 47516 27132 47572 27134
rect 45724 27074 45780 27076
rect 45724 27022 45726 27074
rect 45726 27022 45778 27074
rect 45778 27022 45780 27074
rect 45724 27020 45780 27022
rect 49196 31106 49252 31108
rect 49196 31054 49198 31106
rect 49198 31054 49250 31106
rect 49250 31054 49252 31106
rect 49196 31052 49252 31054
rect 49308 30994 49364 30996
rect 49308 30942 49310 30994
rect 49310 30942 49362 30994
rect 49362 30942 49364 30994
rect 49308 30940 49364 30942
rect 49980 33346 50036 33348
rect 49980 33294 49982 33346
rect 49982 33294 50034 33346
rect 50034 33294 50036 33346
rect 49980 33292 50036 33294
rect 50092 33234 50148 33236
rect 50092 33182 50094 33234
rect 50094 33182 50146 33234
rect 50146 33182 50148 33234
rect 50092 33180 50148 33182
rect 50316 37100 50372 37156
rect 50556 37658 50612 37660
rect 50556 37606 50558 37658
rect 50558 37606 50610 37658
rect 50610 37606 50612 37658
rect 50556 37604 50612 37606
rect 50660 37658 50716 37660
rect 50660 37606 50662 37658
rect 50662 37606 50714 37658
rect 50714 37606 50716 37658
rect 50660 37604 50716 37606
rect 50764 37658 50820 37660
rect 50764 37606 50766 37658
rect 50766 37606 50818 37658
rect 50818 37606 50820 37658
rect 50764 37604 50820 37606
rect 50652 37266 50708 37268
rect 50652 37214 50654 37266
rect 50654 37214 50706 37266
rect 50706 37214 50708 37266
rect 50652 37212 50708 37214
rect 50316 36092 50372 36148
rect 53228 45218 53284 45220
rect 53228 45166 53230 45218
rect 53230 45166 53282 45218
rect 53282 45166 53284 45218
rect 53228 45164 53284 45166
rect 52780 44828 52836 44884
rect 52892 44716 52948 44772
rect 52668 44492 52724 44548
rect 53564 43596 53620 43652
rect 52556 43372 52612 43428
rect 52892 42866 52948 42868
rect 52892 42814 52894 42866
rect 52894 42814 52946 42866
rect 52946 42814 52948 42866
rect 52892 42812 52948 42814
rect 52444 42700 52500 42756
rect 53900 42812 53956 42868
rect 54348 42754 54404 42756
rect 54348 42702 54350 42754
rect 54350 42702 54402 42754
rect 54402 42702 54404 42754
rect 54348 42700 54404 42702
rect 53452 41916 53508 41972
rect 53004 41410 53060 41412
rect 53004 41358 53006 41410
rect 53006 41358 53058 41410
rect 53058 41358 53060 41410
rect 53004 41356 53060 41358
rect 53788 41970 53844 41972
rect 53788 41918 53790 41970
rect 53790 41918 53842 41970
rect 53842 41918 53844 41970
rect 53788 41916 53844 41918
rect 54236 41804 54292 41860
rect 53564 41356 53620 41412
rect 52668 41186 52724 41188
rect 52668 41134 52670 41186
rect 52670 41134 52722 41186
rect 52722 41134 52724 41186
rect 52668 41132 52724 41134
rect 52108 39004 52164 39060
rect 51436 38722 51492 38724
rect 51436 38670 51438 38722
rect 51438 38670 51490 38722
rect 51490 38670 51492 38722
rect 51436 38668 51492 38670
rect 52892 40962 52948 40964
rect 52892 40910 52894 40962
rect 52894 40910 52946 40962
rect 52946 40910 52948 40962
rect 52892 40908 52948 40910
rect 52892 40402 52948 40404
rect 52892 40350 52894 40402
rect 52894 40350 52946 40402
rect 52946 40350 52948 40402
rect 52892 40348 52948 40350
rect 54684 41804 54740 41860
rect 51884 38668 51940 38724
rect 53788 38332 53844 38388
rect 50556 36090 50612 36092
rect 50556 36038 50558 36090
rect 50558 36038 50610 36090
rect 50610 36038 50612 36090
rect 50556 36036 50612 36038
rect 50660 36090 50716 36092
rect 50660 36038 50662 36090
rect 50662 36038 50714 36090
rect 50714 36038 50716 36090
rect 50660 36036 50716 36038
rect 50764 36090 50820 36092
rect 50764 36038 50766 36090
rect 50766 36038 50818 36090
rect 50818 36038 50820 36090
rect 50764 36036 50820 36038
rect 54460 39900 54516 39956
rect 54460 39340 54516 39396
rect 54236 38780 54292 38836
rect 54684 38332 54740 38388
rect 55468 39394 55524 39396
rect 55468 39342 55470 39394
rect 55470 39342 55522 39394
rect 55522 39342 55524 39394
rect 55468 39340 55524 39342
rect 55132 38834 55188 38836
rect 55132 38782 55134 38834
rect 55134 38782 55186 38834
rect 55186 38782 55188 38834
rect 55132 38780 55188 38782
rect 55804 38610 55860 38612
rect 55804 38558 55806 38610
rect 55806 38558 55858 38610
rect 55858 38558 55860 38610
rect 55804 38556 55860 38558
rect 55132 38220 55188 38276
rect 51772 36988 51828 37044
rect 51884 36764 51940 36820
rect 50988 35922 51044 35924
rect 50988 35870 50990 35922
rect 50990 35870 51042 35922
rect 51042 35870 51044 35922
rect 50988 35868 51044 35870
rect 50652 35698 50708 35700
rect 50652 35646 50654 35698
rect 50654 35646 50706 35698
rect 50706 35646 50708 35698
rect 50652 35644 50708 35646
rect 51996 35756 52052 35812
rect 51212 35532 51268 35588
rect 52444 36988 52500 37044
rect 53004 36764 53060 36820
rect 53228 36988 53284 37044
rect 52220 35868 52276 35924
rect 54460 37436 54516 37492
rect 54348 37100 54404 37156
rect 54572 37324 54628 37380
rect 56028 38220 56084 38276
rect 57036 38556 57092 38612
rect 54572 36988 54628 37044
rect 54908 36988 54964 37044
rect 53788 35644 53844 35700
rect 54236 35644 54292 35700
rect 51548 34748 51604 34804
rect 50556 34522 50612 34524
rect 50556 34470 50558 34522
rect 50558 34470 50610 34522
rect 50610 34470 50612 34522
rect 50556 34468 50612 34470
rect 50660 34522 50716 34524
rect 50660 34470 50662 34522
rect 50662 34470 50714 34522
rect 50714 34470 50716 34522
rect 50660 34468 50716 34470
rect 50764 34522 50820 34524
rect 50764 34470 50766 34522
rect 50766 34470 50818 34522
rect 50818 34470 50820 34522
rect 50764 34468 50820 34470
rect 50316 34188 50372 34244
rect 50652 34130 50708 34132
rect 50652 34078 50654 34130
rect 50654 34078 50706 34130
rect 50706 34078 50708 34130
rect 50652 34076 50708 34078
rect 50316 33458 50372 33460
rect 50316 33406 50318 33458
rect 50318 33406 50370 33458
rect 50370 33406 50372 33458
rect 50316 33404 50372 33406
rect 51660 34188 51716 34244
rect 51660 33292 51716 33348
rect 52780 35308 52836 35364
rect 52556 34636 52612 34692
rect 50556 32954 50612 32956
rect 50556 32902 50558 32954
rect 50558 32902 50610 32954
rect 50610 32902 50612 32954
rect 50556 32900 50612 32902
rect 50660 32954 50716 32956
rect 50660 32902 50662 32954
rect 50662 32902 50714 32954
rect 50714 32902 50716 32954
rect 50660 32900 50716 32902
rect 50764 32954 50820 32956
rect 50764 32902 50766 32954
rect 50766 32902 50818 32954
rect 50818 32902 50820 32954
rect 50764 32900 50820 32902
rect 50204 32060 50260 32116
rect 50988 32562 51044 32564
rect 50988 32510 50990 32562
rect 50990 32510 51042 32562
rect 51042 32510 51044 32562
rect 50988 32508 51044 32510
rect 51996 33346 52052 33348
rect 51996 33294 51998 33346
rect 51998 33294 52050 33346
rect 52050 33294 52052 33346
rect 51996 33292 52052 33294
rect 51884 33068 51940 33124
rect 51884 32562 51940 32564
rect 51884 32510 51886 32562
rect 51886 32510 51938 32562
rect 51938 32510 51940 32562
rect 51884 32508 51940 32510
rect 50764 31778 50820 31780
rect 50764 31726 50766 31778
rect 50766 31726 50818 31778
rect 50818 31726 50820 31778
rect 50764 31724 50820 31726
rect 50556 31386 50612 31388
rect 50556 31334 50558 31386
rect 50558 31334 50610 31386
rect 50610 31334 50612 31386
rect 50556 31332 50612 31334
rect 50660 31386 50716 31388
rect 50660 31334 50662 31386
rect 50662 31334 50714 31386
rect 50714 31334 50716 31386
rect 50660 31332 50716 31334
rect 50764 31386 50820 31388
rect 50764 31334 50766 31386
rect 50766 31334 50818 31386
rect 50818 31334 50820 31386
rect 50764 31332 50820 31334
rect 50092 30940 50148 30996
rect 50092 30770 50148 30772
rect 50092 30718 50094 30770
rect 50094 30718 50146 30770
rect 50146 30718 50148 30770
rect 50092 30716 50148 30718
rect 52444 31106 52500 31108
rect 52444 31054 52446 31106
rect 52446 31054 52498 31106
rect 52498 31054 52500 31106
rect 52444 31052 52500 31054
rect 51100 30882 51156 30884
rect 51100 30830 51102 30882
rect 51102 30830 51154 30882
rect 51154 30830 51156 30882
rect 51100 30828 51156 30830
rect 50540 30716 50596 30772
rect 51324 30716 51380 30772
rect 52332 30716 52388 30772
rect 50556 29818 50612 29820
rect 50556 29766 50558 29818
rect 50558 29766 50610 29818
rect 50610 29766 50612 29818
rect 50556 29764 50612 29766
rect 50660 29818 50716 29820
rect 50660 29766 50662 29818
rect 50662 29766 50714 29818
rect 50714 29766 50716 29818
rect 50660 29764 50716 29766
rect 50764 29818 50820 29820
rect 50764 29766 50766 29818
rect 50766 29766 50818 29818
rect 50818 29766 50820 29818
rect 50764 29764 50820 29766
rect 52108 29484 52164 29540
rect 53004 34802 53060 34804
rect 53004 34750 53006 34802
rect 53006 34750 53058 34802
rect 53058 34750 53060 34802
rect 53004 34748 53060 34750
rect 52668 33234 52724 33236
rect 52668 33182 52670 33234
rect 52670 33182 52722 33234
rect 52722 33182 52724 33234
rect 52668 33180 52724 33182
rect 52892 33292 52948 33348
rect 53004 33122 53060 33124
rect 53004 33070 53006 33122
rect 53006 33070 53058 33122
rect 53058 33070 53060 33122
rect 53004 33068 53060 33070
rect 53788 34802 53844 34804
rect 53788 34750 53790 34802
rect 53790 34750 53842 34802
rect 53842 34750 53844 34802
rect 53788 34748 53844 34750
rect 54796 33906 54852 33908
rect 54796 33854 54798 33906
rect 54798 33854 54850 33906
rect 54850 33854 54852 33906
rect 54796 33852 54852 33854
rect 53340 31666 53396 31668
rect 53340 31614 53342 31666
rect 53342 31614 53394 31666
rect 53394 31614 53396 31666
rect 53340 31612 53396 31614
rect 52556 28700 52612 28756
rect 53676 31500 53732 31556
rect 54796 31724 54852 31780
rect 52668 31052 52724 31108
rect 52108 28476 52164 28532
rect 50556 28250 50612 28252
rect 50556 28198 50558 28250
rect 50558 28198 50610 28250
rect 50610 28198 50612 28250
rect 50556 28196 50612 28198
rect 50660 28250 50716 28252
rect 50660 28198 50662 28250
rect 50662 28198 50714 28250
rect 50714 28198 50716 28250
rect 50660 28196 50716 28198
rect 50764 28250 50820 28252
rect 50764 28198 50766 28250
rect 50766 28198 50818 28250
rect 50818 28198 50820 28250
rect 50764 28196 50820 28198
rect 49644 27580 49700 27636
rect 44492 25228 44548 25284
rect 44940 25116 44996 25172
rect 45388 25340 45444 25396
rect 45836 25394 45892 25396
rect 45836 25342 45838 25394
rect 45838 25342 45890 25394
rect 45890 25342 45892 25394
rect 45836 25340 45892 25342
rect 46060 25116 46116 25172
rect 46172 25340 46228 25396
rect 45164 24668 45220 24724
rect 45612 23938 45668 23940
rect 45612 23886 45614 23938
rect 45614 23886 45666 23938
rect 45666 23886 45668 23938
rect 45612 23884 45668 23886
rect 44604 23154 44660 23156
rect 44604 23102 44606 23154
rect 44606 23102 44658 23154
rect 44658 23102 44660 23154
rect 44604 23100 44660 23102
rect 45724 23100 45780 23156
rect 44156 22540 44212 22596
rect 45164 22316 45220 22372
rect 42588 22204 42644 22260
rect 44156 22204 44212 22260
rect 42588 21868 42644 21924
rect 42476 19852 42532 19908
rect 42252 19292 42308 19348
rect 42140 18450 42196 18452
rect 42140 18398 42142 18450
rect 42142 18398 42194 18450
rect 42194 18398 42196 18450
rect 42140 18396 42196 18398
rect 41468 17500 41524 17556
rect 41356 17276 41412 17332
rect 41132 16268 41188 16324
rect 41804 17106 41860 17108
rect 41804 17054 41806 17106
rect 41806 17054 41858 17106
rect 41858 17054 41860 17106
rect 41804 17052 41860 17054
rect 41580 16882 41636 16884
rect 41580 16830 41582 16882
rect 41582 16830 41634 16882
rect 41634 16830 41636 16882
rect 41580 16828 41636 16830
rect 41692 16770 41748 16772
rect 41692 16718 41694 16770
rect 41694 16718 41746 16770
rect 41746 16718 41748 16770
rect 41692 16716 41748 16718
rect 41804 16044 41860 16100
rect 41244 15874 41300 15876
rect 41244 15822 41246 15874
rect 41246 15822 41298 15874
rect 41298 15822 41300 15874
rect 41244 15820 41300 15822
rect 42140 16828 42196 16884
rect 42364 18284 42420 18340
rect 42588 16210 42644 16212
rect 42588 16158 42590 16210
rect 42590 16158 42642 16210
rect 42642 16158 42644 16210
rect 42588 16156 42644 16158
rect 42028 15484 42084 15540
rect 42476 16098 42532 16100
rect 42476 16046 42478 16098
rect 42478 16046 42530 16098
rect 42530 16046 42532 16098
rect 42476 16044 42532 16046
rect 43596 21868 43652 21924
rect 43820 21532 43876 21588
rect 43036 21308 43092 21364
rect 43148 20636 43204 20692
rect 42924 19906 42980 19908
rect 42924 19854 42926 19906
rect 42926 19854 42978 19906
rect 42978 19854 42980 19906
rect 42924 19852 42980 19854
rect 42812 19346 42868 19348
rect 42812 19294 42814 19346
rect 42814 19294 42866 19346
rect 42866 19294 42868 19346
rect 42812 19292 42868 19294
rect 45500 22258 45556 22260
rect 45500 22206 45502 22258
rect 45502 22206 45554 22258
rect 45554 22206 45556 22258
rect 45500 22204 45556 22206
rect 44268 21868 44324 21924
rect 44828 21868 44884 21924
rect 48188 26236 48244 26292
rect 46284 25228 46340 25284
rect 46508 25116 46564 25172
rect 46508 24892 46564 24948
rect 47852 24946 47908 24948
rect 47852 24894 47854 24946
rect 47854 24894 47906 24946
rect 47906 24894 47908 24946
rect 47852 24892 47908 24894
rect 47516 24834 47572 24836
rect 47516 24782 47518 24834
rect 47518 24782 47570 24834
rect 47570 24782 47572 24834
rect 47516 24780 47572 24782
rect 50556 26682 50612 26684
rect 50556 26630 50558 26682
rect 50558 26630 50610 26682
rect 50610 26630 50612 26682
rect 50556 26628 50612 26630
rect 50660 26682 50716 26684
rect 50660 26630 50662 26682
rect 50662 26630 50714 26682
rect 50714 26630 50716 26682
rect 50660 26628 50716 26630
rect 50764 26682 50820 26684
rect 50764 26630 50766 26682
rect 50766 26630 50818 26682
rect 50818 26630 50820 26682
rect 50764 26628 50820 26630
rect 49084 26514 49140 26516
rect 49084 26462 49086 26514
rect 49086 26462 49138 26514
rect 49138 26462 49140 26514
rect 49084 26460 49140 26462
rect 48860 26290 48916 26292
rect 48860 26238 48862 26290
rect 48862 26238 48914 26290
rect 48914 26238 48916 26290
rect 48860 26236 48916 26238
rect 52108 26236 52164 26292
rect 50556 25114 50612 25116
rect 50556 25062 50558 25114
rect 50558 25062 50610 25114
rect 50610 25062 50612 25114
rect 50556 25060 50612 25062
rect 50660 25114 50716 25116
rect 50660 25062 50662 25114
rect 50662 25062 50714 25114
rect 50714 25062 50716 25114
rect 50660 25060 50716 25062
rect 50764 25114 50820 25116
rect 50764 25062 50766 25114
rect 50766 25062 50818 25114
rect 50818 25062 50820 25114
rect 50764 25060 50820 25062
rect 48636 24780 48692 24836
rect 46956 24722 47012 24724
rect 46956 24670 46958 24722
rect 46958 24670 47010 24722
rect 47010 24670 47012 24722
rect 46956 24668 47012 24670
rect 46396 23826 46452 23828
rect 46396 23774 46398 23826
rect 46398 23774 46450 23826
rect 46450 23774 46452 23826
rect 46396 23772 46452 23774
rect 46620 23826 46676 23828
rect 46620 23774 46622 23826
rect 46622 23774 46674 23826
rect 46674 23774 46676 23826
rect 46620 23772 46676 23774
rect 46172 23100 46228 23156
rect 46284 22988 46340 23044
rect 46396 22370 46452 22372
rect 46396 22318 46398 22370
rect 46398 22318 46450 22370
rect 46450 22318 46452 22370
rect 46396 22316 46452 22318
rect 43596 19292 43652 19348
rect 44268 19346 44324 19348
rect 44268 19294 44270 19346
rect 44270 19294 44322 19346
rect 44322 19294 44324 19346
rect 44268 19292 44324 19294
rect 44828 19292 44884 19348
rect 43820 18508 43876 18564
rect 44940 18450 44996 18452
rect 44940 18398 44942 18450
rect 44942 18398 44994 18450
rect 44994 18398 44996 18450
rect 44940 18396 44996 18398
rect 49756 23772 49812 23828
rect 47516 23042 47572 23044
rect 47516 22990 47518 23042
rect 47518 22990 47570 23042
rect 47570 22990 47572 23042
rect 47516 22988 47572 22990
rect 47964 23154 48020 23156
rect 47964 23102 47966 23154
rect 47966 23102 48018 23154
rect 48018 23102 48020 23154
rect 47964 23100 48020 23102
rect 50556 23546 50612 23548
rect 50556 23494 50558 23546
rect 50558 23494 50610 23546
rect 50610 23494 50612 23546
rect 50556 23492 50612 23494
rect 50660 23546 50716 23548
rect 50660 23494 50662 23546
rect 50662 23494 50714 23546
rect 50714 23494 50716 23546
rect 50660 23492 50716 23494
rect 50764 23546 50820 23548
rect 50764 23494 50766 23546
rect 50766 23494 50818 23546
rect 50818 23494 50820 23546
rect 50764 23492 50820 23494
rect 49756 22482 49812 22484
rect 49756 22430 49758 22482
rect 49758 22430 49810 22482
rect 49810 22430 49812 22482
rect 49756 22428 49812 22430
rect 46956 22316 47012 22372
rect 52892 30828 52948 30884
rect 54236 31666 54292 31668
rect 54236 31614 54238 31666
rect 54238 31614 54290 31666
rect 54290 31614 54292 31666
rect 54236 31612 54292 31614
rect 53564 30044 53620 30100
rect 54012 30156 54068 30212
rect 54012 29932 54068 29988
rect 55020 36876 55076 36932
rect 55020 35644 55076 35700
rect 55804 37324 55860 37380
rect 55356 37100 55412 37156
rect 56588 37378 56644 37380
rect 56588 37326 56590 37378
rect 56590 37326 56642 37378
rect 56642 37326 56644 37378
rect 56588 37324 56644 37326
rect 56924 37826 56980 37828
rect 56924 37774 56926 37826
rect 56926 37774 56978 37826
rect 56978 37774 56980 37826
rect 56924 37772 56980 37774
rect 57820 37938 57876 37940
rect 57820 37886 57822 37938
rect 57822 37886 57874 37938
rect 57874 37886 57876 37938
rect 57820 37884 57876 37886
rect 57484 37660 57540 37716
rect 58044 37772 58100 37828
rect 57148 37436 57204 37492
rect 57820 37548 57876 37604
rect 55244 34860 55300 34916
rect 55692 34860 55748 34916
rect 55356 34076 55412 34132
rect 55692 34130 55748 34132
rect 55692 34078 55694 34130
rect 55694 34078 55746 34130
rect 55746 34078 55748 34130
rect 55692 34076 55748 34078
rect 55468 33906 55524 33908
rect 55468 33854 55470 33906
rect 55470 33854 55522 33906
rect 55522 33854 55524 33906
rect 55468 33852 55524 33854
rect 55132 31778 55188 31780
rect 55132 31726 55134 31778
rect 55134 31726 55186 31778
rect 55186 31726 55188 31778
rect 55132 31724 55188 31726
rect 55020 31554 55076 31556
rect 55020 31502 55022 31554
rect 55022 31502 55074 31554
rect 55074 31502 55076 31554
rect 55020 31500 55076 31502
rect 56252 36204 56308 36260
rect 55804 31388 55860 31444
rect 55916 34188 55972 34244
rect 55580 30210 55636 30212
rect 55580 30158 55582 30210
rect 55582 30158 55634 30210
rect 55634 30158 55636 30210
rect 55580 30156 55636 30158
rect 55916 29596 55972 29652
rect 55244 28642 55300 28644
rect 55244 28590 55246 28642
rect 55246 28590 55298 28642
rect 55298 28590 55300 28642
rect 55244 28588 55300 28590
rect 55580 28642 55636 28644
rect 55580 28590 55582 28642
rect 55582 28590 55634 28642
rect 55634 28590 55636 28642
rect 55580 28588 55636 28590
rect 54908 27804 54964 27860
rect 56588 35756 56644 35812
rect 58044 36988 58100 37044
rect 57820 36258 57876 36260
rect 57820 36206 57822 36258
rect 57822 36206 57874 36258
rect 57874 36206 57876 36258
rect 57820 36204 57876 36206
rect 57820 35810 57876 35812
rect 57820 35758 57822 35810
rect 57822 35758 57874 35810
rect 57874 35758 57876 35810
rect 57820 35756 57876 35758
rect 57148 35698 57204 35700
rect 57148 35646 57150 35698
rect 57150 35646 57202 35698
rect 57202 35646 57204 35698
rect 57148 35644 57204 35646
rect 58380 36316 58436 36372
rect 58268 35644 58324 35700
rect 58156 34972 58212 35028
rect 57820 34690 57876 34692
rect 57820 34638 57822 34690
rect 57822 34638 57874 34690
rect 57874 34638 57876 34690
rect 57820 34636 57876 34638
rect 57596 34300 57652 34356
rect 58156 34300 58212 34356
rect 57820 34242 57876 34244
rect 57820 34190 57822 34242
rect 57822 34190 57874 34242
rect 57874 34190 57876 34242
rect 57820 34188 57876 34190
rect 56700 33852 56756 33908
rect 58156 33628 58212 33684
rect 57596 32956 57652 33012
rect 57148 32284 57204 32340
rect 58156 32956 58212 33012
rect 57820 32674 57876 32676
rect 57820 32622 57822 32674
rect 57822 32622 57874 32674
rect 57874 32622 57876 32674
rect 57820 32620 57876 32622
rect 58156 32284 58212 32340
rect 57708 31948 57764 32004
rect 56924 31666 56980 31668
rect 56924 31614 56926 31666
rect 56926 31614 56978 31666
rect 56978 31614 56980 31666
rect 56924 31612 56980 31614
rect 57484 31666 57540 31668
rect 57484 31614 57486 31666
rect 57486 31614 57538 31666
rect 57538 31614 57540 31666
rect 57484 31612 57540 31614
rect 57820 31554 57876 31556
rect 57820 31502 57822 31554
rect 57822 31502 57874 31554
rect 57874 31502 57876 31554
rect 57820 31500 57876 31502
rect 57820 31106 57876 31108
rect 57820 31054 57822 31106
rect 57822 31054 57874 31106
rect 57874 31054 57876 31106
rect 57820 31052 57876 31054
rect 58380 30940 58436 30996
rect 57148 30268 57204 30324
rect 58156 30268 58212 30324
rect 57596 29650 57652 29652
rect 57596 29598 57598 29650
rect 57598 29598 57650 29650
rect 57650 29598 57652 29650
rect 57596 29596 57652 29598
rect 58156 29596 58212 29652
rect 57820 29538 57876 29540
rect 57820 29486 57822 29538
rect 57822 29486 57874 29538
rect 57874 29486 57876 29538
rect 57820 29484 57876 29486
rect 57260 28924 57316 28980
rect 57932 28252 57988 28308
rect 57596 27580 57652 27636
rect 56588 27468 56644 27524
rect 58156 27580 58212 27636
rect 57820 27244 57876 27300
rect 56252 27132 56308 27188
rect 55580 26460 55636 26516
rect 57596 26796 57652 26852
rect 55580 25900 55636 25956
rect 52668 24892 52724 24948
rect 55132 25564 55188 25620
rect 53452 24332 53508 24388
rect 58156 26796 58212 26852
rect 57932 26236 57988 26292
rect 57932 25618 57988 25620
rect 57932 25566 57934 25618
rect 57934 25566 57986 25618
rect 57986 25566 57988 25618
rect 57932 25564 57988 25566
rect 57820 25228 57876 25284
rect 57932 24892 57988 24948
rect 55356 24498 55412 24500
rect 55356 24446 55358 24498
rect 55358 24446 55410 24498
rect 55410 24446 55412 24498
rect 55356 24444 55412 24446
rect 57932 23436 57988 23492
rect 53452 22988 53508 23044
rect 55356 22930 55412 22932
rect 55356 22878 55358 22930
rect 55358 22878 55410 22930
rect 55410 22878 55412 22930
rect 55356 22876 55412 22878
rect 52108 22316 52164 22372
rect 52668 22652 52724 22708
rect 53564 22428 53620 22484
rect 50556 21978 50612 21980
rect 50556 21926 50558 21978
rect 50558 21926 50610 21978
rect 50610 21926 50612 21978
rect 50556 21924 50612 21926
rect 50660 21978 50716 21980
rect 50660 21926 50662 21978
rect 50662 21926 50714 21978
rect 50714 21926 50716 21978
rect 50660 21924 50716 21926
rect 50764 21978 50820 21980
rect 50764 21926 50766 21978
rect 50766 21926 50818 21978
rect 50818 21926 50820 21978
rect 50764 21924 50820 21926
rect 53452 21586 53508 21588
rect 53452 21534 53454 21586
rect 53454 21534 53506 21586
rect 53506 21534 53508 21586
rect 53452 21532 53508 21534
rect 46508 19292 46564 19348
rect 45164 18060 45220 18116
rect 45612 17724 45668 17780
rect 45276 17666 45332 17668
rect 45276 17614 45278 17666
rect 45278 17614 45330 17666
rect 45330 17614 45332 17666
rect 45276 17612 45332 17614
rect 43820 16828 43876 16884
rect 46732 18450 46788 18452
rect 46732 18398 46734 18450
rect 46734 18398 46786 18450
rect 46786 18398 46788 18450
rect 46732 18396 46788 18398
rect 46396 18338 46452 18340
rect 46396 18286 46398 18338
rect 46398 18286 46450 18338
rect 46450 18286 46452 18338
rect 46396 18284 46452 18286
rect 45948 18060 46004 18116
rect 47964 20018 48020 20020
rect 47964 19966 47966 20018
rect 47966 19966 48018 20018
rect 48018 19966 48020 20018
rect 47964 19964 48020 19966
rect 48188 19852 48244 19908
rect 47740 18396 47796 18452
rect 46956 17778 47012 17780
rect 46956 17726 46958 17778
rect 46958 17726 47010 17778
rect 47010 17726 47012 17778
rect 46956 17724 47012 17726
rect 48076 17778 48132 17780
rect 48076 17726 48078 17778
rect 48078 17726 48130 17778
rect 48130 17726 48132 17778
rect 48076 17724 48132 17726
rect 45836 17554 45892 17556
rect 45836 17502 45838 17554
rect 45838 17502 45890 17554
rect 45890 17502 45892 17554
rect 45836 17500 45892 17502
rect 45724 16716 45780 16772
rect 46508 17164 46564 17220
rect 43820 16604 43876 16660
rect 43708 16156 43764 16212
rect 42700 16098 42756 16100
rect 42700 16046 42702 16098
rect 42702 16046 42754 16098
rect 42754 16046 42756 16098
rect 42700 16044 42756 16046
rect 43708 15820 43764 15876
rect 41132 15426 41188 15428
rect 41132 15374 41134 15426
rect 41134 15374 41186 15426
rect 41186 15374 41188 15426
rect 41132 15372 41188 15374
rect 41580 15314 41636 15316
rect 41580 15262 41582 15314
rect 41582 15262 41634 15314
rect 41634 15262 41636 15314
rect 41580 15260 41636 15262
rect 41356 15148 41412 15204
rect 40908 14812 40964 14868
rect 42476 15260 42532 15316
rect 42252 15148 42308 15204
rect 40572 14140 40628 14196
rect 45052 15260 45108 15316
rect 44380 14476 44436 14532
rect 45276 15202 45332 15204
rect 45276 15150 45278 15202
rect 45278 15150 45330 15202
rect 45330 15150 45332 15202
rect 45276 15148 45332 15150
rect 45388 15314 45444 15316
rect 45388 15262 45390 15314
rect 45390 15262 45442 15314
rect 45442 15262 45444 15314
rect 45388 15260 45444 15262
rect 45724 15148 45780 15204
rect 40908 13746 40964 13748
rect 40908 13694 40910 13746
rect 40910 13694 40962 13746
rect 40962 13694 40964 13746
rect 40908 13692 40964 13694
rect 45612 14530 45668 14532
rect 45612 14478 45614 14530
rect 45614 14478 45666 14530
rect 45666 14478 45668 14530
rect 45612 14476 45668 14478
rect 41020 13580 41076 13636
rect 41580 13634 41636 13636
rect 41580 13582 41582 13634
rect 41582 13582 41634 13634
rect 41634 13582 41636 13634
rect 41580 13580 41636 13582
rect 43036 12908 43092 12964
rect 41468 12572 41524 12628
rect 41580 12012 41636 12068
rect 42476 12572 42532 12628
rect 41692 12236 41748 12292
rect 39676 11282 39732 11284
rect 39676 11230 39678 11282
rect 39678 11230 39730 11282
rect 39730 11230 39732 11282
rect 39676 11228 39732 11230
rect 39116 10722 39172 10724
rect 39116 10670 39118 10722
rect 39118 10670 39170 10722
rect 39170 10670 39172 10722
rect 39116 10668 39172 10670
rect 39340 10610 39396 10612
rect 39340 10558 39342 10610
rect 39342 10558 39394 10610
rect 39394 10558 39396 10610
rect 39340 10556 39396 10558
rect 38220 8204 38276 8260
rect 38444 8764 38500 8820
rect 38332 7420 38388 7476
rect 37772 6636 37828 6692
rect 38108 6690 38164 6692
rect 38108 6638 38110 6690
rect 38110 6638 38162 6690
rect 38162 6638 38164 6690
rect 38108 6636 38164 6638
rect 37660 6076 37716 6132
rect 37996 6524 38052 6580
rect 37212 6018 37268 6020
rect 37212 5966 37214 6018
rect 37214 5966 37266 6018
rect 37266 5966 37268 6018
rect 37212 5964 37268 5966
rect 37100 5292 37156 5348
rect 37772 5906 37828 5908
rect 37772 5854 37774 5906
rect 37774 5854 37826 5906
rect 37826 5854 37828 5906
rect 37772 5852 37828 5854
rect 37548 5404 37604 5460
rect 37660 5516 37716 5572
rect 37212 5122 37268 5124
rect 37212 5070 37214 5122
rect 37214 5070 37266 5122
rect 37266 5070 37268 5122
rect 37212 5068 37268 5070
rect 37660 5122 37716 5124
rect 37660 5070 37662 5122
rect 37662 5070 37714 5122
rect 37714 5070 37716 5122
rect 37660 5068 37716 5070
rect 37772 4956 37828 5012
rect 37884 5292 37940 5348
rect 37548 4844 37604 4900
rect 36764 4732 36820 4788
rect 36988 4338 37044 4340
rect 36988 4286 36990 4338
rect 36990 4286 37042 4338
rect 37042 4286 37044 4338
rect 36988 4284 37044 4286
rect 36316 3948 36372 4004
rect 36204 3666 36260 3668
rect 36204 3614 36206 3666
rect 36206 3614 36258 3666
rect 36258 3614 36260 3666
rect 36204 3612 36260 3614
rect 37212 3724 37268 3780
rect 38332 6748 38388 6804
rect 38108 6412 38164 6468
rect 37436 3724 37492 3780
rect 36988 3500 37044 3556
rect 38220 5180 38276 5236
rect 38220 4508 38276 4564
rect 39452 9996 39508 10052
rect 38892 9266 38948 9268
rect 38892 9214 38894 9266
rect 38894 9214 38946 9266
rect 38946 9214 38948 9266
rect 38892 9212 38948 9214
rect 40124 11170 40180 11172
rect 40124 11118 40126 11170
rect 40126 11118 40178 11170
rect 40178 11118 40180 11170
rect 40124 11116 40180 11118
rect 40236 11004 40292 11060
rect 40572 10668 40628 10724
rect 39900 9826 39956 9828
rect 39900 9774 39902 9826
rect 39902 9774 39954 9826
rect 39954 9774 39956 9826
rect 39900 9772 39956 9774
rect 40124 10332 40180 10388
rect 41020 10556 41076 10612
rect 40908 10332 40964 10388
rect 41580 10220 41636 10276
rect 40908 9884 40964 9940
rect 39340 9212 39396 9268
rect 40236 9548 40292 9604
rect 38780 8988 38836 9044
rect 40124 9212 40180 9268
rect 40348 9436 40404 9492
rect 42476 12124 42532 12180
rect 43148 13468 43204 13524
rect 42924 11954 42980 11956
rect 42924 11902 42926 11954
rect 42926 11902 42978 11954
rect 42978 11902 42980 11954
rect 42924 11900 42980 11902
rect 42588 10892 42644 10948
rect 43260 12124 43316 12180
rect 43708 12796 43764 12852
rect 45276 13580 45332 13636
rect 44044 12572 44100 12628
rect 44828 12850 44884 12852
rect 44828 12798 44830 12850
rect 44830 12798 44882 12850
rect 44882 12798 44884 12850
rect 44828 12796 44884 12798
rect 44268 12124 44324 12180
rect 45164 12962 45220 12964
rect 45164 12910 45166 12962
rect 45166 12910 45218 12962
rect 45218 12910 45220 12962
rect 45164 12908 45220 12910
rect 45052 12348 45108 12404
rect 43708 12012 43764 12068
rect 45164 12178 45220 12180
rect 45164 12126 45166 12178
rect 45166 12126 45218 12178
rect 45218 12126 45220 12178
rect 45164 12124 45220 12126
rect 43148 11116 43204 11172
rect 41356 9602 41412 9604
rect 41356 9550 41358 9602
rect 41358 9550 41410 9602
rect 41410 9550 41412 9602
rect 41356 9548 41412 9550
rect 41692 9436 41748 9492
rect 39004 8316 39060 8372
rect 38780 8258 38836 8260
rect 38780 8206 38782 8258
rect 38782 8206 38834 8258
rect 38834 8206 38836 8258
rect 38780 8204 38836 8206
rect 38668 7308 38724 7364
rect 38444 6524 38500 6580
rect 38444 6300 38500 6356
rect 39116 7420 39172 7476
rect 39900 7756 39956 7812
rect 40124 7586 40180 7588
rect 40124 7534 40126 7586
rect 40126 7534 40178 7586
rect 40178 7534 40180 7586
rect 40124 7532 40180 7534
rect 40796 7474 40852 7476
rect 40796 7422 40798 7474
rect 40798 7422 40850 7474
rect 40850 7422 40852 7474
rect 40796 7420 40852 7422
rect 41020 7756 41076 7812
rect 41132 7308 41188 7364
rect 40908 7084 40964 7140
rect 39228 6748 39284 6804
rect 39116 6466 39172 6468
rect 39116 6414 39118 6466
rect 39118 6414 39170 6466
rect 39170 6414 39172 6466
rect 39116 6412 39172 6414
rect 39676 6300 39732 6356
rect 38892 5964 38948 6020
rect 39228 6188 39284 6244
rect 38892 5794 38948 5796
rect 38892 5742 38894 5794
rect 38894 5742 38946 5794
rect 38946 5742 38948 5794
rect 38892 5740 38948 5742
rect 38444 5180 38500 5236
rect 38668 5292 38724 5348
rect 39564 6076 39620 6132
rect 39340 5682 39396 5684
rect 39340 5630 39342 5682
rect 39342 5630 39394 5682
rect 39394 5630 39396 5682
rect 39340 5628 39396 5630
rect 39340 5234 39396 5236
rect 39340 5182 39342 5234
rect 39342 5182 39394 5234
rect 39394 5182 39396 5234
rect 39340 5180 39396 5182
rect 40012 5852 40068 5908
rect 39788 5628 39844 5684
rect 41020 6412 41076 6468
rect 41244 6636 41300 6692
rect 40908 5628 40964 5684
rect 41580 7586 41636 7588
rect 41580 7534 41582 7586
rect 41582 7534 41634 7586
rect 41634 7534 41636 7586
rect 41580 7532 41636 7534
rect 42924 9436 42980 9492
rect 43260 10444 43316 10500
rect 45612 11282 45668 11284
rect 45612 11230 45614 11282
rect 45614 11230 45666 11282
rect 45666 11230 45668 11282
rect 45612 11228 45668 11230
rect 43484 11116 43540 11172
rect 44492 11116 44548 11172
rect 45276 11004 45332 11060
rect 43372 10108 43428 10164
rect 43036 9154 43092 9156
rect 43036 9102 43038 9154
rect 43038 9102 43090 9154
rect 43090 9102 43092 9154
rect 43036 9100 43092 9102
rect 43148 8988 43204 9044
rect 46060 14642 46116 14644
rect 46060 14590 46062 14642
rect 46062 14590 46114 14642
rect 46114 14590 46116 14642
rect 46060 14588 46116 14590
rect 46396 15260 46452 15316
rect 46508 15148 46564 15204
rect 47068 15314 47124 15316
rect 47068 15262 47070 15314
rect 47070 15262 47122 15314
rect 47122 15262 47124 15314
rect 47068 15260 47124 15262
rect 46956 14588 47012 14644
rect 46956 13804 47012 13860
rect 47516 15260 47572 15316
rect 48748 17724 48804 17780
rect 50556 20410 50612 20412
rect 50556 20358 50558 20410
rect 50558 20358 50610 20410
rect 50610 20358 50612 20410
rect 50556 20356 50612 20358
rect 50660 20410 50716 20412
rect 50660 20358 50662 20410
rect 50662 20358 50714 20410
rect 50714 20358 50716 20410
rect 50660 20356 50716 20358
rect 50764 20410 50820 20412
rect 50764 20358 50766 20410
rect 50766 20358 50818 20410
rect 50818 20358 50820 20410
rect 50764 20356 50820 20358
rect 49980 20018 50036 20020
rect 49980 19966 49982 20018
rect 49982 19966 50034 20018
rect 50034 19966 50036 20018
rect 49980 19964 50036 19966
rect 49644 19180 49700 19236
rect 52108 19628 52164 19684
rect 50556 18842 50612 18844
rect 50556 18790 50558 18842
rect 50558 18790 50610 18842
rect 50610 18790 50612 18842
rect 50556 18788 50612 18790
rect 50660 18842 50716 18844
rect 50660 18790 50662 18842
rect 50662 18790 50714 18842
rect 50714 18790 50716 18842
rect 50660 18788 50716 18790
rect 50764 18842 50820 18844
rect 50764 18790 50766 18842
rect 50766 18790 50818 18842
rect 50818 18790 50820 18842
rect 50764 18788 50820 18790
rect 48972 18508 49028 18564
rect 48860 18060 48916 18116
rect 49084 17388 49140 17444
rect 51212 18284 51268 18340
rect 51100 17948 51156 18004
rect 50764 17890 50820 17892
rect 50764 17838 50766 17890
rect 50766 17838 50818 17890
rect 50818 17838 50820 17890
rect 50764 17836 50820 17838
rect 51548 18226 51604 18228
rect 51548 18174 51550 18226
rect 51550 18174 51602 18226
rect 51602 18174 51604 18226
rect 51548 18172 51604 18174
rect 48188 15372 48244 15428
rect 48412 14642 48468 14644
rect 48412 14590 48414 14642
rect 48414 14590 48466 14642
rect 48466 14590 48468 14642
rect 48412 14588 48468 14590
rect 48748 16044 48804 16100
rect 49644 16044 49700 16100
rect 53228 19628 53284 19684
rect 51996 18338 52052 18340
rect 51996 18286 51998 18338
rect 51998 18286 52050 18338
rect 52050 18286 52052 18338
rect 51996 18284 52052 18286
rect 51772 17948 51828 18004
rect 52220 17836 52276 17892
rect 52668 17666 52724 17668
rect 52668 17614 52670 17666
rect 52670 17614 52722 17666
rect 52722 17614 52724 17666
rect 52668 17612 52724 17614
rect 50556 17274 50612 17276
rect 50556 17222 50558 17274
rect 50558 17222 50610 17274
rect 50610 17222 50612 17274
rect 50556 17220 50612 17222
rect 50660 17274 50716 17276
rect 50660 17222 50662 17274
rect 50662 17222 50714 17274
rect 50714 17222 50716 17274
rect 50660 17220 50716 17222
rect 50764 17274 50820 17276
rect 50764 17222 50766 17274
rect 50766 17222 50818 17274
rect 50818 17222 50820 17274
rect 50764 17220 50820 17222
rect 50652 16994 50708 16996
rect 50652 16942 50654 16994
rect 50654 16942 50706 16994
rect 50706 16942 50708 16994
rect 50652 16940 50708 16942
rect 51324 16882 51380 16884
rect 51324 16830 51326 16882
rect 51326 16830 51378 16882
rect 51378 16830 51380 16882
rect 51324 16828 51380 16830
rect 50204 16044 50260 16100
rect 50556 15706 50612 15708
rect 50556 15654 50558 15706
rect 50558 15654 50610 15706
rect 50610 15654 50612 15706
rect 50556 15652 50612 15654
rect 50660 15706 50716 15708
rect 50660 15654 50662 15706
rect 50662 15654 50714 15706
rect 50714 15654 50716 15706
rect 50660 15652 50716 15654
rect 50764 15706 50820 15708
rect 50764 15654 50766 15706
rect 50766 15654 50818 15706
rect 50818 15654 50820 15706
rect 50764 15652 50820 15654
rect 49196 14476 49252 14532
rect 50540 14530 50596 14532
rect 50540 14478 50542 14530
rect 50542 14478 50594 14530
rect 50594 14478 50596 14530
rect 50540 14476 50596 14478
rect 47852 13858 47908 13860
rect 47852 13806 47854 13858
rect 47854 13806 47906 13858
rect 47906 13806 47908 13858
rect 47852 13804 47908 13806
rect 46508 13634 46564 13636
rect 46508 13582 46510 13634
rect 46510 13582 46562 13634
rect 46562 13582 46564 13634
rect 46508 13580 46564 13582
rect 47516 13692 47572 13748
rect 46284 12962 46340 12964
rect 46284 12910 46286 12962
rect 46286 12910 46338 12962
rect 46338 12910 46340 12962
rect 46284 12908 46340 12910
rect 47068 12962 47124 12964
rect 47068 12910 47070 12962
rect 47070 12910 47122 12962
rect 47122 12910 47124 12962
rect 47068 12908 47124 12910
rect 46172 12348 46228 12404
rect 47292 12850 47348 12852
rect 47292 12798 47294 12850
rect 47294 12798 47346 12850
rect 47346 12798 47348 12850
rect 47292 12796 47348 12798
rect 47292 12402 47348 12404
rect 47292 12350 47294 12402
rect 47294 12350 47346 12402
rect 47346 12350 47348 12402
rect 47292 12348 47348 12350
rect 48076 13746 48132 13748
rect 48076 13694 48078 13746
rect 48078 13694 48130 13746
rect 48130 13694 48132 13746
rect 48076 13692 48132 13694
rect 47740 13580 47796 13636
rect 48300 12850 48356 12852
rect 48300 12798 48302 12850
rect 48302 12798 48354 12850
rect 48354 12798 48356 12850
rect 48300 12796 48356 12798
rect 47180 11900 47236 11956
rect 48412 12348 48468 12404
rect 47628 11676 47684 11732
rect 47740 11900 47796 11956
rect 47068 11228 47124 11284
rect 42588 8930 42644 8932
rect 42588 8878 42590 8930
rect 42590 8878 42642 8930
rect 42642 8878 42644 8930
rect 42588 8876 42644 8878
rect 42028 7420 42084 7476
rect 42588 7532 42644 7588
rect 42252 7308 42308 7364
rect 41356 5964 41412 6020
rect 41804 5906 41860 5908
rect 41804 5854 41806 5906
rect 41806 5854 41858 5906
rect 41858 5854 41860 5906
rect 41804 5852 41860 5854
rect 41132 5180 41188 5236
rect 39788 5122 39844 5124
rect 39788 5070 39790 5122
rect 39790 5070 39842 5122
rect 39842 5070 39844 5122
rect 39788 5068 39844 5070
rect 40684 4732 40740 4788
rect 38892 3612 38948 3668
rect 39676 3612 39732 3668
rect 39116 3388 39172 3444
rect 39004 3164 39060 3220
rect 40012 4338 40068 4340
rect 40012 4286 40014 4338
rect 40014 4286 40066 4338
rect 40066 4286 40068 4338
rect 40012 4284 40068 4286
rect 40348 3836 40404 3892
rect 40908 4562 40964 4564
rect 40908 4510 40910 4562
rect 40910 4510 40962 4562
rect 40962 4510 40964 4562
rect 40908 4508 40964 4510
rect 40908 3948 40964 4004
rect 41356 5068 41412 5124
rect 42252 6860 42308 6916
rect 42588 6748 42644 6804
rect 42364 6690 42420 6692
rect 42364 6638 42366 6690
rect 42366 6638 42418 6690
rect 42418 6638 42420 6690
rect 42364 6636 42420 6638
rect 43820 9042 43876 9044
rect 43820 8990 43822 9042
rect 43822 8990 43874 9042
rect 43874 8990 43876 9042
rect 43820 8988 43876 8990
rect 45612 9548 45668 9604
rect 44492 9100 44548 9156
rect 44044 8428 44100 8484
rect 43484 7756 43540 7812
rect 42924 5682 42980 5684
rect 42924 5630 42926 5682
rect 42926 5630 42978 5682
rect 42978 5630 42980 5682
rect 42924 5628 42980 5630
rect 43148 5292 43204 5348
rect 43036 5068 43092 5124
rect 42252 4898 42308 4900
rect 42252 4846 42254 4898
rect 42254 4846 42306 4898
rect 42306 4846 42308 4898
rect 42252 4844 42308 4846
rect 42364 4508 42420 4564
rect 42028 4284 42084 4340
rect 42364 4338 42420 4340
rect 42364 4286 42366 4338
rect 42366 4286 42418 4338
rect 42418 4286 42420 4338
rect 42364 4284 42420 4286
rect 42140 4172 42196 4228
rect 42364 3778 42420 3780
rect 42364 3726 42366 3778
rect 42366 3726 42418 3778
rect 42418 3726 42420 3778
rect 42364 3724 42420 3726
rect 42812 4898 42868 4900
rect 42812 4846 42814 4898
rect 42814 4846 42866 4898
rect 42866 4846 42868 4898
rect 42812 4844 42868 4846
rect 42700 3724 42756 3780
rect 43148 4284 43204 4340
rect 43372 3948 43428 4004
rect 41580 3554 41636 3556
rect 41580 3502 41582 3554
rect 41582 3502 41634 3554
rect 41634 3502 41636 3554
rect 41580 3500 41636 3502
rect 43148 3388 43204 3444
rect 43708 7362 43764 7364
rect 43708 7310 43710 7362
rect 43710 7310 43762 7362
rect 43762 7310 43764 7362
rect 43708 7308 43764 7310
rect 44044 6636 44100 6692
rect 44156 7474 44212 7476
rect 44156 7422 44158 7474
rect 44158 7422 44210 7474
rect 44210 7422 44212 7474
rect 44156 7420 44212 7422
rect 44156 5852 44212 5908
rect 43708 5122 43764 5124
rect 43708 5070 43710 5122
rect 43710 5070 43762 5122
rect 43762 5070 43764 5122
rect 43708 5068 43764 5070
rect 44268 5628 44324 5684
rect 44044 5292 44100 5348
rect 44156 4226 44212 4228
rect 44156 4174 44158 4226
rect 44158 4174 44210 4226
rect 44210 4174 44212 4226
rect 44156 4172 44212 4174
rect 43820 3612 43876 3668
rect 40012 3164 40068 3220
rect 45612 9100 45668 9156
rect 45388 8930 45444 8932
rect 45388 8878 45390 8930
rect 45390 8878 45442 8930
rect 45442 8878 45444 8930
rect 45388 8876 45444 8878
rect 45276 8818 45332 8820
rect 45276 8766 45278 8818
rect 45278 8766 45330 8818
rect 45330 8766 45332 8818
rect 45276 8764 45332 8766
rect 45500 6524 45556 6580
rect 45276 6412 45332 6468
rect 45948 9100 46004 9156
rect 46284 10108 46340 10164
rect 46172 9602 46228 9604
rect 46172 9550 46174 9602
rect 46174 9550 46226 9602
rect 46226 9550 46228 9602
rect 46172 9548 46228 9550
rect 46508 8876 46564 8932
rect 46060 8764 46116 8820
rect 48300 11170 48356 11172
rect 48300 11118 48302 11170
rect 48302 11118 48354 11170
rect 48354 11118 48356 11170
rect 48300 11116 48356 11118
rect 50556 14138 50612 14140
rect 50556 14086 50558 14138
rect 50558 14086 50610 14138
rect 50610 14086 50612 14138
rect 50556 14084 50612 14086
rect 50660 14138 50716 14140
rect 50660 14086 50662 14138
rect 50662 14086 50714 14138
rect 50714 14086 50716 14138
rect 50660 14084 50716 14086
rect 50764 14138 50820 14140
rect 50764 14086 50766 14138
rect 50766 14086 50818 14138
rect 50818 14086 50820 14138
rect 50764 14084 50820 14086
rect 49084 13858 49140 13860
rect 49084 13806 49086 13858
rect 49086 13806 49138 13858
rect 49138 13806 49140 13858
rect 49084 13804 49140 13806
rect 49756 13858 49812 13860
rect 49756 13806 49758 13858
rect 49758 13806 49810 13858
rect 49810 13806 49812 13858
rect 49756 13804 49812 13806
rect 50652 13804 50708 13860
rect 48748 13746 48804 13748
rect 48748 13694 48750 13746
rect 48750 13694 48802 13746
rect 48802 13694 48804 13746
rect 48748 13692 48804 13694
rect 49980 13746 50036 13748
rect 49980 13694 49982 13746
rect 49982 13694 50034 13746
rect 50034 13694 50036 13746
rect 49980 13692 50036 13694
rect 51212 14306 51268 14308
rect 51212 14254 51214 14306
rect 51214 14254 51266 14306
rect 51266 14254 51268 14306
rect 51212 14252 51268 14254
rect 51772 14476 51828 14532
rect 52108 16828 52164 16884
rect 51996 15538 52052 15540
rect 51996 15486 51998 15538
rect 51998 15486 52050 15538
rect 52050 15486 52052 15538
rect 51996 15484 52052 15486
rect 53452 18450 53508 18452
rect 53452 18398 53454 18450
rect 53454 18398 53506 18450
rect 53506 18398 53508 18450
rect 53452 18396 53508 18398
rect 52780 16828 52836 16884
rect 55580 22370 55636 22372
rect 55580 22318 55582 22370
rect 55582 22318 55634 22370
rect 55634 22318 55636 22370
rect 55580 22316 55636 22318
rect 57932 22204 57988 22260
rect 55020 21532 55076 21588
rect 55468 21644 55524 21700
rect 53676 20860 53732 20916
rect 55356 20860 55412 20916
rect 57932 20076 57988 20132
rect 55356 19794 55412 19796
rect 55356 19742 55358 19794
rect 55358 19742 55410 19794
rect 55410 19742 55412 19794
rect 55356 19740 55412 19742
rect 55580 19234 55636 19236
rect 55580 19182 55582 19234
rect 55582 19182 55634 19234
rect 55634 19182 55636 19234
rect 55580 19180 55636 19182
rect 57932 18844 57988 18900
rect 55356 18226 55412 18228
rect 55356 18174 55358 18226
rect 55358 18174 55410 18226
rect 55410 18174 55412 18226
rect 55356 18172 55412 18174
rect 55580 17666 55636 17668
rect 55580 17614 55582 17666
rect 55582 17614 55634 17666
rect 55634 17614 55636 17666
rect 55580 17612 55636 17614
rect 55020 16828 55076 16884
rect 55356 17500 55412 17556
rect 52780 16604 52836 16660
rect 52332 15484 52388 15540
rect 51996 14588 52052 14644
rect 51884 13916 51940 13972
rect 50652 13468 50708 13524
rect 49308 11954 49364 11956
rect 49308 11902 49310 11954
rect 49310 11902 49362 11954
rect 49362 11902 49364 11954
rect 49308 11900 49364 11902
rect 49196 11116 49252 11172
rect 50092 12684 50148 12740
rect 49868 12124 49924 12180
rect 49980 12012 50036 12068
rect 51884 12962 51940 12964
rect 51884 12910 51886 12962
rect 51886 12910 51938 12962
rect 51938 12910 51940 12962
rect 51884 12908 51940 12910
rect 50556 12570 50612 12572
rect 50556 12518 50558 12570
rect 50558 12518 50610 12570
rect 50610 12518 50612 12570
rect 50556 12516 50612 12518
rect 50660 12570 50716 12572
rect 50660 12518 50662 12570
rect 50662 12518 50714 12570
rect 50714 12518 50716 12570
rect 50660 12516 50716 12518
rect 50764 12570 50820 12572
rect 50764 12518 50766 12570
rect 50766 12518 50818 12570
rect 50818 12518 50820 12570
rect 50764 12516 50820 12518
rect 50988 12124 51044 12180
rect 50652 11788 50708 11844
rect 51100 11676 51156 11732
rect 50316 11282 50372 11284
rect 50316 11230 50318 11282
rect 50318 11230 50370 11282
rect 50370 11230 50372 11282
rect 50316 11228 50372 11230
rect 47180 9548 47236 9604
rect 47852 9154 47908 9156
rect 47852 9102 47854 9154
rect 47854 9102 47906 9154
rect 47906 9102 47908 9154
rect 47852 9100 47908 9102
rect 46956 8764 47012 8820
rect 46396 7420 46452 7476
rect 47180 7474 47236 7476
rect 47180 7422 47182 7474
rect 47182 7422 47234 7474
rect 47234 7422 47236 7474
rect 47180 7420 47236 7422
rect 44828 5906 44884 5908
rect 44828 5854 44830 5906
rect 44830 5854 44882 5906
rect 44882 5854 44884 5906
rect 44828 5852 44884 5854
rect 45276 5628 45332 5684
rect 45164 5292 45220 5348
rect 44716 5122 44772 5124
rect 44716 5070 44718 5122
rect 44718 5070 44770 5122
rect 44770 5070 44772 5122
rect 44716 5068 44772 5070
rect 44940 4338 44996 4340
rect 44940 4286 44942 4338
rect 44942 4286 44994 4338
rect 44994 4286 44996 4338
rect 44940 4284 44996 4286
rect 44716 4226 44772 4228
rect 44716 4174 44718 4226
rect 44718 4174 44770 4226
rect 44770 4174 44772 4226
rect 44716 4172 44772 4174
rect 44604 3724 44660 3780
rect 44604 3442 44660 3444
rect 44604 3390 44606 3442
rect 44606 3390 44658 3442
rect 44658 3390 44660 3442
rect 44604 3388 44660 3390
rect 45724 5122 45780 5124
rect 45724 5070 45726 5122
rect 45726 5070 45778 5122
rect 45778 5070 45780 5122
rect 45724 5068 45780 5070
rect 45164 4508 45220 4564
rect 46060 6748 46116 6804
rect 46284 6636 46340 6692
rect 48188 10444 48244 10500
rect 49644 10498 49700 10500
rect 49644 10446 49646 10498
rect 49646 10446 49698 10498
rect 49698 10446 49700 10498
rect 49644 10444 49700 10446
rect 48524 9660 48580 9716
rect 50556 11002 50612 11004
rect 50556 10950 50558 11002
rect 50558 10950 50610 11002
rect 50610 10950 50612 11002
rect 50556 10948 50612 10950
rect 50660 11002 50716 11004
rect 50660 10950 50662 11002
rect 50662 10950 50714 11002
rect 50714 10950 50716 11002
rect 50660 10948 50716 10950
rect 50764 11002 50820 11004
rect 50764 10950 50766 11002
rect 50766 10950 50818 11002
rect 50818 10950 50820 11002
rect 50764 10948 50820 10950
rect 51996 12850 52052 12852
rect 51996 12798 51998 12850
rect 51998 12798 52050 12850
rect 52050 12798 52052 12850
rect 51996 12796 52052 12798
rect 52444 15090 52500 15092
rect 52444 15038 52446 15090
rect 52446 15038 52498 15090
rect 52498 15038 52500 15090
rect 52444 15036 52500 15038
rect 52892 14812 52948 14868
rect 57932 17500 57988 17556
rect 55356 16156 55412 16212
rect 55580 16098 55636 16100
rect 55580 16046 55582 16098
rect 55582 16046 55634 16098
rect 55634 16046 55636 16098
rect 55580 16044 55636 16046
rect 54236 15484 54292 15540
rect 57932 15484 57988 15540
rect 53004 14754 53060 14756
rect 53004 14702 53006 14754
rect 53006 14702 53058 14754
rect 53058 14702 53060 14754
rect 53004 14700 53060 14702
rect 52668 14588 52724 14644
rect 52892 14530 52948 14532
rect 52892 14478 52894 14530
rect 52894 14478 52946 14530
rect 52946 14478 52948 14530
rect 52892 14476 52948 14478
rect 53452 15314 53508 15316
rect 53452 15262 53454 15314
rect 53454 15262 53506 15314
rect 53506 15262 53508 15314
rect 53452 15260 53508 15262
rect 53116 14252 53172 14308
rect 53340 15036 53396 15092
rect 54124 14812 54180 14868
rect 55356 14812 55412 14868
rect 55580 15036 55636 15092
rect 54908 14642 54964 14644
rect 54908 14590 54910 14642
rect 54910 14590 54962 14642
rect 54962 14590 54964 14642
rect 54908 14588 54964 14590
rect 54124 14476 54180 14532
rect 53004 13916 53060 13972
rect 53788 14252 53844 14308
rect 53564 13858 53620 13860
rect 53564 13806 53566 13858
rect 53566 13806 53618 13858
rect 53618 13806 53620 13858
rect 53564 13804 53620 13806
rect 54236 13804 54292 13860
rect 52668 12962 52724 12964
rect 52668 12910 52670 12962
rect 52670 12910 52722 12962
rect 52722 12910 52724 12962
rect 52668 12908 52724 12910
rect 56588 14476 56644 14532
rect 53116 12850 53172 12852
rect 53116 12798 53118 12850
rect 53118 12798 53170 12850
rect 53170 12798 53172 12850
rect 53116 12796 53172 12798
rect 51996 12236 52052 12292
rect 51884 12178 51940 12180
rect 51884 12126 51886 12178
rect 51886 12126 51938 12178
rect 51938 12126 51940 12178
rect 51884 12124 51940 12126
rect 51100 10722 51156 10724
rect 51100 10670 51102 10722
rect 51102 10670 51154 10722
rect 51154 10670 51156 10722
rect 51100 10668 51156 10670
rect 49868 9772 49924 9828
rect 50540 9826 50596 9828
rect 50540 9774 50542 9826
rect 50542 9774 50594 9826
rect 50594 9774 50596 9826
rect 50540 9772 50596 9774
rect 49644 9324 49700 9380
rect 49532 8428 49588 8484
rect 47292 6412 47348 6468
rect 46284 6076 46340 6132
rect 47740 6130 47796 6132
rect 47740 6078 47742 6130
rect 47742 6078 47794 6130
rect 47794 6078 47796 6130
rect 47740 6076 47796 6078
rect 46508 5628 46564 5684
rect 45724 3836 45780 3892
rect 46284 3554 46340 3556
rect 46284 3502 46286 3554
rect 46286 3502 46338 3554
rect 46338 3502 46340 3554
rect 46284 3500 46340 3502
rect 46956 5292 47012 5348
rect 47068 5234 47124 5236
rect 47068 5182 47070 5234
rect 47070 5182 47122 5234
rect 47122 5182 47124 5234
rect 47068 5180 47124 5182
rect 47852 5794 47908 5796
rect 47852 5742 47854 5794
rect 47854 5742 47906 5794
rect 47906 5742 47908 5794
rect 47852 5740 47908 5742
rect 47516 5682 47572 5684
rect 47516 5630 47518 5682
rect 47518 5630 47570 5682
rect 47570 5630 47572 5682
rect 47516 5628 47572 5630
rect 46620 3836 46676 3892
rect 47404 3836 47460 3892
rect 49308 8092 49364 8148
rect 48748 7868 48804 7924
rect 48972 7250 49028 7252
rect 48972 7198 48974 7250
rect 48974 7198 49026 7250
rect 49026 7198 49028 7250
rect 48972 7196 49028 7198
rect 50988 9660 51044 9716
rect 50556 9434 50612 9436
rect 50556 9382 50558 9434
rect 50558 9382 50610 9434
rect 50610 9382 50612 9434
rect 50556 9380 50612 9382
rect 50660 9434 50716 9436
rect 50660 9382 50662 9434
rect 50662 9382 50714 9434
rect 50714 9382 50716 9434
rect 50660 9380 50716 9382
rect 50764 9434 50820 9436
rect 50764 9382 50766 9434
rect 50766 9382 50818 9434
rect 50818 9382 50820 9434
rect 50764 9380 50820 9382
rect 52220 11282 52276 11284
rect 52220 11230 52222 11282
rect 52222 11230 52274 11282
rect 52274 11230 52276 11282
rect 52220 11228 52276 11230
rect 51548 10332 51604 10388
rect 51772 9996 51828 10052
rect 51436 9212 51492 9268
rect 50988 8764 51044 8820
rect 49868 8540 49924 8596
rect 49644 8370 49700 8372
rect 49644 8318 49646 8370
rect 49646 8318 49698 8370
rect 49698 8318 49700 8370
rect 49644 8316 49700 8318
rect 55468 12796 55524 12852
rect 55244 12684 55300 12740
rect 54460 12572 54516 12628
rect 53452 12236 53508 12292
rect 55132 12290 55188 12292
rect 55132 12238 55134 12290
rect 55134 12238 55186 12290
rect 55186 12238 55188 12290
rect 55132 12236 55188 12238
rect 53116 10892 53172 10948
rect 53564 11394 53620 11396
rect 53564 11342 53566 11394
rect 53566 11342 53618 11394
rect 53618 11342 53620 11394
rect 53564 11340 53620 11342
rect 55356 11788 55412 11844
rect 52332 10722 52388 10724
rect 52332 10670 52334 10722
rect 52334 10670 52386 10722
rect 52386 10670 52388 10722
rect 52332 10668 52388 10670
rect 52220 10610 52276 10612
rect 52220 10558 52222 10610
rect 52222 10558 52274 10610
rect 52274 10558 52276 10610
rect 52220 10556 52276 10558
rect 52668 9996 52724 10052
rect 52108 9826 52164 9828
rect 52108 9774 52110 9826
rect 52110 9774 52162 9826
rect 52162 9774 52164 9826
rect 52108 9772 52164 9774
rect 52892 10556 52948 10612
rect 53676 10892 53732 10948
rect 53900 10610 53956 10612
rect 53900 10558 53902 10610
rect 53902 10558 53954 10610
rect 53954 10558 53956 10610
rect 53900 10556 53956 10558
rect 54236 10498 54292 10500
rect 54236 10446 54238 10498
rect 54238 10446 54290 10498
rect 54290 10446 54292 10498
rect 54236 10444 54292 10446
rect 54684 10444 54740 10500
rect 54908 10668 54964 10724
rect 53452 9884 53508 9940
rect 51660 9042 51716 9044
rect 51660 8990 51662 9042
rect 51662 8990 51714 9042
rect 51714 8990 51716 9042
rect 51660 8988 51716 8990
rect 51660 8764 51716 8820
rect 51212 8370 51268 8372
rect 51212 8318 51214 8370
rect 51214 8318 51266 8370
rect 51266 8318 51268 8370
rect 51212 8316 51268 8318
rect 50204 8204 50260 8260
rect 50988 8258 51044 8260
rect 50988 8206 50990 8258
rect 50990 8206 51042 8258
rect 51042 8206 51044 8258
rect 50988 8204 51044 8206
rect 50556 7866 50612 7868
rect 50556 7814 50558 7866
rect 50558 7814 50610 7866
rect 50610 7814 50612 7866
rect 50556 7812 50612 7814
rect 50660 7866 50716 7868
rect 50660 7814 50662 7866
rect 50662 7814 50714 7866
rect 50714 7814 50716 7866
rect 50660 7812 50716 7814
rect 50764 7866 50820 7868
rect 50764 7814 50766 7866
rect 50766 7814 50818 7866
rect 50818 7814 50820 7866
rect 50764 7812 50820 7814
rect 49868 6748 49924 6804
rect 50428 6748 50484 6804
rect 50204 6636 50260 6692
rect 50876 6690 50932 6692
rect 50876 6638 50878 6690
rect 50878 6638 50930 6690
rect 50930 6638 50932 6690
rect 50876 6636 50932 6638
rect 49756 6578 49812 6580
rect 49756 6526 49758 6578
rect 49758 6526 49810 6578
rect 49810 6526 49812 6578
rect 49756 6524 49812 6526
rect 50428 6524 50484 6580
rect 50204 6466 50260 6468
rect 50204 6414 50206 6466
rect 50206 6414 50258 6466
rect 50258 6414 50260 6466
rect 50204 6412 50260 6414
rect 49196 5740 49252 5796
rect 49308 5852 49364 5908
rect 48412 5234 48468 5236
rect 48412 5182 48414 5234
rect 48414 5182 48466 5234
rect 48466 5182 48468 5234
rect 48412 5180 48468 5182
rect 48972 5180 49028 5236
rect 49756 5180 49812 5236
rect 50556 6298 50612 6300
rect 50556 6246 50558 6298
rect 50558 6246 50610 6298
rect 50610 6246 50612 6298
rect 50556 6244 50612 6246
rect 50660 6298 50716 6300
rect 50660 6246 50662 6298
rect 50662 6246 50714 6298
rect 50714 6246 50716 6298
rect 50660 6244 50716 6246
rect 50764 6298 50820 6300
rect 50764 6246 50766 6298
rect 50766 6246 50818 6298
rect 50818 6246 50820 6298
rect 50764 6244 50820 6246
rect 49868 5740 49924 5796
rect 51772 8652 51828 8708
rect 51772 8428 51828 8484
rect 52892 9212 52948 9268
rect 54124 9938 54180 9940
rect 54124 9886 54126 9938
rect 54126 9886 54178 9938
rect 54178 9886 54180 9938
rect 54124 9884 54180 9886
rect 53676 9660 53732 9716
rect 52892 8428 52948 8484
rect 54124 9042 54180 9044
rect 54124 8990 54126 9042
rect 54126 8990 54178 9042
rect 54178 8990 54180 9042
rect 54124 8988 54180 8990
rect 54572 9826 54628 9828
rect 54572 9774 54574 9826
rect 54574 9774 54626 9826
rect 54626 9774 54628 9826
rect 54572 9772 54628 9774
rect 55020 10556 55076 10612
rect 54684 8988 54740 9044
rect 52780 8204 52836 8260
rect 53452 8204 53508 8260
rect 52892 8092 52948 8148
rect 51772 7644 51828 7700
rect 51996 7644 52052 7700
rect 51324 6578 51380 6580
rect 51324 6526 51326 6578
rect 51326 6526 51378 6578
rect 51378 6526 51380 6578
rect 51324 6524 51380 6526
rect 51100 5906 51156 5908
rect 51100 5854 51102 5906
rect 51102 5854 51154 5906
rect 51154 5854 51156 5906
rect 51100 5852 51156 5854
rect 52556 6748 52612 6804
rect 52780 6412 52836 6468
rect 54460 8258 54516 8260
rect 54460 8206 54462 8258
rect 54462 8206 54514 8258
rect 54514 8206 54516 8258
rect 54460 8204 54516 8206
rect 56924 12796 56980 12852
rect 56588 12684 56644 12740
rect 55580 12124 55636 12180
rect 55692 11340 55748 11396
rect 56028 12572 56084 12628
rect 57036 12178 57092 12180
rect 57036 12126 57038 12178
rect 57038 12126 57090 12178
rect 57090 12126 57092 12178
rect 57036 12124 57092 12126
rect 55804 11282 55860 11284
rect 55804 11230 55806 11282
rect 55806 11230 55858 11282
rect 55858 11230 55860 11282
rect 55804 11228 55860 11230
rect 56812 10668 56868 10724
rect 56476 10610 56532 10612
rect 56476 10558 56478 10610
rect 56478 10558 56530 10610
rect 56530 10558 56532 10610
rect 56476 10556 56532 10558
rect 56028 10444 56084 10500
rect 55580 9772 55636 9828
rect 57036 10444 57092 10500
rect 57148 9660 57204 9716
rect 55916 8652 55972 8708
rect 53228 6972 53284 7028
rect 53004 6748 53060 6804
rect 53900 6972 53956 7028
rect 57484 8652 57540 8708
rect 55916 7586 55972 7588
rect 55916 7534 55918 7586
rect 55918 7534 55970 7586
rect 55970 7534 55972 7586
rect 55916 7532 55972 7534
rect 57148 7532 57204 7588
rect 54572 7420 54628 7476
rect 56588 7474 56644 7476
rect 56588 7422 56590 7474
rect 56590 7422 56642 7474
rect 56642 7422 56644 7474
rect 56588 7420 56644 7422
rect 57260 7644 57316 7700
rect 54684 6972 54740 7028
rect 50092 5234 50148 5236
rect 50092 5182 50094 5234
rect 50094 5182 50146 5234
rect 50146 5182 50148 5234
rect 50092 5180 50148 5182
rect 48188 5122 48244 5124
rect 48188 5070 48190 5122
rect 48190 5070 48242 5122
rect 48242 5070 48244 5122
rect 48188 5068 48244 5070
rect 50556 4730 50612 4732
rect 50556 4678 50558 4730
rect 50558 4678 50610 4730
rect 50610 4678 50612 4730
rect 50556 4676 50612 4678
rect 50660 4730 50716 4732
rect 50660 4678 50662 4730
rect 50662 4678 50714 4730
rect 50714 4678 50716 4730
rect 50660 4676 50716 4678
rect 50764 4730 50820 4732
rect 50764 4678 50766 4730
rect 50766 4678 50818 4730
rect 50818 4678 50820 4730
rect 50764 4676 50820 4678
rect 46732 3442 46788 3444
rect 46732 3390 46734 3442
rect 46734 3390 46786 3442
rect 46786 3390 46788 3442
rect 46732 3388 46788 3390
rect 46508 3276 46564 3332
rect 50556 3162 50612 3164
rect 50556 3110 50558 3162
rect 50558 3110 50610 3162
rect 50610 3110 50612 3162
rect 50556 3108 50612 3110
rect 50660 3162 50716 3164
rect 50660 3110 50662 3162
rect 50662 3110 50714 3162
rect 50714 3110 50716 3162
rect 50660 3108 50716 3110
rect 50764 3162 50820 3164
rect 50764 3110 50766 3162
rect 50766 3110 50818 3162
rect 50818 3110 50820 3162
rect 50764 3108 50820 3110
<< metal3 >>
rect 44370 46844 44380 46900
rect 44436 46844 51436 46900
rect 51492 46844 51502 46900
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 42242 46172 42252 46228
rect 42308 46172 47404 46228
rect 47460 46172 47470 46228
rect 26226 46060 26236 46116
rect 26292 46060 29372 46116
rect 29428 46060 29438 46116
rect 41346 46060 41356 46116
rect 41412 46060 42588 46116
rect 42644 46060 44604 46116
rect 44660 46060 44670 46116
rect 9650 45948 9660 46004
rect 9716 45948 11900 46004
rect 11956 45948 11966 46004
rect 12338 45948 12348 46004
rect 12404 45948 14476 46004
rect 14532 45948 14542 46004
rect 16034 45948 16044 46004
rect 16100 45948 16828 46004
rect 16884 45948 16894 46004
rect 26786 45948 26796 46004
rect 26852 45948 27580 46004
rect 27636 45948 27646 46004
rect 35074 45948 35084 46004
rect 35140 45948 36988 46004
rect 37044 45948 37054 46004
rect 51426 45948 51436 46004
rect 51492 45948 53788 46004
rect 53844 45948 53854 46004
rect 8372 45836 10780 45892
rect 10836 45836 10846 45892
rect 11554 45836 11564 45892
rect 11620 45836 13132 45892
rect 13188 45836 13198 45892
rect 16482 45836 16492 45892
rect 16548 45836 17500 45892
rect 17556 45836 17566 45892
rect 27122 45836 27132 45892
rect 27188 45836 28364 45892
rect 28420 45836 28430 45892
rect 36530 45836 36540 45892
rect 36596 45836 38108 45892
rect 38164 45836 38174 45892
rect 41010 45836 41020 45892
rect 41076 45836 46228 45892
rect 46386 45836 46396 45892
rect 46452 45836 52780 45892
rect 52836 45836 54236 45892
rect 54292 45836 54302 45892
rect 8372 45780 8428 45836
rect 46172 45780 46228 45836
rect 8194 45724 8204 45780
rect 8260 45724 8428 45780
rect 12562 45724 12572 45780
rect 12628 45724 13244 45780
rect 13300 45724 13916 45780
rect 13972 45724 13982 45780
rect 35522 45724 35532 45780
rect 35588 45724 39004 45780
rect 39060 45724 40012 45780
rect 40068 45724 40078 45780
rect 42354 45724 42364 45780
rect 42420 45724 43036 45780
rect 43092 45724 43596 45780
rect 43652 45724 43662 45780
rect 46172 45724 46732 45780
rect 46788 45724 53340 45780
rect 53396 45724 53406 45780
rect 10098 45612 10108 45668
rect 10164 45612 10556 45668
rect 10612 45612 10622 45668
rect 19618 45612 19628 45668
rect 19684 45612 21084 45668
rect 21140 45612 21150 45668
rect 37202 45612 37212 45668
rect 37268 45612 38668 45668
rect 38724 45612 38734 45668
rect 43138 45612 43148 45668
rect 43204 45612 46284 45668
rect 46340 45612 48748 45668
rect 48804 45612 48814 45668
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 50546 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50830 45500
rect 16044 45388 16828 45444
rect 16884 45388 16894 45444
rect 16044 45332 16100 45388
rect 10434 45276 10444 45332
rect 10500 45276 12124 45332
rect 12180 45276 13804 45332
rect 13860 45276 14364 45332
rect 14420 45276 14430 45332
rect 14802 45276 14812 45332
rect 14868 45276 16100 45332
rect 16258 45276 16268 45332
rect 16324 45276 18172 45332
rect 18228 45276 20748 45332
rect 20804 45276 20814 45332
rect 41010 45276 41020 45332
rect 41076 45276 46396 45332
rect 46452 45276 46462 45332
rect 49074 45276 49084 45332
rect 49140 45276 52220 45332
rect 52276 45276 52286 45332
rect 9874 45164 9884 45220
rect 9940 45164 11116 45220
rect 11172 45164 12236 45220
rect 12292 45164 13468 45220
rect 13524 45164 14140 45220
rect 14196 45164 14206 45220
rect 16594 45164 16604 45220
rect 16660 45164 17724 45220
rect 17780 45164 17790 45220
rect 40674 45164 40684 45220
rect 40740 45164 42252 45220
rect 42308 45164 42318 45220
rect 44258 45164 44268 45220
rect 44324 45164 44940 45220
rect 44996 45164 45006 45220
rect 45714 45164 45724 45220
rect 45780 45164 52108 45220
rect 52164 45164 53228 45220
rect 53284 45164 53294 45220
rect 15586 45052 15596 45108
rect 15652 45052 18956 45108
rect 19012 45052 19022 45108
rect 19282 45052 19292 45108
rect 19348 45052 20188 45108
rect 20244 45052 20748 45108
rect 20804 45052 21980 45108
rect 22036 45052 22046 45108
rect 26786 45052 26796 45108
rect 26852 45052 29260 45108
rect 29316 45052 30436 45108
rect 36306 45052 36316 45108
rect 36372 45052 39564 45108
rect 39620 45052 39630 45108
rect 39788 45052 40236 45108
rect 40292 45052 41580 45108
rect 41636 45052 41646 45108
rect 41794 45052 41804 45108
rect 41860 45052 42588 45108
rect 42644 45052 42924 45108
rect 42980 45052 42990 45108
rect 44146 45052 44156 45108
rect 44212 45052 51212 45108
rect 51268 45052 51278 45108
rect 51762 45052 51772 45108
rect 51828 45052 51996 45108
rect 52052 45052 52062 45108
rect 30380 44996 30436 45052
rect 39788 44996 39844 45052
rect 11554 44940 11564 44996
rect 11620 44940 12460 44996
rect 12516 44940 15708 44996
rect 15764 44940 20636 44996
rect 20692 44940 21308 44996
rect 21364 44940 21374 44996
rect 30370 44940 30380 44996
rect 30436 44940 30446 44996
rect 36194 44940 36204 44996
rect 36260 44940 37548 44996
rect 37604 44940 38108 44996
rect 38164 44940 39844 44996
rect 40338 44940 40348 44996
rect 40404 44940 41356 44996
rect 41412 44940 41422 44996
rect 43362 44940 43372 44996
rect 43428 44940 47628 44996
rect 47684 44940 47694 44996
rect 51538 44940 51548 44996
rect 51604 44940 52108 44996
rect 52164 44940 52174 44996
rect 14242 44828 14252 44884
rect 14308 44828 16492 44884
rect 16548 44828 18956 44884
rect 19012 44828 19022 44884
rect 20402 44828 20412 44884
rect 20468 44828 21532 44884
rect 21588 44828 21598 44884
rect 40226 44828 40236 44884
rect 40292 44828 43708 44884
rect 44370 44828 44380 44884
rect 44436 44828 48412 44884
rect 48468 44828 52780 44884
rect 52836 44828 52846 44884
rect 20412 44772 20468 44828
rect 43652 44772 43708 44828
rect 15586 44716 15596 44772
rect 15652 44716 20468 44772
rect 40338 44716 40348 44772
rect 40404 44716 41020 44772
rect 41076 44716 41086 44772
rect 43652 44716 49980 44772
rect 50036 44716 52892 44772
rect 52948 44716 52958 44772
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 13794 44604 13804 44660
rect 13860 44604 17612 44660
rect 17668 44604 18060 44660
rect 18116 44604 18126 44660
rect 41682 44604 41692 44660
rect 41748 44604 47740 44660
rect 47796 44604 48188 44660
rect 48244 44604 48254 44660
rect 16818 44492 16828 44548
rect 16884 44492 19964 44548
rect 20020 44492 20524 44548
rect 20580 44492 21308 44548
rect 21364 44492 21374 44548
rect 43698 44492 43708 44548
rect 43764 44492 50092 44548
rect 50148 44492 52668 44548
rect 52724 44492 52734 44548
rect 7970 44380 7980 44436
rect 8036 44380 8652 44436
rect 8708 44380 9660 44436
rect 9716 44380 10220 44436
rect 10276 44380 10286 44436
rect 10546 44380 10556 44436
rect 10612 44380 12124 44436
rect 12180 44380 13244 44436
rect 13300 44380 15372 44436
rect 15428 44380 15438 44436
rect 45266 44380 45276 44436
rect 45332 44380 48860 44436
rect 48916 44380 49532 44436
rect 49588 44380 51772 44436
rect 51828 44380 51838 44436
rect 14914 44268 14924 44324
rect 14980 44268 15484 44324
rect 15540 44268 15550 44324
rect 16370 44268 16380 44324
rect 16436 44268 17052 44324
rect 17108 44268 17118 44324
rect 19618 44268 19628 44324
rect 19684 44268 20412 44324
rect 20468 44268 21868 44324
rect 21924 44268 21934 44324
rect 39666 44268 39676 44324
rect 39732 44268 40572 44324
rect 40628 44268 40638 44324
rect 49746 44268 49756 44324
rect 49812 44268 50204 44324
rect 50260 44268 50270 44324
rect 9762 44156 9772 44212
rect 9828 44156 11340 44212
rect 11396 44156 11406 44212
rect 12114 44156 12124 44212
rect 12180 44156 13356 44212
rect 13412 44156 13422 44212
rect 17826 44156 17836 44212
rect 17892 44156 22092 44212
rect 22148 44156 23436 44212
rect 23492 44156 23502 44212
rect 36306 44156 36316 44212
rect 36372 44156 37548 44212
rect 37604 44156 37614 44212
rect 38210 44156 38220 44212
rect 38276 44156 39116 44212
rect 39172 44156 40236 44212
rect 40292 44156 40302 44212
rect 42802 44156 42812 44212
rect 42868 44156 44156 44212
rect 44212 44156 44222 44212
rect 2034 44044 2044 44100
rect 2100 44044 7084 44100
rect 7140 44044 7644 44100
rect 7700 44044 7710 44100
rect 8306 44044 8316 44100
rect 8372 44044 8764 44100
rect 8820 44044 10108 44100
rect 10164 44044 10174 44100
rect 12674 44044 12684 44100
rect 12740 44044 13468 44100
rect 13524 44044 16268 44100
rect 16324 44044 16334 44100
rect 20738 44044 20748 44100
rect 20804 44044 22204 44100
rect 22260 44044 22270 44100
rect 41346 44044 41356 44100
rect 41412 44044 41916 44100
rect 41972 44044 42924 44100
rect 42980 44044 42990 44100
rect 49074 44044 49084 44100
rect 49140 44044 50988 44100
rect 51044 44044 51054 44100
rect 41468 43932 42028 43988
rect 42084 43932 42094 43988
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 0 43764 800 43792
rect 0 43708 1708 43764
rect 1764 43708 2492 43764
rect 2548 43708 2558 43764
rect 9986 43708 9996 43764
rect 10052 43708 10062 43764
rect 13458 43708 13468 43764
rect 13524 43708 15036 43764
rect 15092 43708 15102 43764
rect 21634 43708 21644 43764
rect 21700 43708 22540 43764
rect 22596 43708 24332 43764
rect 24388 43708 24398 43764
rect 40674 43708 40684 43764
rect 40740 43708 40908 43764
rect 40964 43708 40974 43764
rect 0 43680 800 43708
rect 9996 43540 10052 43708
rect 41468 43652 41524 43932
rect 50546 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50830 43932
rect 43026 43708 43036 43764
rect 43092 43708 43102 43764
rect 44594 43708 44604 43764
rect 44660 43708 45052 43764
rect 45108 43708 45118 43764
rect 49522 43708 49532 43764
rect 49588 43708 50092 43764
rect 50148 43708 50158 43764
rect 42690 43652 42700 43708
rect 42756 43652 42766 43708
rect 43036 43652 43092 43708
rect 44146 43652 44156 43708
rect 44212 43652 44222 43708
rect 11330 43596 11340 43652
rect 11396 43596 12124 43652
rect 12180 43596 12684 43652
rect 12740 43596 12750 43652
rect 40114 43596 40124 43652
rect 40180 43596 40348 43652
rect 40404 43596 40414 43652
rect 40572 43596 41244 43652
rect 41300 43596 41524 43652
rect 41580 43596 42756 43652
rect 43036 43596 44212 43652
rect 45826 43596 45836 43652
rect 45892 43596 46956 43652
rect 47012 43596 47022 43652
rect 49970 43596 49980 43652
rect 50036 43596 51548 43652
rect 51604 43596 53564 43652
rect 53620 43596 53630 43652
rect 40572 43540 40628 43596
rect 41580 43540 41636 43596
rect 43036 43540 43092 43596
rect 7186 43484 7196 43540
rect 7252 43484 8428 43540
rect 8484 43484 8876 43540
rect 8932 43484 10052 43540
rect 35858 43484 35868 43540
rect 35924 43484 37324 43540
rect 37380 43484 37390 43540
rect 37650 43484 37660 43540
rect 37716 43484 40628 43540
rect 41346 43484 41356 43540
rect 41412 43484 41580 43540
rect 41636 43484 41646 43540
rect 41794 43484 41804 43540
rect 41860 43484 43092 43540
rect 44258 43484 44268 43540
rect 44324 43484 45612 43540
rect 45668 43484 46060 43540
rect 46116 43484 46126 43540
rect 47954 43484 47964 43540
rect 48020 43484 49308 43540
rect 49364 43484 49374 43540
rect 51202 43484 51212 43540
rect 51268 43484 51884 43540
rect 51940 43484 51950 43540
rect 8530 43372 8540 43428
rect 8596 43372 12796 43428
rect 12852 43372 14140 43428
rect 14196 43372 15260 43428
rect 15316 43372 15326 43428
rect 16258 43372 16268 43428
rect 16324 43372 19516 43428
rect 19572 43372 19582 43428
rect 33506 43372 33516 43428
rect 33572 43372 34300 43428
rect 34356 43372 34366 43428
rect 39778 43372 39788 43428
rect 39844 43372 45948 43428
rect 46004 43372 46014 43428
rect 46498 43372 46508 43428
rect 46564 43372 48748 43428
rect 48804 43372 52556 43428
rect 52612 43372 52622 43428
rect 7074 43260 7084 43316
rect 7140 43260 7868 43316
rect 7924 43260 7934 43316
rect 21410 43260 21420 43316
rect 21476 43260 22764 43316
rect 22820 43260 23436 43316
rect 23492 43260 23502 43316
rect 34626 43260 34636 43316
rect 34692 43260 37436 43316
rect 37492 43260 37502 43316
rect 39106 43260 39116 43316
rect 39172 43260 40012 43316
rect 40068 43260 40078 43316
rect 44044 43260 50428 43316
rect 50484 43260 51548 43316
rect 51604 43260 51614 43316
rect 10322 43148 10332 43204
rect 10388 43148 10668 43204
rect 10724 43148 10734 43204
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 44044 43092 44100 43260
rect 46274 43148 46284 43204
rect 46340 43148 48748 43204
rect 48804 43148 48814 43204
rect 32162 43036 32172 43092
rect 32228 43036 34748 43092
rect 34804 43036 34814 43092
rect 42130 43036 42140 43092
rect 42196 43036 44100 43092
rect 44156 43036 50876 43092
rect 50932 43036 51324 43092
rect 51380 43036 51390 43092
rect 44156 42980 44212 43036
rect 33618 42924 33628 42980
rect 33684 42924 34412 42980
rect 34468 42924 34478 42980
rect 37202 42924 37212 42980
rect 37268 42924 39004 42980
rect 39060 42924 39070 42980
rect 41122 42924 41132 42980
rect 41188 42924 44212 42980
rect 44370 42924 44380 42980
rect 44436 42924 45388 42980
rect 45444 42924 45454 42980
rect 11442 42812 11452 42868
rect 11508 42812 20972 42868
rect 21028 42812 21038 42868
rect 52882 42812 52892 42868
rect 52948 42812 53900 42868
rect 53956 42812 53966 42868
rect 9090 42700 9100 42756
rect 9156 42700 9436 42756
rect 9492 42700 10108 42756
rect 10164 42700 11676 42756
rect 11732 42700 11742 42756
rect 37202 42700 37212 42756
rect 37268 42700 37772 42756
rect 37828 42700 37838 42756
rect 41794 42700 41804 42756
rect 41860 42700 42812 42756
rect 42868 42700 42878 42756
rect 47170 42700 47180 42756
rect 47236 42700 49532 42756
rect 49588 42700 49598 42756
rect 51874 42700 51884 42756
rect 51940 42700 52444 42756
rect 52500 42700 54348 42756
rect 54404 42700 54414 42756
rect 7298 42588 7308 42644
rect 7364 42588 8204 42644
rect 8260 42588 8270 42644
rect 10434 42588 10444 42644
rect 10500 42588 10892 42644
rect 10948 42588 11732 42644
rect 30146 42588 30156 42644
rect 30212 42588 30492 42644
rect 30548 42588 31276 42644
rect 31332 42588 31342 42644
rect 31714 42588 31724 42644
rect 31780 42588 33292 42644
rect 33348 42588 35308 42644
rect 35364 42588 35374 42644
rect 39330 42588 39340 42644
rect 39396 42588 40348 42644
rect 40404 42588 41132 42644
rect 41188 42588 41198 42644
rect 42018 42588 42028 42644
rect 42084 42588 42700 42644
rect 42756 42588 42766 42644
rect 11676 42532 11732 42588
rect 2706 42476 2716 42532
rect 2772 42476 7532 42532
rect 7588 42476 7598 42532
rect 9202 42476 9212 42532
rect 9268 42476 10332 42532
rect 10388 42476 10398 42532
rect 11666 42476 11676 42532
rect 11732 42476 13692 42532
rect 13748 42476 13758 42532
rect 30370 42476 30380 42532
rect 30436 42476 31948 42532
rect 32004 42476 32014 42532
rect 33394 42476 33404 42532
rect 33460 42476 35196 42532
rect 35252 42476 35262 42532
rect 41682 42476 41692 42532
rect 41748 42476 43820 42532
rect 43876 42476 43886 42532
rect 45154 42476 45164 42532
rect 45220 42476 45836 42532
rect 45892 42476 47964 42532
rect 48020 42476 48860 42532
rect 48916 42476 48926 42532
rect 0 42420 800 42448
rect 0 42364 2380 42420
rect 2436 42364 2446 42420
rect 28690 42364 28700 42420
rect 28756 42364 30044 42420
rect 30100 42364 30716 42420
rect 30772 42364 31948 42420
rect 33618 42364 33628 42420
rect 33684 42364 34188 42420
rect 34244 42364 37548 42420
rect 37604 42364 37614 42420
rect 39666 42364 39676 42420
rect 39732 42364 40124 42420
rect 40180 42364 40190 42420
rect 42690 42364 42700 42420
rect 42756 42364 48972 42420
rect 49028 42364 49038 42420
rect 0 42336 800 42364
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 31892 42308 31948 42364
rect 50546 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50830 42364
rect 2034 42252 2044 42308
rect 2100 42252 4396 42308
rect 4452 42252 4462 42308
rect 8530 42252 8540 42308
rect 8596 42252 13468 42308
rect 13524 42252 14588 42308
rect 14644 42252 14654 42308
rect 19506 42252 19516 42308
rect 19572 42252 19582 42308
rect 31892 42252 39900 42308
rect 39956 42252 39966 42308
rect 19516 42196 19572 42252
rect 12908 42140 13580 42196
rect 13636 42140 16604 42196
rect 16660 42140 16670 42196
rect 19516 42140 19964 42196
rect 20020 42140 20030 42196
rect 40226 42140 40236 42196
rect 40292 42140 41244 42196
rect 41300 42140 43708 42196
rect 44818 42140 44828 42196
rect 44884 42140 45724 42196
rect 45780 42140 45790 42196
rect 12908 42084 12964 42140
rect 43652 42084 43708 42140
rect 10994 42028 11004 42084
rect 11060 42028 11900 42084
rect 11956 42028 11966 42084
rect 12898 42028 12908 42084
rect 12964 42028 12974 42084
rect 13234 42028 13244 42084
rect 13300 42028 14476 42084
rect 14532 42028 15372 42084
rect 15428 42028 16268 42084
rect 16324 42028 16334 42084
rect 41010 42028 41020 42084
rect 41076 42028 41804 42084
rect 41860 42028 42476 42084
rect 42532 42028 42542 42084
rect 42802 42028 42812 42084
rect 42868 42028 43372 42084
rect 43428 42028 43438 42084
rect 43652 42028 48076 42084
rect 48132 42028 48142 42084
rect 1698 41916 1708 41972
rect 1764 41916 3612 41972
rect 3668 41916 3678 41972
rect 8372 41916 8988 41972
rect 9044 41916 9996 41972
rect 10052 41916 10062 41972
rect 11442 41916 11452 41972
rect 11508 41916 15596 41972
rect 15652 41916 16492 41972
rect 16548 41916 16558 41972
rect 20626 41916 20636 41972
rect 20692 41916 22204 41972
rect 22260 41916 23324 41972
rect 23380 41916 23390 41972
rect 23650 41916 23660 41972
rect 23716 41916 23726 41972
rect 32498 41916 32508 41972
rect 32564 41916 35084 41972
rect 35140 41916 35150 41972
rect 43138 41916 43148 41972
rect 43204 41916 43820 41972
rect 43876 41916 43886 41972
rect 45266 41916 45276 41972
rect 45332 41916 45948 41972
rect 46004 41916 46508 41972
rect 46564 41916 46574 41972
rect 48290 41916 48300 41972
rect 48356 41916 53452 41972
rect 53508 41916 53788 41972
rect 53844 41916 53854 41972
rect 2370 41804 2380 41860
rect 2436 41804 3164 41860
rect 3220 41804 3230 41860
rect 0 41748 800 41776
rect 8372 41748 8428 41916
rect 23660 41860 23716 41916
rect 13122 41804 13132 41860
rect 13188 41804 13468 41860
rect 13524 41804 13534 41860
rect 21186 41804 21196 41860
rect 21252 41804 21980 41860
rect 22036 41804 22046 41860
rect 22642 41804 22652 41860
rect 22708 41804 23716 41860
rect 36530 41804 36540 41860
rect 36596 41804 42364 41860
rect 42420 41804 42430 41860
rect 43698 41804 43708 41860
rect 43764 41804 45052 41860
rect 45108 41804 45118 41860
rect 49634 41804 49644 41860
rect 49700 41804 50092 41860
rect 50148 41804 50158 41860
rect 50754 41804 50764 41860
rect 50820 41804 54236 41860
rect 54292 41804 54684 41860
rect 54740 41804 54750 41860
rect 0 41692 1708 41748
rect 1764 41692 2940 41748
rect 2996 41692 3006 41748
rect 3378 41692 3388 41748
rect 3444 41692 4396 41748
rect 4452 41692 4462 41748
rect 5954 41692 5964 41748
rect 6020 41692 7644 41748
rect 7700 41692 8428 41748
rect 42466 41692 42476 41748
rect 42532 41692 43596 41748
rect 43652 41692 43662 41748
rect 0 41664 800 41692
rect 2034 41580 2044 41636
rect 2100 41580 4284 41636
rect 4340 41580 4350 41636
rect 37874 41580 37884 41636
rect 37940 41580 39788 41636
rect 39844 41580 39854 41636
rect 44706 41580 44716 41636
rect 44772 41580 48412 41636
rect 48468 41580 48478 41636
rect 4284 41412 4340 41580
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 12786 41468 12796 41524
rect 12852 41468 13244 41524
rect 13300 41468 13310 41524
rect 4284 41356 5292 41412
rect 5348 41356 5358 41412
rect 16594 41356 16604 41412
rect 16660 41356 19964 41412
rect 20020 41356 20030 41412
rect 29810 41356 29820 41412
rect 29876 41356 32508 41412
rect 32564 41356 32574 41412
rect 42354 41356 42364 41412
rect 42420 41356 43708 41412
rect 44146 41356 44156 41412
rect 44212 41356 45724 41412
rect 45780 41356 46620 41412
rect 46676 41356 46686 41412
rect 51650 41356 51660 41412
rect 51716 41356 53004 41412
rect 53060 41356 53564 41412
rect 53620 41356 53630 41412
rect 43652 41300 43708 41356
rect 5058 41244 5068 41300
rect 5124 41244 6412 41300
rect 6468 41244 8876 41300
rect 8932 41244 9548 41300
rect 9604 41244 9614 41300
rect 10658 41244 10668 41300
rect 10724 41244 13580 41300
rect 13636 41244 14028 41300
rect 14084 41244 14094 41300
rect 16370 41244 16380 41300
rect 16436 41244 18060 41300
rect 18116 41244 18126 41300
rect 31042 41244 31052 41300
rect 31108 41244 36540 41300
rect 36596 41244 36606 41300
rect 37762 41244 37772 41300
rect 37828 41244 39452 41300
rect 39508 41244 39518 41300
rect 43652 41244 45836 41300
rect 45892 41244 45902 41300
rect 2258 41132 2268 41188
rect 2324 41132 6972 41188
rect 7028 41132 7038 41188
rect 17490 41132 17500 41188
rect 17556 41132 18732 41188
rect 18788 41132 19292 41188
rect 19348 41132 19358 41188
rect 19506 41132 19516 41188
rect 19572 41132 23100 41188
rect 23156 41132 23166 41188
rect 29698 41132 29708 41188
rect 29764 41132 32172 41188
rect 32228 41132 32238 41188
rect 36194 41132 36204 41188
rect 36260 41132 37324 41188
rect 37380 41132 38332 41188
rect 38388 41132 38398 41188
rect 51426 41132 51436 41188
rect 51492 41132 52668 41188
rect 52724 41132 52734 41188
rect 0 41076 800 41104
rect 0 41020 2380 41076
rect 2436 41020 2446 41076
rect 2706 41020 2716 41076
rect 2772 41020 7196 41076
rect 7252 41020 7262 41076
rect 12562 41020 12572 41076
rect 12628 41020 13804 41076
rect 13860 41020 14588 41076
rect 14644 41020 14654 41076
rect 16370 41020 16380 41076
rect 16436 41020 17948 41076
rect 18004 41020 21420 41076
rect 21476 41020 21486 41076
rect 22306 41020 22316 41076
rect 22372 41020 23660 41076
rect 23716 41020 23726 41076
rect 37538 41020 37548 41076
rect 37604 41020 38556 41076
rect 38612 41020 38622 41076
rect 41356 41020 43708 41076
rect 49298 41020 49308 41076
rect 49364 41020 50652 41076
rect 50708 41020 50718 41076
rect 0 40992 800 41020
rect 21420 40964 21476 41020
rect 41356 40964 41412 41020
rect 43652 40964 43708 41020
rect 7970 40908 7980 40964
rect 8036 40908 12796 40964
rect 12852 40908 12862 40964
rect 14242 40908 14252 40964
rect 14308 40908 16156 40964
rect 16212 40908 16716 40964
rect 16772 40908 16782 40964
rect 19068 40908 19852 40964
rect 19908 40908 19918 40964
rect 21420 40908 22428 40964
rect 22484 40908 22494 40964
rect 36418 40908 36428 40964
rect 36484 40908 36764 40964
rect 36820 40908 36830 40964
rect 37874 40908 37884 40964
rect 37940 40908 39004 40964
rect 39060 40908 40124 40964
rect 40180 40908 40190 40964
rect 41346 40908 41356 40964
rect 41412 40908 41422 40964
rect 42578 40908 42588 40964
rect 42644 40908 42654 40964
rect 43652 40908 48468 40964
rect 49074 40908 49084 40964
rect 49140 40908 51660 40964
rect 51716 40908 51726 40964
rect 51986 40908 51996 40964
rect 52052 40908 52892 40964
rect 52948 40908 52958 40964
rect 19068 40852 19124 40908
rect 40124 40852 40180 40908
rect 42588 40852 42644 40908
rect 48412 40852 48468 40908
rect 18274 40796 18284 40852
rect 18340 40796 19068 40852
rect 19124 40796 19134 40852
rect 28354 40796 28364 40852
rect 28420 40796 29708 40852
rect 29764 40796 29774 40852
rect 40124 40796 41580 40852
rect 41636 40796 41646 40852
rect 42588 40796 44268 40852
rect 44324 40796 44334 40852
rect 48412 40796 49532 40852
rect 49588 40796 49598 40852
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 50546 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50830 40796
rect 31154 40684 31164 40740
rect 31220 40684 31836 40740
rect 31892 40684 40348 40740
rect 40404 40684 40414 40740
rect 41682 40684 41692 40740
rect 41748 40684 43036 40740
rect 43092 40684 43102 40740
rect 43362 40684 43372 40740
rect 43428 40684 44716 40740
rect 44772 40684 44782 40740
rect 5282 40572 5292 40628
rect 5348 40572 5852 40628
rect 5908 40572 5918 40628
rect 9762 40572 9772 40628
rect 9828 40572 11004 40628
rect 11060 40572 11070 40628
rect 11890 40572 11900 40628
rect 11956 40572 16604 40628
rect 16660 40572 16670 40628
rect 18386 40572 18396 40628
rect 18452 40572 20972 40628
rect 21028 40572 21644 40628
rect 21700 40572 21710 40628
rect 39778 40572 39788 40628
rect 39844 40572 40460 40628
rect 40516 40572 40526 40628
rect 43586 40572 43596 40628
rect 43652 40572 44156 40628
rect 44212 40572 44222 40628
rect 45938 40572 45948 40628
rect 46004 40572 47404 40628
rect 47460 40572 49308 40628
rect 49364 40572 49374 40628
rect 7186 40460 7196 40516
rect 7252 40460 7868 40516
rect 7924 40460 7934 40516
rect 10098 40460 10108 40516
rect 10164 40460 13020 40516
rect 13076 40460 13086 40516
rect 13244 40460 19628 40516
rect 19684 40460 19694 40516
rect 19842 40460 19852 40516
rect 19908 40460 21532 40516
rect 21588 40460 23548 40516
rect 23604 40460 23614 40516
rect 31042 40460 31052 40516
rect 31108 40460 35084 40516
rect 35140 40460 35150 40516
rect 36428 40460 46284 40516
rect 46340 40460 46350 40516
rect 0 40404 800 40432
rect 13244 40404 13300 40460
rect 19628 40404 19684 40460
rect 36428 40404 36484 40460
rect 0 40348 1708 40404
rect 1764 40348 1774 40404
rect 10322 40348 10332 40404
rect 10388 40348 11452 40404
rect 11508 40348 11900 40404
rect 11956 40348 11966 40404
rect 12226 40348 12236 40404
rect 12292 40348 13300 40404
rect 14690 40348 14700 40404
rect 14756 40348 17388 40404
rect 17444 40348 17454 40404
rect 19058 40348 19068 40404
rect 19124 40348 19404 40404
rect 19460 40348 19470 40404
rect 19628 40348 20188 40404
rect 20244 40348 20254 40404
rect 22642 40348 22652 40404
rect 22708 40348 23436 40404
rect 23492 40348 23502 40404
rect 30370 40348 30380 40404
rect 30436 40348 31500 40404
rect 31556 40348 31566 40404
rect 33954 40348 33964 40404
rect 34020 40348 36484 40404
rect 37650 40348 37660 40404
rect 37716 40348 37726 40404
rect 42354 40348 42364 40404
rect 42420 40348 43260 40404
rect 43316 40348 44604 40404
rect 44660 40348 44670 40404
rect 50194 40348 50204 40404
rect 50260 40348 51100 40404
rect 51156 40348 51772 40404
rect 51828 40348 52892 40404
rect 52948 40348 52958 40404
rect 0 40320 800 40348
rect 2594 40236 2604 40292
rect 2660 40236 3276 40292
rect 3332 40236 3342 40292
rect 28018 40236 28028 40292
rect 28084 40236 28812 40292
rect 28868 40236 37100 40292
rect 37156 40236 37166 40292
rect 37660 40180 37716 40348
rect 40338 40236 40348 40292
rect 40404 40236 44044 40292
rect 44100 40236 44110 40292
rect 44930 40236 44940 40292
rect 44996 40236 49308 40292
rect 49364 40236 49868 40292
rect 49924 40236 49934 40292
rect 5058 40124 5068 40180
rect 5124 40124 5628 40180
rect 5684 40124 5694 40180
rect 28690 40124 28700 40180
rect 28756 40124 30380 40180
rect 30436 40124 30446 40180
rect 37660 40124 41132 40180
rect 41188 40124 41198 40180
rect 42130 40124 42140 40180
rect 42196 40124 42700 40180
rect 42756 40124 42766 40180
rect 37660 40068 37716 40124
rect 36530 40012 36540 40068
rect 36596 40012 37716 40068
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 46946 39900 46956 39956
rect 47012 39900 54460 39956
rect 54516 39900 54526 39956
rect 2930 39788 2940 39844
rect 2996 39788 4060 39844
rect 4116 39788 4396 39844
rect 4452 39788 11116 39844
rect 11172 39788 11182 39844
rect 18722 39788 18732 39844
rect 18788 39788 19180 39844
rect 19236 39788 19246 39844
rect 37090 39788 37100 39844
rect 37156 39788 40124 39844
rect 40180 39788 40190 39844
rect 0 39732 800 39760
rect 0 39676 1708 39732
rect 1764 39676 1774 39732
rect 4722 39676 4732 39732
rect 4788 39676 5740 39732
rect 5796 39676 5806 39732
rect 6514 39676 6524 39732
rect 6580 39676 7644 39732
rect 7700 39676 7710 39732
rect 17714 39676 17724 39732
rect 17780 39676 18844 39732
rect 18900 39676 18910 39732
rect 36642 39676 36652 39732
rect 36708 39676 40684 39732
rect 40740 39676 41244 39732
rect 41300 39676 41310 39732
rect 0 39648 800 39676
rect 2258 39564 2268 39620
rect 2324 39564 3724 39620
rect 3780 39564 7140 39620
rect 7084 39508 7140 39564
rect 8372 39564 8652 39620
rect 8708 39564 9660 39620
rect 9716 39564 9726 39620
rect 13010 39564 13020 39620
rect 13076 39564 14588 39620
rect 14644 39564 14654 39620
rect 21970 39564 21980 39620
rect 22036 39564 23324 39620
rect 23380 39564 23390 39620
rect 28690 39564 28700 39620
rect 28756 39564 29484 39620
rect 29540 39564 29550 39620
rect 31938 39564 31948 39620
rect 32004 39564 32620 39620
rect 32676 39564 32686 39620
rect 36978 39564 36988 39620
rect 37044 39564 39676 39620
rect 39732 39564 46284 39620
rect 46340 39564 48860 39620
rect 48916 39564 48926 39620
rect 8372 39508 8428 39564
rect 4834 39452 4844 39508
rect 4900 39452 5852 39508
rect 5908 39452 6412 39508
rect 6468 39452 6860 39508
rect 6916 39452 6926 39508
rect 7074 39452 7084 39508
rect 7140 39452 8428 39508
rect 10770 39452 10780 39508
rect 10836 39452 12012 39508
rect 12068 39452 12078 39508
rect 16818 39452 16828 39508
rect 16884 39452 18620 39508
rect 18676 39452 18686 39508
rect 21858 39452 21868 39508
rect 21924 39452 22540 39508
rect 22596 39452 23660 39508
rect 23716 39452 23726 39508
rect 35858 39452 35868 39508
rect 35924 39452 36540 39508
rect 36596 39452 36606 39508
rect 42242 39452 42252 39508
rect 42308 39452 43148 39508
rect 43204 39452 43214 39508
rect 8306 39340 8316 39396
rect 8372 39340 8988 39396
rect 9044 39340 10556 39396
rect 10612 39340 10622 39396
rect 14690 39340 14700 39396
rect 14756 39340 15372 39396
rect 15428 39340 15438 39396
rect 18834 39340 18844 39396
rect 18900 39340 22316 39396
rect 22372 39340 23100 39396
rect 23156 39340 23166 39396
rect 35186 39340 35196 39396
rect 35252 39340 39116 39396
rect 39172 39340 39182 39396
rect 39778 39340 39788 39396
rect 39844 39340 41468 39396
rect 41524 39340 41534 39396
rect 45714 39340 45724 39396
rect 45780 39340 45948 39396
rect 46004 39340 51100 39396
rect 51156 39340 51166 39396
rect 54450 39340 54460 39396
rect 54516 39340 55468 39396
rect 55524 39340 55534 39396
rect 3042 39228 3052 39284
rect 3108 39228 7308 39284
rect 7364 39228 7374 39284
rect 8754 39228 8764 39284
rect 8820 39228 18172 39284
rect 18228 39228 19180 39284
rect 19236 39228 19246 39284
rect 33394 39228 33404 39284
rect 33460 39228 46732 39284
rect 46788 39228 47292 39284
rect 47348 39228 47358 39284
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 50546 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50830 39228
rect 2706 39116 2716 39172
rect 2772 39116 9884 39172
rect 9940 39116 9950 39172
rect 17938 39116 17948 39172
rect 18004 39116 18620 39172
rect 18676 39116 18686 39172
rect 29922 39116 29932 39172
rect 29988 39116 30380 39172
rect 30436 39116 30446 39172
rect 42242 39116 42252 39172
rect 42308 39116 42318 39172
rect 0 39060 800 39088
rect 42252 39060 42308 39116
rect 0 39004 1708 39060
rect 1764 39004 1774 39060
rect 2034 39004 2044 39060
rect 2100 39004 3724 39060
rect 3780 39004 3790 39060
rect 4946 39004 4956 39060
rect 5012 39004 5022 39060
rect 13682 39004 13692 39060
rect 13748 39004 14364 39060
rect 14420 39004 14430 39060
rect 28690 39004 28700 39060
rect 28756 39004 29372 39060
rect 29428 39004 42924 39060
rect 42980 39004 44828 39060
rect 44884 39004 46060 39060
rect 46116 39004 46126 39060
rect 46722 39004 46732 39060
rect 46788 39004 52108 39060
rect 52164 39004 52174 39060
rect 0 38976 800 39004
rect 4956 38836 5012 39004
rect 24322 38892 24332 38948
rect 24388 38892 25452 38948
rect 25508 38892 25518 38948
rect 28802 38892 28812 38948
rect 28868 38892 29820 38948
rect 29876 38892 36652 38948
rect 36708 38892 36718 38948
rect 46498 38892 46508 38948
rect 46564 38892 47068 38948
rect 47124 38892 47134 38948
rect 49410 38892 49420 38948
rect 49476 38892 51548 38948
rect 51604 38892 51614 38948
rect 4050 38780 4060 38836
rect 4116 38780 4284 38836
rect 4340 38780 5852 38836
rect 5908 38780 5918 38836
rect 12002 38780 12012 38836
rect 12068 38780 12796 38836
rect 12852 38780 13916 38836
rect 13972 38780 14588 38836
rect 14644 38780 14654 38836
rect 40002 38780 40012 38836
rect 40068 38780 40908 38836
rect 40964 38780 41916 38836
rect 41972 38780 41982 38836
rect 45826 38780 45836 38836
rect 45892 38780 46732 38836
rect 46788 38780 46798 38836
rect 54226 38780 54236 38836
rect 54292 38780 55132 38836
rect 55188 38780 55198 38836
rect 3490 38668 3500 38724
rect 3556 38668 4844 38724
rect 4900 38668 4910 38724
rect 5058 38668 5068 38724
rect 5124 38668 5740 38724
rect 5796 38668 6748 38724
rect 6804 38668 6814 38724
rect 10882 38668 10892 38724
rect 10948 38668 11900 38724
rect 11956 38668 11966 38724
rect 13794 38668 13804 38724
rect 13860 38668 13870 38724
rect 16034 38668 16044 38724
rect 16100 38668 18508 38724
rect 18564 38668 19852 38724
rect 19908 38668 19918 38724
rect 20402 38668 20412 38724
rect 20468 38668 23548 38724
rect 23604 38668 23614 38724
rect 36530 38668 36540 38724
rect 36596 38668 37772 38724
rect 37828 38668 37838 38724
rect 41570 38668 41580 38724
rect 41636 38668 42252 38724
rect 42308 38668 42318 38724
rect 47730 38668 47740 38724
rect 47796 38668 48748 38724
rect 48804 38668 48814 38724
rect 51090 38668 51100 38724
rect 51156 38668 51436 38724
rect 51492 38668 51884 38724
rect 51940 38668 51950 38724
rect 13804 38612 13860 38668
rect 3154 38556 3164 38612
rect 3220 38556 4732 38612
rect 4788 38556 4798 38612
rect 9986 38556 9996 38612
rect 10052 38556 13860 38612
rect 55794 38556 55804 38612
rect 55860 38556 57036 38612
rect 57092 38556 57102 38612
rect 16258 38444 16268 38500
rect 16324 38444 19292 38500
rect 19348 38444 20076 38500
rect 20132 38444 20142 38500
rect 46386 38444 46396 38500
rect 46452 38444 48300 38500
rect 48356 38444 48366 38500
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 40226 38332 40236 38388
rect 40292 38332 43596 38388
rect 43652 38332 43662 38388
rect 46610 38332 46620 38388
rect 46676 38332 53788 38388
rect 53844 38332 54684 38388
rect 54740 38332 54750 38388
rect 33506 38220 33516 38276
rect 33572 38220 33796 38276
rect 39330 38220 39340 38276
rect 39396 38220 39900 38276
rect 39956 38220 45724 38276
rect 45780 38220 45790 38276
rect 50194 38220 50204 38276
rect 50260 38220 51212 38276
rect 51268 38220 51278 38276
rect 55122 38220 55132 38276
rect 55188 38220 56028 38276
rect 56084 38220 56094 38276
rect 33740 38164 33796 38220
rect 2146 38108 2156 38164
rect 2212 38108 2828 38164
rect 2884 38108 2894 38164
rect 10098 38108 10108 38164
rect 10164 38108 11116 38164
rect 11172 38108 11182 38164
rect 20850 38108 20860 38164
rect 20916 38108 21980 38164
rect 22036 38108 22046 38164
rect 33730 38108 33740 38164
rect 33796 38108 33806 38164
rect 37090 38108 37100 38164
rect 37156 38108 38444 38164
rect 38500 38108 40348 38164
rect 40404 38108 40414 38164
rect 49634 38108 49644 38164
rect 49700 38108 50316 38164
rect 50372 38108 50382 38164
rect 9650 37996 9660 38052
rect 9716 37996 24108 38052
rect 24164 37996 25004 38052
rect 25060 37996 25070 38052
rect 30930 37996 30940 38052
rect 30996 37996 33404 38052
rect 33460 37996 33470 38052
rect 40002 37996 40012 38052
rect 40068 37996 41580 38052
rect 41636 37996 41646 38052
rect 41794 37996 41804 38052
rect 41860 37996 42700 38052
rect 42756 37996 43484 38052
rect 43540 37996 43550 38052
rect 5058 37884 5068 37940
rect 5124 37884 9996 37940
rect 10052 37884 10062 37940
rect 33282 37884 33292 37940
rect 33348 37884 33964 37940
rect 34020 37884 34030 37940
rect 40226 37884 40236 37940
rect 40292 37884 40460 37940
rect 40516 37884 42476 37940
rect 42532 37884 42542 37940
rect 47394 37884 47404 37940
rect 47460 37884 49196 37940
rect 49252 37884 49262 37940
rect 49410 37884 49420 37940
rect 49476 37884 57820 37940
rect 57876 37884 57886 37940
rect 5068 37828 5124 37884
rect 2370 37772 2380 37828
rect 2436 37772 2940 37828
rect 2996 37772 5124 37828
rect 11106 37772 11116 37828
rect 11172 37772 15148 37828
rect 17378 37772 17388 37828
rect 17444 37772 23884 37828
rect 23940 37772 25228 37828
rect 25284 37772 25294 37828
rect 28578 37772 28588 37828
rect 28644 37772 29708 37828
rect 29764 37772 29774 37828
rect 33842 37772 33852 37828
rect 33908 37772 37212 37828
rect 37268 37772 37278 37828
rect 38612 37772 43820 37828
rect 43876 37772 43886 37828
rect 44034 37772 44044 37828
rect 44100 37772 44940 37828
rect 44996 37772 45500 37828
rect 45556 37772 45566 37828
rect 48514 37772 48524 37828
rect 48580 37772 50316 37828
rect 50372 37772 50382 37828
rect 56914 37772 56924 37828
rect 56980 37772 58044 37828
rect 58100 37772 58110 37828
rect 15092 37716 15148 37772
rect 38612 37716 38668 37772
rect 59200 37716 60000 37744
rect 2258 37660 2268 37716
rect 2324 37660 2716 37716
rect 2772 37660 2782 37716
rect 6514 37660 6524 37716
rect 6580 37660 7084 37716
rect 7140 37660 14756 37716
rect 15092 37660 17500 37716
rect 17556 37660 19628 37716
rect 19684 37660 19694 37716
rect 31938 37660 31948 37716
rect 32004 37660 38668 37716
rect 57474 37660 57484 37716
rect 57540 37660 60000 37716
rect 14700 37604 14756 37660
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 50546 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50830 37660
rect 59200 37632 60000 37660
rect 12226 37548 12236 37604
rect 12292 37548 14476 37604
rect 14532 37548 14542 37604
rect 14700 37548 16492 37604
rect 16548 37548 18060 37604
rect 18116 37548 18126 37604
rect 43362 37548 43372 37604
rect 43428 37548 44156 37604
rect 44212 37548 44828 37604
rect 44884 37548 44894 37604
rect 50988 37548 57820 37604
rect 57876 37548 57886 37604
rect 50988 37492 51044 37548
rect 13458 37436 13468 37492
rect 13524 37436 14588 37492
rect 14644 37436 14654 37492
rect 15092 37436 23212 37492
rect 23268 37436 23548 37492
rect 23604 37436 23614 37492
rect 29362 37436 29372 37492
rect 29428 37436 29932 37492
rect 29988 37436 30492 37492
rect 30548 37436 30940 37492
rect 30996 37436 31006 37492
rect 32050 37436 32060 37492
rect 32116 37436 32508 37492
rect 32564 37436 39788 37492
rect 39844 37436 39854 37492
rect 50194 37436 50204 37492
rect 50260 37436 51044 37492
rect 54450 37436 54460 37492
rect 54516 37436 55468 37492
rect 57138 37436 57148 37492
rect 57204 37436 57214 37492
rect 15092 37380 15148 37436
rect 55412 37380 55468 37436
rect 9650 37324 9660 37380
rect 9716 37324 9726 37380
rect 12450 37324 12460 37380
rect 12516 37324 15148 37380
rect 15810 37324 15820 37380
rect 15876 37324 16716 37380
rect 16772 37324 16782 37380
rect 28466 37324 28476 37380
rect 28532 37324 29260 37380
rect 29316 37324 29326 37380
rect 30818 37324 30828 37380
rect 30884 37324 32396 37380
rect 32452 37324 32462 37380
rect 33282 37324 33292 37380
rect 33348 37324 33628 37380
rect 33684 37324 34300 37380
rect 34356 37324 38332 37380
rect 38388 37324 39452 37380
rect 39508 37324 39518 37380
rect 47282 37324 47292 37380
rect 47348 37324 54572 37380
rect 54628 37324 54638 37380
rect 55412 37324 55804 37380
rect 55860 37324 56588 37380
rect 56644 37324 56654 37380
rect 9660 37156 9716 37324
rect 12338 37212 12348 37268
rect 12404 37212 13244 37268
rect 13300 37212 14028 37268
rect 14084 37212 16268 37268
rect 16324 37212 17612 37268
rect 17668 37212 17678 37268
rect 18162 37212 18172 37268
rect 18228 37212 19068 37268
rect 19124 37212 19134 37268
rect 20290 37212 20300 37268
rect 20356 37212 23324 37268
rect 23380 37212 23390 37268
rect 24434 37212 24444 37268
rect 24500 37212 25228 37268
rect 25284 37212 25294 37268
rect 33394 37212 33404 37268
rect 33460 37212 34524 37268
rect 34580 37212 34590 37268
rect 36306 37212 36316 37268
rect 36372 37212 37100 37268
rect 37156 37212 37166 37268
rect 46722 37212 46732 37268
rect 46788 37212 47180 37268
rect 47236 37212 47246 37268
rect 48290 37212 48300 37268
rect 48356 37212 50652 37268
rect 50708 37212 50718 37268
rect 9660 37100 9772 37156
rect 9828 37100 9838 37156
rect 11442 37100 11452 37156
rect 11508 37100 15820 37156
rect 15876 37100 15886 37156
rect 16370 37100 16380 37156
rect 16436 37100 17948 37156
rect 18004 37100 18014 37156
rect 43698 37100 43708 37156
rect 43764 37100 44716 37156
rect 44772 37100 44782 37156
rect 50306 37100 50316 37156
rect 50372 37100 54348 37156
rect 54404 37100 55356 37156
rect 55412 37100 55422 37156
rect 57148 37044 57204 37436
rect 59200 37044 60000 37072
rect 9650 36988 9660 37044
rect 9716 36988 10220 37044
rect 10276 36988 10286 37044
rect 15026 36988 15036 37044
rect 15092 36988 16156 37044
rect 16212 36988 17388 37044
rect 17444 36988 17454 37044
rect 23986 36988 23996 37044
rect 24052 36988 24556 37044
rect 24612 36988 25340 37044
rect 25396 36988 25788 37044
rect 25844 36988 25854 37044
rect 32722 36988 32732 37044
rect 32788 36988 34076 37044
rect 34132 36988 34142 37044
rect 42476 36988 46396 37044
rect 46452 36988 46462 37044
rect 51762 36988 51772 37044
rect 51828 36988 52444 37044
rect 52500 36988 53228 37044
rect 53284 36988 53294 37044
rect 54562 36988 54572 37044
rect 54628 36988 54740 37044
rect 54898 36988 54908 37044
rect 54964 36988 57204 37044
rect 58034 36988 58044 37044
rect 58100 36988 60000 37044
rect 37762 36876 37772 36932
rect 37828 36876 41580 36932
rect 41636 36876 41646 36932
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 42476 36820 42532 36988
rect 54684 36932 54740 36988
rect 59200 36960 60000 36988
rect 54684 36876 55020 36932
rect 55076 36876 55086 36932
rect 35634 36764 35644 36820
rect 35700 36764 42532 36820
rect 45602 36764 45612 36820
rect 45668 36764 51884 36820
rect 51940 36764 53004 36820
rect 53060 36764 53070 36820
rect 19170 36652 19180 36708
rect 19236 36652 21308 36708
rect 21364 36652 22092 36708
rect 22148 36652 22158 36708
rect 30034 36652 30044 36708
rect 30100 36652 30268 36708
rect 30324 36652 30334 36708
rect 41122 36652 41132 36708
rect 41188 36652 43260 36708
rect 43316 36652 44156 36708
rect 44212 36652 44222 36708
rect 18610 36540 18620 36596
rect 18676 36540 19516 36596
rect 19572 36540 19582 36596
rect 20738 36540 20748 36596
rect 20804 36540 21756 36596
rect 21812 36540 21822 36596
rect 28242 36540 28252 36596
rect 28308 36540 29484 36596
rect 29540 36540 29550 36596
rect 41458 36540 41468 36596
rect 41524 36540 42028 36596
rect 42084 36540 42094 36596
rect 7410 36428 7420 36484
rect 7476 36428 7980 36484
rect 8036 36428 10220 36484
rect 10276 36428 10286 36484
rect 11554 36428 11564 36484
rect 11620 36428 12460 36484
rect 12516 36428 14140 36484
rect 14196 36428 15148 36484
rect 15204 36428 15214 36484
rect 21522 36428 21532 36484
rect 21588 36428 21980 36484
rect 22036 36428 22046 36484
rect 44370 36428 44380 36484
rect 44436 36428 45052 36484
rect 45108 36428 45724 36484
rect 45780 36428 45790 36484
rect 46274 36428 46284 36484
rect 46340 36428 47068 36484
rect 47124 36428 47134 36484
rect 59200 36372 60000 36400
rect 6402 36316 6412 36372
rect 6468 36316 10332 36372
rect 10388 36316 10780 36372
rect 10836 36316 10846 36372
rect 18274 36316 18284 36372
rect 18340 36316 18956 36372
rect 19012 36316 20636 36372
rect 20692 36316 20702 36372
rect 26226 36316 26236 36372
rect 26292 36316 27020 36372
rect 27076 36316 27086 36372
rect 43586 36316 43596 36372
rect 43652 36316 43932 36372
rect 43988 36316 45276 36372
rect 45332 36316 45342 36372
rect 58370 36316 58380 36372
rect 58436 36316 60000 36372
rect 59200 36288 60000 36316
rect 9762 36204 9772 36260
rect 9828 36204 10892 36260
rect 10948 36204 11900 36260
rect 11956 36204 11966 36260
rect 12898 36204 12908 36260
rect 12964 36204 14476 36260
rect 14532 36204 14542 36260
rect 31042 36204 31052 36260
rect 31108 36204 31948 36260
rect 32004 36204 32014 36260
rect 45826 36204 45836 36260
rect 45892 36204 47292 36260
rect 47348 36204 48524 36260
rect 48580 36204 49084 36260
rect 49140 36204 49150 36260
rect 56242 36204 56252 36260
rect 56308 36204 57820 36260
rect 57876 36204 57886 36260
rect 41346 36092 41356 36148
rect 41412 36092 50316 36148
rect 50372 36092 50382 36148
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 50546 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50830 36092
rect 2034 35980 2044 36036
rect 2100 35980 6636 36036
rect 6692 35980 6972 36036
rect 7028 35980 7308 36036
rect 7364 35980 7374 36036
rect 34962 35980 34972 36036
rect 35028 35980 37660 36036
rect 37716 35980 38164 36036
rect 3938 35868 3948 35924
rect 4004 35868 7420 35924
rect 7476 35868 7486 35924
rect 13906 35868 13916 35924
rect 13972 35868 14700 35924
rect 14756 35868 14766 35924
rect 38108 35812 38164 35980
rect 47394 35868 47404 35924
rect 47460 35868 48188 35924
rect 48244 35868 48254 35924
rect 50978 35868 50988 35924
rect 51044 35868 52220 35924
rect 52276 35868 52286 35924
rect 2482 35756 2492 35812
rect 2548 35756 4956 35812
rect 5012 35756 6076 35812
rect 6132 35756 6142 35812
rect 7074 35756 7084 35812
rect 7140 35756 7364 35812
rect 8194 35756 8204 35812
rect 8260 35756 8652 35812
rect 8708 35756 8718 35812
rect 16594 35756 16604 35812
rect 16660 35756 17948 35812
rect 18004 35756 18508 35812
rect 18564 35756 18574 35812
rect 29810 35756 29820 35812
rect 29876 35756 36092 35812
rect 36148 35756 36540 35812
rect 36596 35756 37324 35812
rect 37380 35756 37390 35812
rect 38098 35756 38108 35812
rect 38164 35756 38174 35812
rect 40002 35756 40012 35812
rect 40068 35756 41244 35812
rect 41300 35756 41310 35812
rect 47618 35756 47628 35812
rect 47684 35756 48300 35812
rect 48356 35756 49308 35812
rect 49364 35756 51996 35812
rect 52052 35756 52062 35812
rect 56578 35756 56588 35812
rect 56644 35756 57820 35812
rect 57876 35756 57886 35812
rect 0 35700 800 35728
rect 7308 35700 7364 35756
rect 29820 35700 29876 35756
rect 59200 35700 60000 35728
rect 0 35644 1708 35700
rect 1764 35644 1774 35700
rect 3154 35644 3164 35700
rect 3220 35644 4396 35700
rect 4452 35644 4462 35700
rect 7298 35644 7308 35700
rect 7364 35644 7374 35700
rect 14354 35644 14364 35700
rect 14420 35644 16268 35700
rect 16324 35644 16334 35700
rect 18050 35644 18060 35700
rect 18116 35644 18620 35700
rect 18676 35644 18686 35700
rect 20178 35644 20188 35700
rect 20244 35644 20524 35700
rect 20580 35644 20590 35700
rect 24770 35644 24780 35700
rect 24836 35644 25340 35700
rect 25396 35644 25406 35700
rect 28578 35644 28588 35700
rect 28644 35644 29876 35700
rect 36866 35644 36876 35700
rect 36932 35644 37436 35700
rect 37492 35644 37502 35700
rect 37986 35644 37996 35700
rect 38052 35644 38780 35700
rect 38836 35644 39228 35700
rect 39284 35644 39294 35700
rect 40114 35644 40124 35700
rect 40180 35644 40908 35700
rect 40964 35644 40974 35700
rect 45602 35644 45612 35700
rect 45668 35644 47516 35700
rect 47572 35644 47852 35700
rect 47908 35644 48636 35700
rect 48692 35644 48702 35700
rect 49970 35644 49980 35700
rect 50036 35644 50652 35700
rect 50708 35644 50718 35700
rect 53778 35644 53788 35700
rect 53844 35644 54236 35700
rect 54292 35644 55020 35700
rect 55076 35644 55086 35700
rect 57138 35644 57148 35700
rect 57204 35644 58268 35700
rect 58324 35644 60000 35700
rect 0 35616 800 35644
rect 59200 35616 60000 35644
rect 6850 35532 6860 35588
rect 6916 35532 7196 35588
rect 7252 35532 7262 35588
rect 7410 35532 7420 35588
rect 7476 35532 8540 35588
rect 8596 35532 8606 35588
rect 30034 35532 30044 35588
rect 30100 35532 30492 35588
rect 30548 35532 30558 35588
rect 33618 35532 33628 35588
rect 33684 35532 34412 35588
rect 34468 35532 35420 35588
rect 35476 35532 35486 35588
rect 36306 35532 36316 35588
rect 36372 35532 37100 35588
rect 37156 35532 38556 35588
rect 38612 35476 38668 35588
rect 48178 35532 48188 35588
rect 48244 35532 51212 35588
rect 51268 35532 51278 35588
rect 4172 35420 8876 35476
rect 8932 35420 8942 35476
rect 14018 35420 14028 35476
rect 14084 35420 14812 35476
rect 14868 35420 14878 35476
rect 16482 35420 16492 35476
rect 16548 35420 17948 35476
rect 18004 35420 19292 35476
rect 19348 35420 20076 35476
rect 20132 35420 20142 35476
rect 29250 35420 29260 35476
rect 29316 35420 30380 35476
rect 30436 35420 31836 35476
rect 31892 35420 32396 35476
rect 32452 35420 35588 35476
rect 36642 35420 36652 35476
rect 36708 35420 37436 35476
rect 37492 35420 38444 35476
rect 38500 35420 38510 35476
rect 38612 35420 49980 35476
rect 50036 35420 50428 35476
rect 4172 35364 4228 35420
rect 35532 35364 35588 35420
rect 50372 35364 50428 35420
rect 4162 35308 4172 35364
rect 4228 35308 4238 35364
rect 20514 35308 20524 35364
rect 20580 35308 21868 35364
rect 21924 35308 21934 35364
rect 35532 35308 44044 35364
rect 44100 35308 45836 35364
rect 45892 35308 45902 35364
rect 50372 35308 52780 35364
rect 52836 35308 52846 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 9090 35196 9100 35252
rect 9156 35196 9660 35252
rect 9716 35196 9726 35252
rect 17826 35196 17836 35252
rect 17892 35196 18844 35252
rect 18900 35196 18910 35252
rect 27906 35196 27916 35252
rect 27972 35196 28364 35252
rect 28420 35196 29148 35252
rect 29204 35196 29214 35252
rect 29362 35196 29372 35252
rect 29428 35196 29820 35252
rect 29876 35196 29886 35252
rect 31938 35196 31948 35252
rect 32004 35196 34244 35252
rect 34188 35140 34244 35196
rect 9202 35084 9212 35140
rect 9268 35084 24444 35140
rect 24500 35084 25116 35140
rect 25172 35084 25182 35140
rect 32162 35084 32172 35140
rect 32228 35084 33404 35140
rect 33460 35084 33964 35140
rect 34020 35084 34030 35140
rect 34188 35084 36316 35140
rect 36372 35084 36382 35140
rect 59200 35028 60000 35056
rect 5068 34972 22316 35028
rect 22372 34972 22988 35028
rect 23044 34972 23548 35028
rect 23604 34972 23614 35028
rect 24882 34972 24892 35028
rect 24948 34972 26908 35028
rect 26964 34972 27804 35028
rect 27860 34972 33628 35028
rect 33684 34972 33694 35028
rect 58146 34972 58156 35028
rect 58212 34972 60000 35028
rect 5068 34916 5124 34972
rect 59200 34944 60000 34972
rect 5058 34860 5068 34916
rect 5124 34860 5134 34916
rect 9762 34860 9772 34916
rect 9828 34860 10668 34916
rect 10724 34860 10734 34916
rect 15026 34860 15036 34916
rect 15092 34860 17388 34916
rect 17444 34860 17454 34916
rect 22754 34860 22764 34916
rect 22820 34860 23772 34916
rect 23828 34860 23838 34916
rect 24546 34860 24556 34916
rect 24612 34860 25340 34916
rect 25396 34860 25406 34916
rect 26114 34860 26124 34916
rect 26180 34860 26684 34916
rect 26740 34860 26750 34916
rect 30146 34860 30156 34916
rect 30212 34860 31500 34916
rect 31556 34860 32396 34916
rect 32452 34860 32462 34916
rect 34738 34860 34748 34916
rect 34804 34860 36092 34916
rect 36148 34860 36158 34916
rect 38322 34860 38332 34916
rect 38388 34860 39900 34916
rect 39956 34860 39966 34916
rect 44930 34860 44940 34916
rect 44996 34860 45836 34916
rect 45892 34860 45902 34916
rect 55234 34860 55244 34916
rect 55300 34860 55692 34916
rect 55748 34860 55758 34916
rect 6850 34748 6860 34804
rect 6916 34748 9100 34804
rect 9156 34748 9166 34804
rect 9622 34748 9660 34804
rect 9716 34748 9726 34804
rect 9874 34748 9884 34804
rect 9940 34748 10556 34804
rect 10612 34748 11004 34804
rect 11060 34748 11070 34804
rect 18386 34748 18396 34804
rect 18452 34748 19516 34804
rect 19572 34748 19582 34804
rect 20066 34748 20076 34804
rect 20132 34748 21644 34804
rect 21700 34748 21710 34804
rect 22642 34748 22652 34804
rect 22708 34748 23324 34804
rect 23380 34748 23390 34804
rect 24322 34748 24332 34804
rect 24388 34748 25564 34804
rect 25620 34748 25630 34804
rect 31938 34748 31948 34804
rect 32004 34748 32284 34804
rect 32340 34748 32350 34804
rect 34514 34748 34524 34804
rect 34580 34748 35980 34804
rect 36036 34748 36046 34804
rect 51538 34748 51548 34804
rect 51604 34748 53004 34804
rect 53060 34748 53788 34804
rect 53844 34748 53854 34804
rect 7410 34636 7420 34692
rect 7476 34636 14252 34692
rect 14308 34636 18956 34692
rect 19012 34636 19022 34692
rect 28466 34636 28476 34692
rect 28532 34636 29484 34692
rect 29540 34636 29550 34692
rect 31266 34636 31276 34692
rect 31332 34636 32172 34692
rect 32228 34636 32238 34692
rect 39890 34636 39900 34692
rect 39956 34636 41132 34692
rect 41188 34636 41198 34692
rect 52546 34636 52556 34692
rect 52612 34636 57820 34692
rect 57876 34636 57886 34692
rect 28914 34524 28924 34580
rect 28980 34524 29596 34580
rect 29652 34524 29662 34580
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 50546 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50830 34524
rect 9874 34412 9884 34468
rect 9940 34412 11452 34468
rect 11508 34412 11518 34468
rect 25890 34412 25900 34468
rect 25956 34412 26348 34468
rect 26404 34412 26414 34468
rect 47852 34412 48748 34468
rect 48804 34412 48814 34468
rect 47852 34356 47908 34412
rect 59200 34356 60000 34384
rect 2034 34300 2044 34356
rect 2100 34300 6188 34356
rect 6244 34300 6254 34356
rect 8978 34300 8988 34356
rect 9044 34300 9436 34356
rect 9492 34300 9772 34356
rect 9828 34300 9838 34356
rect 11218 34300 11228 34356
rect 11284 34300 13132 34356
rect 13188 34300 14364 34356
rect 14420 34300 14430 34356
rect 28802 34300 28812 34356
rect 28868 34300 29596 34356
rect 29652 34300 29662 34356
rect 41570 34300 41580 34356
rect 41636 34300 42812 34356
rect 42868 34300 42878 34356
rect 45826 34300 45836 34356
rect 45892 34300 47852 34356
rect 47908 34300 47918 34356
rect 48066 34300 48076 34356
rect 48132 34300 48972 34356
rect 49028 34300 49644 34356
rect 49700 34300 49710 34356
rect 57586 34300 57596 34356
rect 57652 34300 58156 34356
rect 58212 34300 60000 34356
rect 59200 34272 60000 34300
rect 10658 34188 10668 34244
rect 10724 34188 11788 34244
rect 11844 34188 11854 34244
rect 20850 34188 20860 34244
rect 20916 34188 21532 34244
rect 21588 34188 22316 34244
rect 22372 34188 22382 34244
rect 27682 34188 27692 34244
rect 27748 34188 28924 34244
rect 28980 34188 28990 34244
rect 33730 34188 33740 34244
rect 33796 34188 34748 34244
rect 34804 34188 34814 34244
rect 42578 34188 42588 34244
rect 42644 34188 45500 34244
rect 45556 34188 45566 34244
rect 47506 34188 47516 34244
rect 47572 34188 49196 34244
rect 49252 34188 49262 34244
rect 50306 34188 50316 34244
rect 50372 34188 51660 34244
rect 51716 34188 51726 34244
rect 55906 34188 55916 34244
rect 55972 34188 57820 34244
rect 57876 34188 57886 34244
rect 9538 34076 9548 34132
rect 9604 34076 11116 34132
rect 11172 34076 11182 34132
rect 13570 34076 13580 34132
rect 13636 34076 14700 34132
rect 14756 34076 14766 34132
rect 15250 34076 15260 34132
rect 15316 34076 20300 34132
rect 20356 34076 20366 34132
rect 24322 34076 24332 34132
rect 24388 34076 24892 34132
rect 24948 34076 25228 34132
rect 25284 34076 25294 34132
rect 25890 34076 25900 34132
rect 25956 34076 27468 34132
rect 27524 34076 27534 34132
rect 28578 34076 28588 34132
rect 28644 34076 29372 34132
rect 29428 34076 29438 34132
rect 29810 34076 29820 34132
rect 29876 34076 30828 34132
rect 30884 34076 31612 34132
rect 31668 34076 31678 34132
rect 33954 34076 33964 34132
rect 34020 34076 34636 34132
rect 34692 34076 34702 34132
rect 36866 34076 36876 34132
rect 36932 34076 39004 34132
rect 39060 34076 39070 34132
rect 41234 34076 41244 34132
rect 41300 34076 42252 34132
rect 42308 34076 42318 34132
rect 43138 34076 43148 34132
rect 43204 34076 45052 34132
rect 45108 34076 45388 34132
rect 45444 34076 45454 34132
rect 48290 34076 48300 34132
rect 48356 34076 49308 34132
rect 49364 34076 49374 34132
rect 49746 34076 49756 34132
rect 49812 34076 50652 34132
rect 50708 34076 50718 34132
rect 55346 34076 55356 34132
rect 55412 34076 55692 34132
rect 55748 34076 55758 34132
rect 8642 33964 8652 34020
rect 8708 33964 11228 34020
rect 11284 33964 11294 34020
rect 17938 33964 17948 34020
rect 18004 33964 18844 34020
rect 18900 33964 18910 34020
rect 30370 33964 30380 34020
rect 30436 33964 31388 34020
rect 31444 33964 31454 34020
rect 37090 33964 37100 34020
rect 37156 33964 37660 34020
rect 37716 33964 38780 34020
rect 38836 33964 38846 34020
rect 36306 33852 36316 33908
rect 36372 33852 43932 33908
rect 43988 33852 45724 33908
rect 45780 33852 45790 33908
rect 46722 33852 46732 33908
rect 46788 33852 54796 33908
rect 54852 33852 54862 33908
rect 55458 33852 55468 33908
rect 55524 33852 56700 33908
rect 56756 33852 56766 33908
rect 16706 33740 16716 33796
rect 16772 33740 18508 33796
rect 18564 33740 18844 33796
rect 18900 33740 18910 33796
rect 31042 33740 31052 33796
rect 31108 33740 33628 33796
rect 33684 33740 33694 33796
rect 40114 33740 40124 33796
rect 40180 33740 41020 33796
rect 41076 33740 43036 33796
rect 43092 33740 43102 33796
rect 0 33684 800 33712
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 59200 33684 60000 33712
rect 0 33628 1708 33684
rect 1764 33628 2492 33684
rect 2548 33628 2558 33684
rect 5058 33628 5068 33684
rect 5124 33628 7196 33684
rect 7252 33628 7262 33684
rect 38210 33628 38220 33684
rect 38276 33628 38668 33684
rect 38724 33628 38734 33684
rect 58146 33628 58156 33684
rect 58212 33628 60000 33684
rect 0 33600 800 33628
rect 59200 33600 60000 33628
rect 15698 33516 15708 33572
rect 15764 33516 17500 33572
rect 17556 33516 17948 33572
rect 18004 33516 18014 33572
rect 31042 33516 31052 33572
rect 31108 33516 32060 33572
rect 32116 33516 32732 33572
rect 32788 33516 33516 33572
rect 33572 33516 33582 33572
rect 44370 33516 44380 33572
rect 44436 33516 45276 33572
rect 45332 33516 45342 33572
rect 3714 33404 3724 33460
rect 3780 33404 5964 33460
rect 6020 33404 6030 33460
rect 12674 33404 12684 33460
rect 12740 33404 13132 33460
rect 13188 33404 13580 33460
rect 13636 33404 13646 33460
rect 13906 33404 13916 33460
rect 13972 33404 16492 33460
rect 16548 33404 16558 33460
rect 31826 33404 31836 33460
rect 31892 33404 32844 33460
rect 32900 33404 32910 33460
rect 34738 33404 34748 33460
rect 34804 33404 35532 33460
rect 35588 33404 35598 33460
rect 36530 33404 36540 33460
rect 36596 33404 37100 33460
rect 37156 33404 39676 33460
rect 39732 33404 39742 33460
rect 47170 33404 47180 33460
rect 47236 33404 48748 33460
rect 48804 33404 50316 33460
rect 50372 33404 50382 33460
rect 6402 33292 6412 33348
rect 6468 33292 6860 33348
rect 6916 33292 7588 33348
rect 7970 33292 7980 33348
rect 8036 33292 8988 33348
rect 9044 33292 9054 33348
rect 14018 33292 14028 33348
rect 14084 33292 16828 33348
rect 16884 33292 16894 33348
rect 17266 33292 17276 33348
rect 17332 33292 19404 33348
rect 19460 33292 19470 33348
rect 20962 33292 20972 33348
rect 21028 33292 21420 33348
rect 21476 33292 22540 33348
rect 22596 33292 22606 33348
rect 34290 33292 34300 33348
rect 34356 33292 35644 33348
rect 35700 33292 35710 33348
rect 48962 33292 48972 33348
rect 49028 33292 49980 33348
rect 50036 33292 50046 33348
rect 51650 33292 51660 33348
rect 51716 33292 51996 33348
rect 52052 33292 52892 33348
rect 52948 33292 52958 33348
rect 7532 33124 7588 33292
rect 17836 33236 17892 33292
rect 8642 33180 8652 33236
rect 8708 33180 16380 33236
rect 16436 33180 16446 33236
rect 17826 33180 17836 33236
rect 17892 33180 17902 33236
rect 26674 33180 26684 33236
rect 26740 33180 27580 33236
rect 27636 33180 27646 33236
rect 34962 33180 34972 33236
rect 35028 33180 35756 33236
rect 35812 33180 35822 33236
rect 44258 33180 44268 33236
rect 44324 33180 45052 33236
rect 45108 33180 47404 33236
rect 47460 33180 48412 33236
rect 48468 33180 50092 33236
rect 50148 33180 50158 33236
rect 50372 33180 52668 33236
rect 52724 33180 52734 33236
rect 50372 33124 50428 33180
rect 2706 33068 2716 33124
rect 2772 33068 3276 33124
rect 3332 33068 6188 33124
rect 6244 33068 7308 33124
rect 7364 33068 7374 33124
rect 7522 33068 7532 33124
rect 7588 33068 7598 33124
rect 9622 33068 9660 33124
rect 9716 33068 9726 33124
rect 9986 33068 9996 33124
rect 10052 33068 10556 33124
rect 10612 33068 10622 33124
rect 17714 33068 17724 33124
rect 17780 33068 19068 33124
rect 19124 33068 19134 33124
rect 19292 33068 20412 33124
rect 20468 33068 20478 33124
rect 48178 33068 48188 33124
rect 48244 33068 49532 33124
rect 49588 33068 50428 33124
rect 51874 33068 51884 33124
rect 51940 33068 53004 33124
rect 53060 33068 53070 33124
rect 19292 33012 19348 33068
rect 59200 33012 60000 33040
rect 5954 32956 5964 33012
rect 6020 32956 6412 33012
rect 6468 32956 10332 33012
rect 10388 32956 10398 33012
rect 15138 32956 15148 33012
rect 15204 32956 19348 33012
rect 57586 32956 57596 33012
rect 57652 32956 58156 33012
rect 58212 32956 60000 33012
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 50546 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50830 32956
rect 59200 32928 60000 32956
rect 16482 32844 16492 32900
rect 16548 32844 18620 32900
rect 18676 32844 18686 32900
rect 38882 32844 38892 32900
rect 38948 32844 39676 32900
rect 39732 32844 40236 32900
rect 40292 32844 47628 32900
rect 47684 32844 47694 32900
rect 6850 32732 6860 32788
rect 6916 32732 7980 32788
rect 8036 32732 9436 32788
rect 9492 32732 9502 32788
rect 11218 32732 11228 32788
rect 11284 32732 11788 32788
rect 11844 32732 15148 32788
rect 18386 32732 18396 32788
rect 18452 32732 23212 32788
rect 23268 32732 23278 32788
rect 45154 32732 45164 32788
rect 45220 32732 46732 32788
rect 46788 32732 46798 32788
rect 15092 32676 15148 32732
rect 14914 32620 14924 32676
rect 14980 32620 14990 32676
rect 15092 32620 16380 32676
rect 16436 32620 18284 32676
rect 18340 32620 19180 32676
rect 19236 32620 19246 32676
rect 26898 32620 26908 32676
rect 26964 32620 29372 32676
rect 29428 32620 29438 32676
rect 41570 32620 41580 32676
rect 41636 32620 43260 32676
rect 43316 32620 43326 32676
rect 43586 32620 43596 32676
rect 43652 32620 57820 32676
rect 57876 32620 57886 32676
rect 14924 32564 14980 32620
rect 5954 32508 5964 32564
rect 6020 32508 7084 32564
rect 7140 32508 7150 32564
rect 14924 32508 15708 32564
rect 15764 32508 15774 32564
rect 16706 32508 16716 32564
rect 16772 32508 17836 32564
rect 17892 32508 17902 32564
rect 19954 32508 19964 32564
rect 20020 32508 20030 32564
rect 29810 32508 29820 32564
rect 29876 32508 30380 32564
rect 30436 32508 31836 32564
rect 31892 32508 31902 32564
rect 37650 32508 37660 32564
rect 37716 32508 41468 32564
rect 41524 32508 42924 32564
rect 42980 32508 42990 32564
rect 43138 32508 43148 32564
rect 43204 32508 45388 32564
rect 45444 32508 46508 32564
rect 46564 32508 46574 32564
rect 50978 32508 50988 32564
rect 51044 32508 51884 32564
rect 51940 32508 51950 32564
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 7298 31948 7308 32004
rect 7364 31948 8204 32004
rect 8260 31948 8270 32004
rect 19964 31892 20020 32508
rect 23314 32396 23324 32452
rect 23380 32396 23772 32452
rect 23828 32396 23838 32452
rect 30930 32396 30940 32452
rect 30996 32396 31724 32452
rect 31780 32396 31790 32452
rect 32050 32396 32060 32452
rect 32116 32396 37884 32452
rect 37940 32396 37950 32452
rect 59200 32340 60000 32368
rect 33618 32284 33628 32340
rect 33684 32284 35084 32340
rect 35140 32284 35150 32340
rect 57138 32284 57148 32340
rect 57204 32284 58156 32340
rect 58212 32284 60000 32340
rect 59200 32256 60000 32284
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 22978 32060 22988 32116
rect 23044 32060 28700 32116
rect 28756 32060 28766 32116
rect 46722 32060 46732 32116
rect 46788 32060 50204 32116
rect 50260 32060 50270 32116
rect 27682 31948 27692 32004
rect 27748 31948 28140 32004
rect 28196 31948 28588 32004
rect 28644 31948 28654 32004
rect 30594 31948 30604 32004
rect 30660 31948 33292 32004
rect 33348 31948 33358 32004
rect 47058 31948 47068 32004
rect 47124 31948 57708 32004
rect 57764 31948 57774 32004
rect 4498 31836 4508 31892
rect 4564 31836 5068 31892
rect 5124 31836 5134 31892
rect 7186 31836 7196 31892
rect 7252 31836 10556 31892
rect 10612 31836 10622 31892
rect 10994 31836 11004 31892
rect 11060 31836 14924 31892
rect 14980 31836 16268 31892
rect 16324 31836 16334 31892
rect 19292 31836 20020 31892
rect 30034 31836 30044 31892
rect 30100 31836 34524 31892
rect 34580 31836 34590 31892
rect 35186 31836 35196 31892
rect 35252 31836 36092 31892
rect 36148 31836 36158 31892
rect 39218 31836 39228 31892
rect 39284 31836 41356 31892
rect 41412 31836 41422 31892
rect 42354 31836 42364 31892
rect 42420 31836 43708 31892
rect 43764 31836 46844 31892
rect 46900 31836 46910 31892
rect 47954 31836 47964 31892
rect 48020 31836 49308 31892
rect 49364 31836 49374 31892
rect 19292 31780 19348 31836
rect 4834 31724 4844 31780
rect 4900 31724 4910 31780
rect 8754 31724 8764 31780
rect 8820 31724 9660 31780
rect 9716 31724 9726 31780
rect 12114 31724 12124 31780
rect 12180 31724 12572 31780
rect 12628 31724 15092 31780
rect 15586 31724 15596 31780
rect 15652 31724 17164 31780
rect 17220 31724 17230 31780
rect 18162 31724 18172 31780
rect 18228 31724 19348 31780
rect 26562 31724 26572 31780
rect 26628 31724 29708 31780
rect 29764 31724 29774 31780
rect 36194 31724 36204 31780
rect 36260 31724 37100 31780
rect 37156 31724 38556 31780
rect 38612 31724 38622 31780
rect 44930 31724 44940 31780
rect 44996 31724 45836 31780
rect 45892 31724 46396 31780
rect 46452 31724 46462 31780
rect 48626 31724 48636 31780
rect 48692 31724 50764 31780
rect 50820 31724 50830 31780
rect 54786 31724 54796 31780
rect 54852 31724 55132 31780
rect 55188 31724 55198 31780
rect 4844 31668 4900 31724
rect 15036 31668 15092 31724
rect 19292 31668 19348 31724
rect 59200 31668 60000 31696
rect 4162 31612 4172 31668
rect 4228 31612 4900 31668
rect 7858 31612 7868 31668
rect 7924 31612 8428 31668
rect 8484 31612 9884 31668
rect 9940 31612 9950 31668
rect 11554 31612 11564 31668
rect 11620 31612 14140 31668
rect 14196 31612 14476 31668
rect 14532 31612 14542 31668
rect 15026 31612 15036 31668
rect 15092 31612 15484 31668
rect 15540 31612 15550 31668
rect 19282 31612 19292 31668
rect 19348 31612 19358 31668
rect 24434 31612 24444 31668
rect 24500 31612 25340 31668
rect 25396 31612 25406 31668
rect 28354 31612 28364 31668
rect 28420 31612 29148 31668
rect 29204 31612 29214 31668
rect 34738 31612 34748 31668
rect 34804 31612 34814 31668
rect 36418 31612 36428 31668
rect 36484 31612 37212 31668
rect 37268 31612 37278 31668
rect 38994 31612 39004 31668
rect 39060 31612 39676 31668
rect 39732 31612 39742 31668
rect 45154 31612 45164 31668
rect 45220 31612 45948 31668
rect 46004 31612 53340 31668
rect 53396 31612 54236 31668
rect 54292 31612 54302 31668
rect 56914 31612 56924 31668
rect 56980 31612 57484 31668
rect 57540 31612 60000 31668
rect 2706 31500 2716 31556
rect 2772 31500 3164 31556
rect 3220 31500 3724 31556
rect 3780 31500 3790 31556
rect 6402 31500 6412 31556
rect 6468 31500 8540 31556
rect 8596 31500 8606 31556
rect 10882 31500 10892 31556
rect 10948 31500 12012 31556
rect 12068 31500 12078 31556
rect 20066 31500 20076 31556
rect 20132 31500 24220 31556
rect 24276 31500 24286 31556
rect 24658 31500 24668 31556
rect 24724 31500 25900 31556
rect 25956 31500 25966 31556
rect 27122 31500 27132 31556
rect 27188 31500 28252 31556
rect 28308 31500 30044 31556
rect 30100 31500 30110 31556
rect 4946 31388 4956 31444
rect 5012 31388 9100 31444
rect 9156 31388 9548 31444
rect 9604 31388 9614 31444
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 34748 31332 34804 31612
rect 59200 31584 60000 31612
rect 34962 31500 34972 31556
rect 35028 31500 37324 31556
rect 37380 31500 38108 31556
rect 38164 31500 38174 31556
rect 44146 31500 44156 31556
rect 44212 31500 45276 31556
rect 45332 31500 51044 31556
rect 53666 31500 53676 31556
rect 53732 31500 55020 31556
rect 55076 31500 55086 31556
rect 57810 31500 57820 31556
rect 57876 31500 57886 31556
rect 50988 31444 51044 31500
rect 47954 31388 47964 31444
rect 48020 31388 48860 31444
rect 48916 31388 48926 31444
rect 50988 31388 55804 31444
rect 55860 31388 55870 31444
rect 50546 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50830 31388
rect 11218 31276 11228 31332
rect 11284 31276 16828 31332
rect 16884 31276 16894 31332
rect 34748 31276 39900 31332
rect 39956 31276 39966 31332
rect 45714 31276 45724 31332
rect 45780 31276 46060 31332
rect 46116 31276 46126 31332
rect 57820 31220 57876 31500
rect 4274 31164 4284 31220
rect 4340 31164 4676 31220
rect 15922 31164 15932 31220
rect 15988 31164 16604 31220
rect 16660 31164 17164 31220
rect 17220 31164 17612 31220
rect 17668 31164 17678 31220
rect 27346 31164 27356 31220
rect 27412 31164 27916 31220
rect 27972 31164 28364 31220
rect 28420 31164 28430 31220
rect 28914 31164 28924 31220
rect 28980 31164 29820 31220
rect 29876 31164 29886 31220
rect 37202 31164 37212 31220
rect 37268 31164 38108 31220
rect 38164 31164 38174 31220
rect 38658 31164 38668 31220
rect 38724 31164 39788 31220
rect 39844 31164 39854 31220
rect 41906 31164 41916 31220
rect 41972 31164 42812 31220
rect 42868 31164 43148 31220
rect 43204 31164 43214 31220
rect 48850 31164 48860 31220
rect 48916 31164 57876 31220
rect 4620 31108 4676 31164
rect 2818 31052 2828 31108
rect 2884 31052 3276 31108
rect 3332 31052 4172 31108
rect 4228 31052 4238 31108
rect 4610 31052 4620 31108
rect 4676 31052 9716 31108
rect 12450 31052 12460 31108
rect 12516 31052 15596 31108
rect 15652 31052 15662 31108
rect 16258 31052 16268 31108
rect 16324 31052 17388 31108
rect 17444 31052 17454 31108
rect 21410 31052 21420 31108
rect 21476 31052 21868 31108
rect 21924 31052 21934 31108
rect 23538 31052 23548 31108
rect 23604 31052 26908 31108
rect 26964 31052 32508 31108
rect 32564 31052 36092 31108
rect 36148 31052 36158 31108
rect 43362 31052 43372 31108
rect 43428 31052 44604 31108
rect 44660 31052 44670 31108
rect 47282 31052 47292 31108
rect 47348 31052 48524 31108
rect 48580 31052 49196 31108
rect 49252 31052 49262 31108
rect 50372 31052 52444 31108
rect 52500 31052 52510 31108
rect 52658 31052 52668 31108
rect 52724 31052 57820 31108
rect 57876 31052 57886 31108
rect 9660 30996 9716 31052
rect 50372 30996 50428 31052
rect 59200 30996 60000 31024
rect 3490 30940 3500 30996
rect 3556 30940 5404 30996
rect 5460 30940 5470 30996
rect 9650 30940 9660 30996
rect 9716 30940 12348 30996
rect 12404 30940 13468 30996
rect 13524 30940 13534 30996
rect 16482 30940 16492 30996
rect 16548 30940 17836 30996
rect 17892 30940 17902 30996
rect 19282 30940 19292 30996
rect 19348 30940 20972 30996
rect 21028 30940 21038 30996
rect 22642 30940 22652 30996
rect 22708 30940 23324 30996
rect 23380 30940 23390 30996
rect 28242 30940 28252 30996
rect 28308 30940 28924 30996
rect 28980 30940 28990 30996
rect 29698 30940 29708 30996
rect 29764 30940 30044 30996
rect 30100 30940 31388 30996
rect 31444 30940 32284 30996
rect 32340 30940 32350 30996
rect 34178 30940 34188 30996
rect 34244 30940 35868 30996
rect 35924 30940 35934 30996
rect 48178 30940 48188 30996
rect 48244 30940 49308 30996
rect 49364 30940 50092 30996
rect 50148 30940 50428 30996
rect 58370 30940 58380 30996
rect 58436 30940 60000 30996
rect 59200 30912 60000 30940
rect 6178 30828 6188 30884
rect 6244 30828 7196 30884
rect 7252 30828 7262 30884
rect 13794 30828 13804 30884
rect 13860 30828 14364 30884
rect 14420 30828 14430 30884
rect 21634 30828 21644 30884
rect 21700 30828 24332 30884
rect 24388 30828 24398 30884
rect 24658 30828 24668 30884
rect 24724 30828 25676 30884
rect 25732 30828 26236 30884
rect 26292 30828 26572 30884
rect 26628 30828 26638 30884
rect 28466 30828 28476 30884
rect 28532 30828 29596 30884
rect 29652 30828 29662 30884
rect 51090 30828 51100 30884
rect 51156 30828 52892 30884
rect 52948 30828 52958 30884
rect 24332 30772 24388 30828
rect 4162 30716 4172 30772
rect 4228 30716 6972 30772
rect 7028 30716 7756 30772
rect 7812 30716 7822 30772
rect 9874 30716 9884 30772
rect 9940 30716 11676 30772
rect 11732 30716 12684 30772
rect 12740 30716 12750 30772
rect 24332 30716 25228 30772
rect 25284 30716 25294 30772
rect 29250 30716 29260 30772
rect 29316 30716 29932 30772
rect 29988 30716 29998 30772
rect 35186 30716 35196 30772
rect 35252 30716 35868 30772
rect 35924 30716 35934 30772
rect 40450 30716 40460 30772
rect 40516 30716 50092 30772
rect 50148 30716 50158 30772
rect 50530 30716 50540 30772
rect 50596 30716 51324 30772
rect 51380 30716 52332 30772
rect 52388 30716 52398 30772
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 35532 30492 38668 30548
rect 38724 30492 38734 30548
rect 38882 30492 38892 30548
rect 38948 30492 47628 30548
rect 47684 30492 47694 30548
rect 35532 30436 35588 30492
rect 3826 30380 3836 30436
rect 3892 30380 4508 30436
rect 4564 30380 6076 30436
rect 6132 30380 6142 30436
rect 8978 30380 8988 30436
rect 9044 30380 9884 30436
rect 9940 30380 10444 30436
rect 10500 30380 10510 30436
rect 16930 30380 16940 30436
rect 16996 30380 17948 30436
rect 18004 30380 18014 30436
rect 20178 30380 20188 30436
rect 20244 30380 21420 30436
rect 21476 30380 21486 30436
rect 28354 30380 28364 30436
rect 28420 30380 30492 30436
rect 30548 30380 30558 30436
rect 32274 30380 32284 30436
rect 32340 30380 35588 30436
rect 37874 30380 37884 30436
rect 37940 30380 38780 30436
rect 38836 30380 38846 30436
rect 44034 30380 44044 30436
rect 44100 30380 45388 30436
rect 45444 30380 45454 30436
rect 59200 30324 60000 30352
rect 2370 30268 2380 30324
rect 2436 30268 4732 30324
rect 4788 30268 4798 30324
rect 16034 30268 16044 30324
rect 16100 30268 17612 30324
rect 17668 30268 17678 30324
rect 23538 30268 23548 30324
rect 23604 30268 24332 30324
rect 24388 30268 24398 30324
rect 29026 30268 29036 30324
rect 29092 30268 29708 30324
rect 29764 30268 29774 30324
rect 31602 30268 31612 30324
rect 31668 30268 40964 30324
rect 41122 30268 41132 30324
rect 41188 30268 41916 30324
rect 41972 30268 41982 30324
rect 43362 30268 43372 30324
rect 43428 30268 43820 30324
rect 43876 30268 44940 30324
rect 44996 30268 45006 30324
rect 47842 30268 47852 30324
rect 47908 30268 48748 30324
rect 48804 30268 48814 30324
rect 55804 30268 57148 30324
rect 57204 30268 57214 30324
rect 58146 30268 58156 30324
rect 58212 30268 60000 30324
rect 24332 30212 24388 30268
rect 40908 30212 40964 30268
rect 6626 30156 6636 30212
rect 6692 30156 7756 30212
rect 7812 30156 9212 30212
rect 9268 30156 9278 30212
rect 15250 30156 15260 30212
rect 15316 30156 16604 30212
rect 16660 30156 17388 30212
rect 17444 30156 17454 30212
rect 19730 30156 19740 30212
rect 19796 30156 21532 30212
rect 21588 30156 22428 30212
rect 22484 30156 22494 30212
rect 23202 30156 23212 30212
rect 23268 30156 24108 30212
rect 24164 30156 24174 30212
rect 24332 30156 25340 30212
rect 25396 30156 25406 30212
rect 26852 30156 32060 30212
rect 32116 30156 32508 30212
rect 32564 30156 33068 30212
rect 33124 30156 33134 30212
rect 36194 30156 36204 30212
rect 36260 30156 36988 30212
rect 37044 30156 37054 30212
rect 38994 30156 39004 30212
rect 39060 30156 40124 30212
rect 40180 30156 40190 30212
rect 40908 30156 43708 30212
rect 43764 30156 43774 30212
rect 44370 30156 44380 30212
rect 44436 30156 53844 30212
rect 54002 30156 54012 30212
rect 54068 30156 55580 30212
rect 55636 30156 55646 30212
rect 26852 30100 26908 30156
rect 53788 30100 53844 30156
rect 55804 30100 55860 30268
rect 59200 30240 60000 30268
rect 14578 30044 14588 30100
rect 14644 30044 21028 30100
rect 22194 30044 22204 30100
rect 22260 30044 23324 30100
rect 23380 30044 23390 30100
rect 24882 30044 24892 30100
rect 24948 30044 26908 30100
rect 29922 30044 29932 30100
rect 29988 30044 30268 30100
rect 30324 30044 30334 30100
rect 31490 30044 31500 30100
rect 31556 30044 31948 30100
rect 32004 30044 32014 30100
rect 32162 30044 32172 30100
rect 32228 30044 32238 30100
rect 35298 30044 35308 30100
rect 35364 30044 37100 30100
rect 37156 30044 37166 30100
rect 37314 30044 37324 30100
rect 37380 30044 39228 30100
rect 39284 30044 40460 30100
rect 40516 30044 40526 30100
rect 41234 30044 41244 30100
rect 41300 30044 42476 30100
rect 42532 30044 42542 30100
rect 45490 30044 45500 30100
rect 45556 30044 53564 30100
rect 53620 30044 53630 30100
rect 53788 30044 55860 30100
rect 20972 29988 21028 30044
rect 12786 29932 12796 29988
rect 12852 29932 13580 29988
rect 13636 29932 16268 29988
rect 16324 29932 16334 29988
rect 20972 29932 29036 29988
rect 29092 29932 29102 29988
rect 32172 29876 32228 30044
rect 35746 29932 35756 29988
rect 35812 29932 36204 29988
rect 36260 29932 36270 29988
rect 36754 29932 36764 29988
rect 36820 29932 37660 29988
rect 37716 29932 37726 29988
rect 37874 29932 37884 29988
rect 37940 29932 40908 29988
rect 40964 29932 40974 29988
rect 44258 29932 44268 29988
rect 44324 29932 46060 29988
rect 46116 29932 46126 29988
rect 46274 29932 46284 29988
rect 46340 29932 54012 29988
rect 54068 29932 54078 29988
rect 11442 29820 11452 29876
rect 11508 29820 19628 29876
rect 19684 29820 19694 29876
rect 32172 29820 43820 29876
rect 43876 29820 43886 29876
rect 45378 29820 45388 29876
rect 45444 29820 45948 29876
rect 46004 29820 46014 29876
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 50546 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50830 29820
rect 29362 29708 29372 29764
rect 29428 29708 33740 29764
rect 33796 29708 35196 29764
rect 35252 29708 35262 29764
rect 35970 29708 35980 29764
rect 36036 29708 39340 29764
rect 39396 29708 47292 29764
rect 47348 29708 47358 29764
rect 59200 29652 60000 29680
rect 15922 29596 15932 29652
rect 15988 29596 18732 29652
rect 18788 29596 27972 29652
rect 28130 29596 28140 29652
rect 28196 29596 28476 29652
rect 28532 29596 28542 29652
rect 28802 29596 28812 29652
rect 28868 29596 29932 29652
rect 29988 29596 29998 29652
rect 36194 29596 36204 29652
rect 36260 29596 38444 29652
rect 38500 29596 39116 29652
rect 39172 29596 39182 29652
rect 45602 29596 45612 29652
rect 45668 29596 55916 29652
rect 55972 29596 55982 29652
rect 57586 29596 57596 29652
rect 57652 29596 58156 29652
rect 58212 29596 60000 29652
rect 27916 29540 27972 29596
rect 59200 29568 60000 29596
rect 16370 29484 16380 29540
rect 16436 29484 16716 29540
rect 16772 29484 16782 29540
rect 19954 29484 19964 29540
rect 20020 29484 26908 29540
rect 27916 29484 28588 29540
rect 28644 29484 30828 29540
rect 30884 29484 30894 29540
rect 37090 29484 37100 29540
rect 37156 29484 37884 29540
rect 37940 29484 37950 29540
rect 52098 29484 52108 29540
rect 52164 29484 57820 29540
rect 57876 29484 57886 29540
rect 26852 29428 26908 29484
rect 6514 29372 6524 29428
rect 6580 29372 7308 29428
rect 7364 29372 7374 29428
rect 7746 29372 7756 29428
rect 7812 29372 8764 29428
rect 8820 29372 8830 29428
rect 15698 29372 15708 29428
rect 15764 29372 17388 29428
rect 17444 29372 17454 29428
rect 18386 29372 18396 29428
rect 18452 29372 19292 29428
rect 19348 29372 19358 29428
rect 22082 29372 22092 29428
rect 22148 29372 22652 29428
rect 22708 29372 22718 29428
rect 26852 29372 27580 29428
rect 27636 29372 29148 29428
rect 29204 29372 29214 29428
rect 32274 29372 32284 29428
rect 32340 29372 33628 29428
rect 33684 29372 33694 29428
rect 33842 29372 33852 29428
rect 33908 29372 40908 29428
rect 40964 29372 40974 29428
rect 42914 29372 42924 29428
rect 42980 29372 44156 29428
rect 44212 29372 44222 29428
rect 4722 29260 4732 29316
rect 4788 29260 8092 29316
rect 8148 29260 8540 29316
rect 8596 29260 8606 29316
rect 14018 29260 14028 29316
rect 14084 29260 17052 29316
rect 17108 29260 17118 29316
rect 17462 29260 17500 29316
rect 17556 29260 17566 29316
rect 21410 29260 21420 29316
rect 21476 29260 21980 29316
rect 22036 29260 22046 29316
rect 28802 29260 28812 29316
rect 28868 29260 29596 29316
rect 29652 29260 31388 29316
rect 31444 29260 31454 29316
rect 31826 29260 31836 29316
rect 31892 29260 36876 29316
rect 36932 29260 36942 29316
rect 37202 29260 37212 29316
rect 37268 29260 38668 29316
rect 38724 29260 38734 29316
rect 38612 29204 38668 29260
rect 8306 29148 8316 29204
rect 8372 29148 10556 29204
rect 10612 29148 10622 29204
rect 14130 29148 14140 29204
rect 14196 29148 18620 29204
rect 18676 29148 19516 29204
rect 19572 29148 22428 29204
rect 22484 29148 22494 29204
rect 26786 29148 26796 29204
rect 26852 29148 27804 29204
rect 27860 29148 27870 29204
rect 32050 29148 32060 29204
rect 32116 29148 33180 29204
rect 33236 29148 34076 29204
rect 34132 29148 34142 29204
rect 34300 29148 36204 29204
rect 36260 29148 36270 29204
rect 38612 29148 45388 29204
rect 45444 29148 45454 29204
rect 34300 29092 34356 29148
rect 26898 29036 26908 29092
rect 26964 29036 26974 29092
rect 29698 29036 29708 29092
rect 29764 29036 31052 29092
rect 31108 29036 34356 29092
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 18050 28924 18060 28980
rect 18116 28924 20748 28980
rect 20804 28924 20814 28980
rect 26908 28868 26964 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 59200 28980 60000 29008
rect 29474 28924 29484 28980
rect 29540 28924 30716 28980
rect 30772 28924 30782 28980
rect 57250 28924 57260 28980
rect 57316 28924 60000 28980
rect 59200 28896 60000 28924
rect 4946 28812 4956 28868
rect 5012 28812 20188 28868
rect 20244 28812 20254 28868
rect 26908 28812 28028 28868
rect 28084 28812 28094 28868
rect 32386 28812 32396 28868
rect 32452 28812 35308 28868
rect 35364 28812 35374 28868
rect 39564 28812 44604 28868
rect 44660 28812 44670 28868
rect 39564 28756 39620 28812
rect 7074 28700 7084 28756
rect 7140 28700 7868 28756
rect 7924 28700 7934 28756
rect 16370 28700 16380 28756
rect 16436 28700 22764 28756
rect 22820 28700 22830 28756
rect 27794 28700 27804 28756
rect 27860 28700 28476 28756
rect 28532 28700 28542 28756
rect 31714 28700 31724 28756
rect 31780 28700 32732 28756
rect 32788 28700 36148 28756
rect 37538 28700 37548 28756
rect 37604 28700 39004 28756
rect 39060 28700 39070 28756
rect 39554 28700 39564 28756
rect 39620 28700 39630 28756
rect 43698 28700 43708 28756
rect 43764 28700 44940 28756
rect 44996 28700 52556 28756
rect 52612 28700 52622 28756
rect 36092 28644 36148 28700
rect 6962 28588 6972 28644
rect 7028 28588 8652 28644
rect 8708 28588 8718 28644
rect 11218 28588 11228 28644
rect 11284 28588 12124 28644
rect 12180 28588 12572 28644
rect 12628 28588 12638 28644
rect 12786 28588 12796 28644
rect 12852 28588 14364 28644
rect 14420 28588 14430 28644
rect 18284 28588 18732 28644
rect 18788 28588 18798 28644
rect 20402 28588 20412 28644
rect 20468 28588 22876 28644
rect 22932 28588 22942 28644
rect 25666 28588 25676 28644
rect 25732 28588 27020 28644
rect 27076 28588 27086 28644
rect 30370 28588 30380 28644
rect 30436 28588 30828 28644
rect 30884 28588 30894 28644
rect 34738 28588 34748 28644
rect 34804 28588 35532 28644
rect 35588 28588 35868 28644
rect 35924 28588 35934 28644
rect 36082 28588 36092 28644
rect 36148 28588 37660 28644
rect 37716 28588 37726 28644
rect 38098 28588 38108 28644
rect 38164 28588 55244 28644
rect 55300 28588 55580 28644
rect 55636 28588 55646 28644
rect 12338 28476 12348 28532
rect 12404 28476 13580 28532
rect 13636 28476 13646 28532
rect 16706 28476 16716 28532
rect 16772 28476 18060 28532
rect 18116 28476 18126 28532
rect 18284 28420 18340 28588
rect 12002 28364 12012 28420
rect 12068 28364 12908 28420
rect 12964 28364 13804 28420
rect 13860 28364 16772 28420
rect 16930 28364 16940 28420
rect 16996 28364 17276 28420
rect 17332 28364 17342 28420
rect 18162 28364 18172 28420
rect 18228 28364 18340 28420
rect 18396 28476 20076 28532
rect 20132 28476 20142 28532
rect 22530 28476 22540 28532
rect 22596 28476 23660 28532
rect 23716 28476 23726 28532
rect 27234 28476 27244 28532
rect 27300 28476 27804 28532
rect 27860 28476 27870 28532
rect 33506 28476 33516 28532
rect 33572 28476 34524 28532
rect 34580 28476 34590 28532
rect 45938 28476 45948 28532
rect 46004 28476 52108 28532
rect 52164 28476 52174 28532
rect 0 28308 800 28336
rect 16716 28308 16772 28364
rect 18396 28308 18452 28476
rect 21634 28364 21644 28420
rect 21700 28364 22316 28420
rect 22372 28364 22382 28420
rect 30146 28364 30156 28420
rect 30212 28364 31780 28420
rect 31938 28364 31948 28420
rect 32004 28364 34300 28420
rect 34356 28364 34366 28420
rect 34738 28364 34748 28420
rect 34804 28364 38220 28420
rect 38276 28364 38286 28420
rect 38658 28364 38668 28420
rect 38724 28364 39564 28420
rect 39620 28364 39630 28420
rect 41010 28364 41020 28420
rect 41076 28364 42140 28420
rect 42196 28364 46284 28420
rect 46340 28364 46350 28420
rect 31724 28308 31780 28364
rect 59200 28308 60000 28336
rect 0 28252 15260 28308
rect 15316 28252 15326 28308
rect 16716 28252 18452 28308
rect 20188 28252 29484 28308
rect 29540 28252 29550 28308
rect 31724 28252 33628 28308
rect 33684 28252 33694 28308
rect 57922 28252 57932 28308
rect 57988 28252 60000 28308
rect 0 28224 800 28252
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 20188 28084 20244 28252
rect 50546 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50830 28252
rect 59200 28224 60000 28252
rect 17490 28028 17500 28084
rect 17556 28028 20244 28084
rect 24658 28028 24668 28084
rect 24724 28028 25340 28084
rect 25396 28028 25406 28084
rect 27346 28028 27356 28084
rect 27412 28028 27804 28084
rect 27860 28028 30772 28084
rect 30930 28028 30940 28084
rect 30996 28028 32396 28084
rect 32452 28028 32462 28084
rect 32722 28028 32732 28084
rect 32788 28028 33180 28084
rect 33236 28028 33246 28084
rect 43250 28028 43260 28084
rect 43316 28028 44716 28084
rect 44772 28028 44782 28084
rect 45042 28028 45052 28084
rect 45108 28028 46060 28084
rect 46116 28028 46732 28084
rect 46788 28028 46798 28084
rect 30716 27972 30772 28028
rect 15810 27916 15820 27972
rect 15876 27916 18060 27972
rect 18116 27916 18956 27972
rect 19012 27916 19022 27972
rect 20738 27916 20748 27972
rect 20804 27916 28140 27972
rect 28196 27916 28364 27972
rect 28420 27916 28430 27972
rect 30716 27916 34188 27972
rect 34244 27916 34254 27972
rect 34402 27916 34412 27972
rect 34468 27916 35532 27972
rect 35588 27916 35598 27972
rect 36978 27916 36988 27972
rect 37044 27916 38668 27972
rect 38724 27916 39228 27972
rect 39284 27916 39294 27972
rect 39666 27916 39676 27972
rect 39732 27916 40796 27972
rect 40852 27916 40862 27972
rect 43810 27916 43820 27972
rect 43876 27916 44828 27972
rect 44884 27916 44894 27972
rect 34188 27860 34244 27916
rect 8978 27804 8988 27860
rect 9044 27804 14924 27860
rect 14980 27804 14990 27860
rect 17938 27804 17948 27860
rect 18004 27804 18844 27860
rect 18900 27804 18910 27860
rect 21858 27804 21868 27860
rect 21924 27804 22540 27860
rect 22596 27804 22606 27860
rect 34188 27804 37436 27860
rect 37492 27804 37996 27860
rect 38052 27804 38062 27860
rect 42914 27804 42924 27860
rect 42980 27804 54908 27860
rect 54964 27804 54974 27860
rect 18722 27692 18732 27748
rect 18788 27692 20636 27748
rect 20692 27692 20702 27748
rect 21522 27692 21532 27748
rect 21588 27692 22316 27748
rect 22372 27692 22382 27748
rect 44370 27692 44380 27748
rect 44436 27692 45500 27748
rect 45556 27692 45566 27748
rect 59200 27636 60000 27664
rect 22978 27580 22988 27636
rect 23044 27580 30380 27636
rect 30436 27580 30446 27636
rect 43922 27580 43932 27636
rect 43988 27580 45612 27636
rect 45668 27580 49644 27636
rect 49700 27580 49710 27636
rect 57586 27580 57596 27636
rect 57652 27580 58156 27636
rect 58212 27580 60000 27636
rect 59200 27552 60000 27580
rect 14690 27468 14700 27524
rect 14756 27468 22428 27524
rect 22484 27468 22494 27524
rect 43810 27468 43820 27524
rect 43876 27468 45052 27524
rect 45108 27468 56588 27524
rect 56644 27468 56654 27524
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 45490 27356 45500 27412
rect 45556 27356 47068 27412
rect 47124 27356 47134 27412
rect 14130 27244 14140 27300
rect 14196 27244 16268 27300
rect 16324 27244 16334 27300
rect 45724 27244 57820 27300
rect 57876 27244 57886 27300
rect 1922 27132 1932 27188
rect 1988 27132 1998 27188
rect 15474 27132 15484 27188
rect 15540 27132 17948 27188
rect 18004 27132 18014 27188
rect 27122 27132 27132 27188
rect 27188 27132 27580 27188
rect 27636 27132 27646 27188
rect 29474 27132 29484 27188
rect 29540 27132 30156 27188
rect 30212 27132 30222 27188
rect 33730 27132 33740 27188
rect 33796 27132 34748 27188
rect 34804 27132 37100 27188
rect 37156 27132 38220 27188
rect 38276 27132 38286 27188
rect 0 26964 800 26992
rect 1932 26964 1988 27132
rect 38220 27076 38276 27132
rect 45724 27076 45780 27244
rect 46498 27132 46508 27188
rect 46564 27132 47516 27188
rect 47572 27132 56252 27188
rect 56308 27132 56318 27188
rect 19170 27020 19180 27076
rect 19236 27020 19852 27076
rect 19908 27020 19918 27076
rect 20710 27020 20748 27076
rect 20804 27020 20814 27076
rect 23314 27020 23324 27076
rect 23380 27020 24220 27076
rect 24276 27020 24286 27076
rect 28578 27020 28588 27076
rect 28644 27020 29596 27076
rect 29652 27020 29932 27076
rect 29988 27020 30492 27076
rect 30548 27020 30558 27076
rect 38220 27020 39228 27076
rect 39284 27020 39294 27076
rect 45714 27020 45724 27076
rect 45780 27020 45790 27076
rect 59200 26964 60000 26992
rect 0 26908 1988 26964
rect 12338 26908 12348 26964
rect 12404 26908 18732 26964
rect 18788 26908 18798 26964
rect 23090 26908 23100 26964
rect 23156 26908 23772 26964
rect 23828 26908 24332 26964
rect 24388 26908 24398 26964
rect 26450 26908 26460 26964
rect 26516 26908 27356 26964
rect 27412 26908 27422 26964
rect 29810 26908 29820 26964
rect 29876 26908 31612 26964
rect 31668 26908 31678 26964
rect 58156 26908 60000 26964
rect 0 26880 800 26908
rect 58156 26852 58212 26908
rect 59200 26880 60000 26908
rect 12226 26796 12236 26852
rect 12292 26796 13580 26852
rect 13636 26796 13646 26852
rect 28914 26796 28924 26852
rect 28980 26796 32116 26852
rect 34514 26796 34524 26852
rect 34580 26796 35084 26852
rect 35140 26796 35150 26852
rect 37762 26796 37772 26852
rect 37828 26796 38108 26852
rect 38164 26796 38444 26852
rect 38500 26796 38510 26852
rect 57586 26796 57596 26852
rect 57652 26796 58156 26852
rect 58212 26796 58222 26852
rect 22754 26684 22764 26740
rect 22820 26684 31164 26740
rect 31220 26684 31230 26740
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 17154 26572 17164 26628
rect 17220 26572 17500 26628
rect 17556 26572 17566 26628
rect 23426 26572 23436 26628
rect 23492 26572 24108 26628
rect 24164 26572 24174 26628
rect 27682 26572 27692 26628
rect 27748 26572 31836 26628
rect 31892 26572 31902 26628
rect 32060 26516 32116 26796
rect 50546 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50830 26684
rect 33394 26572 33404 26628
rect 33460 26572 44940 26628
rect 44996 26572 45006 26628
rect 4274 26460 4284 26516
rect 4340 26460 8652 26516
rect 8708 26460 8718 26516
rect 26852 26460 29148 26516
rect 29204 26460 30044 26516
rect 30100 26460 31276 26516
rect 31332 26460 31342 26516
rect 32060 26460 40348 26516
rect 40404 26460 40414 26516
rect 49074 26460 49084 26516
rect 49140 26460 55580 26516
rect 55636 26460 55646 26516
rect 26852 26404 26908 26460
rect 12898 26348 12908 26404
rect 12964 26348 16268 26404
rect 16324 26348 16334 26404
rect 16482 26348 16492 26404
rect 16548 26348 16828 26404
rect 16884 26348 26908 26404
rect 28578 26348 28588 26404
rect 28644 26348 29260 26404
rect 29316 26348 29326 26404
rect 30706 26348 30716 26404
rect 30772 26348 32396 26404
rect 32452 26348 32462 26404
rect 32620 26348 38780 26404
rect 38836 26348 41132 26404
rect 41188 26348 41198 26404
rect 43362 26348 43372 26404
rect 43428 26348 44156 26404
rect 44212 26348 44222 26404
rect 0 26292 800 26320
rect 32620 26292 32676 26348
rect 59200 26292 60000 26320
rect 0 26236 1988 26292
rect 11554 26236 11564 26292
rect 11620 26236 12460 26292
rect 12516 26236 15708 26292
rect 15764 26236 17836 26292
rect 17892 26236 17902 26292
rect 31602 26236 31612 26292
rect 31668 26236 32060 26292
rect 32116 26236 32126 26292
rect 32396 26236 32676 26292
rect 35186 26236 35196 26292
rect 35252 26236 36988 26292
rect 37044 26236 37054 26292
rect 38444 26236 39004 26292
rect 39060 26236 39070 26292
rect 41010 26236 41020 26292
rect 41076 26236 42588 26292
rect 42644 26236 42654 26292
rect 48178 26236 48188 26292
rect 48244 26236 48860 26292
rect 48916 26236 52108 26292
rect 52164 26236 52174 26292
rect 57922 26236 57932 26292
rect 57988 26236 60000 26292
rect 0 26208 800 26236
rect 1932 26180 1988 26236
rect 1922 26124 1932 26180
rect 1988 26124 1998 26180
rect 4274 26124 4284 26180
rect 4340 26124 12908 26180
rect 12964 26124 12974 26180
rect 22418 26124 22428 26180
rect 22484 26124 23660 26180
rect 23716 26124 23726 26180
rect 32396 26068 32452 26236
rect 38444 26068 38500 26236
rect 59200 26208 60000 26236
rect 15250 26012 15260 26068
rect 15316 26012 29036 26068
rect 29092 26012 29102 26068
rect 29586 26012 29596 26068
rect 29652 26012 32452 26068
rect 32732 26012 38500 26068
rect 38994 26012 39004 26068
rect 39060 26012 42700 26068
rect 42756 26012 42766 26068
rect 23202 25900 23212 25956
rect 23268 25900 28252 25956
rect 28308 25900 28318 25956
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 32732 25844 32788 26012
rect 42578 25900 42588 25956
rect 42644 25900 43820 25956
rect 43876 25900 55580 25956
rect 55636 25900 55646 25956
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 14242 25788 14252 25844
rect 14308 25788 20300 25844
rect 20356 25788 22876 25844
rect 22932 25788 22942 25844
rect 23100 25788 32788 25844
rect 39900 25788 41356 25844
rect 41412 25788 41422 25844
rect 23100 25732 23156 25788
rect 39900 25732 39956 25788
rect 14130 25676 14140 25732
rect 14196 25676 16716 25732
rect 16772 25676 23156 25732
rect 24994 25676 25004 25732
rect 25060 25676 25900 25732
rect 25956 25676 25966 25732
rect 29698 25676 29708 25732
rect 29764 25676 39956 25732
rect 40114 25676 40124 25732
rect 40180 25676 41132 25732
rect 41188 25676 41198 25732
rect 0 25620 800 25648
rect 59200 25620 60000 25648
rect 0 25564 1932 25620
rect 1988 25564 1998 25620
rect 9548 25564 13468 25620
rect 13524 25564 13534 25620
rect 15092 25564 17388 25620
rect 17444 25564 17454 25620
rect 17826 25564 17836 25620
rect 17892 25564 21868 25620
rect 21924 25564 23100 25620
rect 23156 25564 23166 25620
rect 27906 25564 27916 25620
rect 27972 25564 28924 25620
rect 28980 25564 28990 25620
rect 36418 25564 36428 25620
rect 36484 25564 36764 25620
rect 36820 25564 37212 25620
rect 37268 25564 55132 25620
rect 55188 25564 55198 25620
rect 57922 25564 57932 25620
rect 57988 25564 60000 25620
rect 0 25536 800 25564
rect 9548 25508 9604 25564
rect 15092 25508 15148 25564
rect 59200 25536 60000 25564
rect 4274 25452 4284 25508
rect 4340 25452 9548 25508
rect 9604 25452 9614 25508
rect 12786 25452 12796 25508
rect 12852 25452 15148 25508
rect 16594 25452 16604 25508
rect 16660 25452 17276 25508
rect 17332 25452 17342 25508
rect 18386 25452 18396 25508
rect 18452 25452 19740 25508
rect 19796 25452 19806 25508
rect 20066 25452 20076 25508
rect 20132 25452 22204 25508
rect 22260 25452 22270 25508
rect 29474 25452 29484 25508
rect 29540 25452 30492 25508
rect 30548 25452 32116 25508
rect 38098 25452 38108 25508
rect 38164 25452 39004 25508
rect 39060 25452 39070 25508
rect 19292 25396 19348 25452
rect 32060 25396 32116 25452
rect 10770 25340 10780 25396
rect 10836 25340 12460 25396
rect 12516 25340 12526 25396
rect 19282 25340 19292 25396
rect 19348 25340 19358 25396
rect 22642 25340 22652 25396
rect 22708 25340 25676 25396
rect 25732 25340 25742 25396
rect 26338 25340 26348 25396
rect 26404 25340 28252 25396
rect 28308 25340 28318 25396
rect 30706 25340 30716 25396
rect 30772 25340 31612 25396
rect 31668 25340 31678 25396
rect 32060 25340 38892 25396
rect 38948 25340 38958 25396
rect 39778 25340 39788 25396
rect 39844 25340 43036 25396
rect 43092 25340 43932 25396
rect 43988 25340 43998 25396
rect 45378 25340 45388 25396
rect 45444 25340 45836 25396
rect 45892 25340 46172 25396
rect 46228 25340 46238 25396
rect 8642 25228 8652 25284
rect 8708 25228 12124 25284
rect 12180 25228 12190 25284
rect 12338 25228 12348 25284
rect 12404 25228 13132 25284
rect 13188 25228 13692 25284
rect 13748 25228 13758 25284
rect 26348 25172 26404 25340
rect 28354 25228 28364 25284
rect 28420 25228 28430 25284
rect 28578 25228 28588 25284
rect 28644 25228 29148 25284
rect 29204 25228 30940 25284
rect 30996 25228 31006 25284
rect 32274 25228 32284 25284
rect 32340 25228 32956 25284
rect 33012 25228 33022 25284
rect 44482 25228 44492 25284
rect 44548 25228 46284 25284
rect 46340 25228 46350 25284
rect 50372 25228 57820 25284
rect 57876 25228 57886 25284
rect 28364 25172 28420 25228
rect 50372 25172 50428 25228
rect 19058 25116 19068 25172
rect 19124 25116 19516 25172
rect 19572 25116 19582 25172
rect 23538 25116 23548 25172
rect 23604 25116 24444 25172
rect 24500 25116 26404 25172
rect 27346 25116 27356 25172
rect 27412 25116 28420 25172
rect 34066 25116 34076 25172
rect 34132 25116 36876 25172
rect 36932 25116 36942 25172
rect 41346 25116 41356 25172
rect 41412 25116 44940 25172
rect 44996 25116 46060 25172
rect 46116 25116 46126 25172
rect 46498 25116 46508 25172
rect 46564 25116 50428 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 50546 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50830 25116
rect 20188 25004 28588 25060
rect 28644 25004 28654 25060
rect 30370 25004 30380 25060
rect 30436 25004 32060 25060
rect 32116 25004 33404 25060
rect 33460 25004 33470 25060
rect 33730 25004 33740 25060
rect 33796 25004 34188 25060
rect 34244 25004 34254 25060
rect 0 24948 800 24976
rect 20188 24948 20244 25004
rect 59200 24948 60000 24976
rect 0 24892 1932 24948
rect 1988 24892 1998 24948
rect 4274 24892 4284 24948
rect 4340 24892 4732 24948
rect 4788 24892 14252 24948
rect 14308 24892 14318 24948
rect 18722 24892 18732 24948
rect 18788 24892 19516 24948
rect 19572 24892 20244 24948
rect 23762 24892 23772 24948
rect 23828 24892 24220 24948
rect 24276 24892 25564 24948
rect 25620 24892 26684 24948
rect 26740 24892 26750 24948
rect 27234 24892 27244 24948
rect 27300 24892 27804 24948
rect 27860 24892 27870 24948
rect 28018 24892 28028 24948
rect 28084 24892 31836 24948
rect 31892 24892 31902 24948
rect 32722 24892 32732 24948
rect 32788 24892 33516 24948
rect 33572 24892 33582 24948
rect 35522 24892 35532 24948
rect 35588 24892 38892 24948
rect 38948 24892 38958 24948
rect 46498 24892 46508 24948
rect 46564 24892 47852 24948
rect 47908 24892 52668 24948
rect 52724 24892 52734 24948
rect 57922 24892 57932 24948
rect 57988 24892 60000 24948
rect 0 24864 800 24892
rect 59200 24864 60000 24892
rect 18834 24780 18844 24836
rect 18900 24780 20300 24836
rect 20356 24780 20366 24836
rect 20626 24780 20636 24836
rect 20692 24780 21084 24836
rect 21140 24780 24332 24836
rect 24388 24780 24398 24836
rect 26338 24780 26348 24836
rect 26404 24780 27468 24836
rect 27524 24780 27972 24836
rect 28802 24780 28812 24836
rect 28868 24780 30828 24836
rect 30884 24780 30894 24836
rect 39218 24780 39228 24836
rect 39284 24780 40236 24836
rect 40292 24780 40302 24836
rect 43922 24780 43932 24836
rect 43988 24780 47516 24836
rect 47572 24780 48636 24836
rect 48692 24780 48702 24836
rect 27916 24724 27972 24780
rect 19842 24668 19852 24724
rect 19908 24668 21532 24724
rect 21588 24668 21598 24724
rect 25442 24668 25452 24724
rect 25508 24668 27356 24724
rect 27412 24668 27422 24724
rect 27906 24668 27916 24724
rect 27972 24668 27982 24724
rect 29698 24668 29708 24724
rect 29764 24668 41132 24724
rect 41188 24668 41198 24724
rect 45154 24668 45164 24724
rect 45220 24668 46956 24724
rect 47012 24668 47022 24724
rect 12562 24556 12572 24612
rect 12628 24556 24668 24612
rect 24724 24556 24734 24612
rect 25330 24556 25340 24612
rect 25396 24556 26908 24612
rect 27794 24556 27804 24612
rect 27860 24556 29484 24612
rect 29540 24556 29550 24612
rect 40674 24556 40684 24612
rect 40740 24556 41916 24612
rect 41972 24556 41982 24612
rect 25340 24388 25396 24556
rect 5282 24332 5292 24388
rect 5348 24332 21308 24388
rect 21364 24332 21374 24388
rect 24770 24332 24780 24388
rect 24836 24332 25396 24388
rect 26852 24388 26908 24556
rect 27234 24444 27244 24500
rect 27300 24444 29148 24500
rect 29204 24444 29214 24500
rect 36194 24444 36204 24500
rect 36260 24444 37548 24500
rect 37604 24444 37614 24500
rect 55346 24444 55356 24500
rect 26852 24332 29596 24388
rect 29652 24332 29662 24388
rect 30034 24332 30044 24388
rect 30100 24332 34636 24388
rect 34692 24332 34702 24388
rect 37426 24332 37436 24388
rect 37492 24332 53452 24388
rect 53508 24332 53518 24388
rect 0 24276 800 24304
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 55412 24276 55468 24500
rect 59200 24276 60000 24304
rect 0 24220 1932 24276
rect 1988 24220 1998 24276
rect 33506 24220 33516 24276
rect 33572 24220 34188 24276
rect 34244 24220 34254 24276
rect 55412 24220 60000 24276
rect 0 24192 800 24220
rect 59200 24192 60000 24220
rect 22754 24108 22764 24164
rect 22820 24108 24444 24164
rect 24500 24108 24510 24164
rect 24994 24108 25004 24164
rect 25060 24108 28028 24164
rect 28084 24108 28094 24164
rect 33282 24108 33292 24164
rect 33348 24108 33964 24164
rect 34020 24108 34748 24164
rect 34804 24108 34814 24164
rect 4274 23996 4284 24052
rect 4340 23996 20636 24052
rect 20692 23996 20702 24052
rect 25330 23996 25340 24052
rect 25396 23996 28420 24052
rect 28578 23996 28588 24052
rect 28644 23996 31276 24052
rect 31332 23996 31342 24052
rect 32050 23996 32060 24052
rect 32116 23996 33740 24052
rect 33796 23996 33806 24052
rect 34962 23996 34972 24052
rect 35028 23996 35644 24052
rect 35700 23996 35710 24052
rect 39330 23996 39340 24052
rect 39396 23996 40908 24052
rect 40964 23996 40974 24052
rect 28364 23940 28420 23996
rect 6962 23884 6972 23940
rect 7028 23884 10108 23940
rect 10164 23884 10174 23940
rect 14018 23884 14028 23940
rect 14084 23884 16828 23940
rect 16884 23884 16894 23940
rect 19058 23884 19068 23940
rect 19124 23884 19740 23940
rect 19796 23884 27244 23940
rect 27300 23884 27310 23940
rect 28364 23884 30604 23940
rect 30660 23884 30670 23940
rect 30818 23884 30828 23940
rect 30884 23884 32172 23940
rect 32228 23884 32238 23940
rect 33506 23884 33516 23940
rect 33572 23884 38556 23940
rect 38612 23884 40236 23940
rect 40292 23884 40302 23940
rect 41458 23884 41468 23940
rect 41524 23884 45612 23940
rect 45668 23884 45678 23940
rect 3042 23772 3052 23828
rect 3108 23772 4620 23828
rect 4676 23772 4686 23828
rect 8530 23772 8540 23828
rect 8596 23772 14252 23828
rect 14308 23772 14588 23828
rect 14644 23772 14654 23828
rect 21298 23772 21308 23828
rect 21364 23772 24332 23828
rect 24388 23772 24668 23828
rect 24724 23772 24734 23828
rect 25666 23772 25676 23828
rect 25732 23772 27020 23828
rect 27076 23772 27692 23828
rect 27748 23772 27758 23828
rect 29922 23772 29932 23828
rect 29988 23772 32956 23828
rect 33012 23772 34748 23828
rect 34804 23772 34814 23828
rect 46386 23772 46396 23828
rect 46452 23772 46462 23828
rect 46610 23772 46620 23828
rect 46676 23772 49756 23828
rect 49812 23772 49822 23828
rect 4274 23660 4284 23716
rect 4340 23660 4844 23716
rect 4900 23660 6636 23716
rect 6692 23660 6702 23716
rect 11106 23660 11116 23716
rect 11172 23660 11788 23716
rect 11844 23660 11854 23716
rect 26852 23660 29372 23716
rect 29428 23660 29438 23716
rect 30034 23660 30044 23716
rect 30100 23660 30940 23716
rect 30996 23660 31612 23716
rect 31668 23660 31678 23716
rect 31826 23660 31836 23716
rect 31892 23660 37548 23716
rect 37604 23660 37614 23716
rect 0 23604 800 23632
rect 26852 23604 26908 23660
rect 46396 23604 46452 23772
rect 59200 23604 60000 23632
rect 0 23548 1932 23604
rect 1988 23548 1998 23604
rect 21522 23548 21532 23604
rect 21588 23548 23492 23604
rect 24770 23548 24780 23604
rect 24836 23548 26908 23604
rect 28354 23548 28364 23604
rect 28420 23548 39228 23604
rect 39284 23548 39294 23604
rect 43708 23548 46452 23604
rect 58044 23548 60000 23604
rect 0 23520 800 23548
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 23436 23492 23492 23548
rect 23436 23436 24220 23492
rect 24276 23436 25228 23492
rect 25284 23436 25294 23492
rect 26786 23436 26796 23492
rect 13794 23324 13804 23380
rect 13860 23324 15148 23380
rect 15204 23324 15484 23380
rect 15540 23324 15550 23380
rect 25228 23268 25284 23436
rect 26852 23324 26908 23492
rect 31154 23436 31164 23492
rect 31220 23436 31724 23492
rect 31780 23436 32620 23492
rect 32676 23436 38388 23492
rect 38332 23380 38388 23436
rect 43708 23380 43764 23548
rect 50546 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50830 23548
rect 58044 23492 58100 23548
rect 59200 23520 60000 23548
rect 57922 23436 57932 23492
rect 57988 23436 58100 23492
rect 26964 23324 26974 23380
rect 37650 23324 37660 23380
rect 37716 23324 37726 23380
rect 38322 23324 38332 23380
rect 38388 23324 38398 23380
rect 38546 23324 38556 23380
rect 38612 23324 43764 23380
rect 37660 23268 37716 23324
rect 16146 23212 16156 23268
rect 16212 23212 20412 23268
rect 20468 23212 24444 23268
rect 24500 23212 24510 23268
rect 25228 23212 32172 23268
rect 32228 23212 32238 23268
rect 32386 23212 32396 23268
rect 32452 23212 33516 23268
rect 33572 23212 33582 23268
rect 37660 23212 39452 23268
rect 39508 23212 39518 23268
rect 32396 23156 32452 23212
rect 4274 23100 4284 23156
rect 4340 23100 5292 23156
rect 5348 23100 5358 23156
rect 11218 23100 11228 23156
rect 11284 23100 13468 23156
rect 13524 23100 13534 23156
rect 16706 23100 16716 23156
rect 16772 23100 22428 23156
rect 22484 23100 22494 23156
rect 26786 23100 26796 23156
rect 3378 22988 3388 23044
rect 3444 22988 4732 23044
rect 4788 22988 4798 23044
rect 16482 22988 16492 23044
rect 16548 22988 18508 23044
rect 18564 22988 18574 23044
rect 22530 22988 22540 23044
rect 22596 22988 26124 23044
rect 26180 22988 26190 23044
rect 26852 22988 26908 23156
rect 27132 23100 32452 23156
rect 34626 23100 34636 23156
rect 34692 23100 38108 23156
rect 38164 23100 38174 23156
rect 38770 23100 38780 23156
rect 38836 23100 41244 23156
rect 41300 23100 42252 23156
rect 42308 23100 44604 23156
rect 44660 23100 45724 23156
rect 45780 23100 46172 23156
rect 46228 23100 47964 23156
rect 48020 23100 48030 23156
rect 27132 23044 27188 23100
rect 26964 22988 27188 23044
rect 28914 22988 28924 23044
rect 28980 22988 29596 23044
rect 29652 22988 31948 23044
rect 32004 22988 37324 23044
rect 37380 22988 37390 23044
rect 37874 22988 37884 23044
rect 37940 22988 39004 23044
rect 39060 22988 39070 23044
rect 39666 22988 39676 23044
rect 39732 22988 42140 23044
rect 42196 22988 42206 23044
rect 46274 22988 46284 23044
rect 46340 22988 47516 23044
rect 47572 22988 53452 23044
rect 53508 22988 53518 23044
rect 59200 22932 60000 22960
rect 4834 22876 4844 22932
rect 4900 22876 7868 22932
rect 7924 22876 7934 22932
rect 11106 22876 11116 22932
rect 11172 22876 12124 22932
rect 12180 22876 12190 22932
rect 18610 22876 18620 22932
rect 18676 22876 18686 22932
rect 19282 22876 19292 22932
rect 19348 22876 27244 22932
rect 27300 22876 27310 22932
rect 55346 22876 55356 22932
rect 55412 22876 60000 22932
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 18620 22708 18676 22876
rect 59200 22848 60000 22876
rect 39554 22764 39564 22820
rect 39620 22764 40012 22820
rect 40068 22764 40078 22820
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 18620 22652 28588 22708
rect 28644 22652 28654 22708
rect 35970 22652 35980 22708
rect 36036 22652 52668 22708
rect 52724 22652 52734 22708
rect 3332 22540 4732 22596
rect 4788 22540 5628 22596
rect 5684 22540 5694 22596
rect 7186 22540 7196 22596
rect 7252 22540 8428 22596
rect 8484 22540 8494 22596
rect 22754 22540 22764 22596
rect 22820 22540 24108 22596
rect 24164 22540 24174 22596
rect 35410 22540 35420 22596
rect 35476 22540 37884 22596
rect 37940 22540 37950 22596
rect 38994 22540 39004 22596
rect 39060 22540 40012 22596
rect 40068 22540 40078 22596
rect 42466 22540 42476 22596
rect 42532 22540 44156 22596
rect 44212 22540 44222 22596
rect 3332 22372 3388 22540
rect 4498 22428 4508 22484
rect 4564 22428 5068 22484
rect 5124 22428 6188 22484
rect 6244 22428 6254 22484
rect 12114 22428 12124 22484
rect 12180 22428 13580 22484
rect 13636 22428 13646 22484
rect 14914 22428 14924 22484
rect 14980 22428 15708 22484
rect 15764 22428 15774 22484
rect 16594 22428 16604 22484
rect 16660 22428 22876 22484
rect 22932 22428 22942 22484
rect 26450 22428 26460 22484
rect 26516 22428 33180 22484
rect 33236 22428 33246 22484
rect 36978 22428 36988 22484
rect 37044 22428 38108 22484
rect 38164 22428 38174 22484
rect 38658 22428 38668 22484
rect 38724 22428 39956 22484
rect 40898 22428 40908 22484
rect 40964 22428 41244 22484
rect 41300 22428 43036 22484
rect 43092 22428 43102 22484
rect 49746 22428 49756 22484
rect 49812 22428 53564 22484
rect 53620 22428 53630 22484
rect 39900 22372 39956 22428
rect 2258 22316 2268 22372
rect 2324 22316 2828 22372
rect 2884 22316 3388 22372
rect 12562 22316 12572 22372
rect 12628 22316 14028 22372
rect 14084 22316 14252 22372
rect 14308 22316 14318 22372
rect 14466 22316 14476 22372
rect 14532 22316 23884 22372
rect 23940 22316 25900 22372
rect 25956 22316 30828 22372
rect 30884 22316 30894 22372
rect 35186 22316 35196 22372
rect 35252 22316 37212 22372
rect 37268 22316 37278 22372
rect 37650 22316 37660 22372
rect 37716 22316 39564 22372
rect 39620 22316 39630 22372
rect 39890 22316 39900 22372
rect 39956 22316 39966 22372
rect 40226 22316 40236 22372
rect 40292 22316 42700 22372
rect 42756 22316 45164 22372
rect 45220 22316 46396 22372
rect 46452 22316 46956 22372
rect 47012 22316 47022 22372
rect 52098 22316 52108 22372
rect 52164 22316 55580 22372
rect 55636 22316 55646 22372
rect 59200 22260 60000 22288
rect 2482 22204 2492 22260
rect 2548 22204 4172 22260
rect 4228 22204 4238 22260
rect 6514 22204 6524 22260
rect 6580 22204 8316 22260
rect 8372 22204 8876 22260
rect 8932 22204 8942 22260
rect 17490 22204 17500 22260
rect 17556 22204 18172 22260
rect 18228 22204 18238 22260
rect 28700 22204 41244 22260
rect 41300 22204 41310 22260
rect 41794 22204 41804 22260
rect 41860 22204 42588 22260
rect 42644 22204 42654 22260
rect 44146 22204 44156 22260
rect 44212 22204 45500 22260
rect 45556 22204 45566 22260
rect 57922 22204 57932 22260
rect 57988 22204 60000 22260
rect 28700 22148 28756 22204
rect 59200 22176 60000 22204
rect 10210 22092 10220 22148
rect 10276 22092 12124 22148
rect 12180 22092 12190 22148
rect 17602 22092 17612 22148
rect 17668 22092 17948 22148
rect 18004 22092 18014 22148
rect 28690 22092 28700 22148
rect 28756 22092 28766 22148
rect 34066 22092 34076 22148
rect 34132 22092 35756 22148
rect 35812 22092 35822 22148
rect 36082 22092 36092 22148
rect 36148 22092 37548 22148
rect 37604 22092 38220 22148
rect 38276 22092 38286 22148
rect 38994 22092 39004 22148
rect 39060 22092 41468 22148
rect 41524 22092 41534 22148
rect 6626 21980 6636 22036
rect 6692 21980 11004 22036
rect 11060 21980 11070 22036
rect 34178 21980 34188 22036
rect 34244 21980 35420 22036
rect 35476 21980 35486 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 50546 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50830 21980
rect 17714 21868 17724 21924
rect 17780 21868 18732 21924
rect 18788 21868 18798 21924
rect 25554 21868 25564 21924
rect 25620 21868 26460 21924
rect 26516 21868 26526 21924
rect 35186 21868 35196 21924
rect 35252 21868 36316 21924
rect 36372 21868 36382 21924
rect 39890 21868 39900 21924
rect 39956 21868 39966 21924
rect 42578 21868 42588 21924
rect 42644 21868 43596 21924
rect 43652 21868 44268 21924
rect 44324 21868 44828 21924
rect 44884 21868 44894 21924
rect 39900 21812 39956 21868
rect 3154 21756 3164 21812
rect 3220 21756 5068 21812
rect 5124 21756 5134 21812
rect 14690 21756 14700 21812
rect 14756 21756 15148 21812
rect 15204 21756 15932 21812
rect 15988 21756 15998 21812
rect 25666 21756 25676 21812
rect 25732 21756 27020 21812
rect 27076 21756 27086 21812
rect 30594 21756 30604 21812
rect 30660 21756 34412 21812
rect 34468 21756 34478 21812
rect 39900 21756 40348 21812
rect 40404 21756 40414 21812
rect 2258 21644 2268 21700
rect 2324 21644 3052 21700
rect 3108 21644 3612 21700
rect 3668 21644 3678 21700
rect 8530 21644 8540 21700
rect 8596 21644 12348 21700
rect 12404 21644 12414 21700
rect 13570 21644 13580 21700
rect 13636 21644 20748 21700
rect 20804 21644 21644 21700
rect 21700 21644 21710 21700
rect 23650 21644 23660 21700
rect 23716 21644 25340 21700
rect 25396 21644 28812 21700
rect 28868 21644 29820 21700
rect 29876 21644 30156 21700
rect 30212 21644 32060 21700
rect 32116 21644 32508 21700
rect 32564 21644 33068 21700
rect 33124 21644 33134 21700
rect 38658 21644 38668 21700
rect 38724 21644 39228 21700
rect 39284 21644 39676 21700
rect 39732 21644 55468 21700
rect 55524 21644 55534 21700
rect 59200 21588 60000 21616
rect 2706 21532 2716 21588
rect 2772 21532 3276 21588
rect 3332 21532 4620 21588
rect 4676 21532 4686 21588
rect 4834 21532 4844 21588
rect 4900 21532 4910 21588
rect 43810 21532 43820 21588
rect 43876 21532 53452 21588
rect 53508 21532 53518 21588
rect 55010 21532 55020 21588
rect 55076 21532 60000 21588
rect 4844 21476 4900 21532
rect 59200 21504 60000 21532
rect 2930 21420 2940 21476
rect 2996 21420 4900 21476
rect 8082 21420 8092 21476
rect 8148 21420 8652 21476
rect 8708 21420 10108 21476
rect 10164 21420 10174 21476
rect 4274 21308 4284 21364
rect 4340 21308 5180 21364
rect 5236 21308 6188 21364
rect 6244 21308 6254 21364
rect 41682 21308 41692 21364
rect 41748 21308 43036 21364
rect 43092 21308 43102 21364
rect 14130 21196 14140 21252
rect 14196 21196 16212 21252
rect 24658 21196 24668 21252
rect 24724 21196 26796 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 16156 21028 16212 21196
rect 26852 21140 26908 21252
rect 28130 21196 28140 21252
rect 28196 21196 29260 21252
rect 29316 21196 29326 21252
rect 32050 21196 32060 21252
rect 32116 21196 33964 21252
rect 34020 21196 34030 21252
rect 32060 21140 32116 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 26852 21084 32116 21140
rect 12338 20972 12348 21028
rect 12404 20972 15148 21028
rect 16146 20972 16156 21028
rect 16212 20972 16222 21028
rect 27010 20972 27020 21028
rect 27076 20972 28140 21028
rect 28196 20972 28206 21028
rect 33964 20972 34972 21028
rect 35028 20972 35038 21028
rect 15092 20916 15148 20972
rect 33964 20916 34020 20972
rect 59200 20916 60000 20944
rect 15092 20860 21420 20916
rect 21476 20860 21486 20916
rect 30380 20860 33964 20916
rect 34020 20860 34030 20916
rect 34850 20860 34860 20916
rect 34916 20860 35980 20916
rect 36036 20860 36988 20916
rect 37044 20860 37054 20916
rect 41122 20860 41132 20916
rect 41188 20860 41692 20916
rect 41748 20860 53676 20916
rect 53732 20860 53742 20916
rect 55346 20860 55356 20916
rect 55412 20860 60000 20916
rect 30380 20804 30436 20860
rect 59200 20832 60000 20860
rect 13916 20748 14812 20804
rect 14868 20748 15596 20804
rect 15652 20748 15662 20804
rect 17378 20748 17388 20804
rect 17444 20748 17948 20804
rect 18004 20748 18014 20804
rect 22082 20748 22092 20804
rect 22148 20748 22988 20804
rect 23044 20748 23996 20804
rect 24052 20748 24062 20804
rect 27580 20748 30380 20804
rect 30436 20748 30446 20804
rect 33282 20748 33292 20804
rect 33348 20748 35420 20804
rect 35476 20748 35486 20804
rect 38210 20748 38220 20804
rect 38276 20748 38668 20804
rect 13916 20692 13972 20748
rect 27580 20692 27636 20748
rect 38612 20692 38668 20748
rect 13906 20636 13916 20692
rect 13972 20636 13982 20692
rect 19730 20636 19740 20692
rect 19796 20636 21196 20692
rect 21252 20636 21262 20692
rect 22530 20636 22540 20692
rect 22596 20636 23100 20692
rect 23156 20636 25452 20692
rect 25508 20636 25518 20692
rect 27570 20636 27580 20692
rect 27636 20636 27646 20692
rect 27794 20636 27804 20692
rect 27860 20636 29036 20692
rect 29092 20636 29102 20692
rect 29362 20636 29372 20692
rect 29428 20636 31164 20692
rect 31220 20636 38276 20692
rect 38612 20636 42028 20692
rect 42084 20636 43148 20692
rect 43204 20636 43214 20692
rect 4610 20524 4620 20580
rect 4676 20524 5740 20580
rect 5796 20524 7084 20580
rect 7140 20524 7150 20580
rect 10210 20524 10220 20580
rect 10276 20524 11004 20580
rect 11060 20524 11564 20580
rect 11620 20524 11630 20580
rect 18722 20524 18732 20580
rect 18788 20524 19180 20580
rect 19236 20524 25676 20580
rect 25732 20524 25742 20580
rect 26114 20524 26124 20580
rect 26180 20524 26908 20580
rect 26964 20524 26974 20580
rect 28242 20524 28252 20580
rect 28308 20524 28924 20580
rect 28980 20524 28990 20580
rect 29138 20524 29148 20580
rect 29204 20524 34636 20580
rect 34692 20524 34702 20580
rect 34962 20524 34972 20580
rect 35028 20524 36540 20580
rect 36596 20524 37996 20580
rect 38052 20524 38062 20580
rect 28252 20468 28308 20524
rect 8194 20412 8204 20468
rect 8260 20412 14588 20468
rect 14644 20412 15820 20468
rect 15876 20412 15886 20468
rect 26226 20412 26236 20468
rect 26292 20412 28308 20468
rect 38220 20468 38276 20636
rect 38220 20412 41356 20468
rect 41412 20412 41422 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 50546 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50830 20412
rect 25890 20300 25900 20356
rect 25956 20300 29820 20356
rect 29876 20300 29886 20356
rect 59200 20244 60000 20272
rect 3042 20188 3052 20244
rect 3108 20188 3500 20244
rect 3556 20188 3566 20244
rect 5506 20188 5516 20244
rect 5572 20188 6412 20244
rect 6468 20188 6478 20244
rect 14466 20188 14476 20244
rect 14532 20188 15092 20244
rect 23874 20188 23884 20244
rect 23940 20188 26012 20244
rect 26068 20188 26078 20244
rect 31042 20188 31052 20244
rect 31108 20188 32060 20244
rect 32116 20188 32126 20244
rect 57932 20188 60000 20244
rect 15036 20132 15092 20188
rect 57932 20132 57988 20188
rect 59200 20160 60000 20188
rect 14242 20076 14252 20132
rect 14308 20076 14980 20132
rect 15036 20076 15260 20132
rect 15316 20076 15326 20132
rect 16258 20076 16268 20132
rect 16324 20076 16940 20132
rect 16996 20076 18060 20132
rect 18116 20076 20916 20132
rect 23202 20076 23212 20132
rect 23268 20076 24556 20132
rect 24612 20076 26124 20132
rect 26180 20076 26190 20132
rect 26852 20076 27020 20132
rect 27076 20076 27086 20132
rect 27682 20076 27692 20132
rect 27748 20076 31948 20132
rect 32004 20076 32014 20132
rect 35634 20076 35644 20132
rect 35700 20076 36316 20132
rect 36372 20076 38780 20132
rect 38836 20076 39452 20132
rect 39508 20076 39518 20132
rect 40226 20076 40236 20132
rect 40292 20076 40908 20132
rect 40964 20076 40974 20132
rect 57922 20076 57932 20132
rect 57988 20076 57998 20132
rect 14924 20020 14980 20076
rect 20860 20020 20916 20076
rect 26852 20020 26908 20076
rect 4722 19964 4732 20020
rect 4788 19964 5516 20020
rect 5572 19964 6636 20020
rect 6692 19964 6702 20020
rect 14690 19964 14700 20020
rect 14756 19964 14766 20020
rect 14924 19964 17276 20020
rect 17332 19964 17342 20020
rect 17602 19964 17612 20020
rect 17668 19964 19068 20020
rect 19124 19964 19134 20020
rect 20860 19964 26012 20020
rect 26068 19964 26908 20020
rect 29026 19964 29036 20020
rect 29092 19964 30380 20020
rect 30436 19964 30446 20020
rect 38658 19964 38668 20020
rect 38724 19964 39900 20020
rect 39956 19964 39966 20020
rect 47954 19964 47964 20020
rect 48020 19964 49980 20020
rect 50036 19964 50046 20020
rect 14700 19908 14756 19964
rect 6514 19852 6524 19908
rect 6580 19852 7756 19908
rect 7812 19852 7822 19908
rect 9426 19852 9436 19908
rect 9492 19852 13244 19908
rect 13300 19852 13310 19908
rect 14700 19852 15484 19908
rect 15540 19852 15550 19908
rect 30482 19852 30492 19908
rect 30548 19852 37212 19908
rect 37268 19852 37278 19908
rect 42466 19852 42476 19908
rect 42532 19852 42924 19908
rect 42980 19852 48188 19908
rect 48244 19852 48254 19908
rect 13244 19796 13300 19852
rect 13244 19740 15932 19796
rect 15988 19740 15998 19796
rect 24098 19740 24108 19796
rect 24164 19740 25788 19796
rect 25844 19740 25854 19796
rect 34738 19740 34748 19796
rect 34804 19740 35196 19796
rect 35252 19740 35756 19796
rect 35812 19740 35822 19796
rect 55346 19740 55356 19796
rect 36978 19628 36988 19684
rect 37044 19628 38108 19684
rect 38164 19628 38892 19684
rect 38948 19628 52108 19684
rect 52164 19628 53228 19684
rect 53284 19628 53294 19684
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 55412 19572 55468 19796
rect 59200 19572 60000 19600
rect 55412 19516 60000 19572
rect 59200 19488 60000 19516
rect 11106 19404 11116 19460
rect 11172 19404 12124 19460
rect 12180 19404 12190 19460
rect 15092 19292 20524 19348
rect 20580 19292 21420 19348
rect 21476 19292 21486 19348
rect 23202 19292 23212 19348
rect 23268 19292 27132 19348
rect 27188 19292 27692 19348
rect 27748 19292 28476 19348
rect 28532 19292 28542 19348
rect 39442 19292 39452 19348
rect 39508 19292 42252 19348
rect 42308 19292 42812 19348
rect 42868 19292 43596 19348
rect 43652 19292 44268 19348
rect 44324 19292 44828 19348
rect 44884 19292 46508 19348
rect 46564 19292 46574 19348
rect 4498 19180 4508 19236
rect 4564 19180 5068 19236
rect 5124 19180 5134 19236
rect 11330 19180 11340 19236
rect 11396 19180 12572 19236
rect 12628 19180 12638 19236
rect 15092 19124 15148 19292
rect 18722 19180 18732 19236
rect 18788 19180 19404 19236
rect 19460 19180 19470 19236
rect 20402 19180 20412 19236
rect 20468 19180 21756 19236
rect 21812 19180 21822 19236
rect 28130 19180 28140 19236
rect 28196 19180 29036 19236
rect 29092 19180 29764 19236
rect 49634 19180 49644 19236
rect 49700 19180 55580 19236
rect 55636 19180 55646 19236
rect 29708 19124 29764 19180
rect 2818 19068 2828 19124
rect 2884 19068 3388 19124
rect 3444 19068 3454 19124
rect 4386 19068 4396 19124
rect 4452 19068 5628 19124
rect 5684 19068 5694 19124
rect 7186 19068 7196 19124
rect 7252 19068 7924 19124
rect 11666 19068 11676 19124
rect 11732 19068 15148 19124
rect 19170 19068 19180 19124
rect 19236 19068 19740 19124
rect 19796 19068 19806 19124
rect 25218 19068 25228 19124
rect 25284 19068 25900 19124
rect 25956 19068 25966 19124
rect 27346 19068 27356 19124
rect 27412 19068 28588 19124
rect 28644 19068 28654 19124
rect 29698 19068 29708 19124
rect 29764 19068 29774 19124
rect 36418 19068 36428 19124
rect 36484 19068 37100 19124
rect 37156 19068 37166 19124
rect 4396 19012 4452 19068
rect 7868 19012 7924 19068
rect 2034 18956 2044 19012
rect 2100 18956 4452 19012
rect 5954 18956 5964 19012
rect 6020 18956 7532 19012
rect 7588 18956 7598 19012
rect 7858 18956 7868 19012
rect 7924 18956 12124 19012
rect 12180 18956 18508 19012
rect 18564 18956 19404 19012
rect 19460 18956 19470 19012
rect 28802 18956 28812 19012
rect 28868 18956 29932 19012
rect 29988 18956 30716 19012
rect 30772 18956 30782 19012
rect 0 18900 800 18928
rect 59200 18900 60000 18928
rect 0 18844 1708 18900
rect 1764 18844 1774 18900
rect 4946 18844 4956 18900
rect 5012 18844 9996 18900
rect 10052 18844 11452 18900
rect 11508 18844 11518 18900
rect 13458 18844 13468 18900
rect 13524 18844 17612 18900
rect 17668 18844 17678 18900
rect 57922 18844 57932 18900
rect 57988 18844 60000 18900
rect 0 18816 800 18844
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 50546 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50830 18844
rect 59200 18816 60000 18844
rect 2706 18732 2716 18788
rect 2772 18732 3052 18788
rect 3108 18732 3724 18788
rect 3780 18732 5180 18788
rect 5236 18732 5246 18788
rect 9874 18732 9884 18788
rect 9940 18732 12236 18788
rect 12292 18732 12302 18788
rect 29474 18732 29484 18788
rect 29540 18732 30324 18788
rect 30268 18676 30324 18732
rect 10322 18620 10332 18676
rect 10388 18620 11116 18676
rect 11172 18620 12684 18676
rect 12740 18620 12750 18676
rect 15810 18620 15820 18676
rect 15876 18620 18620 18676
rect 18676 18620 18686 18676
rect 19170 18620 19180 18676
rect 19236 18620 20412 18676
rect 20468 18620 20478 18676
rect 28242 18620 28252 18676
rect 28308 18620 29596 18676
rect 29652 18620 29662 18676
rect 30258 18620 30268 18676
rect 30324 18620 31052 18676
rect 31108 18620 31118 18676
rect 2034 18508 2044 18564
rect 2100 18508 2940 18564
rect 2996 18508 5628 18564
rect 5684 18508 5694 18564
rect 7522 18508 7532 18564
rect 7588 18508 8316 18564
rect 8372 18508 9996 18564
rect 10052 18508 10062 18564
rect 13346 18508 13356 18564
rect 13412 18508 16828 18564
rect 16884 18508 17500 18564
rect 17556 18508 17566 18564
rect 20290 18508 20300 18564
rect 20356 18508 22764 18564
rect 22820 18508 23548 18564
rect 23604 18508 23614 18564
rect 26562 18508 26572 18564
rect 26628 18508 27916 18564
rect 27972 18508 27982 18564
rect 38098 18508 38108 18564
rect 38164 18508 38668 18564
rect 39218 18508 39228 18564
rect 39284 18508 41132 18564
rect 41188 18508 41198 18564
rect 43810 18508 43820 18564
rect 43876 18508 48972 18564
rect 49028 18508 49038 18564
rect 4284 18452 4340 18508
rect 4274 18396 4284 18452
rect 4340 18396 4350 18452
rect 11778 18396 11788 18452
rect 11844 18396 13468 18452
rect 13524 18396 13534 18452
rect 15138 18396 15148 18452
rect 15204 18396 16268 18452
rect 16324 18396 16334 18452
rect 27234 18396 27244 18452
rect 27300 18396 28028 18452
rect 28084 18396 28094 18452
rect 28578 18396 28588 18452
rect 28644 18396 30604 18452
rect 30660 18396 30670 18452
rect 35074 18396 35084 18452
rect 35140 18396 37212 18452
rect 37268 18396 37278 18452
rect 37426 18396 37436 18452
rect 37492 18396 38444 18452
rect 38500 18396 38510 18452
rect 10210 18284 10220 18340
rect 10276 18284 13916 18340
rect 13972 18284 13982 18340
rect 15922 18284 15932 18340
rect 15988 18284 16716 18340
rect 16772 18284 16782 18340
rect 33730 18284 33740 18340
rect 33796 18284 35756 18340
rect 35812 18284 35822 18340
rect 38612 18228 38668 18508
rect 41234 18396 41244 18452
rect 41300 18396 42140 18452
rect 42196 18396 42206 18452
rect 44930 18396 44940 18452
rect 44996 18396 46732 18452
rect 46788 18396 46798 18452
rect 47730 18396 47740 18452
rect 47796 18396 53452 18452
rect 53508 18396 53518 18452
rect 47740 18340 47796 18396
rect 41794 18284 41804 18340
rect 41860 18284 42364 18340
rect 42420 18284 42430 18340
rect 46386 18284 46396 18340
rect 46452 18284 47796 18340
rect 51202 18284 51212 18340
rect 51268 18284 51996 18340
rect 52052 18284 52062 18340
rect 59200 18228 60000 18256
rect 11442 18172 11452 18228
rect 11508 18172 11900 18228
rect 11956 18172 11966 18228
rect 13458 18172 13468 18228
rect 13524 18172 15036 18228
rect 15092 18172 15102 18228
rect 38612 18172 39004 18228
rect 39060 18172 51548 18228
rect 51604 18172 51614 18228
rect 55346 18172 55356 18228
rect 55412 18172 60000 18228
rect 59200 18144 60000 18172
rect 6626 18060 6636 18116
rect 6692 18060 6972 18116
rect 7028 18060 8092 18116
rect 8148 18060 12460 18116
rect 12516 18060 12526 18116
rect 39778 18060 39788 18116
rect 39844 18060 41020 18116
rect 41076 18060 41086 18116
rect 45154 18060 45164 18116
rect 45220 18060 45948 18116
rect 46004 18060 48860 18116
rect 48916 18060 48926 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 51090 17948 51100 18004
rect 51156 17948 51772 18004
rect 51828 17948 51838 18004
rect 3378 17836 3388 17892
rect 3444 17836 3556 17892
rect 4162 17836 4172 17892
rect 4228 17836 4396 17892
rect 4452 17836 6860 17892
rect 6916 17836 7980 17892
rect 8036 17836 8046 17892
rect 22866 17836 22876 17892
rect 22932 17836 23100 17892
rect 23156 17836 23436 17892
rect 23492 17836 23502 17892
rect 29698 17836 29708 17892
rect 29764 17836 37324 17892
rect 37380 17836 37390 17892
rect 38546 17836 38556 17892
rect 38612 17836 50596 17892
rect 50754 17836 50764 17892
rect 50820 17836 52220 17892
rect 52276 17836 52286 17892
rect 3500 17668 3556 17836
rect 50540 17780 50596 17836
rect 26852 17724 27300 17780
rect 31938 17724 31948 17780
rect 32004 17724 34412 17780
rect 34468 17724 34478 17780
rect 36306 17724 36316 17780
rect 36372 17724 38332 17780
rect 38388 17724 38398 17780
rect 45602 17724 45612 17780
rect 45668 17724 46956 17780
rect 47012 17724 47022 17780
rect 48066 17724 48076 17780
rect 48132 17724 48748 17780
rect 48804 17724 48814 17780
rect 50540 17724 55468 17780
rect 3490 17612 3500 17668
rect 3556 17612 3566 17668
rect 5618 17612 5628 17668
rect 5684 17612 7308 17668
rect 7364 17612 7374 17668
rect 10098 17612 10108 17668
rect 10164 17612 13692 17668
rect 13748 17612 13758 17668
rect 16258 17612 16268 17668
rect 16324 17612 17948 17668
rect 18004 17612 18014 17668
rect 22530 17612 22540 17668
rect 22596 17612 23212 17668
rect 23268 17612 23278 17668
rect 26786 17612 26796 17668
rect 26852 17612 26908 17724
rect 27244 17668 27300 17724
rect 55412 17668 55468 17724
rect 27010 17612 27020 17668
rect 27076 17612 27086 17668
rect 27234 17612 27244 17668
rect 27300 17612 27310 17668
rect 37090 17612 37100 17668
rect 37156 17612 39788 17668
rect 39844 17612 39854 17668
rect 45266 17612 45276 17668
rect 45332 17612 52668 17668
rect 52724 17612 52734 17668
rect 55412 17612 55580 17668
rect 55636 17612 55646 17668
rect 0 17556 800 17584
rect 0 17500 1708 17556
rect 1764 17500 1774 17556
rect 9874 17500 9884 17556
rect 9940 17500 10332 17556
rect 10388 17500 10398 17556
rect 19618 17500 19628 17556
rect 19684 17500 20636 17556
rect 20692 17500 21980 17556
rect 22036 17500 22046 17556
rect 24658 17500 24668 17556
rect 24724 17500 26572 17556
rect 26628 17500 26638 17556
rect 0 17472 800 17500
rect 27020 17444 27076 17612
rect 31378 17500 31388 17556
rect 31444 17500 35196 17556
rect 35252 17500 38220 17556
rect 38276 17500 38286 17556
rect 41458 17500 41468 17556
rect 41524 17500 45836 17556
rect 45892 17500 45902 17556
rect 55346 17500 55356 17556
rect 55412 17500 55468 17612
rect 59200 17556 60000 17584
rect 57922 17500 57932 17556
rect 57988 17500 60000 17556
rect 59200 17472 60000 17500
rect 9986 17388 9996 17444
rect 10052 17388 10668 17444
rect 10724 17388 10734 17444
rect 10882 17388 10892 17444
rect 10948 17388 11788 17444
rect 11844 17388 11854 17444
rect 13346 17388 13356 17444
rect 13412 17388 14924 17444
rect 14980 17388 17836 17444
rect 17892 17388 21308 17444
rect 21364 17388 21374 17444
rect 25554 17388 25564 17444
rect 25620 17388 26460 17444
rect 26516 17388 27076 17444
rect 38658 17388 38668 17444
rect 38724 17388 39340 17444
rect 39396 17388 40460 17444
rect 40516 17388 40526 17444
rect 40674 17388 40684 17444
rect 40740 17388 49084 17444
rect 49140 17388 49150 17444
rect 40460 17332 40516 17388
rect 10210 17276 10220 17332
rect 10276 17276 11340 17332
rect 11396 17276 11406 17332
rect 37538 17276 37548 17332
rect 37604 17276 39452 17332
rect 39508 17276 39518 17332
rect 40460 17276 41356 17332
rect 41412 17276 41422 17332
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 50546 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50830 17276
rect 6962 17164 6972 17220
rect 7028 17164 12796 17220
rect 12852 17164 15932 17220
rect 15988 17164 15998 17220
rect 40450 17164 40460 17220
rect 40516 17164 46508 17220
rect 46564 17164 46574 17220
rect 3042 17052 3052 17108
rect 3108 17052 3948 17108
rect 4004 17052 4014 17108
rect 11890 17052 11900 17108
rect 11956 17052 12236 17108
rect 12292 17052 12302 17108
rect 14690 17052 14700 17108
rect 14756 17052 16268 17108
rect 16324 17052 16334 17108
rect 18050 17052 18060 17108
rect 18116 17052 20972 17108
rect 21028 17052 21038 17108
rect 33506 17052 33516 17108
rect 33572 17052 34076 17108
rect 34132 17052 34142 17108
rect 34738 17052 34748 17108
rect 34804 17052 36036 17108
rect 37986 17052 37996 17108
rect 38052 17052 41804 17108
rect 41860 17052 41870 17108
rect 35980 16996 36036 17052
rect 8306 16940 8316 16996
rect 8372 16940 9772 16996
rect 9828 16940 9838 16996
rect 17602 16940 17612 16996
rect 17668 16940 19068 16996
rect 19124 16940 19134 16996
rect 23202 16940 23212 16996
rect 23268 16940 23996 16996
rect 24052 16940 24780 16996
rect 24836 16940 24846 16996
rect 34402 16940 34412 16996
rect 34468 16940 35756 16996
rect 35812 16940 35822 16996
rect 35980 16940 50652 16996
rect 50708 16940 50718 16996
rect 59200 16884 60000 16912
rect 4946 16828 4956 16884
rect 5012 16828 5628 16884
rect 5684 16828 5694 16884
rect 8754 16828 8764 16884
rect 8820 16828 8932 16884
rect 9090 16828 9100 16884
rect 9156 16828 12236 16884
rect 12292 16828 12302 16884
rect 14018 16828 14028 16884
rect 14084 16828 14924 16884
rect 14980 16828 14990 16884
rect 15092 16828 17724 16884
rect 17780 16828 19516 16884
rect 19572 16828 19582 16884
rect 33282 16828 33292 16884
rect 33348 16828 34076 16884
rect 34132 16828 34142 16884
rect 35634 16828 35644 16884
rect 35700 16828 36204 16884
rect 36260 16828 36270 16884
rect 36530 16828 36540 16884
rect 36596 16828 37436 16884
rect 37492 16828 37502 16884
rect 41570 16828 41580 16884
rect 41636 16828 42140 16884
rect 42196 16828 43820 16884
rect 43876 16828 43886 16884
rect 51314 16828 51324 16884
rect 51380 16828 52108 16884
rect 52164 16828 52780 16884
rect 52836 16828 52846 16884
rect 55010 16828 55020 16884
rect 55076 16828 60000 16884
rect 8876 16772 8932 16828
rect 15092 16772 15148 16828
rect 59200 16800 60000 16828
rect 2594 16716 2604 16772
rect 2660 16716 2940 16772
rect 2996 16716 3006 16772
rect 3378 16716 3388 16772
rect 3444 16716 6748 16772
rect 6804 16716 6814 16772
rect 8876 16716 9996 16772
rect 10052 16716 10062 16772
rect 14466 16716 14476 16772
rect 14532 16716 15148 16772
rect 33058 16716 33068 16772
rect 33124 16716 34748 16772
rect 34804 16716 34814 16772
rect 35746 16716 35756 16772
rect 35812 16716 37324 16772
rect 37380 16716 37390 16772
rect 39778 16716 39788 16772
rect 39844 16716 40796 16772
rect 40852 16716 40862 16772
rect 41682 16716 41692 16772
rect 41748 16716 45724 16772
rect 45780 16716 45790 16772
rect 2940 16660 2996 16716
rect 2940 16604 7868 16660
rect 7924 16604 7934 16660
rect 16258 16604 16268 16660
rect 16324 16604 16716 16660
rect 16772 16604 16782 16660
rect 16930 16604 16940 16660
rect 16996 16604 17836 16660
rect 17892 16604 18284 16660
rect 18340 16604 18350 16660
rect 40114 16604 40124 16660
rect 40180 16604 40908 16660
rect 40964 16604 40974 16660
rect 43810 16604 43820 16660
rect 43876 16604 52780 16660
rect 52836 16604 52846 16660
rect 16482 16492 16492 16548
rect 16548 16492 17724 16548
rect 17780 16492 17790 16548
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 12002 16380 12012 16436
rect 12068 16380 12348 16436
rect 12404 16380 18844 16436
rect 18900 16380 18910 16436
rect 37426 16380 37436 16436
rect 37492 16380 38780 16436
rect 38836 16380 40908 16436
rect 40964 16380 40974 16436
rect 6066 16268 6076 16324
rect 6132 16268 6524 16324
rect 6580 16268 10444 16324
rect 10500 16268 14364 16324
rect 14420 16268 14430 16324
rect 14588 16268 15148 16324
rect 15204 16268 15214 16324
rect 16034 16268 16044 16324
rect 16100 16268 16110 16324
rect 20626 16268 20636 16324
rect 20692 16268 23772 16324
rect 23828 16268 25004 16324
rect 25060 16268 25070 16324
rect 31378 16268 31388 16324
rect 31444 16268 32060 16324
rect 32116 16268 32126 16324
rect 38546 16268 38556 16324
rect 38612 16268 41132 16324
rect 41188 16268 41198 16324
rect 0 16212 800 16240
rect 14588 16212 14644 16268
rect 16044 16212 16100 16268
rect 59200 16212 60000 16240
rect 0 16156 1708 16212
rect 1764 16156 1774 16212
rect 12786 16156 12796 16212
rect 12852 16156 14644 16212
rect 14802 16156 14812 16212
rect 14868 16156 16716 16212
rect 16772 16156 16782 16212
rect 31490 16156 31500 16212
rect 31556 16156 32956 16212
rect 33012 16156 33022 16212
rect 42578 16156 42588 16212
rect 42644 16156 43708 16212
rect 43764 16156 43774 16212
rect 55346 16156 55356 16212
rect 55412 16156 60000 16212
rect 0 16128 800 16156
rect 59200 16128 60000 16156
rect 3378 16044 3388 16100
rect 3444 16044 4620 16100
rect 4676 16044 4686 16100
rect 7298 16044 7308 16100
rect 7364 16044 9212 16100
rect 9268 16044 9278 16100
rect 12674 16044 12684 16100
rect 12740 16044 14588 16100
rect 14644 16044 14654 16100
rect 18386 16044 18396 16100
rect 18452 16044 19180 16100
rect 19236 16044 19246 16100
rect 21858 16044 21868 16100
rect 21924 16044 22428 16100
rect 22484 16044 22494 16100
rect 33170 16044 33180 16100
rect 33236 16044 35420 16100
rect 35476 16044 37100 16100
rect 37156 16044 37166 16100
rect 38770 16044 38780 16100
rect 38836 16044 39340 16100
rect 39396 16044 39900 16100
rect 39956 16044 40236 16100
rect 40292 16044 40302 16100
rect 41794 16044 41804 16100
rect 41860 16044 42476 16100
rect 42532 16044 42542 16100
rect 42690 16044 42700 16100
rect 42756 16044 48748 16100
rect 48804 16044 48814 16100
rect 49634 16044 49644 16100
rect 49700 16044 50204 16100
rect 50260 16044 55580 16100
rect 55636 16044 55646 16100
rect 2034 15932 2044 15988
rect 2100 15932 5460 15988
rect 5618 15932 5628 15988
rect 5684 15932 6300 15988
rect 6356 15932 7420 15988
rect 7476 15932 7486 15988
rect 12114 15932 12124 15988
rect 12180 15932 14476 15988
rect 14532 15932 14542 15988
rect 22754 15932 22764 15988
rect 22820 15932 23996 15988
rect 24052 15932 24062 15988
rect 25666 15932 25676 15988
rect 25732 15932 26236 15988
rect 26292 15932 26302 15988
rect 38994 15932 39004 15988
rect 39060 15932 39564 15988
rect 39620 15932 39630 15988
rect 5404 15876 5460 15932
rect 2146 15820 2156 15876
rect 2212 15820 2716 15876
rect 2772 15820 3836 15876
rect 3892 15820 3902 15876
rect 5404 15820 7868 15876
rect 7924 15820 9380 15876
rect 9538 15820 9548 15876
rect 9604 15820 9884 15876
rect 9940 15820 10220 15876
rect 10276 15820 11788 15876
rect 11844 15820 12796 15876
rect 12852 15820 12862 15876
rect 18834 15820 18844 15876
rect 18900 15820 20244 15876
rect 21522 15820 21532 15876
rect 21588 15820 23100 15876
rect 23156 15820 23660 15876
rect 23716 15820 23726 15876
rect 29362 15820 29372 15876
rect 29428 15820 30380 15876
rect 30436 15820 30446 15876
rect 41234 15820 41244 15876
rect 41300 15820 43708 15876
rect 43764 15820 43774 15876
rect 9324 15764 9380 15820
rect 20188 15764 20244 15820
rect 3602 15708 3612 15764
rect 3668 15708 7532 15764
rect 7588 15708 8092 15764
rect 8148 15708 8158 15764
rect 9324 15708 9660 15764
rect 9716 15708 9726 15764
rect 20188 15708 22540 15764
rect 22596 15708 22606 15764
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 50546 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50830 15708
rect 20300 15596 20636 15652
rect 20692 15596 20702 15652
rect 30594 15596 30604 15652
rect 30660 15596 32844 15652
rect 32900 15596 34972 15652
rect 35028 15596 35038 15652
rect 0 15540 800 15568
rect 20300 15540 20356 15596
rect 59200 15540 60000 15568
rect 0 15484 3388 15540
rect 3444 15484 3454 15540
rect 4946 15484 4956 15540
rect 5012 15484 5628 15540
rect 5684 15484 5694 15540
rect 16146 15484 16156 15540
rect 16212 15484 20356 15540
rect 20514 15484 20524 15540
rect 20580 15484 22428 15540
rect 22484 15484 22494 15540
rect 23874 15484 23884 15540
rect 23940 15484 25900 15540
rect 25956 15484 25966 15540
rect 34066 15484 34076 15540
rect 34132 15484 35084 15540
rect 35140 15484 38556 15540
rect 38612 15484 38622 15540
rect 42018 15484 42028 15540
rect 42084 15484 47796 15540
rect 51986 15484 51996 15540
rect 52052 15484 52332 15540
rect 52388 15484 54236 15540
rect 54292 15484 54302 15540
rect 57922 15484 57932 15540
rect 57988 15484 60000 15540
rect 0 15456 800 15484
rect 8642 15372 8652 15428
rect 8708 15372 15596 15428
rect 15652 15372 15932 15428
rect 15988 15372 21196 15428
rect 21252 15372 21262 15428
rect 22642 15372 22652 15428
rect 22708 15372 23996 15428
rect 24052 15372 24062 15428
rect 30034 15372 30044 15428
rect 30100 15372 36988 15428
rect 37044 15372 37772 15428
rect 37828 15372 37838 15428
rect 38612 15372 41132 15428
rect 41188 15372 41198 15428
rect 38612 15316 38668 15372
rect 47740 15316 47796 15484
rect 59200 15456 60000 15484
rect 48178 15372 48188 15428
rect 48244 15372 55468 15428
rect 2594 15260 2604 15316
rect 2660 15260 7868 15316
rect 7924 15260 7934 15316
rect 12786 15260 12796 15316
rect 12852 15260 13692 15316
rect 13748 15260 13758 15316
rect 15138 15260 15148 15316
rect 15204 15260 18284 15316
rect 18340 15260 18350 15316
rect 21298 15260 21308 15316
rect 21364 15260 22204 15316
rect 22260 15260 23548 15316
rect 23604 15260 23614 15316
rect 31490 15260 31500 15316
rect 31556 15260 33180 15316
rect 33236 15260 33246 15316
rect 34962 15260 34972 15316
rect 35028 15260 36092 15316
rect 36148 15260 38668 15316
rect 39330 15260 39340 15316
rect 39396 15260 39900 15316
rect 39956 15260 39966 15316
rect 41570 15260 41580 15316
rect 41636 15260 42476 15316
rect 42532 15260 42542 15316
rect 45042 15260 45052 15316
rect 45108 15260 45388 15316
rect 45444 15260 46396 15316
rect 46452 15260 46462 15316
rect 47058 15260 47068 15316
rect 47124 15260 47516 15316
rect 47572 15260 47582 15316
rect 47740 15260 53452 15316
rect 53508 15260 53518 15316
rect 17714 15148 17724 15204
rect 17780 15148 19292 15204
rect 19348 15148 19358 15204
rect 26338 15148 26348 15204
rect 26404 15148 27356 15204
rect 27412 15148 27422 15204
rect 32946 15148 32956 15204
rect 33012 15148 34468 15204
rect 34412 15092 34468 15148
rect 40012 15148 41356 15204
rect 41412 15148 42252 15204
rect 42308 15148 42318 15204
rect 45266 15148 45276 15204
rect 45332 15148 45724 15204
rect 45780 15148 46508 15204
rect 46564 15148 46574 15204
rect 40012 15092 40068 15148
rect 55412 15092 55468 15372
rect 4274 15036 4284 15092
rect 4340 15036 6748 15092
rect 6804 15036 6814 15092
rect 11218 15036 11228 15092
rect 11284 15036 12684 15092
rect 12740 15036 12750 15092
rect 34402 15036 34412 15092
rect 34468 15036 34478 15092
rect 40002 15036 40012 15092
rect 40068 15036 40078 15092
rect 52434 15036 52444 15092
rect 52500 15036 53340 15092
rect 53396 15036 53406 15092
rect 55412 15036 55580 15092
rect 55636 15036 55646 15092
rect 38322 14924 38332 14980
rect 38388 14924 39004 14980
rect 39060 14924 39676 14980
rect 39732 14924 39742 14980
rect 0 14868 800 14896
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 59200 14868 60000 14896
rect 0 14812 1820 14868
rect 1876 14812 1886 14868
rect 40898 14812 40908 14868
rect 40964 14812 50428 14868
rect 52882 14812 52892 14868
rect 52948 14812 54124 14868
rect 54180 14812 54190 14868
rect 55346 14812 55356 14868
rect 55412 14812 60000 14868
rect 0 14784 800 14812
rect 50372 14756 50428 14812
rect 59200 14784 60000 14812
rect 50372 14700 53004 14756
rect 53060 14700 53070 14756
rect 15474 14588 15484 14644
rect 15540 14588 16044 14644
rect 16100 14588 16110 14644
rect 18386 14588 18396 14644
rect 18452 14588 19068 14644
rect 19124 14588 19134 14644
rect 46050 14588 46060 14644
rect 46116 14588 46956 14644
rect 47012 14588 48412 14644
rect 48468 14588 48478 14644
rect 51986 14588 51996 14644
rect 52052 14588 52668 14644
rect 52724 14588 54908 14644
rect 54964 14588 54974 14644
rect 4946 14476 4956 14532
rect 5012 14476 6300 14532
rect 6356 14476 6366 14532
rect 14690 14476 14700 14532
rect 14756 14476 17388 14532
rect 17444 14476 17454 14532
rect 24210 14476 24220 14532
rect 24276 14476 25676 14532
rect 25732 14476 25742 14532
rect 26002 14476 26012 14532
rect 26068 14476 27580 14532
rect 27636 14476 27646 14532
rect 28466 14476 28476 14532
rect 28532 14476 30828 14532
rect 30884 14476 30894 14532
rect 31266 14476 31276 14532
rect 31332 14476 33180 14532
rect 33236 14476 33246 14532
rect 36194 14476 36204 14532
rect 36260 14476 37660 14532
rect 37716 14476 37726 14532
rect 43652 14476 44380 14532
rect 44436 14476 45612 14532
rect 45668 14476 45678 14532
rect 49186 14476 49196 14532
rect 49252 14476 50540 14532
rect 50596 14476 50606 14532
rect 51762 14476 51772 14532
rect 51828 14476 52892 14532
rect 52948 14476 52958 14532
rect 54114 14476 54124 14532
rect 54180 14476 56588 14532
rect 56644 14476 56654 14532
rect 30828 14420 30884 14476
rect 43652 14420 43708 14476
rect 14466 14364 14476 14420
rect 14532 14364 15372 14420
rect 15428 14364 15438 14420
rect 21746 14364 21756 14420
rect 21812 14364 22428 14420
rect 22484 14364 22494 14420
rect 28130 14364 28140 14420
rect 28196 14364 29148 14420
rect 29204 14364 29820 14420
rect 29876 14364 29886 14420
rect 30828 14364 32172 14420
rect 32228 14364 32238 14420
rect 35634 14364 35644 14420
rect 35700 14364 36316 14420
rect 36372 14364 36382 14420
rect 38322 14364 38332 14420
rect 38388 14364 43708 14420
rect 2034 14252 2044 14308
rect 2100 14252 3724 14308
rect 3780 14252 4284 14308
rect 4340 14252 4350 14308
rect 7634 14252 7644 14308
rect 7700 14252 8316 14308
rect 8372 14252 10892 14308
rect 10948 14252 10958 14308
rect 19618 14252 19628 14308
rect 19684 14252 20412 14308
rect 20468 14252 20478 14308
rect 20626 14252 20636 14308
rect 20692 14252 24780 14308
rect 24836 14252 25340 14308
rect 25396 14252 25406 14308
rect 28802 14252 28812 14308
rect 28868 14252 29484 14308
rect 29540 14252 29550 14308
rect 31490 14252 31500 14308
rect 31556 14252 32284 14308
rect 32340 14252 32350 14308
rect 35298 14252 35308 14308
rect 35364 14252 36876 14308
rect 36932 14252 36942 14308
rect 51202 14252 51212 14308
rect 51268 14252 53116 14308
rect 53172 14252 53788 14308
rect 53844 14252 53854 14308
rect 0 14196 800 14224
rect 0 14140 2380 14196
rect 2436 14140 3164 14196
rect 3220 14140 3230 14196
rect 10546 14140 10556 14196
rect 10612 14140 12684 14196
rect 12740 14140 13356 14196
rect 13412 14140 13422 14196
rect 15362 14140 15372 14196
rect 15428 14140 15708 14196
rect 15764 14140 15774 14196
rect 39890 14140 39900 14196
rect 39956 14140 40572 14196
rect 40628 14140 40638 14196
rect 0 14112 800 14140
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 50546 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50830 14140
rect 2706 14028 2716 14084
rect 2772 14028 7308 14084
rect 7364 14028 8204 14084
rect 8260 14028 8270 14084
rect 4722 13916 4732 13972
rect 4788 13916 5180 13972
rect 5236 13916 5964 13972
rect 6020 13916 6972 13972
rect 7028 13916 7038 13972
rect 20850 13916 20860 13972
rect 20916 13916 22204 13972
rect 22260 13916 22270 13972
rect 51874 13916 51884 13972
rect 51940 13916 53004 13972
rect 53060 13916 53070 13972
rect 15586 13804 15596 13860
rect 15652 13804 18060 13860
rect 18116 13804 18126 13860
rect 19058 13804 19068 13860
rect 19124 13804 19740 13860
rect 19796 13804 20412 13860
rect 20468 13804 20478 13860
rect 23090 13804 23100 13860
rect 23156 13804 23436 13860
rect 23492 13804 23502 13860
rect 46946 13804 46956 13860
rect 47012 13804 47852 13860
rect 47908 13804 47918 13860
rect 49074 13804 49084 13860
rect 49140 13804 49756 13860
rect 49812 13804 50652 13860
rect 50708 13804 50718 13860
rect 53554 13804 53564 13860
rect 53620 13804 54236 13860
rect 54292 13804 54302 13860
rect 1922 13692 1932 13748
rect 1988 13692 3724 13748
rect 3780 13692 3790 13748
rect 12674 13692 12684 13748
rect 12740 13692 14140 13748
rect 14196 13692 14206 13748
rect 16930 13692 16940 13748
rect 16996 13692 18732 13748
rect 18788 13692 18798 13748
rect 23538 13692 23548 13748
rect 23604 13692 24668 13748
rect 24724 13692 25116 13748
rect 25172 13692 25182 13748
rect 32274 13692 32284 13748
rect 32340 13692 37660 13748
rect 37716 13692 37726 13748
rect 37986 13692 37996 13748
rect 38052 13692 38444 13748
rect 38500 13692 39228 13748
rect 39284 13692 40908 13748
rect 40964 13692 40974 13748
rect 43652 13692 47516 13748
rect 47572 13692 47582 13748
rect 48066 13692 48076 13748
rect 48132 13692 48748 13748
rect 48804 13692 48814 13748
rect 49970 13692 49980 13748
rect 50036 13692 50428 13748
rect 43652 13636 43708 13692
rect 16370 13580 16380 13636
rect 16436 13580 20748 13636
rect 20804 13580 22316 13636
rect 22372 13580 22382 13636
rect 30594 13580 30604 13636
rect 30660 13580 41020 13636
rect 41076 13580 41580 13636
rect 41636 13580 43708 13636
rect 45266 13580 45276 13636
rect 45332 13580 46508 13636
rect 46564 13580 47740 13636
rect 47796 13580 47806 13636
rect 0 13524 800 13552
rect 50372 13524 50428 13692
rect 0 13468 1708 13524
rect 1764 13468 1774 13524
rect 2034 13468 2044 13524
rect 2100 13468 3948 13524
rect 4004 13468 4014 13524
rect 6962 13468 6972 13524
rect 7028 13468 12908 13524
rect 12964 13468 13916 13524
rect 13972 13468 13982 13524
rect 14466 13468 14476 13524
rect 14532 13468 15708 13524
rect 15764 13468 15774 13524
rect 18722 13468 18732 13524
rect 18788 13468 19292 13524
rect 19348 13468 20076 13524
rect 20132 13468 20142 13524
rect 36306 13468 36316 13524
rect 36372 13468 43148 13524
rect 43204 13468 43214 13524
rect 50372 13468 50652 13524
rect 50708 13468 50718 13524
rect 0 13440 800 13468
rect 9202 13356 9212 13412
rect 9268 13356 9996 13412
rect 10052 13356 10062 13412
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 8530 13244 8540 13300
rect 8596 13244 12124 13300
rect 12180 13244 12190 13300
rect 7858 13020 7868 13076
rect 7924 13020 8932 13076
rect 23062 13020 23100 13076
rect 23156 13020 23166 13076
rect 33506 13020 33516 13076
rect 33572 13020 37100 13076
rect 37156 13020 37166 13076
rect 8876 12964 8932 13020
rect 7522 12908 7532 12964
rect 7588 12908 8652 12964
rect 8708 12908 8718 12964
rect 8866 12908 8876 12964
rect 8932 12908 8942 12964
rect 14578 12908 14588 12964
rect 14644 12908 15596 12964
rect 15652 12908 15662 12964
rect 20738 12908 20748 12964
rect 20804 12908 23212 12964
rect 23268 12908 23772 12964
rect 23828 12908 23838 12964
rect 43026 12908 43036 12964
rect 43092 12908 45164 12964
rect 45220 12908 45230 12964
rect 46274 12908 46284 12964
rect 46340 12908 47068 12964
rect 47124 12908 47134 12964
rect 51874 12908 51884 12964
rect 51940 12908 52668 12964
rect 52724 12908 52734 12964
rect 0 12852 800 12880
rect 0 12796 2380 12852
rect 2436 12796 4508 12852
rect 4564 12796 4574 12852
rect 7074 12796 7084 12852
rect 7140 12796 9212 12852
rect 9268 12796 9278 12852
rect 9538 12796 9548 12852
rect 9604 12796 10556 12852
rect 10612 12796 10622 12852
rect 26898 12796 26908 12852
rect 26964 12796 26974 12852
rect 38294 12796 38332 12852
rect 38388 12796 38398 12852
rect 43698 12796 43708 12852
rect 43764 12796 44828 12852
rect 44884 12796 44894 12852
rect 47282 12796 47292 12852
rect 47348 12796 48300 12852
rect 48356 12796 48366 12852
rect 51986 12796 51996 12852
rect 52052 12796 53116 12852
rect 53172 12796 53182 12852
rect 55458 12796 55468 12852
rect 55524 12796 56924 12852
rect 56980 12796 56990 12852
rect 0 12768 800 12796
rect 26908 12740 26964 12796
rect 1698 12684 1708 12740
rect 1764 12684 4956 12740
rect 5012 12684 5022 12740
rect 12114 12684 12124 12740
rect 12180 12684 14700 12740
rect 14756 12684 14766 12740
rect 20738 12684 20748 12740
rect 20804 12684 21420 12740
rect 21476 12684 21486 12740
rect 25890 12684 25900 12740
rect 25956 12684 27132 12740
rect 27188 12684 27198 12740
rect 30706 12684 30716 12740
rect 30772 12684 31948 12740
rect 32004 12684 38108 12740
rect 38164 12684 39116 12740
rect 39172 12684 39182 12740
rect 50082 12684 50092 12740
rect 50148 12684 55244 12740
rect 55300 12684 56588 12740
rect 56644 12684 56654 12740
rect 3378 12572 3388 12628
rect 3444 12572 4284 12628
rect 4340 12572 4350 12628
rect 8866 12572 8876 12628
rect 8932 12572 9548 12628
rect 9604 12572 9614 12628
rect 38210 12572 38220 12628
rect 38276 12572 38892 12628
rect 38948 12572 38958 12628
rect 41458 12572 41468 12628
rect 41524 12572 42476 12628
rect 42532 12572 44044 12628
rect 44100 12572 44110 12628
rect 54450 12572 54460 12628
rect 54516 12572 56028 12628
rect 56084 12572 56094 12628
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 50546 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50830 12572
rect 6290 12460 6300 12516
rect 6356 12460 7420 12516
rect 7476 12460 8540 12516
rect 8596 12460 8606 12516
rect 4610 12348 4620 12404
rect 4676 12348 10724 12404
rect 12002 12348 12012 12404
rect 12068 12348 13804 12404
rect 13860 12348 14812 12404
rect 14868 12348 14878 12404
rect 15362 12348 15372 12404
rect 15428 12348 16268 12404
rect 16324 12348 16334 12404
rect 18386 12348 18396 12404
rect 18452 12348 19964 12404
rect 20020 12348 20030 12404
rect 28354 12348 28364 12404
rect 28420 12348 30156 12404
rect 30212 12348 30222 12404
rect 35970 12348 35980 12404
rect 36036 12348 45052 12404
rect 45108 12348 45118 12404
rect 46162 12348 46172 12404
rect 46228 12348 47292 12404
rect 47348 12348 48412 12404
rect 48468 12348 48478 12404
rect 2034 12236 2044 12292
rect 2100 12236 5516 12292
rect 5572 12236 5582 12292
rect 6402 12236 6412 12292
rect 6468 12236 8204 12292
rect 8260 12236 8270 12292
rect 9874 12236 9884 12292
rect 9940 12236 10332 12292
rect 10388 12236 10398 12292
rect 0 12180 800 12208
rect 10668 12180 10724 12348
rect 19506 12236 19516 12292
rect 19572 12236 20076 12292
rect 20132 12236 20748 12292
rect 20804 12236 20814 12292
rect 29586 12236 29596 12292
rect 29652 12236 31388 12292
rect 31444 12236 31454 12292
rect 32620 12236 35084 12292
rect 35140 12236 35150 12292
rect 41682 12236 41692 12292
rect 41748 12236 51996 12292
rect 52052 12236 52062 12292
rect 53442 12236 53452 12292
rect 53508 12236 55132 12292
rect 55188 12236 55198 12292
rect 32620 12180 32676 12236
rect 0 12124 1708 12180
rect 1764 12124 1774 12180
rect 6290 12124 6300 12180
rect 6356 12124 6636 12180
rect 6692 12124 8764 12180
rect 8820 12124 9772 12180
rect 9828 12124 9838 12180
rect 10658 12124 10668 12180
rect 10724 12124 10734 12180
rect 13906 12124 13916 12180
rect 13972 12124 14588 12180
rect 14644 12124 14654 12180
rect 26898 12124 26908 12180
rect 26964 12124 27356 12180
rect 27412 12124 28252 12180
rect 28308 12124 28318 12180
rect 28466 12124 28476 12180
rect 28532 12124 32676 12180
rect 37202 12124 37212 12180
rect 37268 12124 42476 12180
rect 42532 12124 43260 12180
rect 43316 12124 43708 12180
rect 44258 12124 44268 12180
rect 44324 12124 45164 12180
rect 45220 12124 45230 12180
rect 49858 12124 49868 12180
rect 49924 12124 50988 12180
rect 51044 12124 51884 12180
rect 51940 12124 51950 12180
rect 55570 12124 55580 12180
rect 55636 12124 57036 12180
rect 57092 12124 57102 12180
rect 0 12096 800 12124
rect 2370 12012 2380 12068
rect 2436 12012 5180 12068
rect 5236 12012 5246 12068
rect 5730 12012 5740 12068
rect 5796 12012 6748 12068
rect 6804 12012 6814 12068
rect 7970 12012 7980 12068
rect 8036 12012 8046 12068
rect 8194 12012 8204 12068
rect 8260 12012 12012 12068
rect 12068 12012 12078 12068
rect 33394 12012 33404 12068
rect 33460 12012 33964 12068
rect 34020 12012 34030 12068
rect 38612 12012 41580 12068
rect 41636 12012 41646 12068
rect 43652 12012 43708 12124
rect 43764 12012 43774 12068
rect 49970 12012 49980 12068
rect 50036 12012 50046 12068
rect 7980 11956 8036 12012
rect 38612 11956 38668 12012
rect 49980 11956 50036 12012
rect 3602 11900 3612 11956
rect 3668 11900 3678 11956
rect 7980 11900 9212 11956
rect 9268 11900 9660 11956
rect 9716 11900 9726 11956
rect 15810 11900 15820 11956
rect 15876 11900 16828 11956
rect 16884 11900 17948 11956
rect 18004 11900 18014 11956
rect 27122 11900 27132 11956
rect 27188 11900 28252 11956
rect 28308 11900 28318 11956
rect 29810 11900 29820 11956
rect 29876 11900 30940 11956
rect 30996 11900 33068 11956
rect 33124 11900 38668 11956
rect 42914 11900 42924 11956
rect 42980 11900 47180 11956
rect 47236 11900 47246 11956
rect 47730 11900 47740 11956
rect 47796 11900 49308 11956
rect 49364 11900 50036 11956
rect 3612 11620 3668 11900
rect 4834 11788 4844 11844
rect 4900 11788 6300 11844
rect 6356 11788 6366 11844
rect 7634 11788 7644 11844
rect 7700 11788 8316 11844
rect 8372 11788 8382 11844
rect 11442 11788 11452 11844
rect 11508 11788 12124 11844
rect 12180 11788 12190 11844
rect 18274 11788 18284 11844
rect 18340 11788 19180 11844
rect 19236 11788 19246 11844
rect 33282 11788 33292 11844
rect 33348 11788 33852 11844
rect 33908 11788 34188 11844
rect 34244 11788 34254 11844
rect 50642 11788 50652 11844
rect 50708 11788 55356 11844
rect 55412 11788 55422 11844
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 28578 11676 28588 11732
rect 28644 11676 30380 11732
rect 30436 11676 30446 11732
rect 47618 11676 47628 11732
rect 47684 11676 51100 11732
rect 51156 11676 51166 11732
rect 3612 11564 5740 11620
rect 5796 11564 5806 11620
rect 13570 11564 13580 11620
rect 13636 11564 15988 11620
rect 16370 11564 16380 11620
rect 16436 11564 17164 11620
rect 17220 11564 17724 11620
rect 17780 11564 17790 11620
rect 20290 11564 20300 11620
rect 20356 11564 21532 11620
rect 21588 11564 21598 11620
rect 34514 11564 34524 11620
rect 34580 11564 35420 11620
rect 35476 11564 35486 11620
rect 35634 11564 35644 11620
rect 35700 11564 36428 11620
rect 36484 11564 36494 11620
rect 0 11508 800 11536
rect 3612 11508 3668 11564
rect 15932 11508 15988 11564
rect 35644 11508 35700 11564
rect 0 11452 2380 11508
rect 2436 11452 2446 11508
rect 3602 11452 3612 11508
rect 3668 11452 3678 11508
rect 4946 11452 4956 11508
rect 5012 11452 15148 11508
rect 15922 11452 15932 11508
rect 15988 11452 16940 11508
rect 16996 11452 17006 11508
rect 20178 11452 20188 11508
rect 20244 11452 21420 11508
rect 21476 11452 22876 11508
rect 22932 11452 22942 11508
rect 33170 11452 33180 11508
rect 33236 11452 33628 11508
rect 33684 11452 33694 11508
rect 34962 11452 34972 11508
rect 35028 11452 35700 11508
rect 0 11424 800 11452
rect 15092 11396 15148 11452
rect 6402 11340 6412 11396
rect 6468 11340 6972 11396
rect 7028 11340 7038 11396
rect 12562 11340 12572 11396
rect 12628 11340 13916 11396
rect 13972 11340 13982 11396
rect 15092 11340 15484 11396
rect 15540 11340 16492 11396
rect 16548 11340 16558 11396
rect 17602 11340 17612 11396
rect 17668 11340 19180 11396
rect 19236 11340 19246 11396
rect 27794 11340 27804 11396
rect 27860 11340 29428 11396
rect 32498 11340 32508 11396
rect 32564 11340 37548 11396
rect 37604 11340 37614 11396
rect 38882 11340 38892 11396
rect 38948 11340 39564 11396
rect 39620 11340 39630 11396
rect 53554 11340 53564 11396
rect 53620 11340 55692 11396
rect 55748 11340 55758 11396
rect 29372 11284 29428 11340
rect 3378 11228 3388 11284
rect 3444 11228 5740 11284
rect 5796 11228 6524 11284
rect 6580 11228 6590 11284
rect 10098 11228 10108 11284
rect 10164 11228 11340 11284
rect 11396 11228 13412 11284
rect 25106 11228 25116 11284
rect 25172 11228 29036 11284
rect 29092 11228 29102 11284
rect 29362 11228 29372 11284
rect 29428 11228 29708 11284
rect 29764 11228 29774 11284
rect 33394 11228 33404 11284
rect 33460 11228 35868 11284
rect 35924 11228 35934 11284
rect 38434 11228 38444 11284
rect 38500 11228 39676 11284
rect 39732 11228 45612 11284
rect 45668 11228 47068 11284
rect 47124 11228 50316 11284
rect 50372 11228 50382 11284
rect 52210 11228 52220 11284
rect 52276 11228 55804 11284
rect 55860 11228 55870 11284
rect 13356 11172 13412 11228
rect 2706 11116 2716 11172
rect 2772 11116 3948 11172
rect 4004 11116 4014 11172
rect 10770 11116 10780 11172
rect 10836 11116 12460 11172
rect 12516 11116 12526 11172
rect 13356 11116 14476 11172
rect 14532 11116 14542 11172
rect 27346 11116 27356 11172
rect 27412 11116 33964 11172
rect 34020 11116 34030 11172
rect 39218 11116 39228 11172
rect 39284 11116 40124 11172
rect 40180 11116 40190 11172
rect 43138 11116 43148 11172
rect 43204 11116 43484 11172
rect 43540 11116 44492 11172
rect 44548 11116 44558 11172
rect 48290 11116 48300 11172
rect 48356 11116 49196 11172
rect 49252 11116 49262 11172
rect 38658 11004 38668 11060
rect 38724 11004 39116 11060
rect 39172 11004 40236 11060
rect 40292 11004 45276 11060
rect 45332 11004 45342 11060
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 50546 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50830 11004
rect 12786 10892 12796 10948
rect 12852 10892 13692 10948
rect 13748 10892 13758 10948
rect 30370 10892 30380 10948
rect 30436 10892 42588 10948
rect 42644 10892 42654 10948
rect 53106 10892 53116 10948
rect 53172 10892 53676 10948
rect 53732 10892 53742 10948
rect 0 10836 800 10864
rect 0 10780 1708 10836
rect 1764 10780 1774 10836
rect 2034 10780 2044 10836
rect 2100 10780 2828 10836
rect 2884 10780 3500 10836
rect 3556 10780 3566 10836
rect 26562 10780 26572 10836
rect 26628 10780 28028 10836
rect 28084 10780 28094 10836
rect 28466 10780 28476 10836
rect 28532 10780 29596 10836
rect 29652 10780 29662 10836
rect 33618 10780 33628 10836
rect 33684 10780 33964 10836
rect 34020 10780 34030 10836
rect 34850 10780 34860 10836
rect 34916 10780 38108 10836
rect 38164 10780 38780 10836
rect 38836 10780 38846 10836
rect 0 10752 800 10780
rect 2482 10668 2492 10724
rect 2548 10668 5068 10724
rect 5124 10668 5134 10724
rect 9650 10668 9660 10724
rect 9716 10668 11004 10724
rect 11060 10668 11070 10724
rect 34514 10668 34524 10724
rect 34580 10668 38444 10724
rect 38500 10668 39116 10724
rect 39172 10668 40572 10724
rect 40628 10668 40638 10724
rect 51090 10668 51100 10724
rect 51156 10668 52332 10724
rect 52388 10668 52398 10724
rect 54898 10668 54908 10724
rect 54964 10668 56812 10724
rect 56868 10668 56878 10724
rect 4050 10556 4060 10612
rect 4116 10556 5852 10612
rect 5908 10556 5918 10612
rect 16930 10556 16940 10612
rect 16996 10556 19180 10612
rect 19236 10556 19246 10612
rect 25778 10556 25788 10612
rect 25844 10556 26460 10612
rect 26516 10556 27468 10612
rect 27524 10556 27534 10612
rect 32274 10556 32284 10612
rect 32340 10556 33628 10612
rect 33684 10556 33694 10612
rect 35634 10556 35644 10612
rect 35700 10556 39340 10612
rect 39396 10556 41020 10612
rect 41076 10556 41086 10612
rect 52210 10556 52220 10612
rect 52276 10556 52892 10612
rect 52948 10556 53900 10612
rect 53956 10556 53966 10612
rect 55010 10556 55020 10612
rect 55076 10556 56476 10612
rect 56532 10556 56542 10612
rect 4498 10444 4508 10500
rect 4564 10444 5068 10500
rect 5124 10444 5134 10500
rect 8978 10444 8988 10500
rect 9044 10444 9884 10500
rect 9940 10444 9950 10500
rect 16482 10444 16492 10500
rect 16548 10444 17724 10500
rect 17780 10444 17790 10500
rect 26338 10444 26348 10500
rect 26404 10444 27692 10500
rect 27748 10444 27758 10500
rect 37986 10444 37996 10500
rect 38052 10444 43260 10500
rect 43316 10444 43326 10500
rect 48178 10444 48188 10500
rect 48244 10444 49644 10500
rect 49700 10444 49710 10500
rect 54226 10444 54236 10500
rect 54292 10444 54684 10500
rect 54740 10444 56028 10500
rect 56084 10444 57036 10500
rect 57092 10444 57102 10500
rect 38668 10388 38724 10444
rect 1810 10332 1820 10388
rect 1876 10332 3164 10388
rect 3220 10332 3230 10388
rect 12226 10332 12236 10388
rect 12292 10332 14476 10388
rect 14532 10332 14924 10388
rect 14980 10332 14990 10388
rect 26450 10332 26460 10388
rect 26516 10332 27020 10388
rect 27076 10332 27086 10388
rect 35074 10332 35084 10388
rect 35140 10332 35868 10388
rect 35924 10332 36540 10388
rect 36596 10332 36606 10388
rect 38658 10332 38668 10388
rect 38724 10332 38734 10388
rect 40114 10332 40124 10388
rect 40180 10332 40908 10388
rect 40964 10332 51548 10388
rect 51604 10332 51614 10388
rect 36642 10220 36652 10276
rect 36708 10220 41580 10276
rect 41636 10220 41646 10276
rect 0 10164 800 10192
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 0 10108 1708 10164
rect 1764 10108 2492 10164
rect 2548 10108 2558 10164
rect 3042 10108 3052 10164
rect 3108 10108 3892 10164
rect 5282 10108 5292 10164
rect 5348 10108 6412 10164
rect 6468 10108 6478 10164
rect 43362 10108 43372 10164
rect 43428 10108 46284 10164
rect 46340 10108 46350 10164
rect 0 10080 800 10108
rect 3836 10052 3892 10108
rect 3826 9996 3836 10052
rect 3892 9996 3902 10052
rect 10322 9996 10332 10052
rect 10388 9996 12124 10052
rect 12180 9996 12190 10052
rect 14578 9996 14588 10052
rect 14644 9996 15148 10052
rect 29810 9996 29820 10052
rect 29876 9996 30492 10052
rect 30548 9996 30558 10052
rect 31798 9996 31836 10052
rect 31892 9996 31902 10052
rect 39442 9996 39452 10052
rect 39508 9996 51772 10052
rect 51828 9996 52668 10052
rect 52724 9996 52734 10052
rect 4946 9884 4956 9940
rect 5012 9884 6972 9940
rect 7028 9884 8204 9940
rect 8260 9884 8270 9940
rect 15092 9828 15148 9996
rect 25554 9884 25564 9940
rect 25620 9884 26796 9940
rect 26852 9884 26862 9940
rect 40898 9884 40908 9940
rect 40964 9884 53452 9940
rect 53508 9884 54124 9940
rect 54180 9884 54190 9940
rect 15092 9772 17612 9828
rect 17668 9772 18284 9828
rect 18340 9772 18350 9828
rect 22754 9772 22764 9828
rect 22820 9772 23772 9828
rect 23828 9772 23838 9828
rect 28578 9772 28588 9828
rect 28644 9772 31836 9828
rect 31892 9772 35644 9828
rect 35700 9772 35710 9828
rect 38434 9772 38444 9828
rect 38500 9772 39900 9828
rect 39956 9772 39966 9828
rect 49858 9772 49868 9828
rect 49924 9772 50540 9828
rect 50596 9772 50606 9828
rect 52098 9772 52108 9828
rect 52164 9772 54572 9828
rect 54628 9772 55580 9828
rect 55636 9772 55646 9828
rect 2706 9660 2716 9716
rect 2772 9660 4172 9716
rect 4228 9660 4238 9716
rect 6738 9660 6748 9716
rect 6804 9660 7756 9716
rect 7812 9660 7822 9716
rect 9762 9660 9772 9716
rect 9828 9660 10444 9716
rect 10500 9660 10510 9716
rect 14802 9660 14812 9716
rect 14868 9660 21532 9716
rect 21588 9660 21598 9716
rect 22082 9660 22092 9716
rect 22148 9660 23212 9716
rect 23268 9660 23278 9716
rect 28466 9660 28476 9716
rect 28532 9660 29260 9716
rect 29316 9660 31052 9716
rect 31108 9660 31118 9716
rect 34962 9660 34972 9716
rect 35028 9660 36316 9716
rect 36372 9660 36382 9716
rect 48514 9660 48524 9716
rect 48580 9660 50988 9716
rect 51044 9660 51054 9716
rect 53666 9660 53676 9716
rect 53732 9660 57148 9716
rect 57204 9660 57214 9716
rect 20972 9604 21028 9660
rect 4946 9548 4956 9604
rect 5012 9548 7084 9604
rect 7140 9548 7150 9604
rect 17938 9548 17948 9604
rect 18004 9548 18732 9604
rect 18788 9548 18798 9604
rect 20962 9548 20972 9604
rect 21028 9548 21038 9604
rect 33954 9548 33964 9604
rect 34020 9548 34412 9604
rect 34468 9548 34478 9604
rect 35746 9548 35756 9604
rect 35812 9548 40236 9604
rect 40292 9548 41356 9604
rect 41412 9548 41422 9604
rect 45602 9548 45612 9604
rect 45668 9548 46172 9604
rect 46228 9548 47180 9604
rect 47236 9548 47246 9604
rect 0 9492 800 9520
rect 0 9436 1708 9492
rect 1764 9436 1774 9492
rect 34738 9436 34748 9492
rect 34804 9436 35308 9492
rect 35364 9436 36204 9492
rect 36260 9436 36270 9492
rect 36866 9436 36876 9492
rect 36932 9436 38220 9492
rect 38276 9436 40348 9492
rect 40404 9436 41692 9492
rect 41748 9436 42924 9492
rect 42980 9436 42990 9492
rect 0 9408 800 9436
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 50546 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50830 9436
rect 3266 9324 3276 9380
rect 3332 9324 5180 9380
rect 5236 9324 13580 9380
rect 13636 9324 14868 9380
rect 29698 9324 29708 9380
rect 29764 9324 49644 9380
rect 49700 9324 49710 9380
rect 3490 9212 3500 9268
rect 3556 9212 5404 9268
rect 5460 9212 5470 9268
rect 6626 9212 6636 9268
rect 6692 9212 8092 9268
rect 8148 9212 8158 9268
rect 9874 9212 9884 9268
rect 9940 9212 11452 9268
rect 11508 9212 14644 9268
rect 14588 9156 14644 9212
rect 14812 9156 14868 9324
rect 30706 9212 30716 9268
rect 30772 9212 36428 9268
rect 36484 9212 36494 9268
rect 38882 9212 38892 9268
rect 38948 9212 39340 9268
rect 39396 9212 40124 9268
rect 40180 9212 40190 9268
rect 51426 9212 51436 9268
rect 51492 9212 52892 9268
rect 52948 9212 52958 9268
rect 38892 9156 38948 9212
rect 2034 9100 2044 9156
rect 2100 9100 4284 9156
rect 4340 9100 4350 9156
rect 4620 9100 5292 9156
rect 5348 9100 5358 9156
rect 14578 9100 14588 9156
rect 14644 9100 14654 9156
rect 14802 9100 14812 9156
rect 14868 9100 14878 9156
rect 18834 9100 18844 9156
rect 18900 9100 19964 9156
rect 20020 9100 20030 9156
rect 21186 9100 21196 9156
rect 21252 9100 21980 9156
rect 22036 9100 22046 9156
rect 27570 9100 27580 9156
rect 27636 9100 31388 9156
rect 31444 9100 31948 9156
rect 32004 9100 32014 9156
rect 35298 9100 35308 9156
rect 35364 9100 35980 9156
rect 36036 9100 36046 9156
rect 36306 9100 36316 9156
rect 36372 9100 38948 9156
rect 43026 9100 43036 9156
rect 43092 9100 44492 9156
rect 44548 9100 45612 9156
rect 45668 9100 45678 9156
rect 45938 9100 45948 9156
rect 46004 9100 47852 9156
rect 47908 9100 47918 9156
rect 4620 9044 4676 9100
rect 3826 8988 3836 9044
rect 3892 8988 4620 9044
rect 4676 8988 4686 9044
rect 5058 8988 5068 9044
rect 5124 8988 6412 9044
rect 6468 8988 7196 9044
rect 7252 8988 7262 9044
rect 16482 8988 16492 9044
rect 16548 8988 17948 9044
rect 18004 8988 18014 9044
rect 22082 8988 22092 9044
rect 22148 8988 23436 9044
rect 23492 8988 23502 9044
rect 27458 8988 27468 9044
rect 27524 8988 28588 9044
rect 28644 8988 28654 9044
rect 31154 8988 31164 9044
rect 31220 8988 36092 9044
rect 36148 8988 38780 9044
rect 38836 8988 38846 9044
rect 43138 8988 43148 9044
rect 43204 8988 43820 9044
rect 43876 8988 43886 9044
rect 51650 8988 51660 9044
rect 51716 8988 51726 9044
rect 54114 8988 54124 9044
rect 54180 8988 54684 9044
rect 54740 8988 54750 9044
rect 51660 8932 51716 8988
rect 29026 8876 29036 8932
rect 29092 8876 30268 8932
rect 30324 8876 31612 8932
rect 31668 8876 31678 8932
rect 42578 8876 42588 8932
rect 42644 8876 45388 8932
rect 45444 8876 45454 8932
rect 46498 8876 46508 8932
rect 46564 8876 51716 8932
rect 0 8820 800 8848
rect 0 8764 2380 8820
rect 2436 8764 3612 8820
rect 3668 8764 3678 8820
rect 26898 8764 26908 8820
rect 26964 8764 27916 8820
rect 27972 8764 28812 8820
rect 28868 8764 38444 8820
rect 38500 8764 38510 8820
rect 45266 8764 45276 8820
rect 45332 8764 46060 8820
rect 46116 8764 46956 8820
rect 47012 8764 47022 8820
rect 50978 8764 50988 8820
rect 51044 8764 51660 8820
rect 51716 8764 51726 8820
rect 0 8736 800 8764
rect 51762 8652 51772 8708
rect 51828 8652 55916 8708
rect 55972 8652 57484 8708
rect 57540 8652 57550 8708
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 33954 8540 33964 8596
rect 34020 8540 34636 8596
rect 34692 8540 34702 8596
rect 49858 8540 49868 8596
rect 49924 8540 49934 8596
rect 49868 8484 49924 8540
rect 20178 8428 20188 8484
rect 20244 8428 22092 8484
rect 22148 8428 22158 8484
rect 24658 8428 24668 8484
rect 24724 8428 25788 8484
rect 25844 8428 25854 8484
rect 31826 8428 31836 8484
rect 31892 8428 31902 8484
rect 33506 8428 33516 8484
rect 33572 8428 44044 8484
rect 44100 8428 44110 8484
rect 49522 8428 49532 8484
rect 49588 8428 49924 8484
rect 51762 8428 51772 8484
rect 51828 8428 52892 8484
rect 52948 8428 52958 8484
rect 7410 8316 7420 8372
rect 7476 8316 9548 8372
rect 9604 8316 9614 8372
rect 10210 8316 10220 8372
rect 10276 8316 13244 8372
rect 13300 8316 13580 8372
rect 13636 8316 13646 8372
rect 18162 8316 18172 8372
rect 18228 8316 19404 8372
rect 19460 8316 19470 8372
rect 24994 8316 25004 8372
rect 25060 8316 25900 8372
rect 25956 8316 28140 8372
rect 28196 8316 28206 8372
rect 31836 8260 31892 8428
rect 33282 8316 33292 8372
rect 33348 8316 33852 8372
rect 33908 8316 39004 8372
rect 39060 8316 39070 8372
rect 49634 8316 49644 8372
rect 49700 8316 51212 8372
rect 51268 8316 51278 8372
rect 4722 8204 4732 8260
rect 4788 8204 5404 8260
rect 5460 8204 5964 8260
rect 6020 8204 6030 8260
rect 6626 8204 6636 8260
rect 6692 8204 7084 8260
rect 7140 8204 8428 8260
rect 8484 8204 9436 8260
rect 9492 8204 9502 8260
rect 12562 8204 12572 8260
rect 12628 8204 13804 8260
rect 13860 8204 13870 8260
rect 27234 8204 27244 8260
rect 27300 8204 28252 8260
rect 28308 8204 28318 8260
rect 31836 8204 33628 8260
rect 33684 8204 33694 8260
rect 34402 8204 34412 8260
rect 34468 8204 34748 8260
rect 34804 8204 34814 8260
rect 36642 8204 36652 8260
rect 36708 8204 38220 8260
rect 38276 8204 38780 8260
rect 38836 8204 38846 8260
rect 50194 8204 50204 8260
rect 50260 8204 50988 8260
rect 51044 8204 52780 8260
rect 52836 8204 52846 8260
rect 53442 8204 53452 8260
rect 53508 8204 54460 8260
rect 54516 8204 54526 8260
rect 0 8148 800 8176
rect 0 8092 1708 8148
rect 1764 8092 2940 8148
rect 2996 8092 3006 8148
rect 8306 8092 8316 8148
rect 8372 8092 10108 8148
rect 10164 8092 11676 8148
rect 11732 8092 11742 8148
rect 14914 8092 14924 8148
rect 14980 8092 15820 8148
rect 15876 8092 15886 8148
rect 30482 8092 30492 8148
rect 30548 8092 30940 8148
rect 30996 8092 31006 8148
rect 31826 8092 31836 8148
rect 31892 8092 34076 8148
rect 34132 8092 35084 8148
rect 35140 8092 35980 8148
rect 36036 8092 36046 8148
rect 49298 8092 49308 8148
rect 49364 8092 52892 8148
rect 52948 8092 52958 8148
rect 0 8064 800 8092
rect 7410 7980 7420 8036
rect 7476 7980 13916 8036
rect 13972 7980 13982 8036
rect 22866 7980 22876 8036
rect 22932 7980 24668 8036
rect 24724 7980 26236 8036
rect 26292 7980 26302 8036
rect 27458 7980 27468 8036
rect 27524 7980 28028 8036
rect 28084 7980 29036 8036
rect 29092 7980 29102 8036
rect 30370 7980 30380 8036
rect 30436 7980 33068 8036
rect 33124 7980 33134 8036
rect 33618 7980 33628 8036
rect 33684 7980 34300 8036
rect 34356 7980 34366 8036
rect 36194 7980 36204 8036
rect 36260 7980 43708 8036
rect 43652 7924 43708 7980
rect 11218 7868 11228 7924
rect 11284 7868 14812 7924
rect 14868 7868 16268 7924
rect 16324 7868 16828 7924
rect 16884 7868 16894 7924
rect 43652 7868 48748 7924
rect 48804 7868 48814 7924
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 50546 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50830 7868
rect 34626 7756 34636 7812
rect 34692 7756 38668 7812
rect 39890 7756 39900 7812
rect 39956 7756 41020 7812
rect 41076 7756 43484 7812
rect 43540 7756 43550 7812
rect 38612 7700 38668 7756
rect 8866 7644 8876 7700
rect 8932 7644 11116 7700
rect 11172 7644 11182 7700
rect 14578 7644 14588 7700
rect 14644 7644 15484 7700
rect 15540 7644 15550 7700
rect 35298 7644 35308 7700
rect 35364 7644 35868 7700
rect 35924 7644 36652 7700
rect 36708 7644 36718 7700
rect 38612 7644 51772 7700
rect 51828 7644 51838 7700
rect 51986 7644 51996 7700
rect 52052 7644 57260 7700
rect 57316 7644 57326 7700
rect 11442 7532 11452 7588
rect 11508 7532 13580 7588
rect 13636 7532 14700 7588
rect 14756 7532 15148 7588
rect 15204 7532 15214 7588
rect 30594 7532 30604 7588
rect 30660 7532 32284 7588
rect 32340 7532 35420 7588
rect 35476 7532 36764 7588
rect 36820 7532 36830 7588
rect 40114 7532 40124 7588
rect 40180 7532 41580 7588
rect 41636 7532 42588 7588
rect 42644 7532 42654 7588
rect 55906 7532 55916 7588
rect 55972 7532 57148 7588
rect 57204 7532 57214 7588
rect 2034 7420 2044 7476
rect 2100 7420 9772 7476
rect 9828 7420 9838 7476
rect 10994 7420 11004 7476
rect 11060 7420 12572 7476
rect 12628 7420 12638 7476
rect 23202 7420 23212 7476
rect 23268 7420 24444 7476
rect 24500 7420 30380 7476
rect 30436 7420 30446 7476
rect 31724 7420 34188 7476
rect 34244 7420 34254 7476
rect 38322 7420 38332 7476
rect 38388 7420 39116 7476
rect 39172 7420 40796 7476
rect 40852 7420 40862 7476
rect 42018 7420 42028 7476
rect 42084 7420 44156 7476
rect 44212 7420 44222 7476
rect 46386 7420 46396 7476
rect 46452 7420 47180 7476
rect 47236 7420 47246 7476
rect 54562 7420 54572 7476
rect 54628 7420 56588 7476
rect 56644 7420 56654 7476
rect 31724 7364 31780 7420
rect 8372 7308 14476 7364
rect 14532 7308 14542 7364
rect 15250 7308 15260 7364
rect 15316 7308 15708 7364
rect 15764 7308 15774 7364
rect 29810 7308 29820 7364
rect 29876 7308 31724 7364
rect 31780 7308 31790 7364
rect 32498 7308 32508 7364
rect 32564 7308 33628 7364
rect 33684 7308 33694 7364
rect 34402 7308 34412 7364
rect 34468 7308 38668 7364
rect 38724 7308 41132 7364
rect 41188 7308 41198 7364
rect 42242 7308 42252 7364
rect 42308 7308 43708 7364
rect 43764 7308 43774 7364
rect 8372 7252 8428 7308
rect 5954 7196 5964 7252
rect 6020 7196 8428 7252
rect 14018 7196 14028 7252
rect 14084 7196 18844 7252
rect 18900 7196 18910 7252
rect 27010 7196 27020 7252
rect 27076 7196 27086 7252
rect 37202 7196 37212 7252
rect 37268 7196 48972 7252
rect 49028 7196 49038 7252
rect 27020 7140 27076 7196
rect 26450 7084 26460 7140
rect 26516 7084 27580 7140
rect 27636 7084 27646 7140
rect 33058 7084 33068 7140
rect 33124 7084 33740 7140
rect 33796 7084 33806 7140
rect 40898 7084 40908 7140
rect 40964 7084 43708 7140
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 43652 7028 43708 7084
rect 43652 6972 53228 7028
rect 53284 6972 53900 7028
rect 53956 6972 54684 7028
rect 54740 6972 54750 7028
rect 27122 6860 27132 6916
rect 27188 6860 28364 6916
rect 28420 6860 29372 6916
rect 29428 6860 29438 6916
rect 34290 6860 34300 6916
rect 34356 6860 42252 6916
rect 42308 6860 42318 6916
rect 13906 6748 13916 6804
rect 13972 6748 14700 6804
rect 14756 6748 14766 6804
rect 27458 6748 27468 6804
rect 27524 6748 28028 6804
rect 28084 6748 28094 6804
rect 35746 6748 35756 6804
rect 35812 6748 37436 6804
rect 37492 6748 37502 6804
rect 38322 6748 38332 6804
rect 38388 6748 39228 6804
rect 39284 6748 39294 6804
rect 42578 6748 42588 6804
rect 42644 6748 46060 6804
rect 46116 6748 49868 6804
rect 49924 6748 49934 6804
rect 50418 6748 50428 6804
rect 50484 6748 52556 6804
rect 52612 6748 53004 6804
rect 53060 6748 53070 6804
rect 24210 6636 24220 6692
rect 24276 6636 24668 6692
rect 24724 6636 25340 6692
rect 25396 6636 25406 6692
rect 26114 6636 26124 6692
rect 26180 6636 26908 6692
rect 26964 6636 27972 6692
rect 29586 6636 29596 6692
rect 29652 6636 31388 6692
rect 31444 6636 31454 6692
rect 36530 6636 36540 6692
rect 36596 6636 37772 6692
rect 37828 6636 38108 6692
rect 38164 6636 38174 6692
rect 41234 6636 41244 6692
rect 41300 6636 42364 6692
rect 42420 6636 42430 6692
rect 44034 6636 44044 6692
rect 44100 6636 46284 6692
rect 46340 6636 46350 6692
rect 50194 6636 50204 6692
rect 50260 6636 50876 6692
rect 50932 6636 50942 6692
rect 27916 6580 27972 6636
rect 51324 6580 51380 6748
rect 27906 6524 27916 6580
rect 27972 6524 32172 6580
rect 32228 6524 32238 6580
rect 35410 6524 35420 6580
rect 35476 6524 36428 6580
rect 36484 6524 36494 6580
rect 37538 6524 37548 6580
rect 37604 6524 37614 6580
rect 37986 6524 37996 6580
rect 38052 6524 38444 6580
rect 38500 6524 45500 6580
rect 45556 6524 45566 6580
rect 49746 6524 49756 6580
rect 49812 6524 50428 6580
rect 50484 6524 50494 6580
rect 51314 6524 51324 6580
rect 51380 6524 51390 6580
rect 37548 6468 37604 6524
rect 26786 6412 26796 6468
rect 26852 6412 27244 6468
rect 27300 6412 27310 6468
rect 28242 6412 28252 6468
rect 28308 6412 29596 6468
rect 29652 6412 29662 6468
rect 33030 6412 33068 6468
rect 33124 6412 33134 6468
rect 34626 6412 34636 6468
rect 34692 6412 35644 6468
rect 35700 6412 36988 6468
rect 37044 6412 37054 6468
rect 37548 6412 38108 6468
rect 38164 6412 38668 6468
rect 39106 6412 39116 6468
rect 39172 6412 41020 6468
rect 41076 6412 41086 6468
rect 45266 6412 45276 6468
rect 45332 6412 47292 6468
rect 47348 6412 47358 6468
rect 50194 6412 50204 6468
rect 50260 6412 52780 6468
rect 52836 6412 52846 6468
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 28252 6244 28308 6412
rect 38612 6356 38668 6412
rect 35522 6300 35532 6356
rect 35588 6300 36204 6356
rect 36260 6300 37212 6356
rect 37268 6300 38444 6356
rect 38500 6300 38510 6356
rect 38612 6300 39676 6356
rect 39732 6300 39742 6356
rect 50546 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50830 6300
rect 26562 6188 26572 6244
rect 26628 6188 27132 6244
rect 27188 6188 27198 6244
rect 27346 6188 27356 6244
rect 27412 6188 28308 6244
rect 32274 6188 32284 6244
rect 32340 6188 33292 6244
rect 33348 6188 35196 6244
rect 35252 6188 35262 6244
rect 37314 6188 37324 6244
rect 37380 6188 39228 6244
rect 39284 6188 39294 6244
rect 26450 6076 26460 6132
rect 26516 6076 31500 6132
rect 31556 6076 32844 6132
rect 32900 6076 32910 6132
rect 36306 6076 36316 6132
rect 36372 6076 37100 6132
rect 37156 6076 37660 6132
rect 37716 6076 39564 6132
rect 39620 6076 39630 6132
rect 46274 6076 46284 6132
rect 46340 6076 47740 6132
rect 47796 6076 47806 6132
rect 37202 5964 37212 6020
rect 37268 5964 38892 6020
rect 38948 5964 38958 6020
rect 39788 5964 41356 6020
rect 41412 5964 41422 6020
rect 39788 5908 39844 5964
rect 25666 5852 25676 5908
rect 25732 5852 26460 5908
rect 26516 5852 26526 5908
rect 31042 5852 31052 5908
rect 31108 5852 31500 5908
rect 31556 5852 31566 5908
rect 33730 5852 33740 5908
rect 33796 5852 34524 5908
rect 34580 5852 35644 5908
rect 35700 5852 35710 5908
rect 36082 5852 36092 5908
rect 36148 5852 36764 5908
rect 36820 5852 36830 5908
rect 37762 5852 37772 5908
rect 37828 5852 39844 5908
rect 40002 5852 40012 5908
rect 40068 5852 41804 5908
rect 41860 5852 41870 5908
rect 44146 5852 44156 5908
rect 44212 5852 44828 5908
rect 44884 5852 44894 5908
rect 49298 5852 49308 5908
rect 49364 5852 51100 5908
rect 51156 5852 51166 5908
rect 36092 5796 36148 5852
rect 30930 5740 30940 5796
rect 30996 5740 31612 5796
rect 31668 5740 31678 5796
rect 31938 5740 31948 5796
rect 32004 5740 36148 5796
rect 37884 5740 38892 5796
rect 38948 5740 38958 5796
rect 47842 5740 47852 5796
rect 47908 5740 49196 5796
rect 49252 5740 49868 5796
rect 49924 5740 49934 5796
rect 27234 5628 27244 5684
rect 27300 5628 31388 5684
rect 31444 5628 33404 5684
rect 33460 5628 33470 5684
rect 33618 5628 33628 5684
rect 33684 5628 35196 5684
rect 35252 5628 35262 5684
rect 33170 5516 33180 5572
rect 33236 5516 33964 5572
rect 34020 5516 34030 5572
rect 36418 5516 36428 5572
rect 36484 5516 36876 5572
rect 36932 5516 37660 5572
rect 37716 5516 37726 5572
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 32946 5404 32956 5460
rect 33012 5404 33516 5460
rect 33572 5404 35028 5460
rect 34972 5348 35028 5404
rect 35532 5404 37548 5460
rect 37604 5404 37614 5460
rect 35532 5348 35588 5404
rect 37884 5348 37940 5740
rect 39330 5628 39340 5684
rect 39396 5628 39788 5684
rect 39844 5628 40908 5684
rect 40964 5628 40974 5684
rect 42914 5628 42924 5684
rect 42980 5628 44268 5684
rect 44324 5628 45276 5684
rect 45332 5628 45342 5684
rect 46498 5628 46508 5684
rect 46564 5628 47516 5684
rect 47572 5628 47582 5684
rect 31714 5292 31724 5348
rect 31780 5292 32732 5348
rect 32788 5292 33964 5348
rect 34020 5292 34748 5348
rect 34804 5292 34814 5348
rect 34962 5292 34972 5348
rect 35028 5292 35588 5348
rect 37090 5292 37100 5348
rect 37156 5292 37884 5348
rect 37940 5292 37950 5348
rect 38658 5292 38668 5348
rect 38724 5292 43148 5348
rect 43204 5292 43214 5348
rect 44034 5292 44044 5348
rect 44100 5292 45164 5348
rect 45220 5292 46956 5348
rect 47012 5292 47022 5348
rect 30594 5180 30604 5236
rect 30660 5180 31836 5236
rect 31892 5180 31902 5236
rect 33506 5180 33516 5236
rect 33572 5180 38220 5236
rect 38276 5180 38286 5236
rect 38434 5180 38444 5236
rect 38500 5180 39340 5236
rect 39396 5180 39406 5236
rect 39564 5180 41132 5236
rect 41188 5180 41198 5236
rect 47058 5180 47068 5236
rect 47124 5180 48412 5236
rect 48468 5180 48972 5236
rect 49028 5180 49756 5236
rect 49812 5180 50092 5236
rect 50148 5180 50158 5236
rect 39564 5124 39620 5180
rect 28812 5068 30940 5124
rect 30996 5068 31006 5124
rect 32610 5068 32620 5124
rect 32676 5068 34636 5124
rect 34692 5068 34702 5124
rect 34860 5068 35868 5124
rect 35924 5068 35934 5124
rect 36306 5068 36316 5124
rect 36372 5068 37212 5124
rect 37268 5068 37278 5124
rect 37650 5068 37660 5124
rect 37716 5068 39620 5124
rect 39778 5068 39788 5124
rect 39844 5068 41356 5124
rect 41412 5068 41422 5124
rect 43026 5068 43036 5124
rect 43092 5068 43708 5124
rect 43764 5068 44716 5124
rect 44772 5068 44782 5124
rect 45714 5068 45724 5124
rect 45780 5068 48188 5124
rect 48244 5068 48254 5124
rect 28812 5012 28868 5068
rect 29372 5012 29428 5068
rect 34860 5012 34916 5068
rect 28802 4956 28812 5012
rect 28868 4956 28878 5012
rect 29362 4956 29372 5012
rect 29428 4956 29438 5012
rect 32722 4956 32732 5012
rect 32788 4956 34300 5012
rect 34356 4956 34916 5012
rect 35634 4956 35644 5012
rect 35700 4956 37772 5012
rect 37828 4956 37838 5012
rect 33058 4844 33068 4900
rect 33124 4844 33628 4900
rect 33684 4844 33694 4900
rect 35410 4844 35420 4900
rect 35476 4844 37548 4900
rect 37604 4844 42252 4900
rect 42308 4844 42812 4900
rect 42868 4844 42878 4900
rect 36754 4732 36764 4788
rect 36820 4732 40684 4788
rect 40740 4732 40750 4788
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 50546 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50830 4732
rect 33170 4620 33180 4676
rect 33236 4620 34748 4676
rect 34804 4620 34814 4676
rect 29474 4508 29484 4564
rect 29540 4508 31388 4564
rect 31444 4508 32060 4564
rect 32116 4508 32126 4564
rect 38210 4508 38220 4564
rect 38276 4508 40908 4564
rect 40964 4508 40974 4564
rect 42354 4508 42364 4564
rect 42420 4508 45164 4564
rect 45220 4508 45230 4564
rect 35186 4284 35196 4340
rect 35252 4284 36988 4340
rect 37044 4284 37054 4340
rect 40002 4284 40012 4340
rect 40068 4284 42028 4340
rect 42084 4284 42364 4340
rect 42420 4284 42430 4340
rect 43138 4284 43148 4340
rect 43204 4284 44940 4340
rect 44996 4284 45006 4340
rect 43148 4228 43204 4284
rect 42130 4172 42140 4228
rect 42196 4172 43204 4228
rect 44146 4172 44156 4228
rect 44212 4172 44716 4228
rect 44772 4172 44782 4228
rect 33618 4060 33628 4116
rect 33684 4060 34860 4116
rect 34916 4060 34926 4116
rect 36306 3948 36316 4004
rect 36372 3948 40908 4004
rect 40964 3948 43372 4004
rect 43428 3948 43438 4004
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 40338 3836 40348 3892
rect 40404 3836 45724 3892
rect 45780 3836 46620 3892
rect 46676 3836 47404 3892
rect 47460 3836 47470 3892
rect 35074 3724 35084 3780
rect 35140 3724 37212 3780
rect 37268 3724 37278 3780
rect 37426 3724 37436 3780
rect 37492 3724 42364 3780
rect 42420 3724 42700 3780
rect 42756 3724 44604 3780
rect 44660 3724 44670 3780
rect 34962 3612 34972 3668
rect 35028 3612 36204 3668
rect 36260 3612 36270 3668
rect 36428 3612 38892 3668
rect 38948 3612 38958 3668
rect 39666 3612 39676 3668
rect 39732 3612 43820 3668
rect 43876 3612 43886 3668
rect 36428 3556 36484 3612
rect 25106 3500 25116 3556
rect 25172 3500 26012 3556
rect 26068 3500 26078 3556
rect 33506 3500 33516 3556
rect 33572 3500 34636 3556
rect 34692 3500 34702 3556
rect 34850 3500 34860 3556
rect 34916 3500 36484 3556
rect 36978 3500 36988 3556
rect 37044 3500 41580 3556
rect 41636 3500 46284 3556
rect 46340 3500 46350 3556
rect 28354 3388 28364 3444
rect 28420 3388 30268 3444
rect 30324 3388 30334 3444
rect 33292 3388 33964 3444
rect 34020 3388 34030 3444
rect 34402 3388 34412 3444
rect 34468 3388 35532 3444
rect 35588 3388 39116 3444
rect 39172 3388 39182 3444
rect 43138 3388 43148 3444
rect 43204 3388 44604 3444
rect 44660 3388 46732 3444
rect 46788 3388 46798 3444
rect 33292 3332 33348 3388
rect 33282 3276 33292 3332
rect 33348 3276 33358 3332
rect 43652 3276 46508 3332
rect 46564 3276 46574 3332
rect 29362 3164 29372 3220
rect 29428 3164 39004 3220
rect 39060 3164 40012 3220
rect 40068 3164 40078 3220
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 43652 3108 43708 3276
rect 50546 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50830 3164
rect 33058 3052 33068 3108
rect 33124 3052 43708 3108
<< via3 >>
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 50556 45444 50612 45500
rect 50660 45444 50716 45500
rect 50764 45444 50820 45500
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 50556 43876 50612 43932
rect 50660 43876 50716 43932
rect 50764 43876 50820 43932
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 50556 42308 50612 42364
rect 50660 42308 50716 42364
rect 50764 42308 50820 42364
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 50556 40740 50612 40796
rect 50660 40740 50716 40796
rect 50764 40740 50820 40796
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 50556 39172 50612 39228
rect 50660 39172 50716 39228
rect 50764 39172 50820 39228
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 50556 37604 50612 37660
rect 50660 37604 50716 37660
rect 50764 37604 50820 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 50556 36036 50612 36092
rect 50660 36036 50716 36092
rect 50764 36036 50820 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 9660 34748 9716 34804
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 50556 34468 50612 34524
rect 50660 34468 50716 34524
rect 50764 34468 50820 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 9660 33068 9716 33124
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 50556 32900 50612 32956
rect 50660 32900 50716 32956
rect 50764 32900 50820 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 50556 31332 50612 31388
rect 50660 31332 50716 31388
rect 50764 31332 50820 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 50556 29764 50612 29820
rect 50660 29764 50716 29820
rect 50764 29764 50820 29820
rect 17500 29260 17556 29316
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 20748 28924 20804 28980
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 50556 28196 50612 28252
rect 50660 28196 50716 28252
rect 50764 28196 50820 28252
rect 20748 27916 20804 27972
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 20748 27020 20804 27076
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 17500 26572 17556 26628
rect 50556 26628 50612 26684
rect 50660 26628 50716 26684
rect 50764 26628 50820 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 50556 25060 50612 25116
rect 50660 25060 50716 25116
rect 50764 25060 50820 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 50556 23492 50612 23548
rect 50660 23492 50716 23548
rect 50764 23492 50820 23548
rect 26908 23324 26964 23380
rect 26908 22988 26964 23044
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 50556 21924 50612 21980
rect 50660 21924 50716 21980
rect 50764 21924 50820 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 50556 20356 50612 20412
rect 50660 20356 50716 20412
rect 50764 20356 50820 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 50556 18788 50612 18844
rect 50660 18788 50716 18844
rect 50764 18788 50820 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 23100 17836 23156 17892
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 50556 17220 50612 17276
rect 50660 17220 50716 17276
rect 50764 17220 50820 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 50556 15652 50612 15708
rect 50660 15652 50716 15708
rect 50764 15652 50820 15708
rect 38332 14924 38388 14980
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 50556 14084 50612 14140
rect 50660 14084 50716 14140
rect 50764 14084 50820 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 23100 13020 23156 13076
rect 38332 12796 38388 12852
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 50556 12516 50612 12572
rect 50660 12516 50716 12572
rect 50764 12516 50820 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 50556 10948 50612 11004
rect 50660 10948 50716 11004
rect 50764 10948 50820 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 31836 9996 31892 10052
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 50556 9380 50612 9436
rect 50660 9380 50716 9436
rect 50764 9380 50820 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 50556 7812 50612 7868
rect 50660 7812 50716 7868
rect 50764 7812 50820 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 33068 6412 33124 6468
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 50556 6244 50612 6300
rect 50660 6244 50716 6300
rect 50764 6244 50820 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 31836 5180 31892 5236
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 50556 4676 50612 4732
rect 50660 4676 50716 4732
rect 50764 4676 50820 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
rect 50556 3108 50612 3164
rect 50660 3108 50716 3164
rect 50764 3108 50820 3164
rect 33068 3052 33124 3108
<< metal4 >>
rect 4448 46284 4768 46316
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 19808 45500 20128 46316
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 19808 43932 20128 45444
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 19808 42364 20128 43876
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 9660 34804 9716 34814
rect 9660 33124 9716 34748
rect 9660 33058 9716 33068
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 17500 29316 17556 29326
rect 17500 26628 17556 29260
rect 17500 26562 17556 26572
rect 19808 28252 20128 29764
rect 35168 46284 35488 46316
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 20748 28980 20804 28990
rect 20748 27972 20804 28924
rect 20748 27076 20804 27916
rect 20748 27010 20804 27020
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 26908 23380 26964 23390
rect 26908 23044 26964 23324
rect 26908 22978 26964 22988
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 23100 17892 23156 17902
rect 23100 13076 23156 17836
rect 23100 13010 23156 13020
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 50528 45500 50848 46316
rect 50528 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50848 45500
rect 50528 43932 50848 45444
rect 50528 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50848 43932
rect 50528 42364 50848 43876
rect 50528 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50848 42364
rect 50528 40796 50848 42308
rect 50528 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50848 40796
rect 50528 39228 50848 40740
rect 50528 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50848 39228
rect 50528 37660 50848 39172
rect 50528 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50848 37660
rect 50528 36092 50848 37604
rect 50528 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50848 36092
rect 50528 34524 50848 36036
rect 50528 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50848 34524
rect 50528 32956 50848 34468
rect 50528 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50848 32956
rect 50528 31388 50848 32900
rect 50528 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50848 31388
rect 50528 29820 50848 31332
rect 50528 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50848 29820
rect 50528 28252 50848 29764
rect 50528 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50848 28252
rect 50528 26684 50848 28196
rect 50528 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50848 26684
rect 50528 25116 50848 26628
rect 50528 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50848 25116
rect 50528 23548 50848 25060
rect 50528 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50848 23548
rect 50528 21980 50848 23492
rect 50528 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50848 21980
rect 50528 20412 50848 21924
rect 50528 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50848 20412
rect 50528 18844 50848 20356
rect 50528 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50848 18844
rect 50528 17276 50848 18788
rect 50528 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50848 17276
rect 50528 15708 50848 17220
rect 50528 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50848 15708
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 35168 11788 35488 13300
rect 38332 14980 38388 14990
rect 38332 12852 38388 14924
rect 38332 12786 38388 12796
rect 50528 14140 50848 15652
rect 50528 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50848 14140
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 31836 10052 31892 10062
rect 31836 5236 31892 9996
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 31836 5170 31892 5180
rect 33068 6468 33124 6478
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 33068 3108 33124 6412
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
rect 50528 12572 50848 14084
rect 50528 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50848 12572
rect 50528 11004 50848 12516
rect 50528 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50848 11004
rect 50528 9436 50848 10948
rect 50528 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50848 9436
rect 50528 7868 50848 9380
rect 50528 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50848 7868
rect 50528 6300 50848 7812
rect 50528 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50848 6300
rect 50528 4732 50848 6244
rect 50528 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50848 4732
rect 50528 3164 50848 4676
rect 50528 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50848 3164
rect 50528 3076 50848 3108
rect 33068 3042 33124 3052
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1482_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 44240 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1483_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 42784 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1484_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 44576 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1485_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 44576 0 -1 28224
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1486_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 44688 0 1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1487_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 46704 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1488_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 46704 0 -1 25088
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1489_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 44016 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1490_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 45472 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1491_
timestamp 1698431365
transform 1 0 28000 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1492_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 30128 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1493_
timestamp 1698431365
transform 1 0 30576 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1494_
timestamp 1698431365
transform 1 0 28336 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1495_
timestamp 1698431365
transform 1 0 28672 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1496_
timestamp 1698431365
transform 1 0 29904 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1497_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 38192 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1498_
timestamp 1698431365
transform 1 0 30688 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1499_
timestamp 1698431365
transform 1 0 38416 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1500_
timestamp 1698431365
transform 1 0 33936 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1501_
timestamp 1698431365
transform 1 0 37744 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1502_
timestamp 1698431365
transform -1 0 39536 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1503_
timestamp 1698431365
transform 1 0 38640 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1504_
timestamp 1698431365
transform -1 0 30128 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1505_
timestamp 1698431365
transform 1 0 30800 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1506_
timestamp 1698431365
transform 1 0 26992 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1507_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29008 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1508_
timestamp 1698431365
transform -1 0 29568 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1509_
timestamp 1698431365
transform 1 0 26320 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1510_
timestamp 1698431365
transform 1 0 26992 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1511_
timestamp 1698431365
transform -1 0 30688 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1512_
timestamp 1698431365
transform 1 0 30912 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1513_
timestamp 1698431365
transform 1 0 31360 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1514_
timestamp 1698431365
transform 1 0 25648 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1515_
timestamp 1698431365
transform 1 0 32032 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1516_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 32816 0 1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1517_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 29344 0 -1 9408
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1518_
timestamp 1698431365
transform -1 0 26768 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1519_
timestamp 1698431365
transform -1 0 30912 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1520_
timestamp 1698431365
transform -1 0 25872 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1521_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 25200 0 1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1522_
timestamp 1698431365
transform 1 0 24192 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1523_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 27664 0 1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1524_
timestamp 1698431365
transform 1 0 37520 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1525_
timestamp 1698431365
transform 1 0 26768 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1526_
timestamp 1698431365
transform -1 0 32256 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1527_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29008 0 1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1528_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 27888 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1529_
timestamp 1698431365
transform 1 0 22176 0 -1 7840
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1530_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 24864 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1531_
timestamp 1698431365
transform 1 0 27328 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1532_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 24416 0 1 10976
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1533_
timestamp 1698431365
transform 1 0 29344 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1534_
timestamp 1698431365
transform -1 0 37520 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1535_
timestamp 1698431365
transform -1 0 34832 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1536_
timestamp 1698431365
transform -1 0 31472 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1537_
timestamp 1698431365
transform 1 0 27104 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1538_
timestamp 1698431365
transform 1 0 26544 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1539_
timestamp 1698431365
transform 1 0 27328 0 -1 7840
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1540_
timestamp 1698431365
transform -1 0 31136 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1541_
timestamp 1698431365
transform -1 0 28784 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1542_
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1543_
timestamp 1698431365
transform 1 0 25648 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1544_
timestamp 1698431365
transform 1 0 26656 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1545_
timestamp 1698431365
transform 1 0 26880 0 1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1546_
timestamp 1698431365
transform -1 0 31248 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1547_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25648 0 -1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1548_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25424 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1549_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 28784 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1550_
timestamp 1698431365
transform 1 0 27440 0 -1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1551_
timestamp 1698431365
transform 1 0 33936 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1552_
timestamp 1698431365
transform -1 0 33824 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1553_
timestamp 1698431365
transform 1 0 28112 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1554_
timestamp 1698431365
transform -1 0 39648 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1555_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 31136 0 -1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1556_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 34944 0 -1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1557_
timestamp 1698431365
transform -1 0 33600 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1558_
timestamp 1698431365
transform 1 0 35056 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1559_
timestamp 1698431365
transform 1 0 35504 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1560_
timestamp 1698431365
transform -1 0 36288 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1561_
timestamp 1698431365
transform 1 0 34944 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1562_
timestamp 1698431365
transform 1 0 32816 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1563_
timestamp 1698431365
transform 1 0 34048 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1564_
timestamp 1698431365
transform 1 0 33488 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1565_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 35504 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1566_
timestamp 1698431365
transform -1 0 36400 0 -1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1567_
timestamp 1698431365
transform 1 0 32704 0 1 12544
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1568_
timestamp 1698431365
transform 1 0 34496 0 -1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1569_
timestamp 1698431365
transform 1 0 46032 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1570_
timestamp 1698431365
transform 1 0 43120 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1571_
timestamp 1698431365
transform -1 0 44688 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1572_
timestamp 1698431365
transform 1 0 32704 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1573_
timestamp 1698431365
transform 1 0 31920 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1574_
timestamp 1698431365
transform 1 0 32368 0 1 4704
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1575_
timestamp 1698431365
transform 1 0 40768 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1576_
timestamp 1698431365
transform 1 0 31248 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1577_
timestamp 1698431365
transform -1 0 33600 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1578_
timestamp 1698431365
transform 1 0 34272 0 -1 6272
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1579_
timestamp 1698431365
transform 1 0 34832 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1580_
timestamp 1698431365
transform -1 0 32704 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1581_
timestamp 1698431365
transform 1 0 31696 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1582_
timestamp 1698431365
transform 1 0 35056 0 1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1583_
timestamp 1698431365
transform 1 0 36848 0 1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1584_
timestamp 1698431365
transform 1 0 36064 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1585_
timestamp 1698431365
transform -1 0 41328 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1586_
timestamp 1698431365
transform -1 0 39424 0 1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1587_
timestamp 1698431365
transform 1 0 39648 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1588_
timestamp 1698431365
transform 1 0 36400 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1589_
timestamp 1698431365
transform -1 0 41888 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1590_
timestamp 1698431365
transform -1 0 36624 0 1 4704
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1591_
timestamp 1698431365
transform 1 0 42672 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1592_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 35616 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _1593_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 38192 0 1 4704
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _1594_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 38080 0 -1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1595_
timestamp 1698431365
transform 1 0 40544 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1596_
timestamp 1698431365
transform 1 0 40656 0 1 6272
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1597_
timestamp 1698431365
transform 1 0 43792 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1598_
timestamp 1698431365
transform 1 0 42784 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1599_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 39872 0 1 6272
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1600_
timestamp 1698431365
transform 1 0 39648 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1601_
timestamp 1698431365
transform -1 0 42224 0 -1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1602_
timestamp 1698431365
transform 1 0 42224 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1603_
timestamp 1698431365
transform 1 0 33376 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1604_
timestamp 1698431365
transform 1 0 33600 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1605_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 36624 0 -1 4704
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1606_
timestamp 1698431365
transform 1 0 44464 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1607_
timestamp 1698431365
transform 1 0 36848 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1608_
timestamp 1698431365
transform -1 0 29680 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1609_
timestamp 1698431365
transform 1 0 38864 0 -1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1610_
timestamp 1698431365
transform -1 0 44464 0 -1 4704
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1611_
timestamp 1698431365
transform 1 0 41888 0 1 7840
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1612_
timestamp 1698431365
transform -1 0 44240 0 -1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1613_
timestamp 1698431365
transform -1 0 43792 0 1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1614_
timestamp 1698431365
transform 1 0 26880 0 -1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1615_
timestamp 1698431365
transform 1 0 29680 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1616_
timestamp 1698431365
transform -1 0 31696 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1617_
timestamp 1698431365
transform 1 0 30128 0 1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1618_
timestamp 1698431365
transform 1 0 37968 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1619_
timestamp 1698431365
transform 1 0 35616 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1620_
timestamp 1698431365
transform -1 0 39088 0 1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1621_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 38080 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1622_
timestamp 1698431365
transform -1 0 46144 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1623_
timestamp 1698431365
transform -1 0 38416 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1624_
timestamp 1698431365
transform -1 0 30912 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1625_
timestamp 1698431365
transform 1 0 30912 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1626_
timestamp 1698431365
transform 1 0 31584 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1627_
timestamp 1698431365
transform 1 0 30128 0 -1 10976
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1628_
timestamp 1698431365
transform 1 0 37296 0 1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1629_
timestamp 1698431365
transform -1 0 39536 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1630_
timestamp 1698431365
transform 1 0 32704 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1631_
timestamp 1698431365
transform -1 0 35280 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1632_
timestamp 1698431365
transform -1 0 34384 0 -1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1633_
timestamp 1698431365
transform 1 0 26208 0 1 12544
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1634_
timestamp 1698431365
transform 1 0 37632 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1635_
timestamp 1698431365
transform -1 0 38752 0 -1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1636_
timestamp 1698431365
transform 1 0 30464 0 1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1637_
timestamp 1698431365
transform -1 0 32480 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1638_
timestamp 1698431365
transform -1 0 32480 0 -1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1639_
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1640_
timestamp 1698431365
transform 1 0 29232 0 -1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1641_
timestamp 1698431365
transform 1 0 35280 0 -1 15680
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1642_
timestamp 1698431365
transform 1 0 28336 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1643_
timestamp 1698431365
transform 1 0 31248 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1644_
timestamp 1698431365
transform 1 0 35952 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1645_
timestamp 1698431365
transform -1 0 37520 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1646_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 39984 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1647_
timestamp 1698431365
transform 1 0 43008 0 1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1648_
timestamp 1698431365
transform 1 0 43792 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1649_
timestamp 1698431365
transform -1 0 43792 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1650_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 42448 0 -1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1651_
timestamp 1698431365
transform -1 0 41440 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1652_
timestamp 1698431365
transform -1 0 40432 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1653_
timestamp 1698431365
transform 1 0 38640 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1654_
timestamp 1698431365
transform 1 0 39312 0 -1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1655_
timestamp 1698431365
transform 1 0 39200 0 1 15680
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1656_
timestamp 1698431365
transform -1 0 35280 0 1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1657_
timestamp 1698431365
transform 1 0 33600 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1658_
timestamp 1698431365
transform 1 0 35280 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1659_
timestamp 1698431365
transform -1 0 36288 0 -1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1660_
timestamp 1698431365
transform 1 0 41216 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1661_
timestamp 1698431365
transform -1 0 41888 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1662_
timestamp 1698431365
transform 1 0 40432 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1663_
timestamp 1698431365
transform 1 0 36064 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1664_
timestamp 1698431365
transform 1 0 39088 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1665_
timestamp 1698431365
transform 1 0 40768 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1666_
timestamp 1698431365
transform 1 0 41328 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1667_
timestamp 1698431365
transform -1 0 42560 0 1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1668_
timestamp 1698431365
transform 1 0 36400 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1669_
timestamp 1698431365
transform 1 0 36288 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1670_
timestamp 1698431365
transform 1 0 41888 0 1 12544
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1671_
timestamp 1698431365
transform 1 0 43792 0 -1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1672_
timestamp 1698431365
transform 1 0 43456 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1673_
timestamp 1698431365
transform 1 0 42336 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _1674_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 43456 0 -1 9408
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1675_
timestamp 1698431365
transform 1 0 45472 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1676_
timestamp 1698431365
transform -1 0 42672 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1677_
timestamp 1698431365
transform -1 0 45472 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1678_
timestamp 1698431365
transform 1 0 42000 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1679_
timestamp 1698431365
transform 1 0 44688 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1680_
timestamp 1698431365
transform 1 0 43680 0 1 4704
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1681_
timestamp 1698431365
transform 1 0 44016 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1682_
timestamp 1698431365
transform -1 0 46256 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1683_
timestamp 1698431365
transform 1 0 39648 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1684_
timestamp 1698431365
transform 1 0 45472 0 1 3136
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1685_
timestamp 1698431365
transform 1 0 33152 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1686_
timestamp 1698431365
transform 1 0 32592 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1687_
timestamp 1698431365
transform 1 0 45920 0 -1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _1688_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 45136 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1689_
timestamp 1698431365
transform 1 0 45360 0 1 7840
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1690_
timestamp 1698431365
transform -1 0 46928 0 -1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1691_
timestamp 1698431365
transform -1 0 36512 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1692_
timestamp 1698431365
transform -1 0 35840 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1693_
timestamp 1698431365
transform 1 0 36848 0 1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1694_
timestamp 1698431365
transform -1 0 46144 0 -1 15680
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1695_
timestamp 1698431365
transform 1 0 37520 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _1696_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 40432 0 1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1697_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 44688 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1698_
timestamp 1698431365
transform 1 0 44688 0 1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1699_
timestamp 1698431365
transform -1 0 44016 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1700_
timestamp 1698431365
transform -1 0 39312 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1701_
timestamp 1698431365
transform -1 0 38752 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1702_
timestamp 1698431365
transform -1 0 40096 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1703_
timestamp 1698431365
transform 1 0 37856 0 -1 14112
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1704_
timestamp 1698431365
transform -1 0 48272 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1705_
timestamp 1698431365
transform -1 0 51856 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1706_
timestamp 1698431365
transform -1 0 47824 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1707_
timestamp 1698431365
transform 1 0 46032 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1708_
timestamp 1698431365
transform 1 0 41776 0 -1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1709_
timestamp 1698431365
transform 1 0 46480 0 1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1710_
timestamp 1698431365
transform 1 0 44688 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1711_
timestamp 1698431365
transform 1 0 42896 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _1712_
timestamp 1698431365
transform 1 0 43456 0 -1 12544
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1713_
timestamp 1698431365
transform 1 0 46256 0 -1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1714_
timestamp 1698431365
transform 1 0 46480 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1715_
timestamp 1698431365
transform 1 0 47600 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1716_
timestamp 1698431365
transform 1 0 46704 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1717_
timestamp 1698431365
transform 1 0 47824 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1718_
timestamp 1698431365
transform 1 0 47040 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1719_
timestamp 1698431365
transform -1 0 47936 0 1 4704
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1720_
timestamp 1698431365
transform 1 0 47264 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1721_
timestamp 1698431365
transform -1 0 48832 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1722_
timestamp 1698431365
transform -1 0 48608 0 1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1723_
timestamp 1698431365
transform 1 0 49728 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1724_
timestamp 1698431365
transform -1 0 51408 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1725_
timestamp 1698431365
transform 1 0 47376 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1726_
timestamp 1698431365
transform 1 0 48832 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1727_
timestamp 1698431365
transform 1 0 35728 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1728_
timestamp 1698431365
transform 1 0 36512 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1729_
timestamp 1698431365
transform 1 0 48608 0 1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1730_
timestamp 1698431365
transform -1 0 52192 0 -1 6272
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1731_
timestamp 1698431365
transform 1 0 47712 0 1 9408
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1732_
timestamp 1698431365
transform -1 0 50064 0 -1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1733_
timestamp 1698431365
transform -1 0 46704 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1734_
timestamp 1698431365
transform -1 0 45472 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1735_
timestamp 1698431365
transform 1 0 44912 0 1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1736_
timestamp 1698431365
transform -1 0 48944 0 1 15680
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1737_
timestamp 1698431365
transform 1 0 39984 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1738_
timestamp 1698431365
transform -1 0 50288 0 -1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1739_
timestamp 1698431365
transform -1 0 49280 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1740_
timestamp 1698431365
transform 1 0 48160 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1741_
timestamp 1698431365
transform 1 0 47600 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1742_
timestamp 1698431365
transform 1 0 48608 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1743_
timestamp 1698431365
transform -1 0 51632 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1744_
timestamp 1698431365
transform -1 0 51632 0 1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1745_
timestamp 1698431365
transform 1 0 49840 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1746_
timestamp 1698431365
transform 1 0 47488 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1747_
timestamp 1698431365
transform 1 0 49168 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1748_
timestamp 1698431365
transform 1 0 51520 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1749_
timestamp 1698431365
transform 1 0 49952 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1750_
timestamp 1698431365
transform -1 0 53088 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1751_
timestamp 1698431365
transform 1 0 49728 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1752_
timestamp 1698431365
transform 1 0 50848 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1753_
timestamp 1698431365
transform 1 0 50064 0 -1 7840
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1754_
timestamp 1698431365
transform 1 0 50848 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1755_
timestamp 1698431365
transform 1 0 52640 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1756_
timestamp 1698431365
transform 1 0 48608 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1757_
timestamp 1698431365
transform 1 0 53088 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1758_
timestamp 1698431365
transform 1 0 39984 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1759_
timestamp 1698431365
transform 1 0 38640 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1760_
timestamp 1698431365
transform 1 0 39648 0 1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _1761_
timestamp 1698431365
transform 1 0 52976 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1762_
timestamp 1698431365
transform -1 0 58352 0 1 7840
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1763_
timestamp 1698431365
transform 1 0 49392 0 1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1764_
timestamp 1698431365
transform 1 0 47488 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1765_
timestamp 1698431365
transform 1 0 46928 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1766_
timestamp 1698431365
transform 1 0 47712 0 1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1767_
timestamp 1698431365
transform -1 0 51296 0 -1 15680
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1768_
timestamp 1698431365
transform -1 0 39872 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1769_
timestamp 1698431365
transform -1 0 40432 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1770_
timestamp 1698431365
transform 1 0 39088 0 -1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1771_
timestamp 1698431365
transform 1 0 40432 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1772_
timestamp 1698431365
transform 1 0 40768 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1773_
timestamp 1698431365
transform 1 0 40992 0 1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1774_
timestamp 1698431365
transform -1 0 36624 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1775_
timestamp 1698431365
transform -1 0 41888 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1776_
timestamp 1698431365
transform 1 0 41888 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1777_
timestamp 1698431365
transform -1 0 42896 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1778_
timestamp 1698431365
transform -1 0 50288 0 -1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1779_
timestamp 1698431365
transform -1 0 48160 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1780_
timestamp 1698431365
transform -1 0 40432 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1781_
timestamp 1698431365
transform 1 0 49616 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1782_
timestamp 1698431365
transform 1 0 50512 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1783_
timestamp 1698431365
transform -1 0 51632 0 1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1784_
timestamp 1698431365
transform -1 0 57792 0 -1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1785_
timestamp 1698431365
transform -1 0 56224 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1786_
timestamp 1698431365
transform 1 0 49840 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1787_
timestamp 1698431365
transform 1 0 55104 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1788_
timestamp 1698431365
transform 1 0 51744 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1789_
timestamp 1698431365
transform -1 0 54320 0 1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1790_
timestamp 1698431365
transform 1 0 52752 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1791_
timestamp 1698431365
transform 1 0 53872 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1792_
timestamp 1698431365
transform 1 0 56448 0 -1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1793_
timestamp 1698431365
transform 1 0 53536 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1794_
timestamp 1698431365
transform 1 0 51632 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1795_
timestamp 1698431365
transform -1 0 41216 0 1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1796_
timestamp 1698431365
transform -1 0 53872 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1797_
timestamp 1698431365
transform 1 0 55328 0 1 9408
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1798_
timestamp 1698431365
transform 1 0 55328 0 1 10976
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1799_
timestamp 1698431365
transform -1 0 57792 0 -1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1800_
timestamp 1698431365
transform -1 0 53984 0 1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _1801_
timestamp 1698431365
transform 1 0 40768 0 -1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1802_
timestamp 1698431365
transform -1 0 47040 0 -1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1803_
timestamp 1698431365
transform 1 0 44688 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1804_
timestamp 1698431365
transform 1 0 33712 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1805_
timestamp 1698431365
transform -1 0 57904 0 -1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1806_
timestamp 1698431365
transform 1 0 56560 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1807_
timestamp 1698431365
transform 1 0 55664 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1808_
timestamp 1698431365
transform 1 0 51744 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1809_
timestamp 1698431365
transform -1 0 53984 0 1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1810_
timestamp 1698431365
transform -1 0 53536 0 -1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1811_
timestamp 1698431365
transform 1 0 53872 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1812_
timestamp 1698431365
transform 1 0 53984 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1813_
timestamp 1698431365
transform 1 0 56448 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1814_
timestamp 1698431365
transform -1 0 55328 0 1 10976
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1815_
timestamp 1698431365
transform 1 0 54544 0 -1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1816_
timestamp 1698431365
transform 1 0 52528 0 1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1817_
timestamp 1698431365
transform 1 0 52416 0 -1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1818_
timestamp 1698431365
transform 1 0 54656 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1819_
timestamp 1698431365
transform -1 0 54656 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or4_2  _1820_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 53312 0 -1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1821_
timestamp 1698431365
transform -1 0 52304 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _1822_
timestamp 1698431365
transform 1 0 52528 0 1 14112
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1823_
timestamp 1698431365
transform -1 0 36736 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _1824_
timestamp 1698431365
transform 1 0 34384 0 1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1825_
timestamp 1698431365
transform -1 0 42784 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1826_
timestamp 1698431365
transform 1 0 33824 0 -1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1827_
timestamp 1698431365
transform 1 0 33040 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1828_
timestamp 1698431365
transform 1 0 31696 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1829_
timestamp 1698431365
transform 1 0 31248 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1830_
timestamp 1698431365
transform -1 0 53984 0 1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1831_
timestamp 1698431365
transform 1 0 51520 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1832_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 56224 0 -1 12544
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1833_
timestamp 1698431365
transform -1 0 53088 0 -1 17248
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _1834_
timestamp 1698431365
transform 1 0 32144 0 1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1835_
timestamp 1698431365
transform 1 0 30128 0 1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1836_
timestamp 1698431365
transform -1 0 30128 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1837_
timestamp 1698431365
transform -1 0 52976 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1838_
timestamp 1698431365
transform 1 0 50512 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1839_
timestamp 1698431365
transform 1 0 51408 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1840_
timestamp 1698431365
transform 1 0 51296 0 -1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1841_
timestamp 1698431365
transform 1 0 27888 0 -1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1842_
timestamp 1698431365
transform 1 0 29904 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1843_
timestamp 1698431365
transform 1 0 29008 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1844_
timestamp 1698431365
transform -1 0 38192 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1845_
timestamp 1698431365
transform 1 0 36848 0 1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1846_
timestamp 1698431365
transform -1 0 36624 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1847_
timestamp 1698431365
transform 1 0 44688 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1848_
timestamp 1698431365
transform -1 0 46592 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1849_
timestamp 1698431365
transform -1 0 29904 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1850_
timestamp 1698431365
transform -1 0 29680 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1851_
timestamp 1698431365
transform 1 0 31472 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1852_
timestamp 1698431365
transform -1 0 37856 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1853_
timestamp 1698431365
transform 1 0 3808 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1854_
timestamp 1698431365
transform -1 0 14112 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1855_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 14560 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1856_
timestamp 1698431365
transform 1 0 5376 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1857_
timestamp 1698431365
transform 1 0 2688 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1858_
timestamp 1698431365
transform 1 0 3360 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1859_
timestamp 1698431365
transform 1 0 6048 0 -1 12544
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1860_
timestamp 1698431365
transform 1 0 4032 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1861_
timestamp 1698431365
transform 1 0 6048 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1862_
timestamp 1698431365
transform 1 0 5824 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1863_
timestamp 1698431365
transform 1 0 6496 0 1 12544
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1864_
timestamp 1698431365
transform 1 0 6832 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1865_
timestamp 1698431365
transform 1 0 8176 0 -1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1866_
timestamp 1698431365
transform 1 0 8512 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1867_
timestamp 1698431365
transform 1 0 7280 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1868_
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1869_
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1870_
timestamp 1698431365
transform -1 0 12320 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1871_
timestamp 1698431365
transform -1 0 11760 0 1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1872_
timestamp 1698431365
transform 1 0 2016 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1873_
timestamp 1698431365
transform 1 0 2576 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1874_
timestamp 1698431365
transform 1 0 3920 0 -1 9408
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1875_
timestamp 1698431365
transform 1 0 6160 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1876_
timestamp 1698431365
transform 1 0 3472 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _1877_
timestamp 1698431365
transform 1 0 8064 0 1 9408
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__or4_2  _1878_
timestamp 1698431365
transform 1 0 7616 0 -1 10976
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1879_
timestamp 1698431365
transform 1 0 9632 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1880_
timestamp 1698431365
transform -1 0 11648 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1881_
timestamp 1698431365
transform -1 0 11088 0 1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1882_
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1883_
timestamp 1698431365
transform -1 0 12544 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1884_
timestamp 1698431365
transform 1 0 11200 0 -1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1885_
timestamp 1698431365
transform -1 0 13104 0 1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1886_
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1887_
timestamp 1698431365
transform 1 0 7392 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1888_
timestamp 1698431365
transform 1 0 4480 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1889_
timestamp 1698431365
transform 1 0 6160 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1890_
timestamp 1698431365
transform -1 0 7392 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1891_
timestamp 1698431365
transform -1 0 4368 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1892_
timestamp 1698431365
transform -1 0 8400 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1893_
timestamp 1698431365
transform -1 0 4256 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1894_
timestamp 1698431365
transform -1 0 4032 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1895_
timestamp 1698431365
transform 1 0 2016 0 1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1896_
timestamp 1698431365
transform -1 0 3136 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1897_
timestamp 1698431365
transform -1 0 7840 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1898_
timestamp 1698431365
transform 1 0 4256 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1899_
timestamp 1698431365
transform 1 0 4368 0 -1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1900_
timestamp 1698431365
transform 1 0 2576 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1901_
timestamp 1698431365
transform -1 0 5936 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1902_
timestamp 1698431365
transform -1 0 7056 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1903_
timestamp 1698431365
transform -1 0 6384 0 -1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1904_
timestamp 1698431365
transform 1 0 4816 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1905_
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1906_
timestamp 1698431365
transform -1 0 3248 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1907_
timestamp 1698431365
transform -1 0 3248 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1908_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7728 0 1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1909_
timestamp 1698431365
transform -1 0 7504 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1910_
timestamp 1698431365
transform -1 0 7504 0 1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1911_
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1912_
timestamp 1698431365
transform 1 0 4480 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1913_
timestamp 1698431365
transform -1 0 3360 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1914_
timestamp 1698431365
transform 1 0 2688 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1915_
timestamp 1698431365
transform -1 0 4704 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1916_
timestamp 1698431365
transform 1 0 3248 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1917_
timestamp 1698431365
transform 1 0 3024 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1918_
timestamp 1698431365
transform -1 0 7504 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1919_
timestamp 1698431365
transform 1 0 3808 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1920_
timestamp 1698431365
transform -1 0 7056 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1921_
timestamp 1698431365
transform -1 0 6384 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1922_
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1923_
timestamp 1698431365
transform -1 0 7840 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1924_
timestamp 1698431365
transform -1 0 6944 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1925_
timestamp 1698431365
transform 1 0 2240 0 -1 20384
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1926_
timestamp 1698431365
transform -1 0 5712 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1927_
timestamp 1698431365
transform 1 0 4256 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1928_
timestamp 1698431365
transform 1 0 4480 0 -1 23520
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1929_
timestamp 1698431365
transform 1 0 9408 0 1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1930_
timestamp 1698431365
transform 1 0 10864 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1931_
timestamp 1698431365
transform 1 0 6944 0 -1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1932_
timestamp 1698431365
transform 1 0 14672 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1933_
timestamp 1698431365
transform 1 0 9856 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1934_
timestamp 1698431365
transform 1 0 11984 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1935_
timestamp 1698431365
transform 1 0 13776 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1936_
timestamp 1698431365
transform 1 0 14112 0 -1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1937_
timestamp 1698431365
transform 1 0 15456 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1938_
timestamp 1698431365
transform 1 0 15120 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1939_
timestamp 1698431365
transform 1 0 14224 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1940_
timestamp 1698431365
transform 1 0 14896 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1941_
timestamp 1698431365
transform -1 0 16576 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1942_
timestamp 1698431365
transform 1 0 9856 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1943_
timestamp 1698431365
transform 1 0 12544 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1944_
timestamp 1698431365
transform 1 0 4256 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1945_
timestamp 1698431365
transform 1 0 11312 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1946_
timestamp 1698431365
transform 1 0 10752 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1947_
timestamp 1698431365
transform 1 0 13216 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1948_
timestamp 1698431365
transform 1 0 13328 0 1 17248
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1949_
timestamp 1698431365
transform 1 0 14448 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1950_
timestamp 1698431365
transform -1 0 14112 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1951_
timestamp 1698431365
transform 1 0 14112 0 1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1952_
timestamp 1698431365
transform -1 0 15344 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1953_
timestamp 1698431365
transform -1 0 14784 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1954_
timestamp 1698431365
transform 1 0 10192 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1955_
timestamp 1698431365
transform -1 0 11760 0 -1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1956_
timestamp 1698431365
transform 1 0 5600 0 1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1957_
timestamp 1698431365
transform 1 0 9968 0 -1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1958_
timestamp 1698431365
transform 1 0 10864 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1959_
timestamp 1698431365
transform 1 0 11424 0 1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1960_
timestamp 1698431365
transform 1 0 10192 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1961_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11424 0 -1 23520
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1962_
timestamp 1698431365
transform 1 0 2016 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1963_
timestamp 1698431365
transform 1 0 3584 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1964_
timestamp 1698431365
transform 1 0 4480 0 1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1965_
timestamp 1698431365
transform -1 0 5264 0 1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1966_
timestamp 1698431365
transform 1 0 8176 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1967_
timestamp 1698431365
transform -1 0 8624 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1968_
timestamp 1698431365
transform 1 0 2464 0 -1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1969_
timestamp 1698431365
transform -1 0 5376 0 -1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1970_
timestamp 1698431365
transform 1 0 5488 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1971_
timestamp 1698431365
transform 1 0 8400 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1972_
timestamp 1698431365
transform -1 0 12544 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1973_
timestamp 1698431365
transform -1 0 10192 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1974_
timestamp 1698431365
transform -1 0 9184 0 -1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1975_
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1976_
timestamp 1698431365
transform -1 0 10640 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1977_
timestamp 1698431365
transform 1 0 9072 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1978_
timestamp 1698431365
transform -1 0 10304 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1979_
timestamp 1698431365
transform -1 0 9296 0 1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1980_
timestamp 1698431365
transform 1 0 5712 0 1 21952
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1981_
timestamp 1698431365
transform 1 0 7392 0 1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1982_
timestamp 1698431365
transform 1 0 13552 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1983_
timestamp 1698431365
transform -1 0 14784 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1984_
timestamp 1698431365
transform -1 0 11648 0 1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1985_
timestamp 1698431365
transform 1 0 10528 0 -1 10976
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1986_
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1987_
timestamp 1698431365
transform 1 0 4928 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1988_
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1989_
timestamp 1698431365
transform 1 0 5824 0 1 9408
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1990_
timestamp 1698431365
transform 1 0 7616 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1991_
timestamp 1698431365
transform 1 0 4256 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1992_
timestamp 1698431365
transform 1 0 5152 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1993_
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1994_
timestamp 1698431365
transform 1 0 7728 0 1 7840
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1995_
timestamp 1698431365
transform 1 0 11536 0 -1 9408
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1996_
timestamp 1698431365
transform 1 0 13552 0 1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1997_
timestamp 1698431365
transform 1 0 14112 0 -1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1998_
timestamp 1698431365
transform -1 0 15904 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1999_
timestamp 1698431365
transform 1 0 15008 0 -1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2000_
timestamp 1698431365
transform 1 0 24304 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2001_
timestamp 1698431365
transform 1 0 15792 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2002_
timestamp 1698431365
transform 1 0 18256 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2003_
timestamp 1698431365
transform 1 0 29568 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2004_
timestamp 1698431365
transform -1 0 27328 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2005_
timestamp 1698431365
transform -1 0 27552 0 -1 25088
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2006_
timestamp 1698431365
transform 1 0 29008 0 1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2007_
timestamp 1698431365
transform -1 0 30464 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2008_
timestamp 1698431365
transform 1 0 30464 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2009_
timestamp 1698431365
transform 1 0 38752 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2010_
timestamp 1698431365
transform 1 0 38752 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2011_
timestamp 1698431365
transform 1 0 40768 0 -1 25088
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2012_
timestamp 1698431365
transform 1 0 45472 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2013_
timestamp 1698431365
transform -1 0 29904 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2014_
timestamp 1698431365
transform -1 0 29904 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2015_
timestamp 1698431365
transform -1 0 8400 0 -1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2016_
timestamp 1698431365
transform 1 0 6272 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2017_
timestamp 1698431365
transform 1 0 8288 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2018_
timestamp 1698431365
transform -1 0 9184 0 -1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2019_
timestamp 1698431365
transform -1 0 12432 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2020_
timestamp 1698431365
transform 1 0 9744 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2021_
timestamp 1698431365
transform 1 0 11536 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2022_
timestamp 1698431365
transform -1 0 12208 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2023_
timestamp 1698431365
transform -1 0 11648 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2024_
timestamp 1698431365
transform 1 0 10304 0 1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2025_
timestamp 1698431365
transform 1 0 10416 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2026_
timestamp 1698431365
transform -1 0 12880 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2027_
timestamp 1698431365
transform 1 0 9408 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2028_
timestamp 1698431365
transform 1 0 9296 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2029_
timestamp 1698431365
transform 1 0 10304 0 -1 20384
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_2  _2030_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11984 0 -1 21952
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2031_
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2032_
timestamp 1698431365
transform 1 0 14784 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _2033_
timestamp 1698431365
transform 1 0 13440 0 1 9408
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2034_
timestamp 1698431365
transform 1 0 17472 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2035_
timestamp 1698431365
transform -1 0 7728 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2036_
timestamp 1698431365
transform -1 0 14224 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2037_
timestamp 1698431365
transform 1 0 7840 0 -1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2038_
timestamp 1698431365
transform 1 0 10080 0 -1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2039_
timestamp 1698431365
transform -1 0 12432 0 1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _2040_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 14336 0 -1 7840
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2041_
timestamp 1698431365
transform 1 0 14448 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2042_
timestamp 1698431365
transform 1 0 5264 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2043_
timestamp 1698431365
transform 1 0 14560 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2044_
timestamp 1698431365
transform 1 0 3248 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2045_
timestamp 1698431365
transform -1 0 3808 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_2  _2046_
timestamp 1698431365
transform 1 0 3024 0 -1 12544
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2047_
timestamp 1698431365
transform 1 0 15120 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2048_
timestamp 1698431365
transform 1 0 18032 0 1 9408
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_2  _2049_
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2050_
timestamp 1698431365
transform -1 0 14560 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _2051_
timestamp 1698431365
transform 1 0 14560 0 1 23520
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2052_
timestamp 1698431365
transform 1 0 20272 0 -1 21952
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2053_
timestamp 1698431365
transform 1 0 17808 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2054_
timestamp 1698431365
transform -1 0 17920 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2055_
timestamp 1698431365
transform 1 0 17920 0 1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2056_
timestamp 1698431365
transform -1 0 28560 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2057_
timestamp 1698431365
transform -1 0 28784 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _2058_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 28448 0 1 23520
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2059_
timestamp 1698431365
transform -1 0 40544 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2060_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 39984 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2061_
timestamp 1698431365
transform -1 0 42896 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2062_
timestamp 1698431365
transform -1 0 42560 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2063_
timestamp 1698431365
transform 1 0 30352 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2064_
timestamp 1698431365
transform 1 0 10864 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2065_
timestamp 1698431365
transform -1 0 10528 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _2066_
timestamp 1698431365
transform 1 0 10528 0 1 20384
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _2067_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19376 0 1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2068_
timestamp 1698431365
transform -1 0 19712 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2069_
timestamp 1698431365
transform 1 0 10192 0 1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2070_
timestamp 1698431365
transform -1 0 22512 0 1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _2071_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 20720 0 -1 20384
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2072_
timestamp 1698431365
transform 1 0 18368 0 1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2073_
timestamp 1698431365
transform 1 0 19712 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2074_
timestamp 1698431365
transform 1 0 20720 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2075_
timestamp 1698431365
transform 1 0 21840 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2076_
timestamp 1698431365
transform 1 0 19040 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2077_
timestamp 1698431365
transform 1 0 20608 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2078_
timestamp 1698431365
transform -1 0 16464 0 -1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2079_
timestamp 1698431365
transform 1 0 14336 0 -1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2080_
timestamp 1698431365
transform -1 0 17024 0 -1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2081_
timestamp 1698431365
transform -1 0 20496 0 -1 9408
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2082_
timestamp 1698431365
transform 1 0 14560 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2083_
timestamp 1698431365
transform -1 0 18480 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2084_
timestamp 1698431365
transform 1 0 4480 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2085_
timestamp 1698431365
transform 1 0 16016 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2086_
timestamp 1698431365
transform 1 0 6720 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2087_
timestamp 1698431365
transform 1 0 11984 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2088_
timestamp 1698431365
transform 1 0 12432 0 -1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2089_
timestamp 1698431365
transform 1 0 17472 0 -1 10976
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2090_
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_2  _2091_
timestamp 1698431365
transform 1 0 21952 0 -1 10976
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2092_
timestamp 1698431365
transform 1 0 21392 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2093_
timestamp 1698431365
transform 1 0 21280 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2094_
timestamp 1698431365
transform 1 0 22400 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2095_
timestamp 1698431365
transform 1 0 22400 0 1 21952
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2096_
timestamp 1698431365
transform 1 0 16688 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2097_
timestamp 1698431365
transform 1 0 17248 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2098_
timestamp 1698431365
transform 1 0 18928 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2099_
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _2100_
timestamp 1698431365
transform -1 0 30128 0 -1 25088
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2101_
timestamp 1698431365
transform -1 0 38864 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2102_
timestamp 1698431365
transform -1 0 47152 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2103_
timestamp 1698431365
transform 1 0 47152 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2104_
timestamp 1698431365
transform -1 0 20720 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2105_
timestamp 1698431365
transform -1 0 21728 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2106_
timestamp 1698431365
transform 1 0 19712 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2107_
timestamp 1698431365
transform 1 0 21616 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2108_
timestamp 1698431365
transform 1 0 21168 0 -1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2109_
timestamp 1698431365
transform -1 0 22848 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2110_
timestamp 1698431365
transform 1 0 23072 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2111_
timestamp 1698431365
transform 1 0 22960 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2112_
timestamp 1698431365
transform -1 0 20272 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2113_
timestamp 1698431365
transform 1 0 16128 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2114_
timestamp 1698431365
transform 1 0 15232 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2115_
timestamp 1698431365
transform 1 0 15344 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2116_
timestamp 1698431365
transform -1 0 17920 0 1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2117_
timestamp 1698431365
transform -1 0 19040 0 -1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _2118_
timestamp 1698431365
transform -1 0 20944 0 1 10976
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2119_
timestamp 1698431365
transform 1 0 15344 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2120_
timestamp 1698431365
transform 1 0 13776 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2121_
timestamp 1698431365
transform 1 0 15120 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2122_
timestamp 1698431365
transform 1 0 12544 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2123_
timestamp 1698431365
transform 1 0 12544 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _2124_
timestamp 1698431365
transform 1 0 12880 0 -1 15680
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2125_
timestamp 1698431365
transform 1 0 15344 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2126_
timestamp 1698431365
transform 1 0 18368 0 1 12544
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2127_
timestamp 1698431365
transform -1 0 24304 0 1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2128_
timestamp 1698431365
transform -1 0 23520 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _2129_
timestamp 1698431365
transform -1 0 26544 0 1 20384
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2130_
timestamp 1698431365
transform 1 0 25648 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2131_
timestamp 1698431365
transform 1 0 23072 0 1 18816
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2132_
timestamp 1698431365
transform 1 0 18368 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2133_
timestamp 1698431365
transform 1 0 16464 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2134_
timestamp 1698431365
transform -1 0 17808 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2135_
timestamp 1698431365
transform 1 0 17696 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2136_
timestamp 1698431365
transform 1 0 16464 0 1 18816
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2137_
timestamp 1698431365
transform -1 0 20496 0 1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2138_
timestamp 1698431365
transform 1 0 19040 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2139_
timestamp 1698431365
transform 1 0 30240 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _2140_
timestamp 1698431365
transform -1 0 28784 0 1 21952
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2141_
timestamp 1698431365
transform -1 0 42000 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2142_
timestamp 1698431365
transform -1 0 44464 0 1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2143_
timestamp 1698431365
transform 1 0 45360 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2144_
timestamp 1698431365
transform -1 0 39984 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2145_
timestamp 1698431365
transform 1 0 38304 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2146_
timestamp 1698431365
transform -1 0 42896 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2147_
timestamp 1698431365
transform -1 0 30576 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2148_
timestamp 1698431365
transform 1 0 31136 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2149_
timestamp 1698431365
transform 1 0 23408 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2150_
timestamp 1698431365
transform -1 0 23072 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2151_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22736 0 -1 20384
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2152_
timestamp 1698431365
transform 1 0 18816 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2153_
timestamp 1698431365
transform 1 0 20160 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2154_
timestamp 1698431365
transform 1 0 23072 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2155_
timestamp 1698431365
transform 1 0 24528 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2156_
timestamp 1698431365
transform 1 0 21280 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2157_
timestamp 1698431365
transform 1 0 15456 0 1 12544
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2158_
timestamp 1698431365
transform 1 0 14224 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2159_
timestamp 1698431365
transform -1 0 17024 0 -1 14112
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2160_
timestamp 1698431365
transform -1 0 21280 0 -1 14112
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2161_
timestamp 1698431365
transform -1 0 19040 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2162_
timestamp 1698431365
transform -1 0 18032 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2163_
timestamp 1698431365
transform 1 0 13664 0 1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2164_
timestamp 1698431365
transform 1 0 15904 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2165_
timestamp 1698431365
transform 1 0 18816 0 -1 15680
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2166_
timestamp 1698431365
transform 1 0 21840 0 1 14112
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2167_
timestamp 1698431365
transform 1 0 25088 0 1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2168_
timestamp 1698431365
transform 1 0 26320 0 -1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2169_
timestamp 1698431365
transform 1 0 15456 0 1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2170_
timestamp 1698431365
transform 1 0 28112 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2171_
timestamp 1698431365
transform -1 0 31136 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2172_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 28784 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2173_
timestamp 1698431365
transform -1 0 42112 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2174_
timestamp 1698431365
transform -1 0 41776 0 1 25088
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2175_
timestamp 1698431365
transform 1 0 41776 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2176_
timestamp 1698431365
transform -1 0 35728 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2177_
timestamp 1698431365
transform -1 0 32928 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2178_
timestamp 1698431365
transform -1 0 28784 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2179_
timestamp 1698431365
transform 1 0 21952 0 -1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2180_
timestamp 1698431365
transform -1 0 24192 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2181_
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2182_
timestamp 1698431365
transform 1 0 25648 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2183_
timestamp 1698431365
transform 1 0 22288 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2184_
timestamp 1698431365
transform -1 0 22960 0 -1 18816
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2185_
timestamp 1698431365
transform 1 0 20832 0 -1 17248
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2186_
timestamp 1698431365
transform -1 0 17920 0 1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2187_
timestamp 1698431365
transform 1 0 15904 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2188_
timestamp 1698431365
transform -1 0 18816 0 -1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2189_
timestamp 1698431365
transform 1 0 18144 0 -1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _2190_
timestamp 1698431365
transform -1 0 20944 0 1 15680
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2191_
timestamp 1698431365
transform 1 0 23296 0 1 15680
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2192_
timestamp 1698431365
transform 1 0 25872 0 1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2193_
timestamp 1698431365
transform 1 0 26432 0 -1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2194_
timestamp 1698431365
transform 1 0 14784 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2195_
timestamp 1698431365
transform 1 0 15344 0 -1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2196_
timestamp 1698431365
transform 1 0 18368 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2197_
timestamp 1698431365
transform 1 0 30576 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2198_
timestamp 1698431365
transform -1 0 33824 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _2199_
timestamp 1698431365
transform 1 0 30128 0 -1 25088
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2200_
timestamp 1698431365
transform -1 0 38640 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2201_
timestamp 1698431365
transform -1 0 38304 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2202_
timestamp 1698431365
transform 1 0 38080 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2203_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 36848 0 1 21952
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2204_
timestamp 1698431365
transform -1 0 28224 0 1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2205_
timestamp 1698431365
transform 1 0 23520 0 -1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2206_
timestamp 1698431365
transform 1 0 24192 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2207_
timestamp 1698431365
transform 1 0 25536 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2208_
timestamp 1698431365
transform 1 0 26320 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _2209_
timestamp 1698431365
transform -1 0 25648 0 1 17248
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2210_
timestamp 1698431365
transform 1 0 26768 0 1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2211_
timestamp 1698431365
transform 1 0 28560 0 -1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2212_
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _2213_
timestamp 1698431365
transform 1 0 31024 0 1 23520
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2214_
timestamp 1698431365
transform 1 0 35056 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2215_
timestamp 1698431365
transform -1 0 36176 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2216_
timestamp 1698431365
transform -1 0 36288 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2217_
timestamp 1698431365
transform -1 0 34272 0 1 20384
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2218_
timestamp 1698431365
transform 1 0 26320 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2219_
timestamp 1698431365
transform 1 0 27776 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2220_
timestamp 1698431365
transform -1 0 30128 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2221_
timestamp 1698431365
transform 1 0 11424 0 -1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2222_
timestamp 1698431365
transform 1 0 24976 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2223_
timestamp 1698431365
transform 1 0 34272 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2224_
timestamp 1698431365
transform 1 0 32928 0 -1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2225_
timestamp 1698431365
transform -1 0 32256 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2226_
timestamp 1698431365
transform -1 0 18144 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2227_
timestamp 1698431365
transform -1 0 19376 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2228_
timestamp 1698431365
transform 1 0 19040 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2229_
timestamp 1698431365
transform 1 0 9408 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2230_
timestamp 1698431365
transform 1 0 9744 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _2231_
timestamp 1698431365
transform 1 0 13664 0 -1 45472
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _2232_
timestamp 1698431365
transform 1 0 12992 0 1 45472
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2233_
timestamp 1698431365
transform 1 0 18816 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2234_
timestamp 1698431365
transform -1 0 14000 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2235_
timestamp 1698431365
transform -1 0 12432 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2236_
timestamp 1698431365
transform 1 0 8736 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2237_
timestamp 1698431365
transform 1 0 10416 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2238_
timestamp 1698431365
transform 1 0 8624 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2239_
timestamp 1698431365
transform 1 0 9856 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2240_
timestamp 1698431365
transform 1 0 9744 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2241_
timestamp 1698431365
transform 1 0 10752 0 1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2242_
timestamp 1698431365
transform 1 0 20384 0 -1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2243_
timestamp 1698431365
transform 1 0 21168 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2244_
timestamp 1698431365
transform 1 0 22288 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2245_
timestamp 1698431365
transform 1 0 17360 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2246_
timestamp 1698431365
transform 1 0 21952 0 1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2247_
timestamp 1698431365
transform 1 0 16352 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2248_
timestamp 1698431365
transform -1 0 16576 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2249_
timestamp 1698431365
transform 1 0 7504 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _2250_
timestamp 1698431365
transform 1 0 9408 0 1 43904
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _2251_
timestamp 1698431365
transform 1 0 10080 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2252_
timestamp 1698431365
transform -1 0 15904 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2253_
timestamp 1698431365
transform 1 0 17248 0 -1 45472
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2254_
timestamp 1698431365
transform 1 0 21504 0 -1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2255_
timestamp 1698431365
transform 1 0 22736 0 1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2256_
timestamp 1698431365
transform 1 0 3584 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2257_
timestamp 1698431365
transform 1 0 5600 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2258_
timestamp 1698431365
transform 1 0 4592 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2259_
timestamp 1698431365
transform 1 0 6160 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2260_
timestamp 1698431365
transform -1 0 6720 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2261_
timestamp 1698431365
transform 1 0 5712 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2262_
timestamp 1698431365
transform 1 0 7168 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2263_
timestamp 1698431365
transform -1 0 6160 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2264_
timestamp 1698431365
transform 1 0 5600 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2265_
timestamp 1698431365
transform -1 0 8176 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2266_
timestamp 1698431365
transform 1 0 5824 0 1 37632
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2267_
timestamp 1698431365
transform -1 0 7392 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2268_
timestamp 1698431365
transform -1 0 11984 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2269_
timestamp 1698431365
transform 1 0 11760 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2270_
timestamp 1698431365
transform -1 0 9968 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2271_
timestamp 1698431365
transform -1 0 8960 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2272_
timestamp 1698431365
transform -1 0 8512 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2273_
timestamp 1698431365
transform -1 0 7616 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2274_
timestamp 1698431365
transform -1 0 5712 0 -1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2275_
timestamp 1698431365
transform -1 0 4704 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _2276_
timestamp 1698431365
transform 1 0 3472 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2277_
timestamp 1698431365
transform 1 0 5488 0 1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2278_
timestamp 1698431365
transform -1 0 7504 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2279_
timestamp 1698431365
transform -1 0 3808 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2280_
timestamp 1698431365
transform -1 0 4704 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2281_
timestamp 1698431365
transform 1 0 1568 0 1 40768
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2282_
timestamp 1698431365
transform 1 0 2800 0 1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2283_
timestamp 1698431365
transform 1 0 6944 0 -1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2284_
timestamp 1698431365
transform 1 0 9408 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2285_
timestamp 1698431365
transform 1 0 8288 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2286_
timestamp 1698431365
transform -1 0 9072 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2287_
timestamp 1698431365
transform 1 0 7952 0 1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2288_
timestamp 1698431365
transform 1 0 6608 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2289_
timestamp 1698431365
transform -1 0 6832 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2290_
timestamp 1698431365
transform -1 0 7616 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2291_
timestamp 1698431365
transform -1 0 3248 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2292_
timestamp 1698431365
transform 1 0 4592 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2293_
timestamp 1698431365
transform -1 0 3248 0 -1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2294_
timestamp 1698431365
transform 1 0 2016 0 1 37632
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2295_
timestamp 1698431365
transform 1 0 4480 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2296_
timestamp 1698431365
transform -1 0 3024 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2297_
timestamp 1698431365
transform -1 0 3248 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2298_
timestamp 1698431365
transform 1 0 5712 0 -1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2299_
timestamp 1698431365
transform 1 0 6720 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2300_
timestamp 1698431365
transform -1 0 7168 0 1 32928
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2301_
timestamp 1698431365
transform 1 0 1568 0 -1 32928
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2302_
timestamp 1698431365
transform 1 0 1792 0 -1 36064
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2303_
timestamp 1698431365
transform 1 0 3808 0 1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2304_
timestamp 1698431365
transform 1 0 22288 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2305_
timestamp 1698431365
transform 1 0 23184 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2306_
timestamp 1698431365
transform 1 0 22848 0 -1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2307_
timestamp 1698431365
transform 1 0 8064 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2308_
timestamp 1698431365
transform 1 0 24752 0 1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2309_
timestamp 1698431365
transform 1 0 8400 0 1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2310_
timestamp 1698431365
transform 1 0 10864 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2311_
timestamp 1698431365
transform -1 0 10864 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2312_
timestamp 1698431365
transform 1 0 16352 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _2313_
timestamp 1698431365
transform -1 0 17920 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2314_
timestamp 1698431365
transform 1 0 25088 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2315_
timestamp 1698431365
transform 1 0 24640 0 1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2316_
timestamp 1698431365
transform 1 0 5936 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2317_
timestamp 1698431365
transform 1 0 10080 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2318_
timestamp 1698431365
transform -1 0 9968 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2319_
timestamp 1698431365
transform 1 0 9856 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2320_
timestamp 1698431365
transform -1 0 10416 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2321_
timestamp 1698431365
transform 1 0 10416 0 1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2322_
timestamp 1698431365
transform 1 0 9968 0 -1 37632
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2323_
timestamp 1698431365
transform 1 0 19824 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2324_
timestamp 1698431365
transform 1 0 23184 0 -1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2325_
timestamp 1698431365
transform 1 0 23744 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2326_
timestamp 1698431365
transform 1 0 25088 0 -1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2327_
timestamp 1698431365
transform 1 0 24304 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2328_
timestamp 1698431365
transform 1 0 25312 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2329_
timestamp 1698431365
transform -1 0 23744 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2330_
timestamp 1698431365
transform 1 0 22960 0 1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2331_
timestamp 1698431365
transform 1 0 2576 0 -1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2332_
timestamp 1698431365
transform -1 0 4592 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2333_
timestamp 1698431365
transform 1 0 1680 0 1 32928
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2334_
timestamp 1698431365
transform -1 0 4704 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2335_
timestamp 1698431365
transform -1 0 3472 0 1 34496
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2336_
timestamp 1698431365
transform 1 0 4368 0 -1 36064
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2337_
timestamp 1698431365
transform -1 0 5600 0 -1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2338_
timestamp 1698431365
transform 1 0 6720 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2339_
timestamp 1698431365
transform -1 0 5264 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2340_
timestamp 1698431365
transform 1 0 4144 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2341_
timestamp 1698431365
transform 1 0 2576 0 1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2342_
timestamp 1698431365
transform 1 0 3920 0 1 31360
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2343_
timestamp 1698431365
transform -1 0 3024 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2344_
timestamp 1698431365
transform -1 0 8848 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2345_
timestamp 1698431365
transform -1 0 9184 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2346_
timestamp 1698431365
transform -1 0 7392 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2347_
timestamp 1698431365
transform 1 0 7168 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2348_
timestamp 1698431365
transform 1 0 6048 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2349_
timestamp 1698431365
transform -1 0 7392 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2350_
timestamp 1698431365
transform 1 0 7616 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2351_
timestamp 1698431365
transform 1 0 6720 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2352_
timestamp 1698431365
transform -1 0 6720 0 -1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2353_
timestamp 1698431365
transform 1 0 1568 0 1 29792
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2354_
timestamp 1698431365
transform 1 0 3808 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2355_
timestamp 1698431365
transform -1 0 23184 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2356_
timestamp 1698431365
transform -1 0 20160 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2357_
timestamp 1698431365
transform -1 0 15568 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2358_
timestamp 1698431365
transform 1 0 21168 0 -1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _2359_
timestamp 1698431365
transform 1 0 19824 0 -1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2360_
timestamp 1698431365
transform -1 0 21504 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2361_
timestamp 1698431365
transform 1 0 19488 0 1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2362_
timestamp 1698431365
transform -1 0 17248 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2363_
timestamp 1698431365
transform 1 0 13440 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2364_
timestamp 1698431365
transform -1 0 7392 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2365_
timestamp 1698431365
transform -1 0 7840 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2366_
timestamp 1698431365
transform 1 0 7392 0 -1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _2367_
timestamp 1698431365
transform -1 0 13664 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _2368_
timestamp 1698431365
transform 1 0 10416 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2369_
timestamp 1698431365
transform 1 0 11200 0 1 43904
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2370_
timestamp 1698431365
transform 1 0 15120 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2371_
timestamp 1698431365
transform 1 0 13888 0 -1 43904
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2372_
timestamp 1698431365
transform 1 0 18256 0 -1 42336
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2373_
timestamp 1698431365
transform -1 0 23184 0 -1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2374_
timestamp 1698431365
transform -1 0 22176 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2375_
timestamp 1698431365
transform -1 0 21952 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2376_
timestamp 1698431365
transform -1 0 21840 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2377_
timestamp 1698431365
transform 1 0 21840 0 -1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2378_
timestamp 1698431365
transform 1 0 10192 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2379_
timestamp 1698431365
transform -1 0 17024 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2380_
timestamp 1698431365
transform 1 0 16128 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _2381_
timestamp 1698431365
transform -1 0 32704 0 -1 26656
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2382_
timestamp 1698431365
transform 1 0 25536 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2383_
timestamp 1698431365
transform -1 0 31360 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2384_
timestamp 1698431365
transform -1 0 30800 0 1 20384
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2385_
timestamp 1698431365
transform -1 0 13888 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2386_
timestamp 1698431365
transform -1 0 29120 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2387_
timestamp 1698431365
transform -1 0 20944 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2388_
timestamp 1698431365
transform -1 0 4144 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2389_
timestamp 1698431365
transform 1 0 2912 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2390_
timestamp 1698431365
transform 1 0 4144 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2391_
timestamp 1698431365
transform -1 0 5488 0 -1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2392_
timestamp 1698431365
transform -1 0 8176 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2393_
timestamp 1698431365
transform -1 0 9856 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2394_
timestamp 1698431365
transform 1 0 5936 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2395_
timestamp 1698431365
transform 1 0 9520 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2396_
timestamp 1698431365
transform -1 0 9968 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2397_
timestamp 1698431365
transform -1 0 8848 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2398_
timestamp 1698431365
transform 1 0 7504 0 -1 31360
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2399_
timestamp 1698431365
transform -1 0 7392 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2400_
timestamp 1698431365
transform 1 0 5712 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2401_
timestamp 1698431365
transform 1 0 6048 0 1 28224
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2402_
timestamp 1698431365
transform 1 0 7728 0 -1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2403_
timestamp 1698431365
transform 1 0 17472 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2404_
timestamp 1698431365
transform 1 0 18480 0 1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2405_
timestamp 1698431365
transform 1 0 18480 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2406_
timestamp 1698431365
transform 1 0 23184 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2407_
timestamp 1698431365
transform 1 0 19376 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2408_
timestamp 1698431365
transform -1 0 13664 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2409_
timestamp 1698431365
transform 1 0 12208 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2410_
timestamp 1698431365
transform 1 0 14672 0 1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2411_
timestamp 1698431365
transform 1 0 15904 0 1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2412_
timestamp 1698431365
transform -1 0 17248 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _2413_
timestamp 1698431365
transform 1 0 15232 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2414_
timestamp 1698431365
transform 1 0 17360 0 1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2415_
timestamp 1698431365
transform -1 0 13104 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _2416_
timestamp 1698431365
transform 1 0 8624 0 1 40768
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2417_
timestamp 1698431365
transform 1 0 9408 0 -1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2418_
timestamp 1698431365
transform 1 0 9968 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2419_
timestamp 1698431365
transform 1 0 7840 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2420_
timestamp 1698431365
transform 1 0 14336 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2421_
timestamp 1698431365
transform 1 0 13328 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2422_
timestamp 1698431365
transform 1 0 20720 0 -1 40768
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2423_
timestamp 1698431365
transform 1 0 22288 0 1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2424_
timestamp 1698431365
transform 1 0 22176 0 -1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2425_
timestamp 1698431365
transform 1 0 23296 0 -1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2426_
timestamp 1698431365
transform 1 0 14560 0 -1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2427_
timestamp 1698431365
transform 1 0 21392 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2428_
timestamp 1698431365
transform -1 0 21168 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2429_
timestamp 1698431365
transform 1 0 18592 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2430_
timestamp 1698431365
transform -1 0 18592 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2431_
timestamp 1698431365
transform 1 0 10752 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2432_
timestamp 1698431365
transform 1 0 15456 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2433_
timestamp 1698431365
transform 1 0 17248 0 -1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2434_
timestamp 1698431365
transform 1 0 16240 0 -1 29792
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2435_
timestamp 1698431365
transform 1 0 17920 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2436_
timestamp 1698431365
transform -1 0 17920 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2437_
timestamp 1698431365
transform -1 0 20048 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_2  _2438_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17584 0 -1 26656
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2439_
timestamp 1698431365
transform -1 0 12544 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2440_
timestamp 1698431365
transform -1 0 12432 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2441_
timestamp 1698431365
transform -1 0 9296 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2442_
timestamp 1698431365
transform 1 0 6720 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _2443_
timestamp 1698431365
transform 1 0 6608 0 -1 29792
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2444_
timestamp 1698431365
transform 1 0 10304 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2445_
timestamp 1698431365
transform -1 0 11984 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2446_
timestamp 1698431365
transform 1 0 7840 0 1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2447_
timestamp 1698431365
transform 1 0 9632 0 1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2448_
timestamp 1698431365
transform 1 0 10080 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2449_
timestamp 1698431365
transform 1 0 21168 0 1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2450_
timestamp 1698431365
transform -1 0 23856 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2451_
timestamp 1698431365
transform 1 0 21728 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2452_
timestamp 1698431365
transform -1 0 18480 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2453_
timestamp 1698431365
transform -1 0 14336 0 -1 42336
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2454_
timestamp 1698431365
transform 1 0 12880 0 -1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2455_
timestamp 1698431365
transform 1 0 14000 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2456_
timestamp 1698431365
transform 1 0 17248 0 -1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2457_
timestamp 1698431365
transform -1 0 14224 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _2458_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 13104 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2459_
timestamp 1698431365
transform -1 0 12880 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2460_
timestamp 1698431365
transform 1 0 10416 0 -1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2461_
timestamp 1698431365
transform 1 0 11760 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2462_
timestamp 1698431365
transform 1 0 14224 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2463_
timestamp 1698431365
transform 1 0 13664 0 -1 39200
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2464_
timestamp 1698431365
transform 1 0 18144 0 -1 39200
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2465_
timestamp 1698431365
transform -1 0 23072 0 1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2466_
timestamp 1698431365
transform -1 0 14784 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2467_
timestamp 1698431365
transform -1 0 20944 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2468_
timestamp 1698431365
transform 1 0 22176 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2469_
timestamp 1698431365
transform -1 0 15456 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2470_
timestamp 1698431365
transform -1 0 15456 0 1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2471_
timestamp 1698431365
transform 1 0 11760 0 -1 28224
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2472_
timestamp 1698431365
transform 1 0 16128 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2473_
timestamp 1698431365
transform -1 0 15232 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2474_
timestamp 1698431365
transform 1 0 13328 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2475_
timestamp 1698431365
transform 1 0 14112 0 -1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2476_
timestamp 1698431365
transform -1 0 17360 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2477_
timestamp 1698431365
transform 1 0 17360 0 1 29792
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2478_
timestamp 1698431365
transform -1 0 16240 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2479_
timestamp 1698431365
transform 1 0 17248 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_2  _2480_
timestamp 1698431365
transform 1 0 16912 0 1 25088
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2481_
timestamp 1698431365
transform -1 0 12992 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2482_
timestamp 1698431365
transform -1 0 16576 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2483_
timestamp 1698431365
transform 1 0 11872 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2484_
timestamp 1698431365
transform -1 0 13104 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2485_
timestamp 1698431365
transform -1 0 14784 0 1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2486_
timestamp 1698431365
transform 1 0 10192 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2487_
timestamp 1698431365
transform -1 0 11760 0 -1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2488_
timestamp 1698431365
transform 1 0 18256 0 1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2489_
timestamp 1698431365
transform 1 0 18928 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2490_
timestamp 1698431365
transform 1 0 20720 0 -1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2491_
timestamp 1698431365
transform 1 0 17808 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2492_
timestamp 1698431365
transform 1 0 16128 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2493_
timestamp 1698431365
transform -1 0 13664 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2494_
timestamp 1698431365
transform 1 0 13328 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2495_
timestamp 1698431365
transform 1 0 14000 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2496_
timestamp 1698431365
transform 1 0 15904 0 -1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _2497_
timestamp 1698431365
transform -1 0 19040 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2498_
timestamp 1698431365
transform 1 0 17248 0 -1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2499_
timestamp 1698431365
transform -1 0 14560 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2500_
timestamp 1698431365
transform -1 0 14784 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2501_
timestamp 1698431365
transform -1 0 10080 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2502_
timestamp 1698431365
transform -1 0 10080 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2503_
timestamp 1698431365
transform 1 0 10416 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2504_
timestamp 1698431365
transform 1 0 13440 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2505_
timestamp 1698431365
transform 1 0 18368 0 1 36064
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2506_
timestamp 1698431365
transform 1 0 21280 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2507_
timestamp 1698431365
transform 1 0 21168 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2508_
timestamp 1698431365
transform -1 0 22848 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2509_
timestamp 1698431365
transform -1 0 20496 0 1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2510_
timestamp 1698431365
transform 1 0 19152 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2511_
timestamp 1698431365
transform 1 0 18256 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2512_
timestamp 1698431365
transform -1 0 11424 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2513_
timestamp 1698431365
transform -1 0 12320 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2514_
timestamp 1698431365
transform 1 0 10304 0 1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2515_
timestamp 1698431365
transform -1 0 12656 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2516_
timestamp 1698431365
transform 1 0 12544 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2517_
timestamp 1698431365
transform 1 0 12656 0 -1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2518_
timestamp 1698431365
transform -1 0 30128 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2519_
timestamp 1698431365
transform 1 0 13888 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2520_
timestamp 1698431365
transform 1 0 13776 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2521_
timestamp 1698431365
transform 1 0 16912 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_2  _2522_
timestamp 1698431365
transform 1 0 17472 0 1 26656
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2523_
timestamp 1698431365
transform -1 0 15456 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2524_
timestamp 1698431365
transform 1 0 21280 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2525_
timestamp 1698431365
transform 1 0 19040 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2526_
timestamp 1698431365
transform 1 0 20384 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2527_
timestamp 1698431365
transform -1 0 22624 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2528_
timestamp 1698431365
transform 1 0 18704 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2529_
timestamp 1698431365
transform -1 0 14336 0 -1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2530_
timestamp 1698431365
transform 1 0 11984 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2531_
timestamp 1698431365
transform 1 0 14336 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2532_
timestamp 1698431365
transform 1 0 17248 0 1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2533_
timestamp 1698431365
transform -1 0 16912 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2534_
timestamp 1698431365
transform 1 0 11536 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2535_
timestamp 1698431365
transform -1 0 11536 0 -1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2536_
timestamp 1698431365
transform 1 0 14000 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2537_
timestamp 1698431365
transform 1 0 12880 0 -1 32928
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2538_
timestamp 1698431365
transform 1 0 18592 0 -1 34496
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2539_
timestamp 1698431365
transform 1 0 21504 0 1 32928
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2540_
timestamp 1698431365
transform 1 0 21840 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2541_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21952 0 1 29792
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2542_
timestamp 1698431365
transform -1 0 22848 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2543_
timestamp 1698431365
transform 1 0 21616 0 -1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2544_
timestamp 1698431365
transform 1 0 32032 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2545_
timestamp 1698431365
transform 1 0 22848 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2546_
timestamp 1698431365
transform -1 0 29680 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2547_
timestamp 1698431365
transform 1 0 23072 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2548_
timestamp 1698431365
transform 1 0 24192 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2549_
timestamp 1698431365
transform -1 0 32592 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2550_
timestamp 1698431365
transform 1 0 23968 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2551_
timestamp 1698431365
transform -1 0 28784 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2552_
timestamp 1698431365
transform 1 0 25088 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2553_
timestamp 1698431365
transform 1 0 23072 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2554_
timestamp 1698431365
transform -1 0 39312 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2555_
timestamp 1698431365
transform 1 0 22960 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2556_
timestamp 1698431365
transform 1 0 23408 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2557_
timestamp 1698431365
transform 1 0 13328 0 1 32928
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2558_
timestamp 1698431365
transform 1 0 17248 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2559_
timestamp 1698431365
transform -1 0 22064 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2560_
timestamp 1698431365
transform 1 0 19376 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2561_
timestamp 1698431365
transform 1 0 18368 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2562_
timestamp 1698431365
transform 1 0 15568 0 -1 32928
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2563_
timestamp 1698431365
transform 1 0 18816 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2564_
timestamp 1698431365
transform -1 0 14000 0 -1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _2565_
timestamp 1698431365
transform 1 0 16240 0 1 32928
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2566_
timestamp 1698431365
transform 1 0 17024 0 1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2567_
timestamp 1698431365
transform 1 0 19264 0 -1 31360
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2568_
timestamp 1698431365
transform 1 0 25088 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2569_
timestamp 1698431365
transform 1 0 24192 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2570_
timestamp 1698431365
transform 1 0 26432 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2571_
timestamp 1698431365
transform 1 0 25088 0 1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _2572_
timestamp 1698431365
transform -1 0 28336 0 1 29792
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2573_
timestamp 1698431365
transform -1 0 28672 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2574_
timestamp 1698431365
transform -1 0 29568 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2575_
timestamp 1698431365
transform -1 0 28000 0 1 20384
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2576_
timestamp 1698431365
transform 1 0 19152 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2577_
timestamp 1698431365
transform 1 0 19824 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2578_
timestamp 1698431365
transform 1 0 19824 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2579_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 -1 32928
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2580_
timestamp 1698431365
transform 1 0 23072 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2581_
timestamp 1698431365
transform 1 0 23520 0 -1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2582_
timestamp 1698431365
transform 1 0 25536 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2583_
timestamp 1698431365
transform 1 0 25872 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2584_
timestamp 1698431365
transform 1 0 26208 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2585_
timestamp 1698431365
transform 1 0 25984 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _2586_
timestamp 1698431365
transform -1 0 28224 0 -1 32928
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2587_
timestamp 1698431365
transform -1 0 25984 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2588_
timestamp 1698431365
transform -1 0 37968 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2589_
timestamp 1698431365
transform -1 0 27888 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2590_
timestamp 1698431365
transform 1 0 25648 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2591_
timestamp 1698431365
transform 1 0 23968 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2592_
timestamp 1698431365
transform 1 0 23184 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2593_
timestamp 1698431365
transform 1 0 25088 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2594_
timestamp 1698431365
transform 1 0 24864 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2595_
timestamp 1698431365
transform -1 0 25872 0 1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2596_
timestamp 1698431365
transform -1 0 24864 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2597_
timestamp 1698431365
transform -1 0 27552 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2598_
timestamp 1698431365
transform 1 0 25088 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2599_
timestamp 1698431365
transform -1 0 20832 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2600_
timestamp 1698431365
transform -1 0 44352 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2601_
timestamp 1698431365
transform 1 0 45024 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2602_
timestamp 1698431365
transform 1 0 46592 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2603_
timestamp 1698431365
transform 1 0 46144 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2604_
timestamp 1698431365
transform -1 0 44240 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2605_
timestamp 1698431365
transform 1 0 41104 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2606_
timestamp 1698431365
transform 1 0 42896 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2607_
timestamp 1698431365
transform 1 0 40208 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _2608_
timestamp 1698431365
transform -1 0 43680 0 -1 42336
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2609_
timestamp 1698431365
transform 1 0 41552 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2610_
timestamp 1698431365
transform 1 0 41776 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _2611_
timestamp 1698431365
transform 1 0 42560 0 -1 40768
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2612_
timestamp 1698431365
transform 1 0 43680 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2613_
timestamp 1698431365
transform 1 0 41888 0 1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2614_
timestamp 1698431365
transform -1 0 44464 0 1 40768
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2615_
timestamp 1698431365
transform 1 0 40768 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _2616_
timestamp 1698431365
transform 1 0 40880 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _2617_
timestamp 1698431365
transform 1 0 42224 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2618_
timestamp 1698431365
transform -1 0 45584 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2619_
timestamp 1698431365
transform -1 0 46368 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2620_
timestamp 1698431365
transform 1 0 44912 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2621_
timestamp 1698431365
transform 1 0 45808 0 -1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2622_
timestamp 1698431365
transform 1 0 44352 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2623_
timestamp 1698431365
transform 1 0 45808 0 -1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _2624_
timestamp 1698431365
transform 1 0 42000 0 1 45472
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2625_
timestamp 1698431365
transform 1 0 48608 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2626_
timestamp 1698431365
transform -1 0 41552 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _2627_
timestamp 1698431365
transform 1 0 41888 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2628_
timestamp 1698431365
transform 1 0 47488 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2629_
timestamp 1698431365
transform 1 0 45360 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2630_
timestamp 1698431365
transform -1 0 47824 0 1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2631_
timestamp 1698431365
transform 1 0 46928 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2632_
timestamp 1698431365
transform -1 0 43456 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2633_
timestamp 1698431365
transform 1 0 45696 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _2634_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 44352 0 -1 45472
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2635_
timestamp 1698431365
transform -1 0 47488 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  _2636_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 51184 0 1 42336
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2637_
timestamp 1698431365
transform 1 0 48608 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2638_
timestamp 1698431365
transform 1 0 51856 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2639_
timestamp 1698431365
transform 1 0 41216 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2640_
timestamp 1698431365
transform -1 0 40544 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2641_
timestamp 1698431365
transform -1 0 50848 0 1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2642_
timestamp 1698431365
transform -1 0 51856 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2643_
timestamp 1698431365
transform 1 0 47488 0 1 37632
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2644_
timestamp 1698431365
transform -1 0 49952 0 -1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2645_
timestamp 1698431365
transform -1 0 38192 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2646_
timestamp 1698431365
transform 1 0 40992 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2647_
timestamp 1698431365
transform -1 0 38304 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2648_
timestamp 1698431365
transform 1 0 35952 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2649_
timestamp 1698431365
transform -1 0 46480 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2650_
timestamp 1698431365
transform -1 0 39872 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2651_
timestamp 1698431365
transform 1 0 40656 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2652_
timestamp 1698431365
transform 1 0 39872 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2653_
timestamp 1698431365
transform 1 0 38192 0 1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2654_
timestamp 1698431365
transform 1 0 38976 0 1 37632
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2655_
timestamp 1698431365
transform -1 0 39984 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2656_
timestamp 1698431365
transform -1 0 40656 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2657_
timestamp 1698431365
transform -1 0 38976 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2658_
timestamp 1698431365
transform 1 0 37184 0 1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2659_
timestamp 1698431365
transform -1 0 37856 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _2660_
timestamp 1698431365
transform -1 0 39984 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2661_
timestamp 1698431365
transform -1 0 38864 0 -1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2662_
timestamp 1698431365
transform 1 0 36064 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2663_
timestamp 1698431365
transform -1 0 39984 0 -1 45472
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2664_
timestamp 1698431365
transform 1 0 37408 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2665_
timestamp 1698431365
transform -1 0 37632 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2666_
timestamp 1698431365
transform 1 0 40768 0 -1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2667_
timestamp 1698431365
transform 1 0 40096 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2668_
timestamp 1698431365
transform 1 0 40768 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2669_
timestamp 1698431365
transform -1 0 37520 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2670_
timestamp 1698431365
transform 1 0 39984 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2671_
timestamp 1698431365
transform 1 0 39984 0 1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2672_
timestamp 1698431365
transform 1 0 36288 0 -1 39200
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2673_
timestamp 1698431365
transform 1 0 38864 0 -1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2674_
timestamp 1698431365
transform -1 0 38080 0 -1 37632
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2675_
timestamp 1698431365
transform -1 0 40096 0 1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2676_
timestamp 1698431365
transform 1 0 34048 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2677_
timestamp 1698431365
transform 1 0 34272 0 -1 39200
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2678_
timestamp 1698431365
transform -1 0 30240 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2679_
timestamp 1698431365
transform -1 0 32704 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2680_
timestamp 1698431365
transform -1 0 33600 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2681_
timestamp 1698431365
transform -1 0 40432 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2682_
timestamp 1698431365
transform 1 0 29904 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2683_
timestamp 1698431365
transform -1 0 34832 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2684_
timestamp 1698431365
transform -1 0 42896 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2685_
timestamp 1698431365
transform -1 0 47712 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2686_
timestamp 1698431365
transform -1 0 39536 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2687_
timestamp 1698431365
transform -1 0 37408 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2688_
timestamp 1698431365
transform -1 0 37632 0 -1 43904
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2689_
timestamp 1698431365
transform 1 0 32032 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2690_
timestamp 1698431365
transform -1 0 34048 0 1 42336
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2691_
timestamp 1698431365
transform -1 0 35504 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2692_
timestamp 1698431365
transform -1 0 34160 0 1 43904
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2693_
timestamp 1698431365
transform -1 0 34720 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2694_
timestamp 1698431365
transform 1 0 33600 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2695_
timestamp 1698431365
transform 1 0 30576 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2696_
timestamp 1698431365
transform -1 0 50512 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2697_
timestamp 1698431365
transform 1 0 36064 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2698_
timestamp 1698431365
transform -1 0 36624 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2699_
timestamp 1698431365
transform -1 0 38192 0 1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2700_
timestamp 1698431365
transform 1 0 36960 0 -1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2701_
timestamp 1698431365
transform -1 0 43792 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2702_
timestamp 1698431365
transform -1 0 40880 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2703_
timestamp 1698431365
transform -1 0 41776 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2704_
timestamp 1698431365
transform 1 0 41776 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2705_
timestamp 1698431365
transform 1 0 41440 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2706_
timestamp 1698431365
transform 1 0 42336 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2707_
timestamp 1698431365
transform -1 0 42560 0 -1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2708_
timestamp 1698431365
transform -1 0 40768 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2709_
timestamp 1698431365
transform 1 0 38192 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2710_
timestamp 1698431365
transform -1 0 36960 0 -1 36064
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2711_
timestamp 1698431365
transform 1 0 34720 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2712_
timestamp 1698431365
transform -1 0 40544 0 -1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2713_
timestamp 1698431365
transform -1 0 38080 0 1 34496
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2714_
timestamp 1698431365
transform 1 0 37520 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2715_
timestamp 1698431365
transform 1 0 36848 0 1 32928
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2716_
timestamp 1698431365
transform -1 0 39424 0 -1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2717_
timestamp 1698431365
transform -1 0 38864 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2718_
timestamp 1698431365
transform -1 0 36624 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2719_
timestamp 1698431365
transform -1 0 33824 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2720_
timestamp 1698431365
transform 1 0 31696 0 1 36064
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2721_
timestamp 1698431365
transform -1 0 47600 0 -1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2722_
timestamp 1698431365
transform 1 0 33488 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2723_
timestamp 1698431365
transform 1 0 45360 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2724_
timestamp 1698431365
transform -1 0 47040 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2725_
timestamp 1698431365
transform 1 0 32928 0 -1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2726_
timestamp 1698431365
transform -1 0 34272 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2727_
timestamp 1698431365
transform -1 0 30800 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2728_
timestamp 1698431365
transform 1 0 29120 0 -1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2729_
timestamp 1698431365
transform 1 0 42336 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2730_
timestamp 1698431365
transform 1 0 43008 0 1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2731_
timestamp 1698431365
transform 1 0 43792 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2732_
timestamp 1698431365
transform 1 0 29008 0 1 40768
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2733_
timestamp 1698431365
transform 1 0 28560 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2734_
timestamp 1698431365
transform 1 0 28224 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2735_
timestamp 1698431365
transform -1 0 36848 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2736_
timestamp 1698431365
transform -1 0 36176 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2737_
timestamp 1698431365
transform -1 0 36288 0 -1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2738_
timestamp 1698431365
transform 1 0 29008 0 1 39200
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2739_
timestamp 1698431365
transform -1 0 44352 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2740_
timestamp 1698431365
transform -1 0 32256 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2741_
timestamp 1698431365
transform -1 0 32032 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2742_
timestamp 1698431365
transform -1 0 34384 0 -1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2743_
timestamp 1698431365
transform -1 0 32480 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2744_
timestamp 1698431365
transform 1 0 33600 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2745_
timestamp 1698431365
transform -1 0 35616 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2746_
timestamp 1698431365
transform -1 0 35728 0 1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2747_
timestamp 1698431365
transform -1 0 35728 0 1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2748_
timestamp 1698431365
transform -1 0 29008 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2749_
timestamp 1698431365
transform -1 0 29456 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2750_
timestamp 1698431365
transform 1 0 27328 0 -1 34496
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2751_
timestamp 1698431365
transform -1 0 30240 0 -1 32928
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2752_
timestamp 1698431365
transform -1 0 20608 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2753_
timestamp 1698431365
transform -1 0 19152 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2754_
timestamp 1698431365
transform -1 0 24976 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2755_
timestamp 1698431365
transform -1 0 39872 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2756_
timestamp 1698431365
transform -1 0 37520 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2757_
timestamp 1698431365
transform 1 0 38416 0 -1 34496
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2758_
timestamp 1698431365
transform 1 0 37408 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2759_
timestamp 1698431365
transform 1 0 44464 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2760_
timestamp 1698431365
transform -1 0 46032 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2761_
timestamp 1698431365
transform 1 0 42336 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2762_
timestamp 1698431365
transform 1 0 41776 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2763_
timestamp 1698431365
transform 1 0 43792 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2764_
timestamp 1698431365
transform -1 0 43792 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2765_
timestamp 1698431365
transform 1 0 43120 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2766_
timestamp 1698431365
transform -1 0 44464 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2767_
timestamp 1698431365
transform -1 0 41440 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2768_
timestamp 1698431365
transform 1 0 38080 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2769_
timestamp 1698431365
transform 1 0 39872 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2770_
timestamp 1698431365
transform -1 0 43120 0 1 32928
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2771_
timestamp 1698431365
transform 1 0 41104 0 -1 32928
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2772_
timestamp 1698431365
transform 1 0 49952 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2773_
timestamp 1698431365
transform -1 0 50736 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _2774_
timestamp 1698431365
transform -1 0 51520 0 -1 37632
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2775_
timestamp 1698431365
transform 1 0 46480 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2776_
timestamp 1698431365
transform 1 0 48720 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2777_
timestamp 1698431365
transform -1 0 50288 0 1 43904
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2778_
timestamp 1698431365
transform 1 0 49168 0 -1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _2779_
timestamp 1698431365
transform 1 0 49168 0 1 40768
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2780_
timestamp 1698431365
transform -1 0 51072 0 -1 42336
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2781_
timestamp 1698431365
transform 1 0 47824 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2782_
timestamp 1698431365
transform 1 0 52528 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2783_
timestamp 1698431365
transform 1 0 53200 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2784_
timestamp 1698431365
transform 1 0 41664 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2785_
timestamp 1698431365
transform 1 0 40880 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_2  _2786_
timestamp 1698431365
transform 1 0 50288 0 1 43904
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2787_
timestamp 1698431365
transform 1 0 52640 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2788_
timestamp 1698431365
transform 1 0 53984 0 1 40768
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2789_
timestamp 1698431365
transform -1 0 56224 0 -1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2790_
timestamp 1698431365
transform -1 0 43904 0 1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2791_
timestamp 1698431365
transform -1 0 42896 0 1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2792_
timestamp 1698431365
transform -1 0 42784 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2793_
timestamp 1698431365
transform -1 0 41440 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2794_
timestamp 1698431365
transform -1 0 37520 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2795_
timestamp 1698431365
transform 1 0 36848 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2796_
timestamp 1698431365
transform 1 0 37520 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2797_
timestamp 1698431365
transform 1 0 36624 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2798_
timestamp 1698431365
transform 1 0 28112 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2799_
timestamp 1698431365
transform -1 0 29568 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _2800_
timestamp 1698431365
transform -1 0 29344 0 -1 34496
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2801_
timestamp 1698431365
transform 1 0 29008 0 1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2802_
timestamp 1698431365
transform 1 0 27552 0 1 32928
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_2  _2803_
timestamp 1698431365
transform -1 0 28112 0 -1 26656
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2804_
timestamp 1698431365
transform 1 0 22512 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2805_
timestamp 1698431365
transform 1 0 40992 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2806_
timestamp 1698431365
transform 1 0 40768 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2807_
timestamp 1698431365
transform 1 0 41888 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2808_
timestamp 1698431365
transform -1 0 43456 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2809_
timestamp 1698431365
transform -1 0 45584 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2810_
timestamp 1698431365
transform -1 0 44464 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2811_
timestamp 1698431365
transform 1 0 42896 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2812_
timestamp 1698431365
transform 1 0 44688 0 1 32928
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _2813_
timestamp 1698431365
transform -1 0 46144 0 -1 32928
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2814_
timestamp 1698431365
transform 1 0 54432 0 -1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2815_
timestamp 1698431365
transform 1 0 55216 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2816_
timestamp 1698431365
transform -1 0 54768 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2817_
timestamp 1698431365
transform 1 0 55664 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2818_
timestamp 1698431365
transform 1 0 46144 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2819_
timestamp 1698431365
transform -1 0 53200 0 -1 43904
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2820_
timestamp 1698431365
transform 1 0 52304 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _2821_
timestamp 1698431365
transform 1 0 53200 0 -1 42336
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2822_
timestamp 1698431365
transform 1 0 48608 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2823_
timestamp 1698431365
transform 1 0 51184 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2824_
timestamp 1698431365
transform -1 0 53200 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2825_
timestamp 1698431365
transform -1 0 41888 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2826_
timestamp 1698431365
transform 1 0 44464 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2827_
timestamp 1698431365
transform 1 0 49056 0 -1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2828_
timestamp 1698431365
transform 1 0 51184 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2829_
timestamp 1698431365
transform 1 0 53424 0 -1 39200
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_2  _2830_
timestamp 1698431365
transform -1 0 57344 0 1 36064
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2831_
timestamp 1698431365
transform 1 0 39536 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2832_
timestamp 1698431365
transform -1 0 39536 0 1 31360
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2833_
timestamp 1698431365
transform 1 0 41440 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2834_
timestamp 1698431365
transform -1 0 43456 0 -1 29792
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2835_
timestamp 1698431365
transform 1 0 29344 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2836_
timestamp 1698431365
transform -1 0 29568 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2837_
timestamp 1698431365
transform -1 0 28784 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2838_
timestamp 1698431365
transform 1 0 29008 0 1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2839_
timestamp 1698431365
transform 1 0 31248 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2840_
timestamp 1698431365
transform 1 0 30352 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2841_
timestamp 1698431365
transform -1 0 34048 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2842_
timestamp 1698431365
transform 1 0 29792 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2843_
timestamp 1698431365
transform -1 0 33264 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2844_
timestamp 1698431365
transform 1 0 31696 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2845_
timestamp 1698431365
transform 1 0 37856 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2846_
timestamp 1698431365
transform 1 0 34160 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2847_
timestamp 1698431365
transform 1 0 42896 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _2848_
timestamp 1698431365
transform -1 0 45696 0 -1 31360
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2849_
timestamp 1698431365
transform 1 0 53424 0 1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2850_
timestamp 1698431365
transform 1 0 54544 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2851_
timestamp 1698431365
transform 1 0 56448 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2852_
timestamp 1698431365
transform 1 0 46928 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2853_
timestamp 1698431365
transform 1 0 51072 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2854_
timestamp 1698431365
transform 1 0 50624 0 1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2855_
timestamp 1698431365
transform 1 0 51184 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _2856_
timestamp 1698431365
transform 1 0 51296 0 -1 39200
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2857_
timestamp 1698431365
transform 1 0 53088 0 1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2858_
timestamp 1698431365
transform 1 0 50512 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2859_
timestamp 1698431365
transform 1 0 49504 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2860_
timestamp 1698431365
transform 1 0 51072 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2861_
timestamp 1698431365
transform 1 0 43904 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2862_
timestamp 1698431365
transform 1 0 43232 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2863_
timestamp 1698431365
transform 1 0 44464 0 -1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2864_
timestamp 1698431365
transform 1 0 51520 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2865_
timestamp 1698431365
transform 1 0 53312 0 1 34496
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2866_
timestamp 1698431365
transform -1 0 55664 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2867_
timestamp 1698431365
transform -1 0 54768 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2868_
timestamp 1698431365
transform -1 0 55888 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2869_
timestamp 1698431365
transform 1 0 44912 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2870_
timestamp 1698431365
transform 1 0 46144 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2871_
timestamp 1698431365
transform -1 0 46480 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2872_
timestamp 1698431365
transform 1 0 45696 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2873_
timestamp 1698431365
transform -1 0 46816 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2874_
timestamp 1698431365
transform 1 0 43568 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2875_
timestamp 1698431365
transform -1 0 44464 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2876_
timestamp 1698431365
transform -1 0 31808 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2877_
timestamp 1698431365
transform -1 0 30128 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2878_
timestamp 1698431365
transform -1 0 30128 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2879_
timestamp 1698431365
transform 1 0 29008 0 1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2880_
timestamp 1698431365
transform 1 0 29568 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2881_
timestamp 1698431365
transform -1 0 32144 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2882_
timestamp 1698431365
transform 1 0 30128 0 -1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2883_
timestamp 1698431365
transform 1 0 32032 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2884_
timestamp 1698431365
transform 1 0 31136 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2885_
timestamp 1698431365
transform 1 0 31808 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2886_
timestamp 1698431365
transform 1 0 32928 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2887_
timestamp 1698431365
transform -1 0 34384 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2888_
timestamp 1698431365
transform 1 0 32928 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2889_
timestamp 1698431365
transform -1 0 41328 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2890_
timestamp 1698431365
transform -1 0 40544 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2891_
timestamp 1698431365
transform -1 0 45584 0 1 31360
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2892_
timestamp 1698431365
transform 1 0 44688 0 1 29792
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2893_
timestamp 1698431365
transform -1 0 54544 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2894_
timestamp 1698431365
transform -1 0 53312 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2895_
timestamp 1698431365
transform -1 0 55328 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2896_
timestamp 1698431365
transform 1 0 52528 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2897_
timestamp 1698431365
transform -1 0 52304 0 1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2898_
timestamp 1698431365
transform -1 0 53424 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _2899_
timestamp 1698431365
transform 1 0 51632 0 -1 36064
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2900_
timestamp 1698431365
transform -1 0 50176 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2901_
timestamp 1698431365
transform -1 0 48272 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2902_
timestamp 1698431365
transform 1 0 45136 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2903_
timestamp 1698431365
transform -1 0 46144 0 1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2904_
timestamp 1698431365
transform 1 0 48160 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2905_
timestamp 1698431365
transform 1 0 47264 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2906_
timestamp 1698431365
transform 1 0 51184 0 -1 32928
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2907_
timestamp 1698431365
transform -1 0 54768 0 -1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2908_
timestamp 1698431365
transform -1 0 45136 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2909_
timestamp 1698431365
transform -1 0 45696 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2910_
timestamp 1698431365
transform -1 0 38976 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2911_
timestamp 1698431365
transform 1 0 31696 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2912_
timestamp 1698431365
transform -1 0 33152 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2913_
timestamp 1698431365
transform -1 0 32704 0 -1 32928
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2914_
timestamp 1698431365
transform 1 0 38304 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2915_
timestamp 1698431365
transform 1 0 39536 0 -1 26656
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2916_
timestamp 1698431365
transform 1 0 39424 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2917_
timestamp 1698431365
transform -1 0 52304 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2918_
timestamp 1698431365
transform -1 0 51184 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2919_
timestamp 1698431365
transform 1 0 53200 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2920_
timestamp 1698431365
transform -1 0 49728 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2921_
timestamp 1698431365
transform -1 0 49504 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2922_
timestamp 1698431365
transform -1 0 47712 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2923_
timestamp 1698431365
transform -1 0 47824 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2924_
timestamp 1698431365
transform 1 0 47264 0 -1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _2925_
timestamp 1698431365
transform 1 0 48608 0 -1 34496
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2926_
timestamp 1698431365
transform 1 0 50512 0 -1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2927_
timestamp 1698431365
transform 1 0 49056 0 1 31360
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2928_
timestamp 1698431365
transform 1 0 51520 0 -1 31360
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2929_
timestamp 1698431365
transform -1 0 51520 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2930_
timestamp 1698431365
transform -1 0 50400 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2931_
timestamp 1698431365
transform -1 0 37520 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2932_
timestamp 1698431365
transform -1 0 39312 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2933_
timestamp 1698431365
transform 1 0 35616 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2934_
timestamp 1698431365
transform 1 0 32928 0 -1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _2935_
timestamp 1698431365
transform 1 0 33936 0 1 29792
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2936_
timestamp 1698431365
transform 1 0 33600 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2937_
timestamp 1698431365
transform -1 0 37408 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2938_
timestamp 1698431365
transform 1 0 34496 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2939_
timestamp 1698431365
transform 1 0 47600 0 1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2940_
timestamp 1698431365
transform 1 0 48608 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2941_
timestamp 1698431365
transform 1 0 49728 0 1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2942_
timestamp 1698431365
transform 1 0 47824 0 1 32928
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2943_
timestamp 1698431365
transform 1 0 46928 0 -1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2944_
timestamp 1698431365
transform -1 0 49728 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2945_
timestamp 1698431365
transform -1 0 48272 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2946_
timestamp 1698431365
transform -1 0 35616 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2947_
timestamp 1698431365
transform 1 0 35504 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2948_
timestamp 1698431365
transform 1 0 32480 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2949_
timestamp 1698431365
transform 1 0 33040 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2950_
timestamp 1698431365
transform -1 0 35504 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2951_
timestamp 1698431365
transform -1 0 35392 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2952_
timestamp 1698431365
transform -1 0 37856 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2953_
timestamp 1698431365
transform 1 0 35392 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2954_
timestamp 1698431365
transform -1 0 39536 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2955_
timestamp 1698431365
transform 1 0 34496 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2956_
timestamp 1698431365
transform 1 0 34048 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2957_
timestamp 1698431365
transform -1 0 36288 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2958_
timestamp 1698431365
transform -1 0 35952 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2959_
timestamp 1698431365
transform -1 0 35056 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2960_
timestamp 1698431365
transform 1 0 39536 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2961_
timestamp 1698431365
transform -1 0 30800 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2962_
timestamp 1698431365
transform 1 0 36848 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2963_
timestamp 1698431365
transform -1 0 41104 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2964_
timestamp 1698431365
transform -1 0 40544 0 1 21952
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2965_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 39312 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2966_
timestamp 1698431365
transform 1 0 42112 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2967_
timestamp 1698431365
transform 1 0 47152 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2968_
timestamp 1698431365
transform 1 0 46704 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2969_
timestamp 1698431365
transform 1 0 44688 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2970_
timestamp 1698431365
transform -1 0 35056 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2971_
timestamp 1698431365
transform 1 0 28224 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2972_
timestamp 1698431365
transform 1 0 35392 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2973_
timestamp 1698431365
transform 1 0 44464 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2974_
timestamp 1698431365
transform 1 0 41104 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2975_
timestamp 1698431365
transform 1 0 46704 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2976_
timestamp 1698431365
transform -1 0 46816 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2977_
timestamp 1698431365
transform 1 0 40768 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2978_
timestamp 1698431365
transform 1 0 36176 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2979_
timestamp 1698431365
transform 1 0 32928 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2980_
timestamp 1698431365
transform 1 0 30352 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2981_
timestamp 1698431365
transform 1 0 28560 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2982_
timestamp 1698431365
transform -1 0 12656 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2983_
timestamp 1698431365
transform -1 0 11760 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2984_
timestamp 1698431365
transform -1 0 16016 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2985_
timestamp 1698431365
transform -1 0 23408 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2986_
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2987_
timestamp 1698431365
transform 1 0 24080 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2988_
timestamp 1698431365
transform 1 0 23744 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2989_
timestamp 1698431365
transform 1 0 17584 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2990_
timestamp 1698431365
transform -1 0 24416 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2991_
timestamp 1698431365
transform 1 0 34608 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2992_
timestamp 1698431365
transform 1 0 31472 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2993_
timestamp 1698431365
transform 1 0 39088 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2994_
timestamp 1698431365
transform 1 0 33376 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2995_
timestamp 1698431365
transform 1 0 34048 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2996_
timestamp 1698431365
transform 1 0 38640 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2997_
timestamp 1698431365
transform 1 0 45136 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2999_
timestamp 1698431365
transform 1 0 48608 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1482__A1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 44912 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1482__A2
timestamp 1698431365
transform -1 0 45136 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1482__A3
timestamp 1698431365
transform -1 0 45584 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1483__A1
timestamp 1698431365
transform 1 0 43568 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1483__A2
timestamp 1698431365
transform -1 0 42784 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1484__A1
timestamp 1698431365
transform -1 0 46144 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1485__A1
timestamp 1698431365
transform 1 0 45472 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1486__A1
timestamp 1698431365
transform -1 0 47152 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1487__I
timestamp 1698431365
transform -1 0 47600 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1488__A1
timestamp 1698431365
transform -1 0 47600 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1488__A3
timestamp 1698431365
transform 1 0 47824 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1490__I
timestamp 1698431365
transform 1 0 46928 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1492__A2
timestamp 1698431365
transform 1 0 30464 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1494__I
timestamp 1698431365
transform -1 0 28000 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1497__I
timestamp 1698431365
transform -1 0 38192 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1508__A2
timestamp 1698431365
transform 1 0 29792 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1525__A2
timestamp 1698431365
transform -1 0 26992 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1540__A2
timestamp 1698431365
transform 1 0 31920 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1541__A2
timestamp 1698431365
transform 1 0 27888 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1549__A1
timestamp 1698431365
transform -1 0 29232 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1549__A2
timestamp 1698431365
transform 1 0 30240 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1552__A2
timestamp 1698431365
transform -1 0 33264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1556__A2
timestamp 1698431365
transform 1 0 34384 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1615__A1
timestamp 1698431365
transform 1 0 30128 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1620__B2
timestamp 1698431365
transform 1 0 39312 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1622__I
timestamp 1698431365
transform -1 0 45472 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1639__A1
timestamp 1698431365
transform 1 0 29680 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1642__A2
timestamp 1698431365
transform 1 0 28112 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1675__A1
timestamp 1698431365
transform 1 0 45248 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1682__A1
timestamp 1698431365
transform 1 0 45472 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1700__A2
timestamp 1698431365
transform -1 0 38192 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1704__I
timestamp 1698431365
transform 1 0 47600 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1706__A1
timestamp 1698431365
transform 1 0 47040 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1724__A1
timestamp 1698431365
transform -1 0 49728 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1748__A1
timestamp 1698431365
transform 1 0 51296 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1755__A1
timestamp 1698431365
transform -1 0 51856 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1758__A2
timestamp 1698431365
transform 1 0 38864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1769__A2
timestamp 1698431365
transform 1 0 38752 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1772__A1
timestamp 1698431365
transform 1 0 41552 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1774__I
timestamp 1698431365
transform 1 0 35728 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1788__A1
timestamp 1698431365
transform -1 0 51744 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1794__A2
timestamp 1698431365
transform 1 0 52304 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1801__B1
timestamp 1698431365
transform 1 0 42112 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1809__A2
timestamp 1698431365
transform 1 0 52080 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1823__A1
timestamp 1698431365
transform 1 0 36960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1823__A2
timestamp 1698431365
transform 1 0 37408 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1826__I1
timestamp 1698431365
transform 1 0 35728 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1833__A1
timestamp 1698431365
transform 1 0 54208 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1834__B1
timestamp 1698431365
transform -1 0 34496 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1840__A1
timestamp 1698431365
transform 1 0 53200 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1841__A1
timestamp 1698431365
transform 1 0 28560 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1844__A2
timestamp 1698431365
transform 1 0 38976 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1845__I1
timestamp 1698431365
transform 1 0 38528 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1868__A1
timestamp 1698431365
transform 1 0 9184 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1877__A1
timestamp 1698431365
transform -1 0 8736 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1890__A2
timestamp 1698431365
transform 1 0 8064 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1901__A2
timestamp 1698431365
transform 1 0 6160 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1915__A2
timestamp 1698431365
transform -1 0 5152 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1937__A1
timestamp 1698431365
transform 1 0 15904 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1940__I
timestamp 1698431365
transform 1 0 14000 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1943__A2
timestamp 1698431365
transform 1 0 12320 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1950__A1
timestamp 1698431365
transform 1 0 13216 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1967__A2
timestamp 1698431365
transform -1 0 9072 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2000__A1
timestamp 1698431365
transform 1 0 24640 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2041__A1
timestamp 1698431365
transform -1 0 15120 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2060__A1
timestamp 1698431365
transform -1 0 37744 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2061__A1
timestamp 1698431365
transform 1 0 42896 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2083__A1
timestamp 1698431365
transform 1 0 15120 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2112__A1
timestamp 1698431365
transform 1 0 20384 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2119__A1
timestamp 1698431365
transform 1 0 15904 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2140__A1
timestamp 1698431365
transform 1 0 32032 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2140__B2
timestamp 1698431365
transform -1 0 28560 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2146__A2
timestamp 1698431365
transform 1 0 43008 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2156__A1
timestamp 1698431365
transform -1 0 21728 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2172__A1
timestamp 1698431365
transform -1 0 30128 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2172__A2
timestamp 1698431365
transform 1 0 27888 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2172__C
timestamp 1698431365
transform 1 0 30128 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2173__A2
timestamp 1698431365
transform -1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2180__A1
timestamp 1698431365
transform 1 0 23072 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2200__A1
timestamp 1698431365
transform 1 0 38864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2200__A2
timestamp 1698431365
transform 1 0 39872 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2202__A1
timestamp 1698431365
transform 1 0 39648 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2213__B1
timestamp 1698431365
transform 1 0 30800 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2215__A2
timestamp 1698431365
transform 1 0 35168 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2220__C
timestamp 1698431365
transform -1 0 30352 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2223__A2
timestamp 1698431365
transform -1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2270__A2
timestamp 1698431365
transform 1 0 10864 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2304__A2
timestamp 1698431365
transform 1 0 22064 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2329__A2
timestamp 1698431365
transform 1 0 23968 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2374__A1
timestamp 1698431365
transform 1 0 21056 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2375__A1
timestamp 1698431365
transform 1 0 20608 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2381__B1
timestamp 1698431365
transform 1 0 31360 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2383__A1
timestamp 1698431365
transform 1 0 31584 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2385__A2
timestamp 1698431365
transform 1 0 14112 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2407__A1
timestamp 1698431365
transform 1 0 20160 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2426__A2
timestamp 1698431365
transform 1 0 16240 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2434__A3
timestamp 1698431365
transform 1 0 16352 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2435__A1
timestamp 1698431365
transform 1 0 18704 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2436__B
timestamp 1698431365
transform -1 0 17024 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2437__I
timestamp 1698431365
transform 1 0 21504 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2440__A2
timestamp 1698431365
transform -1 0 13216 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2466__A2
timestamp 1698431365
transform 1 0 15008 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2467__A1
timestamp 1698431365
transform 1 0 20160 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2469__A2
timestamp 1698431365
transform 1 0 15680 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2471__A2
timestamp 1698431365
transform -1 0 14000 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2472__A1
timestamp 1698431365
transform 1 0 16800 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2473__A2
timestamp 1698431365
transform 1 0 15456 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2478__A1
timestamp 1698431365
transform -1 0 15680 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2482__A2
timestamp 1698431365
transform 1 0 16576 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2483__A2
timestamp 1698431365
transform -1 0 11872 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2484__A2
timestamp 1698431365
transform 1 0 13104 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2513__A2
timestamp 1698431365
transform 1 0 12544 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2521__A1
timestamp 1698431365
transform 1 0 17472 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2552__I
timestamp 1698431365
transform -1 0 24304 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2555__A1
timestamp 1698431365
transform -1 0 22960 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2555__A2
timestamp 1698431365
transform 1 0 23744 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2586__C
timestamp 1698431365
transform -1 0 29456 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2587__A2
timestamp 1698431365
transform -1 0 23968 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2589__A1
timestamp 1698431365
transform -1 0 27328 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2592__A2
timestamp 1698431365
transform 1 0 22960 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2597__A1
timestamp 1698431365
transform 1 0 27776 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2599__A2
timestamp 1698431365
transform 1 0 21056 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2603__A1
timestamp 1698431365
transform 1 0 45920 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2633__A2
timestamp 1698431365
transform 1 0 44800 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2654__A2
timestamp 1698431365
transform 1 0 39760 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2679__A2
timestamp 1698431365
transform -1 0 32144 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2682__A2
timestamp 1698431365
transform 1 0 30688 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2685__I
timestamp 1698431365
transform 1 0 45920 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2689__A2
timestamp 1698431365
transform 1 0 33376 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2697__A2
timestamp 1698431365
transform -1 0 36064 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2700__A1
timestamp 1698431365
transform 1 0 38304 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2710__A1
timestamp 1698431365
transform 1 0 37072 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2716__A1
timestamp 1698431365
transform 1 0 39648 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2717__A1
timestamp 1698431365
transform 1 0 39760 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2727__A2
timestamp 1698431365
transform 1 0 31024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2730__B2
timestamp 1698431365
transform -1 0 42336 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2733__A2
timestamp 1698431365
transform -1 0 28560 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2734__A2
timestamp 1698431365
transform -1 0 28224 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2736__A2
timestamp 1698431365
transform 1 0 36400 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2739__A1
timestamp 1698431365
transform 1 0 44912 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2749__I
timestamp 1698431365
transform -1 0 30464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2751__A1
timestamp 1698431365
transform -1 0 30464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2754__A1
timestamp 1698431365
transform -1 0 24416 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2754__A2
timestamp 1698431365
transform 1 0 25312 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2775__A1
timestamp 1698431365
transform 1 0 47264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2779__A1
timestamp 1698431365
transform 1 0 50624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2790__A2
timestamp 1698431365
transform -1 0 46928 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2791__A2
timestamp 1698431365
transform 1 0 43680 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2799__I
timestamp 1698431365
transform 1 0 28672 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2818__A1
timestamp 1698431365
transform 1 0 45920 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2831__A1
timestamp 1698431365
transform 1 0 40320 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2834__A2
timestamp 1698431365
transform -1 0 44240 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2836__A2
timestamp 1698431365
transform -1 0 31024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2843__I
timestamp 1698431365
transform -1 0 33488 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2845__A1
timestamp 1698431365
transform 1 0 38080 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2847__A2
timestamp 1698431365
transform 1 0 44128 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2848__B2
timestamp 1698431365
transform 1 0 45920 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2853__A1
timestamp 1698431365
transform -1 0 51072 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2856__A1
timestamp 1698431365
transform 1 0 51072 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2876__A1
timestamp 1698431365
transform 1 0 31808 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2877__A2
timestamp 1698431365
transform 1 0 30352 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2878__A2
timestamp 1698431365
transform -1 0 30576 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2881__A1
timestamp 1698431365
transform 1 0 32368 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2887__A1
timestamp 1698431365
transform -1 0 35168 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2889__A2
timestamp 1698431365
transform 1 0 41552 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2890__A2
timestamp 1698431365
transform 1 0 40768 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2896__A1
timestamp 1698431365
transform 1 0 53312 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2910__A1
timestamp 1698431365
transform 1 0 39200 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2913__A1
timestamp 1698431365
transform 1 0 31696 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2914__C
timestamp 1698431365
transform 1 0 39648 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2935__C
timestamp 1698431365
transform 1 0 33712 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2937__A1
timestamp 1698431365
transform -1 0 36848 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2960__A1
timestamp 1698431365
transform 1 0 39312 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2965__CLK
timestamp 1698431365
transform 1 0 42784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2966__CLK
timestamp 1698431365
transform 1 0 45584 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2967__CLK
timestamp 1698431365
transform 1 0 46928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2968__CLK
timestamp 1698431365
transform 1 0 46480 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2969__CLK
timestamp 1698431365
transform 1 0 44240 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2970__CLK
timestamp 1698431365
transform 1 0 35280 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2971__CLK
timestamp 1698431365
transform -1 0 31248 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2972__CLK
timestamp 1698431365
transform 1 0 38752 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2973__CLK
timestamp 1698431365
transform 1 0 47936 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2974__CLK
timestamp 1698431365
transform 1 0 45808 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2975__CLK
timestamp 1698431365
transform 1 0 46592 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2976__CLK
timestamp 1698431365
transform 1 0 47040 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2977__CLK
timestamp 1698431365
transform 1 0 45808 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2978__CLK
timestamp 1698431365
transform 1 0 39424 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2979__CLK
timestamp 1698431365
transform 1 0 32480 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2980__CLK
timestamp 1698431365
transform 1 0 30576 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2981__CLK
timestamp 1698431365
transform 1 0 32032 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2986__CLK
timestamp 1698431365
transform 1 0 28560 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2990__CLK
timestamp 1698431365
transform 1 0 23632 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2991__CLK
timestamp 1698431365
transform 1 0 38192 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2992__CLK
timestamp 1698431365
transform -1 0 31584 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2993__CLK
timestamp 1698431365
transform 1 0 42560 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2994__CLK
timestamp 1698431365
transform 1 0 37072 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2995__CLK
timestamp 1698431365
transform 1 0 38080 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2996__CLK
timestamp 1698431365
transform -1 0 42112 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2997__CLK
timestamp 1698431365
transform 1 0 46256 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698431365
transform -1 0 29456 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_0__f_clk_I
timestamp 1698431365
transform 1 0 32368 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_1__f_clk_I
timestamp 1698431365
transform 1 0 26992 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_2__f_clk_I
timestamp 1698431365
transform -1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_3__f_clk_I
timestamp 1698431365
transform 1 0 38528 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform -1 0 57904 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform -1 0 26880 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform -1 0 28784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform -1 0 30128 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform -1 0 57232 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform -1 0 57232 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform -1 0 57680 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698431365
transform -1 0 57680 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698431365
transform -1 0 57680 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698431365
transform -1 0 57680 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698431365
transform -1 0 58352 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698431365
transform -1 0 57680 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698431365
transform -1 0 57680 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1698431365
transform -1 0 57680 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1698431365
transform -1 0 57680 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1698431365
transform -1 0 57680 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1698431365
transform -1 0 57008 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1698431365
transform -1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1698431365
transform 1 0 1792 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1698431365
transform 1 0 3584 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1698431365
transform 1 0 4480 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input22_I
timestamp 1698431365
transform 1 0 1792 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input23_I
timestamp 1698431365
transform 1 0 3136 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input24_I
timestamp 1698431365
transform 1 0 1792 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input25_I
timestamp 1698431365
transform -1 0 16576 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input26_I
timestamp 1698431365
transform 1 0 14448 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input27_I
timestamp 1698431365
transform -1 0 9744 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input28_I
timestamp 1698431365
transform 1 0 2464 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input29_I
timestamp 1698431365
transform 1 0 41216 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input30_I
timestamp 1698431365
transform -1 0 2240 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input31_I
timestamp 1698431365
transform 1 0 3136 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input32_I
timestamp 1698431365
transform 1 0 2240 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input33_I
timestamp 1698431365
transform 1 0 2464 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input34_I
timestamp 1698431365
transform 1 0 53760 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input35_I
timestamp 1698431365
transform -1 0 45472 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input36_I
timestamp 1698431365
transform 1 0 44912 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input37_I
timestamp 1698431365
transform 1 0 48048 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input38_I
timestamp 1698431365
transform -1 0 35168 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input39_I
timestamp 1698431365
transform -1 0 40432 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input40_I
timestamp 1698431365
transform 1 0 39424 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input41_I
timestamp 1698431365
transform 1 0 52752 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input42_I
timestamp 1698431365
transform 1 0 40656 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input43_I
timestamp 1698431365
transform 1 0 46256 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input44_I
timestamp 1698431365
transform -1 0 28336 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input45_I
timestamp 1698431365
transform -1 0 25648 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input46_I
timestamp 1698431365
transform 1 0 43344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input47_I
timestamp 1698431365
transform 1 0 34832 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input48_I
timestamp 1698431365
transform 1 0 5152 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input49_I
timestamp 1698431365
transform 1 0 4928 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input50_I
timestamp 1698431365
transform -1 0 31024 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input51_I
timestamp 1698431365
transform 1 0 2240 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input52_I
timestamp 1698431365
transform 1 0 1792 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input53_I
timestamp 1698431365
transform 1 0 3136 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input54_I
timestamp 1698431365
transform 1 0 2464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input55_I
timestamp 1698431365
transform 1 0 2912 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input56_I
timestamp 1698431365
transform -1 0 14224 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input57_I
timestamp 1698431365
transform 1 0 1792 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input58_I
timestamp 1698431365
transform 1 0 3584 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input59_I
timestamp 1698431365
transform 1 0 3136 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input60_I
timestamp 1698431365
transform 1 0 1792 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input61_I
timestamp 1698431365
transform -1 0 25200 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input62_I
timestamp 1698431365
transform -1 0 8288 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input63_I
timestamp 1698431365
transform -1 0 9184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input64_I
timestamp 1698431365
transform -1 0 16128 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input65_I
timestamp 1698431365
transform 1 0 19152 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input66_I
timestamp 1698431365
transform -1 0 35616 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input67_I
timestamp 1698431365
transform -1 0 37296 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input68_I
timestamp 1698431365
transform -1 0 36624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input69_I
timestamp 1698431365
transform -1 0 31136 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input70_I
timestamp 1698431365
transform 1 0 53312 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input71_I
timestamp 1698431365
transform 1 0 44912 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input72_I
timestamp 1698431365
transform -1 0 26992 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input73_I
timestamp 1698431365
transform 1 0 54208 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input74_I
timestamp 1698431365
transform 1 0 53200 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input75_I
timestamp 1698431365
transform -1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input76_I
timestamp 1698431365
transform -1 0 31024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input77_I
timestamp 1698431365
transform 1 0 33152 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input78_I
timestamp 1698431365
transform 1 0 43792 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input79_I
timestamp 1698431365
transform 1 0 46704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input80_I
timestamp 1698431365
transform 1 0 4592 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input81_I
timestamp 1698431365
transform 1 0 4032 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input82_I
timestamp 1698431365
transform -1 0 57008 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output87_I
timestamp 1698431365
transform -1 0 55440 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output90_I
timestamp 1698431365
transform 1 0 30576 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output95_I
timestamp 1698431365
transform 1 0 4704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output97_I
timestamp 1698431365
transform 1 0 30352 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output98_I
timestamp 1698431365
transform 1 0 27104 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output100_I
timestamp 1698431365
transform -1 0 5376 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output101_I
timestamp 1698431365
transform 1 0 55216 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output102_I
timestamp 1698431365
transform 1 0 36848 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output104_I
timestamp 1698431365
transform -1 0 55440 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output110_I
timestamp 1698431365
transform 1 0 39648 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output112_I
timestamp 1698431365
transform -1 0 55440 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output114_I
timestamp 1698431365
transform -1 0 55440 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29456 0 1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1698431365
transform 1 0 25872 0 -1 23520
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1698431365
transform -1 0 26768 0 1 25088
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1698431365
transform 1 0 40768 0 -1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1698431365
transform 1 0 38752 0 1 23520
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_104 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 12992 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_112 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13888 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_121
timestamp 1698431365
transform 1 0 14896 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_129 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15792 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_133 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 16240 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_135
timestamp 1698431365
transform 1 0 16464 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_138
timestamp 1698431365
transform 1 0 16800 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_172
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_180
timestamp 1698431365
transform 1 0 21504 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_185 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22064 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_201
timestamp 1698431365
transform 1 0 23856 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_203
timestamp 1698431365
transform 1 0 24080 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_206
timestamp 1698431365
transform 1 0 24416 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_210
timestamp 1698431365
transform 1 0 24864 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_213
timestamp 1698431365
transform 1 0 25200 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_235
timestamp 1698431365
transform 1 0 27664 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_237
timestamp 1698431365
transform 1 0 27888 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_302
timestamp 1698431365
transform 1 0 35168 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_362
timestamp 1698431365
transform 1 0 41888 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_373
timestamp 1698431365
transform 1 0 43120 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_399
timestamp 1698431365
transform 1 0 46032 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_403
timestamp 1698431365
transform 1 0 46480 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_407
timestamp 1698431365
transform 1 0 46928 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_420
timestamp 1698431365
transform 1 0 48384 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_436
timestamp 1698431365
transform 1 0 50176 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_440
timestamp 1698431365
transform 1 0 50624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_444
timestamp 1698431365
transform 1 0 51072 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_478
timestamp 1698431365
transform 1 0 54880 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_494
timestamp 1698431365
transform 1 0 56672 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_502
timestamp 1698431365
transform 1 0 57568 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_506
timestamp 1698431365
transform 1 0 58016 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_508
timestamp 1698431365
transform 1 0 58240 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698431365
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698431365
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_142
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_206
timestamp 1698431365
transform 1 0 24416 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_212
timestamp 1698431365
transform 1 0 25088 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_220
timestamp 1698431365
transform 1 0 25984 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_224
timestamp 1698431365
transform 1 0 26432 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_226
timestamp 1698431365
transform 1 0 26656 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_229
timestamp 1698431365
transform 1 0 26992 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_237
timestamp 1698431365
transform 1 0 27888 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_279
timestamp 1698431365
transform 1 0 32592 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_288
timestamp 1698431365
transform 1 0 33600 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_332
timestamp 1698431365
transform 1 0 38528 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_334
timestamp 1698431365
transform 1 0 38752 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_347
timestamp 1698431365
transform 1 0 40208 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_349
timestamp 1698431365
transform 1 0 40432 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_360
timestamp 1698431365
transform 1 0 41664 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_422
timestamp 1698431365
transform 1 0 48608 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_486
timestamp 1698431365
transform 1 0 55776 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_492
timestamp 1698431365
transform 1 0 56448 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_508
timestamp 1698431365
transform 1 0 58240 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698431365
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698431365
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698431365
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_241
timestamp 1698431365
transform 1 0 28336 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_247
timestamp 1698431365
transform 1 0 29008 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_259
timestamp 1698431365
transform 1 0 30352 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_269
timestamp 1698431365
transform 1 0 31472 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_348
timestamp 1698431365
transform 1 0 40320 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_358
timestamp 1698431365
transform 1 0 41440 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_360
timestamp 1698431365
transform 1 0 41664 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_375
timestamp 1698431365
transform 1 0 43344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_377
timestamp 1698431365
transform 1 0 43568 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_395
timestamp 1698431365
transform 1 0 45584 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_401
timestamp 1698431365
transform 1 0 46256 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_424
timestamp 1698431365
transform 1 0 48832 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_442
timestamp 1698431365
transform 1 0 50848 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_450
timestamp 1698431365
transform 1 0 51744 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_454
timestamp 1698431365
transform 1 0 52192 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_457
timestamp 1698431365
transform 1 0 52528 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_489
timestamp 1698431365
transform 1 0 56112 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_505
timestamp 1698431365
transform 1 0 57904 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698431365
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698431365
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698431365
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_212
timestamp 1698431365
transform 1 0 25088 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_219
timestamp 1698431365
transform 1 0 25872 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_223
timestamp 1698431365
transform 1 0 26320 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_261
timestamp 1698431365
transform 1 0 30576 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_277
timestamp 1698431365
transform 1 0 32368 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_279
timestamp 1698431365
transform 1 0 32592 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_305
timestamp 1698431365
transform 1 0 35504 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_340
timestamp 1698431365
transform 1 0 39424 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_373
timestamp 1698431365
transform 1 0 43120 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_377
timestamp 1698431365
transform 1 0 43568 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_396
timestamp 1698431365
transform 1 0 45696 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_417
timestamp 1698431365
transform 1 0 48048 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_419
timestamp 1698431365
transform 1 0 48272 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_422
timestamp 1698431365
transform 1 0 48608 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_454
timestamp 1698431365
transform 1 0 52192 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_467
timestamp 1698431365
transform 1 0 53648 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_483
timestamp 1698431365
transform 1 0 55440 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_487
timestamp 1698431365
transform 1 0 55888 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_489
timestamp 1698431365
transform 1 0 56112 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_492
timestamp 1698431365
transform 1 0 56448 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_508
timestamp 1698431365
transform 1 0 58240 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698431365
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_115
timestamp 1698431365
transform 1 0 14224 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_117
timestamp 1698431365
transform 1 0 14448 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_123
timestamp 1698431365
transform 1 0 15120 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_155
timestamp 1698431365
transform 1 0 18704 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698431365
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_177
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_193
timestamp 1698431365
transform 1 0 22960 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_197
timestamp 1698431365
transform 1 0 23408 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_199
timestamp 1698431365
transform 1 0 23632 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_213
timestamp 1698431365
transform 1 0 25200 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_244
timestamp 1698431365
transform 1 0 28672 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_256
timestamp 1698431365
transform 1 0 30016 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_260
timestamp 1698431365
transform 1 0 30464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_262
timestamp 1698431365
transform 1 0 30688 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_265
timestamp 1698431365
transform 1 0 31024 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_267
timestamp 1698431365
transform 1 0 31248 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_289
timestamp 1698431365
transform 1 0 33712 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_297
timestamp 1698431365
transform 1 0 34608 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_340
timestamp 1698431365
transform 1 0 39424 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_375
timestamp 1698431365
transform 1 0 43344 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_383
timestamp 1698431365
transform 1 0 44240 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_387
timestamp 1698431365
transform 1 0 44688 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_391
timestamp 1698431365
transform 1 0 45136 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_393
timestamp 1698431365
transform 1 0 45360 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_396
timestamp 1698431365
transform 1 0 45696 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_404
timestamp 1698431365
transform 1 0 46592 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_408
timestamp 1698431365
transform 1 0 47040 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_450
timestamp 1698431365
transform 1 0 51744 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_454
timestamp 1698431365
transform 1 0 52192 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_457
timestamp 1698431365
transform 1 0 52528 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_459
timestamp 1698431365
transform 1 0 52752 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_473
timestamp 1698431365
transform 1 0 54320 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_505
timestamp 1698431365
transform 1 0 57904 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_6
timestamp 1698431365
transform 1 0 2016 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_22
timestamp 1698431365
transform 1 0 3808 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_30
timestamp 1698431365
transform 1 0 4704 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_34
timestamp 1698431365
transform 1 0 5152 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_43
timestamp 1698431365
transform 1 0 6160 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_51
timestamp 1698431365
transform 1 0 7056 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_55
timestamp 1698431365
transform 1 0 7504 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_57
timestamp 1698431365
transform 1 0 7728 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_68
timestamp 1698431365
transform 1 0 8960 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_80
timestamp 1698431365
transform 1 0 10304 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_88
timestamp 1698431365
transform 1 0 11200 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_142
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_174
timestamp 1698431365
transform 1 0 20832 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_182
timestamp 1698431365
transform 1 0 21728 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_212
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_220
timestamp 1698431365
transform 1 0 25984 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_256
timestamp 1698431365
transform 1 0 30016 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_258
timestamp 1698431365
transform 1 0 30240 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698431365
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_282
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_286
timestamp 1698431365
transform 1 0 33376 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_305
timestamp 1698431365
transform 1 0 35504 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_319
timestamp 1698431365
transform 1 0 37072 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_340
timestamp 1698431365
transform 1 0 39424 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_348
timestamp 1698431365
transform 1 0 40320 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_362
timestamp 1698431365
transform 1 0 41888 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_370
timestamp 1698431365
transform 1 0 42784 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_374
timestamp 1698431365
transform 1 0 43232 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_388
timestamp 1698431365
transform 1 0 44800 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_396
timestamp 1698431365
transform 1 0 45696 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_400
timestamp 1698431365
transform 1 0 46144 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_402
timestamp 1698431365
transform 1 0 46368 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_415
timestamp 1698431365
transform 1 0 47824 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_419
timestamp 1698431365
transform 1 0 48272 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_430
timestamp 1698431365
transform 1 0 49504 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_434
timestamp 1698431365
transform 1 0 49952 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_457
timestamp 1698431365
transform 1 0 52528 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_505
timestamp 1698431365
transform 1 0 57904 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_8
timestamp 1698431365
transform 1 0 2240 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_12
timestamp 1698431365
transform 1 0 2688 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_16
timestamp 1698431365
transform 1 0 3136 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_24
timestamp 1698431365
transform 1 0 4032 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_31
timestamp 1698431365
transform 1 0 4816 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_81
timestamp 1698431365
transform 1 0 10416 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_85
timestamp 1698431365
transform 1 0 10864 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_99
timestamp 1698431365
transform 1 0 12432 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_103
timestamp 1698431365
transform 1 0 12880 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_119
timestamp 1698431365
transform 1 0 14672 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_169
timestamp 1698431365
transform 1 0 20272 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_173
timestamp 1698431365
transform 1 0 20720 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_177
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_193
timestamp 1698431365
transform 1 0 22960 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_201
timestamp 1698431365
transform 1 0 23856 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_203
timestamp 1698431365
transform 1 0 24080 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_218
timestamp 1698431365
transform 1 0 25760 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_226
timestamp 1698431365
transform 1 0 26656 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_234
timestamp 1698431365
transform 1 0 27552 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_236
timestamp 1698431365
transform 1 0 27776 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_247
timestamp 1698431365
transform 1 0 29008 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_255
timestamp 1698431365
transform 1 0 29904 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_287
timestamp 1698431365
transform 1 0 33488 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_299
timestamp 1698431365
transform 1 0 34832 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_312
timestamp 1698431365
transform 1 0 36288 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_314
timestamp 1698431365
transform 1 0 36512 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_322
timestamp 1698431365
transform 1 0 37408 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_329
timestamp 1698431365
transform 1 0 38192 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_338
timestamp 1698431365
transform 1 0 39200 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_354
timestamp 1698431365
transform 1 0 40992 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_358
timestamp 1698431365
transform 1 0 41440 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_387
timestamp 1698431365
transform 1 0 44688 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_391
timestamp 1698431365
transform 1 0 45136 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_416
timestamp 1698431365
transform 1 0 47936 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_424
timestamp 1698431365
transform 1 0 48832 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_428
timestamp 1698431365
transform 1 0 49280 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_438
timestamp 1698431365
transform 1 0 50400 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_447
timestamp 1698431365
transform 1 0 51408 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_451
timestamp 1698431365
transform 1 0 51856 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_457
timestamp 1698431365
transform 1 0 52528 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_477
timestamp 1698431365
transform 1 0 54768 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_485
timestamp 1698431365
transform 1 0 55664 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_14
timestamp 1698431365
transform 1 0 2912 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_18
timestamp 1698431365
transform 1 0 3360 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_22
timestamp 1698431365
transform 1 0 3808 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_39
timestamp 1698431365
transform 1 0 5712 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_55
timestamp 1698431365
transform 1 0 7504 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_62
timestamp 1698431365
transform 1 0 8288 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698431365
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_114
timestamp 1698431365
transform 1 0 14112 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_116
timestamp 1698431365
transform 1 0 14336 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_135
timestamp 1698431365
transform 1 0 16464 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_139
timestamp 1698431365
transform 1 0 16912 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_142
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_146
timestamp 1698431365
transform 1 0 17696 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_171
timestamp 1698431365
transform 1 0 20496 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_178
timestamp 1698431365
transform 1 0 21280 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_182
timestamp 1698431365
transform 1 0 21728 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_188
timestamp 1698431365
transform 1 0 22400 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_204
timestamp 1698431365
transform 1 0 24192 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_208
timestamp 1698431365
transform 1 0 24640 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_225
timestamp 1698431365
transform 1 0 26544 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_250
timestamp 1698431365
transform 1 0 29344 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_278
timestamp 1698431365
transform 1 0 32480 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_282
timestamp 1698431365
transform 1 0 32928 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_290
timestamp 1698431365
transform 1 0 33824 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_312
timestamp 1698431365
transform 1 0 36288 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_319
timestamp 1698431365
transform 1 0 37072 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_333
timestamp 1698431365
transform 1 0 38640 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_352
timestamp 1698431365
transform 1 0 40768 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_360
timestamp 1698431365
transform 1 0 41664 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_364
timestamp 1698431365
transform 1 0 42112 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_375
timestamp 1698431365
transform 1 0 43344 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_399
timestamp 1698431365
transform 1 0 46032 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_407
timestamp 1698431365
transform 1 0 46928 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_418
timestamp 1698431365
transform 1 0 48160 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_422
timestamp 1698431365
transform 1 0 48608 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_438
timestamp 1698431365
transform 1 0 50400 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_453
timestamp 1698431365
transform 1 0 52080 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_457
timestamp 1698431365
transform 1 0 52528 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_477
timestamp 1698431365
transform 1 0 54768 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_504
timestamp 1698431365
transform 1 0 57792 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_508
timestamp 1698431365
transform 1 0 58240 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_8
timestamp 1698431365
transform 1 0 2240 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_10
timestamp 1698431365
transform 1 0 2464 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_39
timestamp 1698431365
transform 1 0 5712 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_57
timestamp 1698431365
transform 1 0 7728 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_59
timestamp 1698431365
transform 1 0 7952 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_100
timestamp 1698431365
transform 1 0 12544 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_104
timestamp 1698431365
transform 1 0 12992 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_131
timestamp 1698431365
transform 1 0 16016 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_139
timestamp 1698431365
transform 1 0 16912 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_143
timestamp 1698431365
transform 1 0 17360 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_172
timestamp 1698431365
transform 1 0 20608 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_174
timestamp 1698431365
transform 1 0 20832 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_202
timestamp 1698431365
transform 1 0 23968 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_210
timestamp 1698431365
transform 1 0 24864 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_214
timestamp 1698431365
transform 1 0 25312 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_225
timestamp 1698431365
transform 1 0 26544 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_233
timestamp 1698431365
transform 1 0 27440 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_255
timestamp 1698431365
transform 1 0 29904 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_269
timestamp 1698431365
transform 1 0 31472 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_275
timestamp 1698431365
transform 1 0 32144 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_291
timestamp 1698431365
transform 1 0 33936 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_317
timestamp 1698431365
transform 1 0 36848 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_337
timestamp 1698431365
transform 1 0 39088 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_341
timestamp 1698431365
transform 1 0 39536 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_362
timestamp 1698431365
transform 1 0 41888 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_366
timestamp 1698431365
transform 1 0 42336 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_387
timestamp 1698431365
transform 1 0 44688 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_391
timestamp 1698431365
transform 1 0 45136 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_410
timestamp 1698431365
transform 1 0 47264 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_454
timestamp 1698431365
transform 1 0 52192 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_480
timestamp 1698431365
transform 1 0 55104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_506
timestamp 1698431365
transform 1 0 58016 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_508
timestamp 1698431365
transform 1 0 58240 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_2
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_30
timestamp 1698431365
transform 1 0 4704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_48
timestamp 1698431365
transform 1 0 6720 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_106
timestamp 1698431365
transform 1 0 13216 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_108
timestamp 1698431365
transform 1 0 13440 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_124
timestamp 1698431365
transform 1 0 15232 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_128
timestamp 1698431365
transform 1 0 15680 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_130
timestamp 1698431365
transform 1 0 15904 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_137
timestamp 1698431365
transform 1 0 16688 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_139
timestamp 1698431365
transform 1 0 16912 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_168
timestamp 1698431365
transform 1 0 20160 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_172
timestamp 1698431365
transform 1 0 20608 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_180
timestamp 1698431365
transform 1 0 21504 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_201
timestamp 1698431365
transform 1 0 23856 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_209
timestamp 1698431365
transform 1 0 24752 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_212
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_216
timestamp 1698431365
transform 1 0 25536 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_245
timestamp 1698431365
transform 1 0 28784 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_249
timestamp 1698431365
transform 1 0 29232 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_282
timestamp 1698431365
transform 1 0 32928 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_286
timestamp 1698431365
transform 1 0 33376 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_319
timestamp 1698431365
transform 1 0 37072 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_323
timestamp 1698431365
transform 1 0 37520 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_325
timestamp 1698431365
transform 1 0 37744 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_331
timestamp 1698431365
transform 1 0 38416 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_333
timestamp 1698431365
transform 1 0 38640 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_342
timestamp 1698431365
transform 1 0 39648 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_349
timestamp 1698431365
transform 1 0 40432 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_362
timestamp 1698431365
transform 1 0 41888 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_387
timestamp 1698431365
transform 1 0 44688 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_391
timestamp 1698431365
transform 1 0 45136 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_393
timestamp 1698431365
transform 1 0 45360 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_407
timestamp 1698431365
transform 1 0 46928 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_411
timestamp 1698431365
transform 1 0 47376 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_435
timestamp 1698431365
transform 1 0 50064 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_451
timestamp 1698431365
transform 1 0 51856 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_474
timestamp 1698431365
transform 1 0 54432 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_500
timestamp 1698431365
transform 1 0 57344 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_508
timestamp 1698431365
transform 1 0 58240 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_8
timestamp 1698431365
transform 1 0 2240 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_10
timestamp 1698431365
transform 1 0 2464 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698431365
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_53
timestamp 1698431365
transform 1 0 7280 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_69
timestamp 1698431365
transform 1 0 9072 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_72
timestamp 1698431365
transform 1 0 9408 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_92
timestamp 1698431365
transform 1 0 11648 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_107
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_122
timestamp 1698431365
transform 1 0 15008 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_124
timestamp 1698431365
transform 1 0 15232 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_200
timestamp 1698431365
transform 1 0 23744 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_204
timestamp 1698431365
transform 1 0 24192 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_252
timestamp 1698431365
transform 1 0 29568 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_256
timestamp 1698431365
transform 1 0 30016 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_260
timestamp 1698431365
transform 1 0 30464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_262
timestamp 1698431365
transform 1 0 30688 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_269
timestamp 1698431365
transform 1 0 31472 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_277
timestamp 1698431365
transform 1 0 32368 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_281
timestamp 1698431365
transform 1 0 32816 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698431365
transform 1 0 36176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_317
timestamp 1698431365
transform 1 0 36848 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_368
timestamp 1698431365
transform 1 0 42560 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_372
timestamp 1698431365
transform 1 0 43008 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_378
timestamp 1698431365
transform 1 0 43680 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_382
timestamp 1698431365
transform 1 0 44128 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_384
timestamp 1698431365
transform 1 0 44352 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_387
timestamp 1698431365
transform 1 0 44688 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_391
timestamp 1698431365
transform 1 0 45136 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_400
timestamp 1698431365
transform 1 0 46144 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_408
timestamp 1698431365
transform 1 0 47040 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_412
timestamp 1698431365
transform 1 0 47488 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_420
timestamp 1698431365
transform 1 0 48384 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_428
timestamp 1698431365
transform 1 0 49280 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_432
timestamp 1698431365
transform 1 0 49728 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_441
timestamp 1698431365
transform 1 0 50736 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_445
timestamp 1698431365
transform 1 0 51184 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_447
timestamp 1698431365
transform 1 0 51408 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_470
timestamp 1698431365
transform 1 0 53984 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_474
timestamp 1698431365
transform 1 0 54432 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_505
timestamp 1698431365
transform 1 0 57904 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_14
timestamp 1698431365
transform 1 0 2912 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_32
timestamp 1698431365
transform 1 0 4928 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_77
timestamp 1698431365
transform 1 0 9968 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_84
timestamp 1698431365
transform 1 0 10752 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_100
timestamp 1698431365
transform 1 0 12544 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_108
timestamp 1698431365
transform 1 0 13440 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_118
timestamp 1698431365
transform 1 0 14560 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_122
timestamp 1698431365
transform 1 0 15008 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_144
timestamp 1698431365
transform 1 0 17472 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_169
timestamp 1698431365
transform 1 0 20272 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_171
timestamp 1698431365
transform 1 0 20496 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_189
timestamp 1698431365
transform 1 0 22512 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_193
timestamp 1698431365
transform 1 0 22960 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_202
timestamp 1698431365
transform 1 0 23968 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_212
timestamp 1698431365
transform 1 0 25088 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_220
timestamp 1698431365
transform 1 0 25984 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_224
timestamp 1698431365
transform 1 0 26432 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_232
timestamp 1698431365
transform 1 0 27328 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_248
timestamp 1698431365
transform 1 0 29120 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_271
timestamp 1698431365
transform 1 0 31696 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_275
timestamp 1698431365
transform 1 0 32144 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_279
timestamp 1698431365
transform 1 0 32592 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_282
timestamp 1698431365
transform 1 0 32928 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_298
timestamp 1698431365
transform 1 0 34720 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_322
timestamp 1698431365
transform 1 0 37408 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_324
timestamp 1698431365
transform 1 0 37632 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_352
timestamp 1698431365
transform 1 0 40768 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_360
timestamp 1698431365
transform 1 0 41664 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_399
timestamp 1698431365
transform 1 0 46032 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_407
timestamp 1698431365
transform 1 0 46928 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_419
timestamp 1698431365
transform 1 0 48272 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_422
timestamp 1698431365
transform 1 0 48608 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_426
timestamp 1698431365
transform 1 0 49056 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_449
timestamp 1698431365
transform 1 0 51632 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_505
timestamp 1698431365
transform 1 0 57904 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_14
timestamp 1698431365
transform 1 0 2912 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_16
timestamp 1698431365
transform 1 0 3136 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_22
timestamp 1698431365
transform 1 0 3808 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_26
timestamp 1698431365
transform 1 0 4256 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_30
timestamp 1698431365
transform 1 0 4704 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698431365
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_37
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_39
timestamp 1698431365
transform 1 0 5712 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_57
timestamp 1698431365
transform 1 0 7728 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_61
timestamp 1698431365
transform 1 0 8176 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_63
timestamp 1698431365
transform 1 0 8400 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_98
timestamp 1698431365
transform 1 0 12320 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_102
timestamp 1698431365
transform 1 0 12768 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_104
timestamp 1698431365
transform 1 0 12992 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_107
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_115
timestamp 1698431365
transform 1 0 14224 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_117
timestamp 1698431365
transform 1 0 14448 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_150
timestamp 1698431365
transform 1 0 18144 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_177
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_189
timestamp 1698431365
transform 1 0 22512 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_205
timestamp 1698431365
transform 1 0 24304 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_213
timestamp 1698431365
transform 1 0 25200 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_247
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_255
timestamp 1698431365
transform 1 0 29904 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_270
timestamp 1698431365
transform 1 0 31584 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_278
timestamp 1698431365
transform 1 0 32480 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_303
timestamp 1698431365
transform 1 0 35280 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698431365
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_317
timestamp 1698431365
transform 1 0 36848 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_325
timestamp 1698431365
transform 1 0 37744 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_339
timestamp 1698431365
transform 1 0 39312 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_346
timestamp 1698431365
transform 1 0 40096 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_354
timestamp 1698431365
transform 1 0 40992 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_356
timestamp 1698431365
transform 1 0 41216 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_393
timestamp 1698431365
transform 1 0 45360 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_397
timestamp 1698431365
transform 1 0 45808 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_423
timestamp 1698431365
transform 1 0 48720 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_427
timestamp 1698431365
transform 1 0 49168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_442
timestamp 1698431365
transform 1 0 50848 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_470
timestamp 1698431365
transform 1 0 53984 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_478
timestamp 1698431365
transform 1 0 54880 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_501
timestamp 1698431365
transform 1 0 57456 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_14
timestamp 1698431365
transform 1 0 2912 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_18
timestamp 1698431365
transform 1 0 3360 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_32
timestamp 1698431365
transform 1 0 4928 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_40
timestamp 1698431365
transform 1 0 5824 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_53
timestamp 1698431365
transform 1 0 7280 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_69
timestamp 1698431365
transform 1 0 9072 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_72
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_93
timestamp 1698431365
transform 1 0 11760 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_97
timestamp 1698431365
transform 1 0 12208 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_125
timestamp 1698431365
transform 1 0 15344 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_142
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_144
timestamp 1698431365
transform 1 0 17472 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_153
timestamp 1698431365
transform 1 0 18480 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_178
timestamp 1698431365
transform 1 0 21280 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_182
timestamp 1698431365
transform 1 0 21728 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_192
timestamp 1698431365
transform 1 0 22848 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_201
timestamp 1698431365
transform 1 0 23856 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_209
timestamp 1698431365
transform 1 0 24752 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_220
timestamp 1698431365
transform 1 0 25984 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_241
timestamp 1698431365
transform 1 0 28336 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_249
timestamp 1698431365
transform 1 0 29232 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_255
timestamp 1698431365
transform 1 0 29904 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_267
timestamp 1698431365
transform 1 0 31248 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_275
timestamp 1698431365
transform 1 0 32144 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_279
timestamp 1698431365
transform 1 0 32592 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_282
timestamp 1698431365
transform 1 0 32928 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_290
timestamp 1698431365
transform 1 0 33824 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_294
timestamp 1698431365
transform 1 0 34272 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_308
timestamp 1698431365
transform 1 0 35840 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_324
timestamp 1698431365
transform 1 0 37632 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_349
timestamp 1698431365
transform 1 0 40432 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_357
timestamp 1698431365
transform 1 0 41328 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_361
timestamp 1698431365
transform 1 0 41776 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_369
timestamp 1698431365
transform 1 0 42672 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_392
timestamp 1698431365
transform 1 0 45248 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_400
timestamp 1698431365
transform 1 0 46144 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_418
timestamp 1698431365
transform 1 0 48160 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_427
timestamp 1698431365
transform 1 0 49168 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_447
timestamp 1698431365
transform 1 0 51408 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_455
timestamp 1698431365
transform 1 0 52304 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_476
timestamp 1698431365
transform 1 0 54656 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_480
timestamp 1698431365
transform 1 0 55104 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_483
timestamp 1698431365
transform 1 0 55440 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_487
timestamp 1698431365
transform 1 0 55888 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_489
timestamp 1698431365
transform 1 0 56112 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_504
timestamp 1698431365
transform 1 0 57792 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_508
timestamp 1698431365
transform 1 0 58240 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_2
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_24
timestamp 1698431365
transform 1 0 4032 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698431365
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_41
timestamp 1698431365
transform 1 0 5936 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_49
timestamp 1698431365
transform 1 0 6832 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_55
timestamp 1698431365
transform 1 0 7504 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_71
timestamp 1698431365
transform 1 0 9296 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_75
timestamp 1698431365
transform 1 0 9744 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_90
timestamp 1698431365
transform 1 0 11424 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_94
timestamp 1698431365
transform 1 0 11872 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_107
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_154
timestamp 1698431365
transform 1 0 18592 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_173
timestamp 1698431365
transform 1 0 20720 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_177
timestamp 1698431365
transform 1 0 21168 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_206
timestamp 1698431365
transform 1 0 24416 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_225
timestamp 1698431365
transform 1 0 26544 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_227
timestamp 1698431365
transform 1 0 26768 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_241
timestamp 1698431365
transform 1 0 28336 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_258
timestamp 1698431365
transform 1 0 30240 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_278
timestamp 1698431365
transform 1 0 32480 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_292
timestamp 1698431365
transform 1 0 34048 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_296
timestamp 1698431365
transform 1 0 34496 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_300
timestamp 1698431365
transform 1 0 34944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_302
timestamp 1698431365
transform 1 0 35168 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_314
timestamp 1698431365
transform 1 0 36512 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_332
timestamp 1698431365
transform 1 0 38528 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_334
timestamp 1698431365
transform 1 0 38752 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_341
timestamp 1698431365
transform 1 0 39536 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_367
timestamp 1698431365
transform 1 0 42448 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_383
timestamp 1698431365
transform 1 0 44240 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_387
timestamp 1698431365
transform 1 0 44688 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_402
timestamp 1698431365
transform 1 0 46368 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_410
timestamp 1698431365
transform 1 0 47264 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_429
timestamp 1698431365
transform 1 0 49392 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_433
timestamp 1698431365
transform 1 0 49840 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_435
timestamp 1698431365
transform 1 0 50064 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_482
timestamp 1698431365
transform 1 0 55328 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_26
timestamp 1698431365
transform 1 0 4256 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_51
timestamp 1698431365
transform 1 0 7056 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_69
timestamp 1698431365
transform 1 0 9072 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_78
timestamp 1698431365
transform 1 0 10080 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_94
timestamp 1698431365
transform 1 0 11872 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_101
timestamp 1698431365
transform 1 0 12656 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_121
timestamp 1698431365
transform 1 0 14896 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_142
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_180
timestamp 1698431365
transform 1 0 21504 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_204
timestamp 1698431365
transform 1 0 24192 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_208
timestamp 1698431365
transform 1 0 24640 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_212
timestamp 1698431365
transform 1 0 25088 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_224
timestamp 1698431365
transform 1 0 26432 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_232
timestamp 1698431365
transform 1 0 27328 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_236
timestamp 1698431365
transform 1 0 27776 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_262
timestamp 1698431365
transform 1 0 30688 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_278
timestamp 1698431365
transform 1 0 32480 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_326
timestamp 1698431365
transform 1 0 37856 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_330
timestamp 1698431365
transform 1 0 38304 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_349
timestamp 1698431365
transform 1 0 40432 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_352
timestamp 1698431365
transform 1 0 40768 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_370
timestamp 1698431365
transform 1 0 42784 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_374
timestamp 1698431365
transform 1 0 43232 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_405
timestamp 1698431365
transform 1 0 46704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_418
timestamp 1698431365
transform 1 0 48160 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_446
timestamp 1698431365
transform 1 0 51296 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_492
timestamp 1698431365
transform 1 0 56448 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_508
timestamp 1698431365
transform 1 0 58240 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_8
timestamp 1698431365
transform 1 0 2240 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_27
timestamp 1698431365
transform 1 0 4368 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_31
timestamp 1698431365
transform 1 0 4816 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_37
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_41
timestamp 1698431365
transform 1 0 5936 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_55
timestamp 1698431365
transform 1 0 7504 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_66
timestamp 1698431365
transform 1 0 8736 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_68
timestamp 1698431365
transform 1 0 8960 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_83
timestamp 1698431365
transform 1 0 10640 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_97
timestamp 1698431365
transform 1 0 12208 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_99
timestamp 1698431365
transform 1 0 12432 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_107
timestamp 1698431365
transform 1 0 13328 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_109
timestamp 1698431365
transform 1 0 13552 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_128
timestamp 1698431365
transform 1 0 15680 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_132
timestamp 1698431365
transform 1 0 16128 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_177
timestamp 1698431365
transform 1 0 21168 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_185
timestamp 1698431365
transform 1 0 22064 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_192
timestamp 1698431365
transform 1 0 22848 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_232
timestamp 1698431365
transform 1 0 27328 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_240
timestamp 1698431365
transform 1 0 28224 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_244
timestamp 1698431365
transform 1 0 28672 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_263
timestamp 1698431365
transform 1 0 30800 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_287
timestamp 1698431365
transform 1 0 33488 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_307
timestamp 1698431365
transform 1 0 35728 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_317
timestamp 1698431365
transform 1 0 36848 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_361
timestamp 1698431365
transform 1 0 41776 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_371
timestamp 1698431365
transform 1 0 42896 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_379
timestamp 1698431365
transform 1 0 43792 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_383
timestamp 1698431365
transform 1 0 44240 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_387
timestamp 1698431365
transform 1 0 44688 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_394
timestamp 1698431365
transform 1 0 45472 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_425
timestamp 1698431365
transform 1 0 48944 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_441
timestamp 1698431365
transform 1 0 50736 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_445
timestamp 1698431365
transform 1 0 51184 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_447
timestamp 1698431365
transform 1 0 51408 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_454
timestamp 1698431365
transform 1 0 52192 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_470
timestamp 1698431365
transform 1 0 53984 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_474
timestamp 1698431365
transform 1 0 54432 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_478
timestamp 1698431365
transform 1 0 54880 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_480
timestamp 1698431365
transform 1 0 55104 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_8
timestamp 1698431365
transform 1 0 2240 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_30
timestamp 1698431365
transform 1 0 4704 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_39
timestamp 1698431365
transform 1 0 5712 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_45
timestamp 1698431365
transform 1 0 6384 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_80
timestamp 1698431365
transform 1 0 10304 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_88
timestamp 1698431365
transform 1 0 11200 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_92
timestamp 1698431365
transform 1 0 11648 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_100
timestamp 1698431365
transform 1 0 12544 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_108
timestamp 1698431365
transform 1 0 13440 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_112
timestamp 1698431365
transform 1 0 13888 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_127
timestamp 1698431365
transform 1 0 15568 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_129
timestamp 1698431365
transform 1 0 15792 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_142
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_149
timestamp 1698431365
transform 1 0 18032 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_163
timestamp 1698431365
transform 1 0 19600 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_171
timestamp 1698431365
transform 1 0 20496 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_173
timestamp 1698431365
transform 1 0 20720 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_212
timestamp 1698431365
transform 1 0 25088 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_216
timestamp 1698431365
transform 1 0 25536 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_228
timestamp 1698431365
transform 1 0 26880 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_236
timestamp 1698431365
transform 1 0 27776 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_269
timestamp 1698431365
transform 1 0 31472 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_277
timestamp 1698431365
transform 1 0 32368 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_279
timestamp 1698431365
transform 1 0 32592 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_282
timestamp 1698431365
transform 1 0 32928 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_289
timestamp 1698431365
transform 1 0 33712 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_305
timestamp 1698431365
transform 1 0 35504 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_309
timestamp 1698431365
transform 1 0 35952 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_316
timestamp 1698431365
transform 1 0 36736 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_320
timestamp 1698431365
transform 1 0 37184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_324
timestamp 1698431365
transform 1 0 37632 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_326
timestamp 1698431365
transform 1 0 37856 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_329
timestamp 1698431365
transform 1 0 38192 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_337
timestamp 1698431365
transform 1 0 39088 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_348
timestamp 1698431365
transform 1 0 40320 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_393
timestamp 1698431365
transform 1 0 45360 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_397
timestamp 1698431365
transform 1 0 45808 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_413
timestamp 1698431365
transform 1 0 47600 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_417
timestamp 1698431365
transform 1 0 48048 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_419
timestamp 1698431365
transform 1 0 48272 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_437
timestamp 1698431365
transform 1 0 50288 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_462
timestamp 1698431365
transform 1 0 53088 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_492
timestamp 1698431365
transform 1 0 56448 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_508
timestamp 1698431365
transform 1 0 58240 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_32
timestamp 1698431365
transform 1 0 4928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698431365
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_60
timestamp 1698431365
transform 1 0 8064 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_67
timestamp 1698431365
transform 1 0 8848 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_97
timestamp 1698431365
transform 1 0 12208 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_99
timestamp 1698431365
transform 1 0 12432 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_136
timestamp 1698431365
transform 1 0 16576 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_144
timestamp 1698431365
transform 1 0 17472 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_148
timestamp 1698431365
transform 1 0 17920 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_158
timestamp 1698431365
transform 1 0 19040 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_160
timestamp 1698431365
transform 1 0 19264 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_217
timestamp 1698431365
transform 1 0 25648 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_221
timestamp 1698431365
transform 1 0 26096 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_239
timestamp 1698431365
transform 1 0 28112 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_243
timestamp 1698431365
transform 1 0 28560 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_247
timestamp 1698431365
transform 1 0 29008 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_301
timestamp 1698431365
transform 1 0 35056 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_305
timestamp 1698431365
transform 1 0 35504 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_355
timestamp 1698431365
transform 1 0 41104 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_363
timestamp 1698431365
transform 1 0 42000 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_366
timestamp 1698431365
transform 1 0 42336 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_374
timestamp 1698431365
transform 1 0 43232 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_381
timestamp 1698431365
transform 1 0 44016 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_402
timestamp 1698431365
transform 1 0 46368 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_406
timestamp 1698431365
transform 1 0 46816 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_438
timestamp 1698431365
transform 1 0 50400 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_2
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_6
timestamp 1698431365
transform 1 0 2016 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_10
timestamp 1698431365
transform 1 0 2464 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_17
timestamp 1698431365
transform 1 0 3248 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_21
timestamp 1698431365
transform 1 0 3696 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_41
timestamp 1698431365
transform 1 0 5936 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_45
timestamp 1698431365
transform 1 0 6384 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_51
timestamp 1698431365
transform 1 0 7056 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_58
timestamp 1698431365
transform 1 0 7840 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_62
timestamp 1698431365
transform 1 0 8288 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_72
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_95
timestamp 1698431365
transform 1 0 11984 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_97
timestamp 1698431365
transform 1 0 12208 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_100
timestamp 1698431365
transform 1 0 12544 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_104
timestamp 1698431365
transform 1 0 12992 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_129
timestamp 1698431365
transform 1 0 15792 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_133
timestamp 1698431365
transform 1 0 16240 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_142
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_151
timestamp 1698431365
transform 1 0 18256 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_157
timestamp 1698431365
transform 1 0 18928 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_193
timestamp 1698431365
transform 1 0 22960 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_203
timestamp 1698431365
transform 1 0 24080 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_209
timestamp 1698431365
transform 1 0 24752 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_212
timestamp 1698431365
transform 1 0 25088 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_220
timestamp 1698431365
transform 1 0 25984 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_222
timestamp 1698431365
transform 1 0 26208 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_241
timestamp 1698431365
transform 1 0 28336 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_245
timestamp 1698431365
transform 1 0 28784 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_253
timestamp 1698431365
transform 1 0 29680 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_259
timestamp 1698431365
transform 1 0 30352 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_263
timestamp 1698431365
transform 1 0 30800 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_279
timestamp 1698431365
transform 1 0 32592 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_282
timestamp 1698431365
transform 1 0 32928 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_314
timestamp 1698431365
transform 1 0 36512 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_318
timestamp 1698431365
transform 1 0 36960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_320
timestamp 1698431365
transform 1 0 37184 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_329
timestamp 1698431365
transform 1 0 38192 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_331
timestamp 1698431365
transform 1 0 38416 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_334
timestamp 1698431365
transform 1 0 38752 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_338
timestamp 1698431365
transform 1 0 39200 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_346
timestamp 1698431365
transform 1 0 40096 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_367
timestamp 1698431365
transform 1 0 42448 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_383
timestamp 1698431365
transform 1 0 44240 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_408
timestamp 1698431365
transform 1 0 47040 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_416
timestamp 1698431365
transform 1 0 47936 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_428
timestamp 1698431365
transform 1 0 49280 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_444
timestamp 1698431365
transform 1 0 51072 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_461
timestamp 1698431365
transform 1 0 52976 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_463
timestamp 1698431365
transform 1 0 53200 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_492
timestamp 1698431365
transform 1 0 56448 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_508
timestamp 1698431365
transform 1 0 58240 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_8
timestamp 1698431365
transform 1 0 2240 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_23
timestamp 1698431365
transform 1 0 3920 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_30
timestamp 1698431365
transform 1 0 4704 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698431365
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_43
timestamp 1698431365
transform 1 0 6160 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_45
timestamp 1698431365
transform 1 0 6384 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_65
timestamp 1698431365
transform 1 0 8624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_69
timestamp 1698431365
transform 1 0 9072 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_73
timestamp 1698431365
transform 1 0 9520 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_103
timestamp 1698431365
transform 1 0 12880 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_107
timestamp 1698431365
transform 1 0 13328 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_123
timestamp 1698431365
transform 1 0 15120 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_127
timestamp 1698431365
transform 1 0 15568 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_171
timestamp 1698431365
transform 1 0 20496 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_223
timestamp 1698431365
transform 1 0 26320 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_257
timestamp 1698431365
transform 1 0 30128 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_288
timestamp 1698431365
transform 1 0 33600 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_304
timestamp 1698431365
transform 1 0 35392 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_308
timestamp 1698431365
transform 1 0 35840 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_332
timestamp 1698431365
transform 1 0 38528 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_336
timestamp 1698431365
transform 1 0 38976 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_338
timestamp 1698431365
transform 1 0 39200 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_368
timestamp 1698431365
transform 1 0 42560 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_372
timestamp 1698431365
transform 1 0 43008 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_380
timestamp 1698431365
transform 1 0 43904 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_382
timestamp 1698431365
transform 1 0 44128 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_416
timestamp 1698431365
transform 1 0 47936 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_448
timestamp 1698431365
transform 1 0 51520 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_452
timestamp 1698431365
transform 1 0 51968 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_454
timestamp 1698431365
transform 1 0 52192 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_461
timestamp 1698431365
transform 1 0 52976 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_465
timestamp 1698431365
transform 1 0 53424 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_481
timestamp 1698431365
transform 1 0 55216 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_2
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_6
timestamp 1698431365
transform 1 0 2016 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_32
timestamp 1698431365
transform 1 0 4928 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_39
timestamp 1698431365
transform 1 0 5712 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_43
timestamp 1698431365
transform 1 0 6160 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_63
timestamp 1698431365
transform 1 0 8400 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_67
timestamp 1698431365
transform 1 0 8848 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_69
timestamp 1698431365
transform 1 0 9072 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_72
timestamp 1698431365
transform 1 0 9408 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_103
timestamp 1698431365
transform 1 0 12880 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_105
timestamp 1698431365
transform 1 0 13104 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_108
timestamp 1698431365
transform 1 0 13440 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_112
timestamp 1698431365
transform 1 0 13888 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_128
timestamp 1698431365
transform 1 0 15680 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_132
timestamp 1698431365
transform 1 0 16128 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_147
timestamp 1698431365
transform 1 0 17808 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_163
timestamp 1698431365
transform 1 0 19600 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_167
timestamp 1698431365
transform 1 0 20048 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_212
timestamp 1698431365
transform 1 0 25088 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_237
timestamp 1698431365
transform 1 0 27888 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_263
timestamp 1698431365
transform 1 0 30800 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_267
timestamp 1698431365
transform 1 0 31248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_269
timestamp 1698431365
transform 1 0 31472 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_276
timestamp 1698431365
transform 1 0 32256 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_297
timestamp 1698431365
transform 1 0 34608 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_301
timestamp 1698431365
transform 1 0 35056 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_333
timestamp 1698431365
transform 1 0 38640 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_337
timestamp 1698431365
transform 1 0 39088 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_339
timestamp 1698431365
transform 1 0 39312 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_342
timestamp 1698431365
transform 1 0 39648 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_346
timestamp 1698431365
transform 1 0 40096 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_358
timestamp 1698431365
transform 1 0 41440 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_364
timestamp 1698431365
transform 1 0 42112 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_368
timestamp 1698431365
transform 1 0 42560 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_370
timestamp 1698431365
transform 1 0 42784 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_373
timestamp 1698431365
transform 1 0 43120 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_406
timestamp 1698431365
transform 1 0 46816 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_410
timestamp 1698431365
transform 1 0 47264 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_418
timestamp 1698431365
transform 1 0 48160 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_437
timestamp 1698431365
transform 1 0 50288 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_453
timestamp 1698431365
transform 1 0 52080 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_461
timestamp 1698431365
transform 1 0 52976 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_463
timestamp 1698431365
transform 1 0 53200 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_492
timestamp 1698431365
transform 1 0 56448 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_508
timestamp 1698431365
transform 1 0 58240 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_2
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_10
timestamp 1698431365
transform 1 0 2464 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_14
timestamp 1698431365
transform 1 0 2912 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_25
timestamp 1698431365
transform 1 0 4144 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698431365
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_50
timestamp 1698431365
transform 1 0 6944 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_81
timestamp 1698431365
transform 1 0 10416 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_107
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_134
timestamp 1698431365
transform 1 0 16352 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_136
timestamp 1698431365
transform 1 0 16576 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_147
timestamp 1698431365
transform 1 0 17808 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_162
timestamp 1698431365
transform 1 0 19488 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_170
timestamp 1698431365
transform 1 0 20384 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_174
timestamp 1698431365
transform 1 0 20832 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_182
timestamp 1698431365
transform 1 0 21728 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_184
timestamp 1698431365
transform 1 0 21952 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_225
timestamp 1698431365
transform 1 0 26544 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_244
timestamp 1698431365
transform 1 0 28672 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_268
timestamp 1698431365
transform 1 0 31360 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_272
timestamp 1698431365
transform 1 0 31808 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_276
timestamp 1698431365
transform 1 0 32256 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_280
timestamp 1698431365
transform 1 0 32704 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_282
timestamp 1698431365
transform 1 0 32928 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_311
timestamp 1698431365
transform 1 0 36176 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_395
timestamp 1698431365
transform 1 0 45584 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_399
timestamp 1698431365
transform 1 0 46032 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_434
timestamp 1698431365
transform 1 0 49952 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_450
timestamp 1698431365
transform 1 0 51744 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_454
timestamp 1698431365
transform 1 0 52192 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_457
timestamp 1698431365
transform 1 0 52528 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_473
timestamp 1698431365
transform 1 0 54320 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_2
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_6
timestamp 1698431365
transform 1 0 2016 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_18
timestamp 1698431365
transform 1 0 3360 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_36
timestamp 1698431365
transform 1 0 5376 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_44
timestamp 1698431365
transform 1 0 6272 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_48
timestamp 1698431365
transform 1 0 6720 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_63
timestamp 1698431365
transform 1 0 8400 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_67
timestamp 1698431365
transform 1 0 8848 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_69
timestamp 1698431365
transform 1 0 9072 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_72
timestamp 1698431365
transform 1 0 9408 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_82
timestamp 1698431365
transform 1 0 10528 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_84
timestamp 1698431365
transform 1 0 10752 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_91
timestamp 1698431365
transform 1 0 11536 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_112
timestamp 1698431365
transform 1 0 13888 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_116
timestamp 1698431365
transform 1 0 14336 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_137
timestamp 1698431365
transform 1 0 16688 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_139
timestamp 1698431365
transform 1 0 16912 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_166
timestamp 1698431365
transform 1 0 19936 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_168
timestamp 1698431365
transform 1 0 20160 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_198
timestamp 1698431365
transform 1 0 23520 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_202
timestamp 1698431365
transform 1 0 23968 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_206
timestamp 1698431365
transform 1 0 24416 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_241
timestamp 1698431365
transform 1 0 28336 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_272
timestamp 1698431365
transform 1 0 31808 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_276
timestamp 1698431365
transform 1 0 32256 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_340
timestamp 1698431365
transform 1 0 39424 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_402
timestamp 1698431365
transform 1 0 46368 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_406
timestamp 1698431365
transform 1 0 46816 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_414
timestamp 1698431365
transform 1 0 47712 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_418
timestamp 1698431365
transform 1 0 48160 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_422
timestamp 1698431365
transform 1 0 48608 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_454
timestamp 1698431365
transform 1 0 52192 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_462
timestamp 1698431365
transform 1 0 53088 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_492
timestamp 1698431365
transform 1 0 56448 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_508
timestamp 1698431365
transform 1 0 58240 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_2
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_37
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_70
timestamp 1698431365
transform 1 0 9184 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_78
timestamp 1698431365
transform 1 0 10080 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_82
timestamp 1698431365
transform 1 0 10528 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_84
timestamp 1698431365
transform 1 0 10752 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_119
timestamp 1698431365
transform 1 0 14672 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_138
timestamp 1698431365
transform 1 0 16800 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_142
timestamp 1698431365
transform 1 0 17248 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_160
timestamp 1698431365
transform 1 0 19264 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_168
timestamp 1698431365
transform 1 0 20160 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_172
timestamp 1698431365
transform 1 0 20608 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_174
timestamp 1698431365
transform 1 0 20832 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_177
timestamp 1698431365
transform 1 0 21168 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_220
timestamp 1698431365
transform 1 0 25984 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_247
timestamp 1698431365
transform 1 0 29008 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_312
timestamp 1698431365
transform 1 0 36288 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_314
timestamp 1698431365
transform 1 0 36512 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_333
timestamp 1698431365
transform 1 0 38640 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_404
timestamp 1698431365
transform 1 0 46592 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_434
timestamp 1698431365
transform 1 0 49952 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_450
timestamp 1698431365
transform 1 0 51744 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_454
timestamp 1698431365
transform 1 0 52192 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_52
timestamp 1698431365
transform 1 0 7168 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_56
timestamp 1698431365
transform 1 0 7616 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_72
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_76
timestamp 1698431365
transform 1 0 9856 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_120
timestamp 1698431365
transform 1 0 14784 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_134
timestamp 1698431365
transform 1 0 16352 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_138
timestamp 1698431365
transform 1 0 16800 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_142
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_146
timestamp 1698431365
transform 1 0 17696 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_156
timestamp 1698431365
transform 1 0 18816 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_162
timestamp 1698431365
transform 1 0 19488 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_178
timestamp 1698431365
transform 1 0 21280 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_196
timestamp 1698431365
transform 1 0 23296 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_198
timestamp 1698431365
transform 1 0 23520 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_201
timestamp 1698431365
transform 1 0 23856 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_218
timestamp 1698431365
transform 1 0 25760 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_275
timestamp 1698431365
transform 1 0 32144 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_279
timestamp 1698431365
transform 1 0 32592 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_282
timestamp 1698431365
transform 1 0 32928 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_314
timestamp 1698431365
transform 1 0 36512 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_322
timestamp 1698431365
transform 1 0 37408 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_345
timestamp 1698431365
transform 1 0 39984 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_349
timestamp 1698431365
transform 1 0 40432 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_352
timestamp 1698431365
transform 1 0 40768 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_354
timestamp 1698431365
transform 1 0 40992 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_384
timestamp 1698431365
transform 1 0 44352 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_414
timestamp 1698431365
transform 1 0 47712 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_418
timestamp 1698431365
transform 1 0 48160 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_422
timestamp 1698431365
transform 1 0 48608 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_454
timestamp 1698431365
transform 1 0 52192 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_462
timestamp 1698431365
transform 1 0 53088 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_492
timestamp 1698431365
transform 1 0 56448 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_508
timestamp 1698431365
transform 1 0 58240 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_42
timestamp 1698431365
transform 1 0 6048 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_66
timestamp 1698431365
transform 1 0 8736 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_70
timestamp 1698431365
transform 1 0 9184 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_89
timestamp 1698431365
transform 1 0 11312 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_107
timestamp 1698431365
transform 1 0 13328 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_111
timestamp 1698431365
transform 1 0 13776 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_174
timestamp 1698431365
transform 1 0 20832 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_242
timestamp 1698431365
transform 1 0 28448 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_244
timestamp 1698431365
transform 1 0 28672 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_260
timestamp 1698431365
transform 1 0 30464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_262
timestamp 1698431365
transform 1 0 30688 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_312
timestamp 1698431365
transform 1 0 36288 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_314
timestamp 1698431365
transform 1 0 36512 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_317
timestamp 1698431365
transform 1 0 36848 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_325
timestamp 1698431365
transform 1 0 37744 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_329
timestamp 1698431365
transform 1 0 38192 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_331
timestamp 1698431365
transform 1 0 38416 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_384
timestamp 1698431365
transform 1 0 44352 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_387
timestamp 1698431365
transform 1 0 44688 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_399
timestamp 1698431365
transform 1 0 46032 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_413
timestamp 1698431365
transform 1 0 47600 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_445
timestamp 1698431365
transform 1 0 51184 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_453
timestamp 1698431365
transform 1 0 52080 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_457
timestamp 1698431365
transform 1 0 52528 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_473
timestamp 1698431365
transform 1 0 54320 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_28
timestamp 1698431365
transform 1 0 4480 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_32
timestamp 1698431365
transform 1 0 4928 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_36
timestamp 1698431365
transform 1 0 5376 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_68
timestamp 1698431365
transform 1 0 8960 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_72
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_76
timestamp 1698431365
transform 1 0 9856 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_78
timestamp 1698431365
transform 1 0 10080 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_87
timestamp 1698431365
transform 1 0 11088 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_89
timestamp 1698431365
transform 1 0 11312 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_102
timestamp 1698431365
transform 1 0 12768 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_106
timestamp 1698431365
transform 1 0 13216 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_130
timestamp 1698431365
transform 1 0 15904 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_138
timestamp 1698431365
transform 1 0 16800 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_142
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_150
timestamp 1698431365
transform 1 0 18144 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_167
timestamp 1698431365
transform 1 0 20048 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_174
timestamp 1698431365
transform 1 0 20832 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_178
timestamp 1698431365
transform 1 0 21280 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_182
timestamp 1698431365
transform 1 0 21728 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_186
timestamp 1698431365
transform 1 0 22176 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_188
timestamp 1698431365
transform 1 0 22400 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_212
timestamp 1698431365
transform 1 0 25088 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_216
timestamp 1698431365
transform 1 0 25536 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_225
timestamp 1698431365
transform 1 0 26544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_290
timestamp 1698431365
transform 1 0 33824 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_326
timestamp 1698431365
transform 1 0 37856 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_330
timestamp 1698431365
transform 1 0 38304 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_340
timestamp 1698431365
transform 1 0 39424 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_405
timestamp 1698431365
transform 1 0 46704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_409
timestamp 1698431365
transform 1 0 47152 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_413
timestamp 1698431365
transform 1 0 47600 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_417
timestamp 1698431365
transform 1 0 48048 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_419
timestamp 1698431365
transform 1 0 48272 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_422
timestamp 1698431365
transform 1 0 48608 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_454
timestamp 1698431365
transform 1 0 52192 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_462
timestamp 1698431365
transform 1 0 53088 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_492
timestamp 1698431365
transform 1 0 56448 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_508
timestamp 1698431365
transform 1 0 58240 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_28
timestamp 1698431365
transform 1 0 4480 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_32
timestamp 1698431365
transform 1 0 4928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698431365
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_37
timestamp 1698431365
transform 1 0 5488 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_53
timestamp 1698431365
transform 1 0 7280 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_61
timestamp 1698431365
transform 1 0 8176 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_63
timestamp 1698431365
transform 1 0 8400 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_93
timestamp 1698431365
transform 1 0 11760 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_104
timestamp 1698431365
transform 1 0 12992 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_112
timestamp 1698431365
transform 1 0 13888 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_116
timestamp 1698431365
transform 1 0 14336 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_120
timestamp 1698431365
transform 1 0 14784 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_126
timestamp 1698431365
transform 1 0 15456 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_134
timestamp 1698431365
transform 1 0 16352 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_138
timestamp 1698431365
transform 1 0 16800 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_172
timestamp 1698431365
transform 1 0 20608 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_174
timestamp 1698431365
transform 1 0 20832 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_227
timestamp 1698431365
transform 1 0 26768 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_231
timestamp 1698431365
transform 1 0 27216 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_235
timestamp 1698431365
transform 1 0 27664 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_253
timestamp 1698431365
transform 1 0 29680 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_257
timestamp 1698431365
transform 1 0 30128 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_266
timestamp 1698431365
transform 1 0 31136 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_270
timestamp 1698431365
transform 1 0 31584 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_285
timestamp 1698431365
transform 1 0 33264 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_322
timestamp 1698431365
transform 1 0 37408 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_330
timestamp 1698431365
transform 1 0 38304 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_332
timestamp 1698431365
transform 1 0 38528 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_350
timestamp 1698431365
transform 1 0 40544 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_371
timestamp 1698431365
transform 1 0 42896 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_387
timestamp 1698431365
transform 1 0 44688 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_391
timestamp 1698431365
transform 1 0 45136 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_395
timestamp 1698431365
transform 1 0 45584 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_399
timestamp 1698431365
transform 1 0 46032 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_403
timestamp 1698431365
transform 1 0 46480 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_435
timestamp 1698431365
transform 1 0 50064 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_451
timestamp 1698431365
transform 1 0 51856 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_457
timestamp 1698431365
transform 1 0 52528 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_473
timestamp 1698431365
transform 1 0 54320 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_481
timestamp 1698431365
transform 1 0 55216 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_28
timestamp 1698431365
transform 1 0 4480 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_60
timestamp 1698431365
transform 1 0 8064 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_68
timestamp 1698431365
transform 1 0 8960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_101
timestamp 1698431365
transform 1 0 12656 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_136
timestamp 1698431365
transform 1 0 16576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_142
timestamp 1698431365
transform 1 0 17248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_144
timestamp 1698431365
transform 1 0 17472 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_205
timestamp 1698431365
transform 1 0 24304 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_209
timestamp 1698431365
transform 1 0 24752 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_212
timestamp 1698431365
transform 1 0 25088 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_244
timestamp 1698431365
transform 1 0 28672 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_255
timestamp 1698431365
transform 1 0 29904 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_282
timestamp 1698431365
transform 1 0 32928 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_284
timestamp 1698431365
transform 1 0 33152 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_287
timestamp 1698431365
transform 1 0 33488 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_295
timestamp 1698431365
transform 1 0 34384 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_304
timestamp 1698431365
transform 1 0 35392 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_312
timestamp 1698431365
transform 1 0 36288 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_314
timestamp 1698431365
transform 1 0 36512 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_317
timestamp 1698431365
transform 1 0 36848 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_321
timestamp 1698431365
transform 1 0 37296 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_329
timestamp 1698431365
transform 1 0 38192 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_338
timestamp 1698431365
transform 1 0 39200 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_340
timestamp 1698431365
transform 1 0 39424 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_348
timestamp 1698431365
transform 1 0 40320 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_428
timestamp 1698431365
transform 1 0 49280 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_460
timestamp 1698431365
transform 1 0 52864 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_476
timestamp 1698431365
transform 1 0 54656 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_484
timestamp 1698431365
transform 1 0 55552 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_488
timestamp 1698431365
transform 1 0 56000 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_492
timestamp 1698431365
transform 1 0 56448 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_500
timestamp 1698431365
transform 1 0 57344 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_28
timestamp 1698431365
transform 1 0 4480 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_32
timestamp 1698431365
transform 1 0 4928 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698431365
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_37
timestamp 1698431365
transform 1 0 5488 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_69
timestamp 1698431365
transform 1 0 9072 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_85
timestamp 1698431365
transform 1 0 10864 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_93
timestamp 1698431365
transform 1 0 11760 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_100
timestamp 1698431365
transform 1 0 12544 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_104
timestamp 1698431365
transform 1 0 12992 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_107
timestamp 1698431365
transform 1 0 13328 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_126
timestamp 1698431365
transform 1 0 15456 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_130
timestamp 1698431365
transform 1 0 15904 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_138
timestamp 1698431365
transform 1 0 16800 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_177
timestamp 1698431365
transform 1 0 21168 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_185
timestamp 1698431365
transform 1 0 22064 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_189
timestamp 1698431365
transform 1 0 22512 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_198
timestamp 1698431365
transform 1 0 23520 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_202
timestamp 1698431365
transform 1 0 23968 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_255
timestamp 1698431365
transform 1 0 29904 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_267
timestamp 1698431365
transform 1 0 31248 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_298
timestamp 1698431365
transform 1 0 34720 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_302
timestamp 1698431365
transform 1 0 35168 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_310
timestamp 1698431365
transform 1 0 36064 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_314
timestamp 1698431365
transform 1 0 36512 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_317
timestamp 1698431365
transform 1 0 36848 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_327
timestamp 1698431365
transform 1 0 37968 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_331
timestamp 1698431365
transform 1 0 38416 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_335
timestamp 1698431365
transform 1 0 38864 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_366
timestamp 1698431365
transform 1 0 42336 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_370
timestamp 1698431365
transform 1 0 42784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_374
timestamp 1698431365
transform 1 0 43232 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_383
timestamp 1698431365
transform 1 0 44240 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_405
timestamp 1698431365
transform 1 0 46704 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_409
timestamp 1698431365
transform 1 0 47152 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_413
timestamp 1698431365
transform 1 0 47600 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_445
timestamp 1698431365
transform 1 0 51184 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_453
timestamp 1698431365
transform 1 0 52080 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_457
timestamp 1698431365
transform 1 0 52528 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_473
timestamp 1698431365
transform 1 0 54320 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_481
timestamp 1698431365
transform 1 0 55216 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_2
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_34
timestamp 1698431365
transform 1 0 5152 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_42
timestamp 1698431365
transform 1 0 6048 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_46
timestamp 1698431365
transform 1 0 6496 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_56
timestamp 1698431365
transform 1 0 7616 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_72
timestamp 1698431365
transform 1 0 9408 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_76
timestamp 1698431365
transform 1 0 9856 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_78
timestamp 1698431365
transform 1 0 10080 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_87
timestamp 1698431365
transform 1 0 11088 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_91
timestamp 1698431365
transform 1 0 11536 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_116
timestamp 1698431365
transform 1 0 14336 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_131
timestamp 1698431365
transform 1 0 16016 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_135
timestamp 1698431365
transform 1 0 16464 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_139
timestamp 1698431365
transform 1 0 16912 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_142
timestamp 1698431365
transform 1 0 17248 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_162
timestamp 1698431365
transform 1 0 19488 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_170
timestamp 1698431365
transform 1 0 20384 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_196
timestamp 1698431365
transform 1 0 23296 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_204
timestamp 1698431365
transform 1 0 24192 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_208
timestamp 1698431365
transform 1 0 24640 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_220
timestamp 1698431365
transform 1 0 25984 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_228
timestamp 1698431365
transform 1 0 26880 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_232
timestamp 1698431365
transform 1 0 27328 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_248
timestamp 1698431365
transform 1 0 29120 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_252
timestamp 1698431365
transform 1 0 29568 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_266
timestamp 1698431365
transform 1 0 31136 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_270
timestamp 1698431365
transform 1 0 31584 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_278
timestamp 1698431365
transform 1 0 32480 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_295
timestamp 1698431365
transform 1 0 34384 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_336
timestamp 1698431365
transform 1 0 38976 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_345
timestamp 1698431365
transform 1 0 39984 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_349
timestamp 1698431365
transform 1 0 40432 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_357
timestamp 1698431365
transform 1 0 41328 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_361
timestamp 1698431365
transform 1 0 41776 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_365
timestamp 1698431365
transform 1 0 42224 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_367
timestamp 1698431365
transform 1 0 42448 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_392
timestamp 1698431365
transform 1 0 45248 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_396
timestamp 1698431365
transform 1 0 45696 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_400
timestamp 1698431365
transform 1 0 46144 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_416
timestamp 1698431365
transform 1 0 47936 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_422
timestamp 1698431365
transform 1 0 48608 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_486
timestamp 1698431365
transform 1 0 55776 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_492
timestamp 1698431365
transform 1 0 56448 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_500
timestamp 1698431365
transform 1 0 57344 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_2
timestamp 1698431365
transform 1 0 1568 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_18
timestamp 1698431365
transform 1 0 3360 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698431365
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_37
timestamp 1698431365
transform 1 0 5488 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_41
timestamp 1698431365
transform 1 0 5936 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_71
timestamp 1698431365
transform 1 0 9296 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_75
timestamp 1698431365
transform 1 0 9744 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_77
timestamp 1698431365
transform 1 0 9968 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_90
timestamp 1698431365
transform 1 0 11424 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_126
timestamp 1698431365
transform 1 0 15456 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_130
timestamp 1698431365
transform 1 0 15904 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_136
timestamp 1698431365
transform 1 0 16576 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_153
timestamp 1698431365
transform 1 0 18480 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_157
timestamp 1698431365
transform 1 0 18928 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_165
timestamp 1698431365
transform 1 0 19824 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_167
timestamp 1698431365
transform 1 0 20048 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_177
timestamp 1698431365
transform 1 0 21168 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_194
timestamp 1698431365
transform 1 0 23072 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_198
timestamp 1698431365
transform 1 0 23520 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_234
timestamp 1698431365
transform 1 0 27552 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_238
timestamp 1698431365
transform 1 0 28000 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_242
timestamp 1698431365
transform 1 0 28448 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_244
timestamp 1698431365
transform 1 0 28672 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_267
timestamp 1698431365
transform 1 0 31248 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_271
timestamp 1698431365
transform 1 0 31696 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_273
timestamp 1698431365
transform 1 0 31920 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_282
timestamp 1698431365
transform 1 0 32928 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_290
timestamp 1698431365
transform 1 0 33824 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_292
timestamp 1698431365
transform 1 0 34048 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_307
timestamp 1698431365
transform 1 0 35728 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_314
timestamp 1698431365
transform 1 0 36512 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_317
timestamp 1698431365
transform 1 0 36848 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_326
timestamp 1698431365
transform 1 0 37856 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_340
timestamp 1698431365
transform 1 0 39424 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_344
timestamp 1698431365
transform 1 0 39872 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_376
timestamp 1698431365
transform 1 0 43456 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_379
timestamp 1698431365
transform 1 0 43792 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_383
timestamp 1698431365
transform 1 0 44240 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_387
timestamp 1698431365
transform 1 0 44688 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_391
timestamp 1698431365
transform 1 0 45136 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_457
timestamp 1698431365
transform 1 0 52528 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_473
timestamp 1698431365
transform 1 0 54320 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_2
timestamp 1698431365
transform 1 0 1568 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_10
timestamp 1698431365
transform 1 0 2464 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_37
timestamp 1698431365
transform 1 0 5488 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_45
timestamp 1698431365
transform 1 0 6384 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_72
timestamp 1698431365
transform 1 0 9408 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_93
timestamp 1698431365
transform 1 0 11760 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_101
timestamp 1698431365
transform 1 0 12656 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_107
timestamp 1698431365
transform 1 0 13328 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_120
timestamp 1698431365
transform 1 0 14784 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_124
timestamp 1698431365
transform 1 0 15232 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_150
timestamp 1698431365
transform 1 0 18144 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_167
timestamp 1698431365
transform 1 0 20048 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_171
timestamp 1698431365
transform 1 0 20496 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_174
timestamp 1698431365
transform 1 0 20832 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_192
timestamp 1698431365
transform 1 0 22848 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_208
timestamp 1698431365
transform 1 0 24640 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_212
timestamp 1698431365
transform 1 0 25088 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_220
timestamp 1698431365
transform 1 0 25984 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_224
timestamp 1698431365
transform 1 0 26432 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_232
timestamp 1698431365
transform 1 0 27328 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_236
timestamp 1698431365
transform 1 0 27776 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_238
timestamp 1698431365
transform 1 0 28000 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_261
timestamp 1698431365
transform 1 0 30576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_265
timestamp 1698431365
transform 1 0 31024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_279
timestamp 1698431365
transform 1 0 32592 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_292
timestamp 1698431365
transform 1 0 34048 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_294
timestamp 1698431365
transform 1 0 34272 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_313
timestamp 1698431365
transform 1 0 36400 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_323
timestamp 1698431365
transform 1 0 37520 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_327
timestamp 1698431365
transform 1 0 37968 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_339
timestamp 1698431365
transform 1 0 39312 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_347
timestamp 1698431365
transform 1 0 40208 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_349
timestamp 1698431365
transform 1 0 40432 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_376
timestamp 1698431365
transform 1 0 43456 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_396
timestamp 1698431365
transform 1 0 45696 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_400
timestamp 1698431365
transform 1 0 46144 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_416
timestamp 1698431365
transform 1 0 47936 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_422
timestamp 1698431365
transform 1 0 48608 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_486
timestamp 1698431365
transform 1 0 55776 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_492
timestamp 1698431365
transform 1 0 56448 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_500
timestamp 1698431365
transform 1 0 57344 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_33
timestamp 1698431365
transform 1 0 5040 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_37
timestamp 1698431365
transform 1 0 5488 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_54
timestamp 1698431365
transform 1 0 7392 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_73
timestamp 1698431365
transform 1 0 9520 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_86
timestamp 1698431365
transform 1 0 10976 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_94
timestamp 1698431365
transform 1 0 11872 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_98
timestamp 1698431365
transform 1 0 12320 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_120
timestamp 1698431365
transform 1 0 14784 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_128
timestamp 1698431365
transform 1 0 15680 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_132
timestamp 1698431365
transform 1 0 16128 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_134
timestamp 1698431365
transform 1 0 16352 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_150
timestamp 1698431365
transform 1 0 18144 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_158
timestamp 1698431365
transform 1 0 19040 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698431365
transform 1 0 20496 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_177
timestamp 1698431365
transform 1 0 21168 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_217
timestamp 1698431365
transform 1 0 25648 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_265
timestamp 1698431365
transform 1 0 31024 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_282
timestamp 1698431365
transform 1 0 32928 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_286
timestamp 1698431365
transform 1 0 33376 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_288
timestamp 1698431365
transform 1 0 33600 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_314
timestamp 1698431365
transform 1 0 36512 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_317
timestamp 1698431365
transform 1 0 36848 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_349
timestamp 1698431365
transform 1 0 40432 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_370
timestamp 1698431365
transform 1 0 42784 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_406
timestamp 1698431365
transform 1 0 46816 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_408
timestamp 1698431365
transform 1 0 47040 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_419
timestamp 1698431365
transform 1 0 48272 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_451
timestamp 1698431365
transform 1 0 51856 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_457
timestamp 1698431365
transform 1 0 52528 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_473
timestamp 1698431365
transform 1 0 54320 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_481
timestamp 1698431365
transform 1 0 55216 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_2
timestamp 1698431365
transform 1 0 1568 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_15
timestamp 1698431365
transform 1 0 3024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_31
timestamp 1698431365
transform 1 0 4816 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_54
timestamp 1698431365
transform 1 0 7392 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_76
timestamp 1698431365
transform 1 0 9856 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_95
timestamp 1698431365
transform 1 0 11984 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_151
timestamp 1698431365
transform 1 0 18256 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_159
timestamp 1698431365
transform 1 0 19152 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_188
timestamp 1698431365
transform 1 0 22400 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_200
timestamp 1698431365
transform 1 0 23744 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_212
timestamp 1698431365
transform 1 0 25088 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_230
timestamp 1698431365
transform 1 0 27104 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_234
timestamp 1698431365
transform 1 0 27552 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_258
timestamp 1698431365
transform 1 0 30240 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_262
timestamp 1698431365
transform 1 0 30688 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_270
timestamp 1698431365
transform 1 0 31584 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_282
timestamp 1698431365
transform 1 0 32928 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_312
timestamp 1698431365
transform 1 0 36288 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_316
timestamp 1698431365
transform 1 0 36736 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_323
timestamp 1698431365
transform 1 0 37520 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_335
timestamp 1698431365
transform 1 0 38864 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_341
timestamp 1698431365
transform 1 0 39536 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_345
timestamp 1698431365
transform 1 0 39984 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_349
timestamp 1698431365
transform 1 0 40432 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_352
timestamp 1698431365
transform 1 0 40768 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_406
timestamp 1698431365
transform 1 0 46816 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_432
timestamp 1698431365
transform 1 0 49728 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_463
timestamp 1698431365
transform 1 0 53200 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_477
timestamp 1698431365
transform 1 0 54768 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_485
timestamp 1698431365
transform 1 0 55664 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_489
timestamp 1698431365
transform 1 0 56112 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_492
timestamp 1698431365
transform 1 0 56448 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_500
timestamp 1698431365
transform 1 0 57344 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_2
timestamp 1698431365
transform 1 0 1568 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_10
timestamp 1698431365
transform 1 0 2464 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_37
timestamp 1698431365
transform 1 0 5488 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_54
timestamp 1698431365
transform 1 0 7392 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_61
timestamp 1698431365
transform 1 0 8176 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_67
timestamp 1698431365
transform 1 0 8848 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_71
timestamp 1698431365
transform 1 0 9296 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_78
timestamp 1698431365
transform 1 0 10080 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_98
timestamp 1698431365
transform 1 0 12320 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_102
timestamp 1698431365
transform 1 0 12768 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_104
timestamp 1698431365
transform 1 0 12992 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_107
timestamp 1698431365
transform 1 0 13328 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_124
timestamp 1698431365
transform 1 0 15232 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_128
timestamp 1698431365
transform 1 0 15680 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_132
timestamp 1698431365
transform 1 0 16128 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_157
timestamp 1698431365
transform 1 0 18928 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_173
timestamp 1698431365
transform 1 0 20720 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_177
timestamp 1698431365
transform 1 0 21168 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_193
timestamp 1698431365
transform 1 0 22960 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_201
timestamp 1698431365
transform 1 0 23856 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_207
timestamp 1698431365
transform 1 0 24528 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_227
timestamp 1698431365
transform 1 0 26768 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_243
timestamp 1698431365
transform 1 0 28560 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_253
timestamp 1698431365
transform 1 0 29680 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_257
timestamp 1698431365
transform 1 0 30128 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_274
timestamp 1698431365
transform 1 0 32032 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_290
timestamp 1698431365
transform 1 0 33824 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_294
timestamp 1698431365
transform 1 0 34272 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_307
timestamp 1698431365
transform 1 0 35728 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_323
timestamp 1698431365
transform 1 0 37520 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_325
timestamp 1698431365
transform 1 0 37744 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_346
timestamp 1698431365
transform 1 0 40096 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_350
timestamp 1698431365
transform 1 0 40544 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_358
timestamp 1698431365
transform 1 0 41440 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_360
timestamp 1698431365
transform 1 0 41664 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_380
timestamp 1698431365
transform 1 0 43904 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_384
timestamp 1698431365
transform 1 0 44352 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_387
timestamp 1698431365
transform 1 0 44688 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_403
timestamp 1698431365
transform 1 0 46480 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_407
timestamp 1698431365
transform 1 0 46928 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_411
timestamp 1698431365
transform 1 0 47376 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_450
timestamp 1698431365
transform 1 0 51744 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_454
timestamp 1698431365
transform 1 0 52192 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_457
timestamp 1698431365
transform 1 0 52528 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_461
timestamp 1698431365
transform 1 0 52976 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_482
timestamp 1698431365
transform 1 0 55328 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_490
timestamp 1698431365
transform 1 0 56224 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_494
timestamp 1698431365
transform 1 0 56672 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_25
timestamp 1698431365
transform 1 0 4144 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_33
timestamp 1698431365
transform 1 0 5040 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_37
timestamp 1698431365
transform 1 0 5488 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_62
timestamp 1698431365
transform 1 0 8288 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_77
timestamp 1698431365
transform 1 0 9968 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_90
timestamp 1698431365
transform 1 0 11424 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_98
timestamp 1698431365
transform 1 0 12320 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_102
timestamp 1698431365
transform 1 0 12768 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_126
timestamp 1698431365
transform 1 0 15456 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_153
timestamp 1698431365
transform 1 0 18480 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_161
timestamp 1698431365
transform 1 0 19376 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_170
timestamp 1698431365
transform 1 0 20384 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_178
timestamp 1698431365
transform 1 0 21280 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_180
timestamp 1698431365
transform 1 0 21504 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_193
timestamp 1698431365
transform 1 0 22960 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_212
timestamp 1698431365
transform 1 0 25088 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_216
timestamp 1698431365
transform 1 0 25536 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_258
timestamp 1698431365
transform 1 0 30240 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_260
timestamp 1698431365
transform 1 0 30464 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_267
timestamp 1698431365
transform 1 0 31248 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_294
timestamp 1698431365
transform 1 0 34272 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_310
timestamp 1698431365
transform 1 0 36064 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_318
timestamp 1698431365
transform 1 0 36960 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_340
timestamp 1698431365
transform 1 0 39424 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_344
timestamp 1698431365
transform 1 0 39872 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_348
timestamp 1698431365
transform 1 0 40320 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_352
timestamp 1698431365
transform 1 0 40768 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_354
timestamp 1698431365
transform 1 0 40992 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_376
timestamp 1698431365
transform 1 0 43456 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_380
timestamp 1698431365
transform 1 0 43904 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_408
timestamp 1698431365
transform 1 0 47040 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_416
timestamp 1698431365
transform 1 0 47936 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_432
timestamp 1698431365
transform 1 0 49728 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_436
timestamp 1698431365
transform 1 0 50176 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_469
timestamp 1698431365
transform 1 0 53872 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_485
timestamp 1698431365
transform 1 0 55664 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_489
timestamp 1698431365
transform 1 0 56112 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_492
timestamp 1698431365
transform 1 0 56448 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_496
timestamp 1698431365
transform 1 0 56896 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_499
timestamp 1698431365
transform 1 0 57232 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_2
timestamp 1698431365
transform 1 0 1568 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_27
timestamp 1698431365
transform 1 0 4368 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_37
timestamp 1698431365
transform 1 0 5488 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_60
timestamp 1698431365
transform 1 0 8064 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_70
timestamp 1698431365
transform 1 0 9184 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_72
timestamp 1698431365
transform 1 0 9408 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_79
timestamp 1698431365
transform 1 0 10192 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_88
timestamp 1698431365
transform 1 0 11200 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_104
timestamp 1698431365
transform 1 0 12992 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_131
timestamp 1698431365
transform 1 0 16016 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_164
timestamp 1698431365
transform 1 0 19712 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_172
timestamp 1698431365
transform 1 0 20608 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_174
timestamp 1698431365
transform 1 0 20832 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_177
timestamp 1698431365
transform 1 0 21168 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_179
timestamp 1698431365
transform 1 0 21392 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_193
timestamp 1698431365
transform 1 0 22960 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_209
timestamp 1698431365
transform 1 0 24752 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_218
timestamp 1698431365
transform 1 0 25760 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_247
timestamp 1698431365
transform 1 0 29008 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_251
timestamp 1698431365
transform 1 0 29456 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_255
timestamp 1698431365
transform 1 0 29904 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_257
timestamp 1698431365
transform 1 0 30128 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_260
timestamp 1698431365
transform 1 0 30464 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_268
timestamp 1698431365
transform 1 0 31360 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_270
timestamp 1698431365
transform 1 0 31584 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_284
timestamp 1698431365
transform 1 0 33152 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_292
timestamp 1698431365
transform 1 0 34048 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_309
timestamp 1698431365
transform 1 0 35952 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_313
timestamp 1698431365
transform 1 0 36400 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_344
timestamp 1698431365
transform 1 0 39872 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_348
timestamp 1698431365
transform 1 0 40320 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_373
timestamp 1698431365
transform 1 0 43120 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_377
timestamp 1698431365
transform 1 0 43568 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_379
timestamp 1698431365
transform 1 0 43792 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_400
timestamp 1698431365
transform 1 0 46144 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_404
timestamp 1698431365
transform 1 0 46592 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_406
timestamp 1698431365
transform 1 0 46816 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_442
timestamp 1698431365
transform 1 0 50848 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_462
timestamp 1698431365
transform 1 0 53088 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_466
timestamp 1698431365
transform 1 0 53536 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_474
timestamp 1698431365
transform 1 0 54432 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_476
timestamp 1698431365
transform 1 0 54656 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_485
timestamp 1698431365
transform 1 0 55664 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_8
timestamp 1698431365
transform 1 0 2240 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_12
timestamp 1698431365
transform 1 0 2688 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_20
timestamp 1698431365
transform 1 0 3584 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_22
timestamp 1698431365
transform 1 0 3808 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_46
timestamp 1698431365
transform 1 0 6496 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_54
timestamp 1698431365
transform 1 0 7392 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_58
timestamp 1698431365
transform 1 0 7840 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_69
timestamp 1698431365
transform 1 0 9072 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_72
timestamp 1698431365
transform 1 0 9408 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_96
timestamp 1698431365
transform 1 0 12096 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_98
timestamp 1698431365
transform 1 0 12320 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_123
timestamp 1698431365
transform 1 0 15120 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_131
timestamp 1698431365
transform 1 0 16016 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_133
timestamp 1698431365
transform 1 0 16240 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_139
timestamp 1698431365
transform 1 0 16912 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_190
timestamp 1698431365
transform 1 0 22624 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_192
timestamp 1698431365
transform 1 0 22848 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_207
timestamp 1698431365
transform 1 0 24528 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_209
timestamp 1698431365
transform 1 0 24752 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_228
timestamp 1698431365
transform 1 0 26880 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_255
timestamp 1698431365
transform 1 0 29904 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_275
timestamp 1698431365
transform 1 0 32144 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_279
timestamp 1698431365
transform 1 0 32592 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_282
timestamp 1698431365
transform 1 0 32928 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_286
timestamp 1698431365
transform 1 0 33376 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_302
timestamp 1698431365
transform 1 0 35168 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_306
timestamp 1698431365
transform 1 0 35616 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_338
timestamp 1698431365
transform 1 0 39200 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_342
timestamp 1698431365
transform 1 0 39648 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_370
timestamp 1698431365
transform 1 0 42784 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_379
timestamp 1698431365
transform 1 0 43792 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_387
timestamp 1698431365
transform 1 0 44688 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_399
timestamp 1698431365
transform 1 0 46032 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_407
timestamp 1698431365
transform 1 0 46928 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_409
timestamp 1698431365
transform 1 0 47152 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_419
timestamp 1698431365
transform 1 0 48272 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_433
timestamp 1698431365
transform 1 0 49840 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_437
timestamp 1698431365
transform 1 0 50288 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_452
timestamp 1698431365
transform 1 0 51968 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_460
timestamp 1698431365
transform 1 0 52864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_462
timestamp 1698431365
transform 1 0 53088 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_475
timestamp 1698431365
transform 1 0 54544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_487
timestamp 1698431365
transform 1 0 55888 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_489
timestamp 1698431365
transform 1 0 56112 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_492
timestamp 1698431365
transform 1 0 56448 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_500
timestamp 1698431365
transform 1 0 57344 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_2
timestamp 1698431365
transform 1 0 1568 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_10
timestamp 1698431365
transform 1 0 2464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_19
timestamp 1698431365
transform 1 0 3472 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_21
timestamp 1698431365
transform 1 0 3696 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_37
timestamp 1698431365
transform 1 0 5488 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_41
timestamp 1698431365
transform 1 0 5936 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_54
timestamp 1698431365
transform 1 0 7392 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_58
timestamp 1698431365
transform 1 0 7840 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_72
timestamp 1698431365
transform 1 0 9408 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_78
timestamp 1698431365
transform 1 0 10080 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_80
timestamp 1698431365
transform 1 0 10304 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_93
timestamp 1698431365
transform 1 0 11760 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698431365
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_107
timestamp 1698431365
transform 1 0 13328 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_111
timestamp 1698431365
transform 1 0 13776 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_118
timestamp 1698431365
transform 1 0 14560 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_134
timestamp 1698431365
transform 1 0 16352 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_160
timestamp 1698431365
transform 1 0 19264 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_169
timestamp 1698431365
transform 1 0 20272 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_173
timestamp 1698431365
transform 1 0 20720 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_177
timestamp 1698431365
transform 1 0 21168 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_208
timestamp 1698431365
transform 1 0 24640 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_230
timestamp 1698431365
transform 1 0 27104 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_238
timestamp 1698431365
transform 1 0 28000 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_242
timestamp 1698431365
transform 1 0 28448 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_244
timestamp 1698431365
transform 1 0 28672 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_256
timestamp 1698431365
transform 1 0 30016 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_260
timestamp 1698431365
transform 1 0 30464 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_264
timestamp 1698431365
transform 1 0 30912 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_282
timestamp 1698431365
transform 1 0 32928 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_291
timestamp 1698431365
transform 1 0 33936 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_293
timestamp 1698431365
transform 1 0 34160 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_312
timestamp 1698431365
transform 1 0 36288 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_314
timestamp 1698431365
transform 1 0 36512 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_317
timestamp 1698431365
transform 1 0 36848 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_328
timestamp 1698431365
transform 1 0 38080 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_332
timestamp 1698431365
transform 1 0 38528 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_352
timestamp 1698431365
transform 1 0 40768 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_362
timestamp 1698431365
transform 1 0 41888 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_370
timestamp 1698431365
transform 1 0 42784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_372
timestamp 1698431365
transform 1 0 43008 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_378
timestamp 1698431365
transform 1 0 43680 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_382
timestamp 1698431365
transform 1 0 44128 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_384
timestamp 1698431365
transform 1 0 44352 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_387
timestamp 1698431365
transform 1 0 44688 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_395
timestamp 1698431365
transform 1 0 45584 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_403
timestamp 1698431365
transform 1 0 46480 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_407
timestamp 1698431365
transform 1 0 46928 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_409
timestamp 1698431365
transform 1 0 47152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_439
timestamp 1698431365
transform 1 0 50512 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_441
timestamp 1698431365
transform 1 0 50736 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_444
timestamp 1698431365
transform 1 0 51072 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_452
timestamp 1698431365
transform 1 0 51968 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_454
timestamp 1698431365
transform 1 0 52192 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_457
timestamp 1698431365
transform 1 0 52528 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_487
timestamp 1698431365
transform 1 0 55888 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_495
timestamp 1698431365
transform 1 0 56784 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_499
timestamp 1698431365
transform 1 0 57232 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_2
timestamp 1698431365
transform 1 0 1568 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_34
timestamp 1698431365
transform 1 0 5152 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_38
timestamp 1698431365
transform 1 0 5600 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_40
timestamp 1698431365
transform 1 0 5824 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_49
timestamp 1698431365
transform 1 0 6832 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_63
timestamp 1698431365
transform 1 0 8400 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_67
timestamp 1698431365
transform 1 0 8848 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_69
timestamp 1698431365
transform 1 0 9072 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_72
timestamp 1698431365
transform 1 0 9408 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_88
timestamp 1698431365
transform 1 0 11200 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_96
timestamp 1698431365
transform 1 0 12096 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_100
timestamp 1698431365
transform 1 0 12544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_102
timestamp 1698431365
transform 1 0 12768 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_124
timestamp 1698431365
transform 1 0 15232 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_138
timestamp 1698431365
transform 1 0 16800 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_175
timestamp 1698431365
transform 1 0 20944 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_177
timestamp 1698431365
transform 1 0 21168 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_193
timestamp 1698431365
transform 1 0 22960 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_200
timestamp 1698431365
transform 1 0 23744 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_204
timestamp 1698431365
transform 1 0 24192 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_212
timestamp 1698431365
transform 1 0 25088 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_229
timestamp 1698431365
transform 1 0 26992 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_237
timestamp 1698431365
transform 1 0 27888 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_239
timestamp 1698431365
transform 1 0 28112 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_251
timestamp 1698431365
transform 1 0 29456 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_275
timestamp 1698431365
transform 1 0 32144 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_279
timestamp 1698431365
transform 1 0 32592 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_282
timestamp 1698431365
transform 1 0 32928 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_286
timestamp 1698431365
transform 1 0 33376 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_306
timestamp 1698431365
transform 1 0 35616 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_310
timestamp 1698431365
transform 1 0 36064 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_336
timestamp 1698431365
transform 1 0 38976 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_358
timestamp 1698431365
transform 1 0 41440 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_396
timestamp 1698431365
transform 1 0 45696 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_400
timestamp 1698431365
transform 1 0 46144 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_408
timestamp 1698431365
transform 1 0 47040 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_436
timestamp 1698431365
transform 1 0 50176 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_438
timestamp 1698431365
transform 1 0 50400 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_472
timestamp 1698431365
transform 1 0 54208 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_488
timestamp 1698431365
transform 1 0 56000 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_492
timestamp 1698431365
transform 1 0 56448 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_496
timestamp 1698431365
transform 1 0 56896 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_499
timestamp 1698431365
transform 1 0 57232 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_8
timestamp 1698431365
transform 1 0 2240 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_30
timestamp 1698431365
transform 1 0 4704 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698431365
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_37
timestamp 1698431365
transform 1 0 5488 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_45
timestamp 1698431365
transform 1 0 6384 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_49
timestamp 1698431365
transform 1 0 6832 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_56
timestamp 1698431365
transform 1 0 7616 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_58
timestamp 1698431365
transform 1 0 7840 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_77
timestamp 1698431365
transform 1 0 9968 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_83
timestamp 1698431365
transform 1 0 10640 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_87
timestamp 1698431365
transform 1 0 11088 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_107
timestamp 1698431365
transform 1 0 13328 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_137
timestamp 1698431365
transform 1 0 16688 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_145
timestamp 1698431365
transform 1 0 17584 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_192
timestamp 1698431365
transform 1 0 22848 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_202
timestamp 1698431365
transform 1 0 23968 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_224
timestamp 1698431365
transform 1 0 26432 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_240
timestamp 1698431365
transform 1 0 28224 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_244
timestamp 1698431365
transform 1 0 28672 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_260
timestamp 1698431365
transform 1 0 30464 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_267
timestamp 1698431365
transform 1 0 31248 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_295
timestamp 1698431365
transform 1 0 34384 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_303
timestamp 1698431365
transform 1 0 35280 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_307
timestamp 1698431365
transform 1 0 35728 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_337
timestamp 1698431365
transform 1 0 39088 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_345
timestamp 1698431365
transform 1 0 39984 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_347
timestamp 1698431365
transform 1 0 40208 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_366
timestamp 1698431365
transform 1 0 42336 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_379
timestamp 1698431365
transform 1 0 43792 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_405
timestamp 1698431365
transform 1 0 46704 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_413
timestamp 1698431365
transform 1 0 47600 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_417
timestamp 1698431365
transform 1 0 48048 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_424
timestamp 1698431365
transform 1 0 48832 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_432
timestamp 1698431365
transform 1 0 49728 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_439
timestamp 1698431365
transform 1 0 50512 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_441
timestamp 1698431365
transform 1 0 50736 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_465
timestamp 1698431365
transform 1 0 53424 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_469
timestamp 1698431365
transform 1 0 53872 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_471
timestamp 1698431365
transform 1 0 54096 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_477
timestamp 1698431365
transform 1 0 54768 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_481
timestamp 1698431365
transform 1 0 55216 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_500
timestamp 1698431365
transform 1 0 57344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_502
timestamp 1698431365
transform 1 0 57568 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_2
timestamp 1698431365
transform 1 0 1568 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_6
timestamp 1698431365
transform 1 0 2016 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_10
timestamp 1698431365
transform 1 0 2464 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_29
timestamp 1698431365
transform 1 0 4592 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_37
timestamp 1698431365
transform 1 0 5488 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_53
timestamp 1698431365
transform 1 0 7280 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_61
timestamp 1698431365
transform 1 0 8176 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_68
timestamp 1698431365
transform 1 0 8960 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_101
timestamp 1698431365
transform 1 0 12656 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_105
timestamp 1698431365
transform 1 0 13104 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_120
timestamp 1698431365
transform 1 0 14784 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_128
timestamp 1698431365
transform 1 0 15680 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_139
timestamp 1698431365
transform 1 0 16912 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_170
timestamp 1698431365
transform 1 0 20384 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_186
timestamp 1698431365
transform 1 0 22176 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_194
timestamp 1698431365
transform 1 0 23072 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_205
timestamp 1698431365
transform 1 0 24304 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698431365
transform 1 0 24752 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_225
timestamp 1698431365
transform 1 0 26544 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_257
timestamp 1698431365
transform 1 0 30128 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_261
timestamp 1698431365
transform 1 0 30576 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_265
timestamp 1698431365
transform 1 0 31024 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_298
timestamp 1698431365
transform 1 0 34720 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_302
timestamp 1698431365
transform 1 0 35168 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_328
timestamp 1698431365
transform 1 0 38080 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_336
timestamp 1698431365
transform 1 0 38976 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_340
timestamp 1698431365
transform 1 0 39424 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_342
timestamp 1698431365
transform 1 0 39648 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_352
timestamp 1698431365
transform 1 0 40768 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_354
timestamp 1698431365
transform 1 0 40992 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_368
timestamp 1698431365
transform 1 0 42560 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_372
timestamp 1698431365
transform 1 0 43008 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_397
timestamp 1698431365
transform 1 0 45808 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_399
timestamp 1698431365
transform 1 0 46032 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_413
timestamp 1698431365
transform 1 0 47600 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_417
timestamp 1698431365
transform 1 0 48048 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_419
timestamp 1698431365
transform 1 0 48272 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_422
timestamp 1698431365
transform 1 0 48608 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_424
timestamp 1698431365
transform 1 0 48832 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_500
timestamp 1698431365
transform 1 0 57344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_502
timestamp 1698431365
transform 1 0 57568 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_2
timestamp 1698431365
transform 1 0 1568 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_25
timestamp 1698431365
transform 1 0 4144 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_37
timestamp 1698431365
transform 1 0 5488 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_39
timestamp 1698431365
transform 1 0 5712 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_93
timestamp 1698431365
transform 1 0 11760 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_101
timestamp 1698431365
transform 1 0 12656 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_107
timestamp 1698431365
transform 1 0 13328 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_111
timestamp 1698431365
transform 1 0 13776 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_123
timestamp 1698431365
transform 1 0 15120 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_131
timestamp 1698431365
transform 1 0 16016 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_148
timestamp 1698431365
transform 1 0 17920 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_150
timestamp 1698431365
transform 1 0 18144 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_163
timestamp 1698431365
transform 1 0 19600 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_171
timestamp 1698431365
transform 1 0 20496 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_177
timestamp 1698431365
transform 1 0 21168 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_194
timestamp 1698431365
transform 1 0 23072 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_198
timestamp 1698431365
transform 1 0 23520 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_221
timestamp 1698431365
transform 1 0 26096 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_237
timestamp 1698431365
transform 1 0 27888 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_260
timestamp 1698431365
transform 1 0 30464 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_276
timestamp 1698431365
transform 1 0 32256 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_296
timestamp 1698431365
transform 1 0 34496 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_306
timestamp 1698431365
transform 1 0 35616 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_314
timestamp 1698431365
transform 1 0 36512 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_317
timestamp 1698431365
transform 1 0 36848 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_333
timestamp 1698431365
transform 1 0 38640 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_335
timestamp 1698431365
transform 1 0 38864 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_343
timestamp 1698431365
transform 1 0 39760 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_372
timestamp 1698431365
transform 1 0 43008 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_384
timestamp 1698431365
transform 1 0 44352 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_387
timestamp 1698431365
transform 1 0 44688 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_391
timestamp 1698431365
transform 1 0 45136 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_395
timestamp 1698431365
transform 1 0 45584 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_397
timestamp 1698431365
transform 1 0 45808 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_405
timestamp 1698431365
transform 1 0 46704 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_441
timestamp 1698431365
transform 1 0 50736 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_443
timestamp 1698431365
transform 1 0 50960 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_452
timestamp 1698431365
transform 1 0 51968 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_454
timestamp 1698431365
transform 1 0 52192 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_457
timestamp 1698431365
transform 1 0 52528 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_461
timestamp 1698431365
transform 1 0 52976 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_483
timestamp 1698431365
transform 1 0 55440 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_490
timestamp 1698431365
transform 1 0 56224 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_494
timestamp 1698431365
transform 1 0 56672 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_8
timestamp 1698431365
transform 1 0 2240 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_10
timestamp 1698431365
transform 1 0 2464 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_17
timestamp 1698431365
transform 1 0 3248 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_19
timestamp 1698431365
transform 1 0 3472 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_33
timestamp 1698431365
transform 1 0 5040 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_37
timestamp 1698431365
transform 1 0 5488 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_53
timestamp 1698431365
transform 1 0 7280 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_61
timestamp 1698431365
transform 1 0 8176 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_68
timestamp 1698431365
transform 1 0 8960 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_72
timestamp 1698431365
transform 1 0 9408 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_90
timestamp 1698431365
transform 1 0 11424 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_92
timestamp 1698431365
transform 1 0 11648 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_99
timestamp 1698431365
transform 1 0 12432 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_101
timestamp 1698431365
transform 1 0 12656 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_133
timestamp 1698431365
transform 1 0 16240 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_142
timestamp 1698431365
transform 1 0 17248 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_205
timestamp 1698431365
transform 1 0 24304 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_209
timestamp 1698431365
transform 1 0 24752 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_218
timestamp 1698431365
transform 1 0 25760 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_234
timestamp 1698431365
transform 1 0 27552 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_242
timestamp 1698431365
transform 1 0 28448 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_257
timestamp 1698431365
transform 1 0 30128 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_261
timestamp 1698431365
transform 1 0 30576 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_265
timestamp 1698431365
transform 1 0 31024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_267
timestamp 1698431365
transform 1 0 31248 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_276
timestamp 1698431365
transform 1 0 32256 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_282
timestamp 1698431365
transform 1 0 32928 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_290
timestamp 1698431365
transform 1 0 33824 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_308
timestamp 1698431365
transform 1 0 35840 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_348
timestamp 1698431365
transform 1 0 40320 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_367
timestamp 1698431365
transform 1 0 42448 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_369
timestamp 1698431365
transform 1 0 42672 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_376
timestamp 1698431365
transform 1 0 43456 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_384
timestamp 1698431365
transform 1 0 44352 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_410
timestamp 1698431365
transform 1 0 47264 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_418
timestamp 1698431365
transform 1 0 48160 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_442
timestamp 1698431365
transform 1 0 50848 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_457
timestamp 1698431365
transform 1 0 52528 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_489
timestamp 1698431365
transform 1 0 56112 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_492
timestamp 1698431365
transform 1 0 56448 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_500
timestamp 1698431365
transform 1 0 57344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_502
timestamp 1698431365
transform 1 0 57568 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_505
timestamp 1698431365
transform 1 0 57904 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_10
timestamp 1698431365
transform 1 0 2464 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_17
timestamp 1698431365
transform 1 0 3248 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_52
timestamp 1698431365
transform 1 0 7168 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_60
timestamp 1698431365
transform 1 0 8064 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_67
timestamp 1698431365
transform 1 0 8848 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_71
timestamp 1698431365
transform 1 0 9296 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_107
timestamp 1698431365
transform 1 0 13328 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_109
timestamp 1698431365
transform 1 0 13552 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_121
timestamp 1698431365
transform 1 0 14896 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_137
timestamp 1698431365
transform 1 0 16688 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_145
timestamp 1698431365
transform 1 0 17584 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_147
timestamp 1698431365
transform 1 0 17808 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_161
timestamp 1698431365
transform 1 0 19376 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_169
timestamp 1698431365
transform 1 0 20272 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_173
timestamp 1698431365
transform 1 0 20720 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_177
timestamp 1698431365
transform 1 0 21168 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_181
timestamp 1698431365
transform 1 0 21616 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_202
timestamp 1698431365
transform 1 0 23968 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_234
timestamp 1698431365
transform 1 0 27552 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_271
timestamp 1698431365
transform 1 0 31696 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_294
timestamp 1698431365
transform 1 0 34272 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_302
timestamp 1698431365
transform 1 0 35168 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_311
timestamp 1698431365
transform 1 0 36176 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_317
timestamp 1698431365
transform 1 0 36848 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_324
timestamp 1698431365
transform 1 0 37632 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_332
timestamp 1698431365
transform 1 0 38528 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_360
timestamp 1698431365
transform 1 0 41664 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_381
timestamp 1698431365
transform 1 0 44016 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_387
timestamp 1698431365
transform 1 0 44688 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_395
timestamp 1698431365
transform 1 0 45584 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_408
timestamp 1698431365
transform 1 0 47040 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_412
timestamp 1698431365
transform 1 0 47488 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_428
timestamp 1698431365
transform 1 0 49280 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_438
timestamp 1698431365
transform 1 0 50400 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_457
timestamp 1698431365
transform 1 0 52528 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_477
timestamp 1698431365
transform 1 0 54768 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_486
timestamp 1698431365
transform 1 0 55776 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_502
timestamp 1698431365
transform 1 0 57568 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_506
timestamp 1698431365
transform 1 0 58016 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_508
timestamp 1698431365
transform 1 0 58240 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_2
timestamp 1698431365
transform 1 0 1568 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_4
timestamp 1698431365
transform 1 0 1792 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_45
timestamp 1698431365
transform 1 0 6384 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_49
timestamp 1698431365
transform 1 0 6832 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_61
timestamp 1698431365
transform 1 0 8176 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_69
timestamp 1698431365
transform 1 0 9072 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_72
timestamp 1698431365
transform 1 0 9408 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_76
timestamp 1698431365
transform 1 0 9856 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_121
timestamp 1698431365
transform 1 0 14896 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_137
timestamp 1698431365
transform 1 0 16688 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_139
timestamp 1698431365
transform 1 0 16912 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_166
timestamp 1698431365
transform 1 0 19936 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_170
timestamp 1698431365
transform 1 0 20384 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_172
timestamp 1698431365
transform 1 0 20608 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_201
timestamp 1698431365
transform 1 0 23856 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_209
timestamp 1698431365
transform 1 0 24752 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_212
timestamp 1698431365
transform 1 0 25088 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_228
timestamp 1698431365
transform 1 0 26880 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_236
timestamp 1698431365
transform 1 0 27776 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_240
timestamp 1698431365
transform 1 0 28224 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_261
timestamp 1698431365
transform 1 0 30576 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_265
timestamp 1698431365
transform 1 0 31024 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_274
timestamp 1698431365
transform 1 0 32032 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_278
timestamp 1698431365
transform 1 0 32480 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_295
timestamp 1698431365
transform 1 0 34384 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_299
timestamp 1698431365
transform 1 0 34832 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_329
timestamp 1698431365
transform 1 0 38192 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_345
timestamp 1698431365
transform 1 0 39984 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_349
timestamp 1698431365
transform 1 0 40432 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_358
timestamp 1698431365
transform 1 0 41440 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_366
timestamp 1698431365
transform 1 0 42336 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_390
timestamp 1698431365
transform 1 0 45024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_394
timestamp 1698431365
transform 1 0 45472 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_414
timestamp 1698431365
transform 1 0 47712 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_418
timestamp 1698431365
transform 1 0 48160 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_422
timestamp 1698431365
transform 1 0 48608 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_438
timestamp 1698431365
transform 1 0 50400 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_442
timestamp 1698431365
transform 1 0 50848 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_444
timestamp 1698431365
transform 1 0 51072 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_486
timestamp 1698431365
transform 1 0 55776 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_492
timestamp 1698431365
transform 1 0 56448 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_508
timestamp 1698431365
transform 1 0 58240 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_26
timestamp 1698431365
transform 1 0 4256 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_28
timestamp 1698431365
transform 1 0 4480 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_49
timestamp 1698431365
transform 1 0 6832 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_55
timestamp 1698431365
transform 1 0 7504 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_57
timestamp 1698431365
transform 1 0 7728 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_64
timestamp 1698431365
transform 1 0 8512 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_76
timestamp 1698431365
transform 1 0 9856 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_85
timestamp 1698431365
transform 1 0 10864 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_93
timestamp 1698431365
transform 1 0 11760 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_97
timestamp 1698431365
transform 1 0 12208 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_99
timestamp 1698431365
transform 1 0 12432 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_142
timestamp 1698431365
transform 1 0 17248 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_168
timestamp 1698431365
transform 1 0 20160 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_172
timestamp 1698431365
transform 1 0 20608 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_174
timestamp 1698431365
transform 1 0 20832 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_189
timestamp 1698431365
transform 1 0 22512 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_204
timestamp 1698431365
transform 1 0 24192 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_236
timestamp 1698431365
transform 1 0 27776 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_244
timestamp 1698431365
transform 1 0 28672 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_270
timestamp 1698431365
transform 1 0 31584 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_284
timestamp 1698431365
transform 1 0 33152 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_288
timestamp 1698431365
transform 1 0 33600 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_304
timestamp 1698431365
transform 1 0 35392 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_308
timestamp 1698431365
transform 1 0 35840 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_317
timestamp 1698431365
transform 1 0 36848 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_319
timestamp 1698431365
transform 1 0 37072 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_387
timestamp 1698431365
transform 1 0 44688 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_391
timestamp 1698431365
transform 1 0 45136 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_415
timestamp 1698431365
transform 1 0 47824 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_419
timestamp 1698431365
transform 1 0 48272 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_421
timestamp 1698431365
transform 1 0 48496 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_438
timestamp 1698431365
transform 1 0 50400 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_442
timestamp 1698431365
transform 1 0 50848 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_444
timestamp 1698431365
transform 1 0 51072 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_463
timestamp 1698431365
transform 1 0 53200 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_467
timestamp 1698431365
transform 1 0 53648 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_469
timestamp 1698431365
transform 1 0 53872 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_493
timestamp 1698431365
transform 1 0 56560 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_14
timestamp 1698431365
transform 1 0 2912 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_18
timestamp 1698431365
transform 1 0 3360 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_22
timestamp 1698431365
transform 1 0 3808 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_24
timestamp 1698431365
transform 1 0 4032 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_30
timestamp 1698431365
transform 1 0 4704 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_46
timestamp 1698431365
transform 1 0 6496 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_50
timestamp 1698431365
transform 1 0 6944 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_58
timestamp 1698431365
transform 1 0 7840 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_66
timestamp 1698431365
transform 1 0 8736 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_95
timestamp 1698431365
transform 1 0 11984 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_121
timestamp 1698431365
transform 1 0 14896 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_123
timestamp 1698431365
transform 1 0 15120 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_142
timestamp 1698431365
transform 1 0 17248 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_150
timestamp 1698431365
transform 1 0 18144 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_174
timestamp 1698431365
transform 1 0 20832 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_182
timestamp 1698431365
transform 1 0 21728 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_201
timestamp 1698431365
transform 1 0 23856 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_209
timestamp 1698431365
transform 1 0 24752 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_212
timestamp 1698431365
transform 1 0 25088 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_244
timestamp 1698431365
transform 1 0 28672 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_263
timestamp 1698431365
transform 1 0 30800 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_267
timestamp 1698431365
transform 1 0 31248 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_275
timestamp 1698431365
transform 1 0 32144 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_279
timestamp 1698431365
transform 1 0 32592 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_294
timestamp 1698431365
transform 1 0 34272 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_310
timestamp 1698431365
transform 1 0 36064 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_318
timestamp 1698431365
transform 1 0 36960 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_335
timestamp 1698431365
transform 1 0 38864 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_345
timestamp 1698431365
transform 1 0 39984 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_349
timestamp 1698431365
transform 1 0 40432 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_352
timestamp 1698431365
transform 1 0 40768 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_412
timestamp 1698431365
transform 1 0 47488 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_414
timestamp 1698431365
transform 1 0 47712 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_422
timestamp 1698431365
transform 1 0 48608 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_429
timestamp 1698431365
transform 1 0 49392 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_444
timestamp 1698431365
transform 1 0 51072 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_452
timestamp 1698431365
transform 1 0 51968 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_454
timestamp 1698431365
transform 1 0 52192 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_486
timestamp 1698431365
transform 1 0 55776 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_492
timestamp 1698431365
transform 1 0 56448 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_508
timestamp 1698431365
transform 1 0 58240 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_14
timestamp 1698431365
transform 1 0 2912 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_18
timestamp 1698431365
transform 1 0 3360 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_34
timestamp 1698431365
transform 1 0 5152 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_37
timestamp 1698431365
transform 1 0 5488 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_72
timestamp 1698431365
transform 1 0 9408 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_99
timestamp 1698431365
transform 1 0 12432 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_103
timestamp 1698431365
transform 1 0 12880 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_107
timestamp 1698431365
transform 1 0 13328 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_113
timestamp 1698431365
transform 1 0 14000 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_117
timestamp 1698431365
transform 1 0 14448 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_129
timestamp 1698431365
transform 1 0 15792 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_139
timestamp 1698431365
transform 1 0 16912 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_147
timestamp 1698431365
transform 1 0 17808 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_151
timestamp 1698431365
transform 1 0 18256 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_165
timestamp 1698431365
transform 1 0 19824 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_173
timestamp 1698431365
transform 1 0 20720 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_177
timestamp 1698431365
transform 1 0 21168 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_185
timestamp 1698431365
transform 1 0 22064 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_189
timestamp 1698431365
transform 1 0 22512 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_200
timestamp 1698431365
transform 1 0 23744 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_232
timestamp 1698431365
transform 1 0 27328 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_240
timestamp 1698431365
transform 1 0 28224 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_244
timestamp 1698431365
transform 1 0 28672 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_247
timestamp 1698431365
transform 1 0 29008 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_260
timestamp 1698431365
transform 1 0 30464 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_264
timestamp 1698431365
transform 1 0 30912 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_305
timestamp 1698431365
transform 1 0 35504 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_313
timestamp 1698431365
transform 1 0 36400 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_327
timestamp 1698431365
transform 1 0 37968 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_335
timestamp 1698431365
transform 1 0 38864 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_341
timestamp 1698431365
transform 1 0 39536 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_349
timestamp 1698431365
transform 1 0 40432 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_358
timestamp 1698431365
transform 1 0 41440 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_383
timestamp 1698431365
transform 1 0 44240 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_387
timestamp 1698431365
transform 1 0 44688 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_395
timestamp 1698431365
transform 1 0 45584 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_451
timestamp 1698431365
transform 1 0 51856 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_457
timestamp 1698431365
transform 1 0 52528 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_487
timestamp 1698431365
transform 1 0 55888 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_503
timestamp 1698431365
transform 1 0 57680 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_507
timestamp 1698431365
transform 1 0 58128 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_2
timestamp 1698431365
transform 1 0 1568 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_51_8
timestamp 1698431365
transform 1 0 2240 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_40
timestamp 1698431365
transform 1 0 5824 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_48
timestamp 1698431365
transform 1 0 6720 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_66
timestamp 1698431365
transform 1 0 8736 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_72
timestamp 1698431365
transform 1 0 9408 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_74
timestamp 1698431365
transform 1 0 9632 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_97
timestamp 1698431365
transform 1 0 12208 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_101
timestamp 1698431365
transform 1 0 12656 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_110
timestamp 1698431365
transform 1 0 13664 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_135
timestamp 1698431365
transform 1 0 16464 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_139
timestamp 1698431365
transform 1 0 16912 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_150
timestamp 1698431365
transform 1 0 18144 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_166
timestamp 1698431365
transform 1 0 19936 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_205
timestamp 1698431365
transform 1 0 24304 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_209
timestamp 1698431365
transform 1 0 24752 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_212
timestamp 1698431365
transform 1 0 25088 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_276
timestamp 1698431365
transform 1 0 32256 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_282
timestamp 1698431365
transform 1 0 32928 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_290
timestamp 1698431365
transform 1 0 33824 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_292
timestamp 1698431365
transform 1 0 34048 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_299
timestamp 1698431365
transform 1 0 34832 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_336
timestamp 1698431365
transform 1 0 38976 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_338
timestamp 1698431365
transform 1 0 39200 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_349
timestamp 1698431365
transform 1 0 40432 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_352
timestamp 1698431365
transform 1 0 40768 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_418
timestamp 1698431365
transform 1 0 48160 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_437
timestamp 1698431365
transform 1 0 50288 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_471
timestamp 1698431365
transform 1 0 54096 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_487
timestamp 1698431365
transform 1 0 55888 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_489
timestamp 1698431365
transform 1 0 56112 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_492
timestamp 1698431365
transform 1 0 56448 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_508
timestamp 1698431365
transform 1 0 58240 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_8
timestamp 1698431365
transform 1 0 2240 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_12
timestamp 1698431365
transform 1 0 2688 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_28
timestamp 1698431365
transform 1 0 4480 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_32
timestamp 1698431365
transform 1 0 4928 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_34
timestamp 1698431365
transform 1 0 5152 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_37
timestamp 1698431365
transform 1 0 5488 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_53
timestamp 1698431365
transform 1 0 7280 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_61
timestamp 1698431365
transform 1 0 8176 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_71
timestamp 1698431365
transform 1 0 9296 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_83
timestamp 1698431365
transform 1 0 10640 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_87
timestamp 1698431365
transform 1 0 11088 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_113
timestamp 1698431365
transform 1 0 14000 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_121
timestamp 1698431365
transform 1 0 14896 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_129
timestamp 1698431365
transform 1 0 15792 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_142
timestamp 1698431365
transform 1 0 17248 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_148
timestamp 1698431365
transform 1 0 17920 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_183
timestamp 1698431365
transform 1 0 21840 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_197
timestamp 1698431365
transform 1 0 23408 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_229
timestamp 1698431365
transform 1 0 26992 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_237
timestamp 1698431365
transform 1 0 27888 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_241
timestamp 1698431365
transform 1 0 28336 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_253
timestamp 1698431365
transform 1 0 29680 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_257
timestamp 1698431365
transform 1 0 30128 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_261
timestamp 1698431365
transform 1 0 30576 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_269
timestamp 1698431365
transform 1 0 31472 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_273
timestamp 1698431365
transform 1 0 31920 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_293
timestamp 1698431365
transform 1 0 34160 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_309
timestamp 1698431365
transform 1 0 35952 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_317
timestamp 1698431365
transform 1 0 36848 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_326
timestamp 1698431365
transform 1 0 37856 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_328
timestamp 1698431365
transform 1 0 38080 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_387
timestamp 1698431365
transform 1 0 44688 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_391
timestamp 1698431365
transform 1 0 45136 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_454
timestamp 1698431365
transform 1 0 52192 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_465
timestamp 1698431365
transform 1 0 53424 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_497
timestamp 1698431365
transform 1 0 57008 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_505
timestamp 1698431365
transform 1 0 57904 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_2
timestamp 1698431365
transform 1 0 1568 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_66
timestamp 1698431365
transform 1 0 8736 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_121
timestamp 1698431365
transform 1 0 14896 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_123
timestamp 1698431365
transform 1 0 15120 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_130
timestamp 1698431365
transform 1 0 15904 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_192
timestamp 1698431365
transform 1 0 22848 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_208
timestamp 1698431365
transform 1 0 24640 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_212
timestamp 1698431365
transform 1 0 25088 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_228
timestamp 1698431365
transform 1 0 26880 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_261
timestamp 1698431365
transform 1 0 30576 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_263
timestamp 1698431365
transform 1 0 30800 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_266
timestamp 1698431365
transform 1 0 31136 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_274
timestamp 1698431365
transform 1 0 32032 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_278
timestamp 1698431365
transform 1 0 32480 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_282
timestamp 1698431365
transform 1 0 32928 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_290
timestamp 1698431365
transform 1 0 33824 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_294
timestamp 1698431365
transform 1 0 34272 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_360
timestamp 1698431365
transform 1 0 41664 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_457
timestamp 1698431365
transform 1 0 52528 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_461
timestamp 1698431365
transform 1 0 52976 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_465
timestamp 1698431365
transform 1 0 53424 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_481
timestamp 1698431365
transform 1 0 55216 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_489
timestamp 1698431365
transform 1 0 56112 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_492
timestamp 1698431365
transform 1 0 56448 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_508
timestamp 1698431365
transform 1 0 58240 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_2
timestamp 1698431365
transform 1 0 1568 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_36
timestamp 1698431365
transform 1 0 5376 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_52
timestamp 1698431365
transform 1 0 7168 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_70
timestamp 1698431365
transform 1 0 9184 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_72
timestamp 1698431365
transform 1 0 9408 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_87
timestamp 1698431365
transform 1 0 11088 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_89
timestamp 1698431365
transform 1 0 11312 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_115
timestamp 1698431365
transform 1 0 14224 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_119
timestamp 1698431365
transform 1 0 14672 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_127
timestamp 1698431365
transform 1 0 15568 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_129
timestamp 1698431365
transform 1 0 15792 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_132
timestamp 1698431365
transform 1 0 16128 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_138
timestamp 1698431365
transform 1 0 16800 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_157
timestamp 1698431365
transform 1 0 18928 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_161
timestamp 1698431365
transform 1 0 19376 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_169
timestamp 1698431365
transform 1 0 20272 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_180
timestamp 1698431365
transform 1 0 21504 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_196
timestamp 1698431365
transform 1 0 23296 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_206
timestamp 1698431365
transform 1 0 24416 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_222
timestamp 1698431365
transform 1 0 26208 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_228
timestamp 1698431365
transform 1 0 26880 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_274
timestamp 1698431365
transform 1 0 32032 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_290
timestamp 1698431365
transform 1 0 33824 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_298
timestamp 1698431365
transform 1 0 34720 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_302
timestamp 1698431365
transform 1 0 35168 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_308
timestamp 1698431365
transform 1 0 35840 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_312
timestamp 1698431365
transform 1 0 36288 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_315
timestamp 1698431365
transform 1 0 36624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_337
timestamp 1698431365
transform 1 0 39088 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_339
timestamp 1698431365
transform 1 0 39312 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_354
timestamp 1698431365
transform 1 0 40992 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_384
timestamp 1698431365
transform 1 0 44352 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_407
timestamp 1698431365
transform 1 0 46928 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_428
timestamp 1698431365
transform 1 0 49280 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_462
timestamp 1698431365
transform 1 0 53088 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_466
timestamp 1698431365
transform 1 0 53536 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_470
timestamp 1698431365
transform 1 0 53984 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_474
timestamp 1698431365
transform 1 0 54432 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_478
timestamp 1698431365
transform 1 0 54880 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_494
timestamp 1698431365
transform 1 0 56672 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_502
timestamp 1698431365
transform 1 0 57568 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_506
timestamp 1698431365
transform 1 0 58016 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_508
timestamp 1698431365
transform 1 0 58240 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1698431365
transform -1 0 57680 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698431365
transform 1 0 27328 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1698431365
transform -1 0 29680 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input4
timestamp 1698431365
transform 1 0 29904 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1698431365
transform -1 0 58352 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1698431365
transform -1 0 58352 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input7
timestamp 1698431365
transform -1 0 58352 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1698431365
transform -1 0 58352 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input9
timestamp 1698431365
transform -1 0 58352 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input10
timestamp 1698431365
transform -1 0 58352 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input11
timestamp 1698431365
transform -1 0 58352 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input12
timestamp 1698431365
transform -1 0 58352 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input13
timestamp 1698431365
transform -1 0 58352 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input14
timestamp 1698431365
transform -1 0 58352 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input15
timestamp 1698431365
transform -1 0 58352 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input16
timestamp 1698431365
transform -1 0 58352 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input17
timestamp 1698431365
transform -1 0 58352 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input18
timestamp 1698431365
transform -1 0 39424 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input19
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input20
timestamp 1698431365
transform 1 0 2240 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input21
timestamp 1698431365
transform 1 0 2240 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input22
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input23
timestamp 1698431365
transform 1 0 2240 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input24
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input25
timestamp 1698431365
transform 1 0 17584 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input26
timestamp 1698431365
transform 1 0 12096 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input27
timestamp 1698431365
transform -1 0 12096 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input28
timestamp 1698431365
transform 1 0 1568 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input29
timestamp 1698431365
transform -1 0 38080 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input30
timestamp 1698431365
transform 1 0 2240 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input31
timestamp 1698431365
transform 1 0 1568 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input32
timestamp 1698431365
transform 1 0 1568 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input33
timestamp 1698431365
transform 1 0 1568 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input34
timestamp 1698431365
transform -1 0 51744 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input35
timestamp 1698431365
transform 1 0 45360 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input36
timestamp 1698431365
transform -1 0 44352 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input37
timestamp 1698431365
transform -1 0 47936 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input38
timestamp 1698431365
transform 1 0 37072 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input39
timestamp 1698431365
transform 1 0 40320 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input40
timestamp 1698431365
transform -1 0 39424 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input41
timestamp 1698431365
transform -1 0 48608 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input42
timestamp 1698431365
transform 1 0 39536 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input43
timestamp 1698431365
transform -1 0 41888 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input44
timestamp 1698431365
transform 1 0 28224 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input45
timestamp 1698431365
transform 1 0 26320 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input46
timestamp 1698431365
transform -1 0 41216 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input47
timestamp 1698431365
transform -1 0 34272 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input48
timestamp 1698431365
transform 1 0 2240 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input49
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input50
timestamp 1698431365
transform -1 0 31696 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input51
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input52
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input53
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input54
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input55
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input56
timestamp 1698431365
transform 1 0 14224 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input57
timestamp 1698431365
transform 1 0 1568 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input58
timestamp 1698431365
transform 1 0 1568 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input59
timestamp 1698431365
transform 1 0 2240 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input60
timestamp 1698431365
transform 1 0 1568 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input61
timestamp 1698431365
transform -1 0 26320 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input62
timestamp 1698431365
transform -1 0 11088 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input63
timestamp 1698431365
transform -1 0 8960 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input64
timestamp 1698431365
transform 1 0 16912 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input65
timestamp 1698431365
transform -1 0 18928 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input66
timestamp 1698431365
transform -1 0 40320 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input67
timestamp 1698431365
transform 1 0 38416 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input68
timestamp 1698431365
transform -1 0 38416 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input69
timestamp 1698431365
transform -1 0 31808 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input70
timestamp 1698431365
transform -1 0 46928 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input71
timestamp 1698431365
transform -1 0 45360 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input72
timestamp 1698431365
transform 1 0 26992 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input73
timestamp 1698431365
transform -1 0 53088 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input74
timestamp 1698431365
transform -1 0 52416 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input75
timestamp 1698431365
transform 1 0 29680 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input76
timestamp 1698431365
transform 1 0 31696 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input77
timestamp 1698431365
transform -1 0 33600 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input78
timestamp 1698431365
transform -1 0 44128 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input79
timestamp 1698431365
transform -1 0 44800 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input80
timestamp 1698431365
transform 1 0 3136 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input81
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input82
timestamp 1698431365
transform -1 0 57680 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output83 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 53312 0 -1 15680
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output84
timestamp 1698431365
transform 1 0 53312 0 -1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output85
timestamp 1698431365
transform 1 0 53312 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output86
timestamp 1698431365
transform 1 0 55440 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output87
timestamp 1698431365
transform 1 0 55440 0 1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output88
timestamp 1698431365
transform 1 0 52528 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output89
timestamp 1698431365
transform 1 0 33712 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output90
timestamp 1698431365
transform -1 0 31248 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output91
timestamp 1698431365
transform -1 0 4480 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output92
timestamp 1698431365
transform -1 0 4480 0 1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output93
timestamp 1698431365
transform -1 0 4480 0 -1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output94
timestamp 1698431365
transform 1 0 52528 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output95
timestamp 1698431365
transform -1 0 4480 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output96
timestamp 1698431365
transform -1 0 30576 0 -1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output97
timestamp 1698431365
transform -1 0 29904 0 -1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output98
timestamp 1698431365
transform 1 0 28224 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output99
timestamp 1698431365
transform -1 0 4480 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output100
timestamp 1698431365
transform -1 0 4480 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output101
timestamp 1698431365
transform 1 0 55440 0 1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output102
timestamp 1698431365
transform -1 0 37296 0 -1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output103
timestamp 1698431365
transform 1 0 55440 0 1 29792
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output104
timestamp 1698431365
transform 1 0 55440 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output105
timestamp 1698431365
transform 1 0 55440 0 1 15680
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output106
timestamp 1698431365
transform 1 0 53312 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output107
timestamp 1698431365
transform 1 0 53312 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output108
timestamp 1698431365
transform 1 0 55440 0 1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output109
timestamp 1698431365
transform 1 0 53312 0 -1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output110
timestamp 1698431365
transform -1 0 38752 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output111
timestamp 1698431365
transform -1 0 31808 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output112
timestamp 1698431365
transform 1 0 55440 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output113
timestamp 1698431365
transform 1 0 53312 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output114
timestamp 1698431365
transform 1 0 55440 0 1 14112
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output115
timestamp 1698431365
transform 1 0 55440 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output116
timestamp 1698431365
transform 1 0 55440 0 1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  pcpi_approx_mul_117 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 22064 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_55 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 58576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_56
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 58576 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_57
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 58576 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_58
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 58576 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_59
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 58576 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_60
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 58576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_61
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 58576 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_62
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 58576 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_63
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 58576 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_64
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 58576 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_65
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 58576 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_66
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 58576 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_67
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 58576 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_68
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 58576 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_69
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 58576 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_70
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 58576 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_71
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 58576 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_72
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 58576 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_73
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 58576 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_74
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 58576 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_75
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 58576 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_76
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 58576 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_77
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 58576 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_78
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 58576 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_79
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 58576 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_80
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 58576 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_81
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 58576 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_82
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 58576 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_83
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 58576 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_84
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 58576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_85
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 58576 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_86
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 58576 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_87
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 58576 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_88
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 58576 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_89
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 58576 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_90
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 58576 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_91
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 58576 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_92
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 58576 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_93
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 58576 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_94
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 58576 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_95
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 58576 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_96
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 58576 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_97
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 58576 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_98
timestamp 1698431365
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698431365
transform -1 0 58576 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_99
timestamp 1698431365
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698431365
transform -1 0 58576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_100
timestamp 1698431365
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698431365
transform -1 0 58576 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_101
timestamp 1698431365
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698431365
transform -1 0 58576 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_102
timestamp 1698431365
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698431365
transform -1 0 58576 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_103
timestamp 1698431365
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698431365
transform -1 0 58576 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_104
timestamp 1698431365
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698431365
transform -1 0 58576 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Left_105
timestamp 1698431365
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1698431365
transform -1 0 58576 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Left_106
timestamp 1698431365
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1698431365
transform -1 0 58576 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Left_107
timestamp 1698431365
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Right_52
timestamp 1698431365
transform -1 0 58576 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Left_108
timestamp 1698431365
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Right_53
timestamp 1698431365
transform -1 0 58576 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Left_109
timestamp 1698431365
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Right_54
timestamp 1698431365
transform -1 0 58576 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_110 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_111
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_112
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_113
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_114
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_115
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_116
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_117
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_118
timestamp 1698431365
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_119
timestamp 1698431365
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_120
timestamp 1698431365
transform 1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_121
timestamp 1698431365
transform 1 0 47040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_122
timestamp 1698431365
transform 1 0 50848 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_123
timestamp 1698431365
transform 1 0 54656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_124
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_125
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_126
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_127
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_128
timestamp 1698431365
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_129
timestamp 1698431365
transform 1 0 48384 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_130
timestamp 1698431365
transform 1 0 56224 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_131
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_132
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_133
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_134
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_135
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_136
timestamp 1698431365
transform 1 0 44464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_137
timestamp 1698431365
transform 1 0 52304 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_138
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_139
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_140
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_141
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_142
timestamp 1698431365
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_143
timestamp 1698431365
transform 1 0 48384 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_144
timestamp 1698431365
transform 1 0 56224 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_145
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_146
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_147
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_148
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_149
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_150
timestamp 1698431365
transform 1 0 44464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_151
timestamp 1698431365
transform 1 0 52304 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_152
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_153
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_154
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_155
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_156
timestamp 1698431365
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_157
timestamp 1698431365
transform 1 0 48384 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_158
timestamp 1698431365
transform 1 0 56224 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_159
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_160
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_161
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_162
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_163
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_164
timestamp 1698431365
transform 1 0 44464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_165
timestamp 1698431365
transform 1 0 52304 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_166
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_167
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_168
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_169
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_170
timestamp 1698431365
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_171
timestamp 1698431365
transform 1 0 48384 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_172
timestamp 1698431365
transform 1 0 56224 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_173
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_174
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_175
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_176
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_177
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_178
timestamp 1698431365
transform 1 0 44464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_179
timestamp 1698431365
transform 1 0 52304 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_180
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_181
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_182
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_183
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_184
timestamp 1698431365
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_185
timestamp 1698431365
transform 1 0 48384 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_186
timestamp 1698431365
transform 1 0 56224 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_187
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_188
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_189
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_190
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_191
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_192
timestamp 1698431365
transform 1 0 44464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_193
timestamp 1698431365
transform 1 0 52304 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_194
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_195
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_196
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_197
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_198
timestamp 1698431365
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_199
timestamp 1698431365
transform 1 0 48384 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_200
timestamp 1698431365
transform 1 0 56224 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_201
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_202
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_203
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_204
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_205
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_206
timestamp 1698431365
transform 1 0 44464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_207
timestamp 1698431365
transform 1 0 52304 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_208
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_209
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_210
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_211
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_212
timestamp 1698431365
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_213
timestamp 1698431365
transform 1 0 48384 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_214
timestamp 1698431365
transform 1 0 56224 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_215
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_216
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_217
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_218
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_219
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_220
timestamp 1698431365
transform 1 0 44464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_221
timestamp 1698431365
transform 1 0 52304 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_222
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_223
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_224
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_225
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_226
timestamp 1698431365
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_227
timestamp 1698431365
transform 1 0 48384 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_228
timestamp 1698431365
transform 1 0 56224 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_229
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_230
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_231
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_232
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_233
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_234
timestamp 1698431365
transform 1 0 44464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_235
timestamp 1698431365
transform 1 0 52304 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_236
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_237
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_238
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_239
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_240
timestamp 1698431365
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_241
timestamp 1698431365
transform 1 0 48384 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_242
timestamp 1698431365
transform 1 0 56224 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_243
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_244
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_245
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_246
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_247
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_248
timestamp 1698431365
transform 1 0 44464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_249
timestamp 1698431365
transform 1 0 52304 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_250
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_251
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_252
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_253
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_254
timestamp 1698431365
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_255
timestamp 1698431365
transform 1 0 48384 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_256
timestamp 1698431365
transform 1 0 56224 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_257
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_258
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_259
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_260
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_261
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_262
timestamp 1698431365
transform 1 0 44464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_263
timestamp 1698431365
transform 1 0 52304 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_264
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_265
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_266
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_267
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_268
timestamp 1698431365
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_269
timestamp 1698431365
transform 1 0 48384 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_270
timestamp 1698431365
transform 1 0 56224 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_271
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_272
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_273
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_274
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_275
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_276
timestamp 1698431365
transform 1 0 44464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_277
timestamp 1698431365
transform 1 0 52304 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_278
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_279
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_280
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_281
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_282
timestamp 1698431365
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_283
timestamp 1698431365
transform 1 0 48384 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_284
timestamp 1698431365
transform 1 0 56224 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_285
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_286
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_287
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_288
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_289
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_290
timestamp 1698431365
transform 1 0 44464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_291
timestamp 1698431365
transform 1 0 52304 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_292
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_293
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_294
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_295
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_296
timestamp 1698431365
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_297
timestamp 1698431365
transform 1 0 48384 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_298
timestamp 1698431365
transform 1 0 56224 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_299
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_300
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_301
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_302
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_303
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_304
timestamp 1698431365
transform 1 0 44464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_305
timestamp 1698431365
transform 1 0 52304 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_306
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_307
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_308
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_309
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_310
timestamp 1698431365
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_311
timestamp 1698431365
transform 1 0 48384 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_312
timestamp 1698431365
transform 1 0 56224 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_313
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_314
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_315
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_316
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_317
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_318
timestamp 1698431365
transform 1 0 44464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_319
timestamp 1698431365
transform 1 0 52304 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_320
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_321
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_322
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_323
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_324
timestamp 1698431365
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_325
timestamp 1698431365
transform 1 0 48384 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_326
timestamp 1698431365
transform 1 0 56224 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_327
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_328
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_329
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_330
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_331
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_332
timestamp 1698431365
transform 1 0 44464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_333
timestamp 1698431365
transform 1 0 52304 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_334
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_335
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_336
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_337
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_338
timestamp 1698431365
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_339
timestamp 1698431365
transform 1 0 48384 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_340
timestamp 1698431365
transform 1 0 56224 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_341
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_342
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_343
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_344
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_345
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_346
timestamp 1698431365
transform 1 0 44464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_347
timestamp 1698431365
transform 1 0 52304 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_348
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_349
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_350
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_351
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_352
timestamp 1698431365
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_353
timestamp 1698431365
transform 1 0 48384 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_354
timestamp 1698431365
transform 1 0 56224 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_355
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_356
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_357
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_358
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_359
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_360
timestamp 1698431365
transform 1 0 44464 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_361
timestamp 1698431365
transform 1 0 52304 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_362
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_363
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_364
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_365
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_366
timestamp 1698431365
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_367
timestamp 1698431365
transform 1 0 48384 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_368
timestamp 1698431365
transform 1 0 56224 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_369
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_370
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_371
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_372
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_373
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_374
timestamp 1698431365
transform 1 0 44464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_375
timestamp 1698431365
transform 1 0 52304 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_376
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_377
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_378
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_379
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_380
timestamp 1698431365
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_381
timestamp 1698431365
transform 1 0 48384 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_382
timestamp 1698431365
transform 1 0 56224 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_383
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_384
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_385
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_386
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_387
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_388
timestamp 1698431365
transform 1 0 44464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_389
timestamp 1698431365
transform 1 0 52304 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_390
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_391
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_392
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_393
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_394
timestamp 1698431365
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_395
timestamp 1698431365
transform 1 0 48384 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_396
timestamp 1698431365
transform 1 0 56224 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_397
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_398
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_399
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_400
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_401
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_402
timestamp 1698431365
transform 1 0 44464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_403
timestamp 1698431365
transform 1 0 52304 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_404
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_405
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_406
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_407
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_408
timestamp 1698431365
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_409
timestamp 1698431365
transform 1 0 48384 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_410
timestamp 1698431365
transform 1 0 56224 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_411
timestamp 1698431365
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_412
timestamp 1698431365
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_413
timestamp 1698431365
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_414
timestamp 1698431365
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_415
timestamp 1698431365
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_416
timestamp 1698431365
transform 1 0 44464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_417
timestamp 1698431365
transform 1 0 52304 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_418
timestamp 1698431365
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_419
timestamp 1698431365
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_420
timestamp 1698431365
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_421
timestamp 1698431365
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_422
timestamp 1698431365
transform 1 0 40544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_423
timestamp 1698431365
transform 1 0 48384 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_424
timestamp 1698431365
transform 1 0 56224 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_425
timestamp 1698431365
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_426
timestamp 1698431365
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_427
timestamp 1698431365
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_428
timestamp 1698431365
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_429
timestamp 1698431365
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_430
timestamp 1698431365
transform 1 0 44464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_431
timestamp 1698431365
transform 1 0 52304 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_432
timestamp 1698431365
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_433
timestamp 1698431365
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_434
timestamp 1698431365
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_435
timestamp 1698431365
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_436
timestamp 1698431365
transform 1 0 40544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_437
timestamp 1698431365
transform 1 0 48384 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_438
timestamp 1698431365
transform 1 0 56224 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_439
timestamp 1698431365
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_440
timestamp 1698431365
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_441
timestamp 1698431365
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_442
timestamp 1698431365
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_443
timestamp 1698431365
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_444
timestamp 1698431365
transform 1 0 44464 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_445
timestamp 1698431365
transform 1 0 52304 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_446
timestamp 1698431365
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_447
timestamp 1698431365
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_448
timestamp 1698431365
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_449
timestamp 1698431365
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_450
timestamp 1698431365
transform 1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_451
timestamp 1698431365
transform 1 0 48384 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_452
timestamp 1698431365
transform 1 0 56224 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_453
timestamp 1698431365
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_454
timestamp 1698431365
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_455
timestamp 1698431365
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_456
timestamp 1698431365
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_457
timestamp 1698431365
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_458
timestamp 1698431365
transform 1 0 44464 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_459
timestamp 1698431365
transform 1 0 52304 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_460
timestamp 1698431365
transform 1 0 9184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_461
timestamp 1698431365
transform 1 0 17024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_462
timestamp 1698431365
transform 1 0 24864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_463
timestamp 1698431365
transform 1 0 32704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_464
timestamp 1698431365
transform 1 0 40544 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_465
timestamp 1698431365
transform 1 0 48384 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_466
timestamp 1698431365
transform 1 0 56224 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_467
timestamp 1698431365
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_468
timestamp 1698431365
transform 1 0 13104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_469
timestamp 1698431365
transform 1 0 20944 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_470
timestamp 1698431365
transform 1 0 28784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_471
timestamp 1698431365
transform 1 0 36624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_472
timestamp 1698431365
transform 1 0 44464 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_473
timestamp 1698431365
transform 1 0 52304 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_474
timestamp 1698431365
transform 1 0 9184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_475
timestamp 1698431365
transform 1 0 17024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_476
timestamp 1698431365
transform 1 0 24864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_477
timestamp 1698431365
transform 1 0 32704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_478
timestamp 1698431365
transform 1 0 40544 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_479
timestamp 1698431365
transform 1 0 48384 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_480
timestamp 1698431365
transform 1 0 56224 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_481
timestamp 1698431365
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_482
timestamp 1698431365
transform 1 0 13104 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_483
timestamp 1698431365
transform 1 0 20944 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_484
timestamp 1698431365
transform 1 0 28784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_485
timestamp 1698431365
transform 1 0 36624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_486
timestamp 1698431365
transform 1 0 44464 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_487
timestamp 1698431365
transform 1 0 52304 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_488
timestamp 1698431365
transform 1 0 9184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_489
timestamp 1698431365
transform 1 0 17024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_490
timestamp 1698431365
transform 1 0 24864 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_491
timestamp 1698431365
transform 1 0 32704 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_492
timestamp 1698431365
transform 1 0 40544 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_493
timestamp 1698431365
transform 1 0 48384 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_494
timestamp 1698431365
transform 1 0 56224 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_495
timestamp 1698431365
transform 1 0 5152 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_496
timestamp 1698431365
transform 1 0 8960 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_497
timestamp 1698431365
transform 1 0 12768 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_498
timestamp 1698431365
transform 1 0 16576 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_499
timestamp 1698431365
transform 1 0 20384 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_500
timestamp 1698431365
transform 1 0 24192 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_501
timestamp 1698431365
transform 1 0 28000 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_502
timestamp 1698431365
transform 1 0 31808 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_503
timestamp 1698431365
transform 1 0 35616 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_504
timestamp 1698431365
transform 1 0 39424 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_505
timestamp 1698431365
transform 1 0 43232 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_506
timestamp 1698431365
transform 1 0 47040 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_507
timestamp 1698431365
transform 1 0 50848 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_508
timestamp 1698431365
transform 1 0 54656 0 1 45472
box -86 -86 310 870
<< labels >>
flabel metal3 s 0 28224 800 28336 0 FreeSans 448 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 59200 37632 60000 37744 0 FreeSans 448 0 0 0 pcpi_insn[0]
port 1 nsew signal input
flabel metal2 s 0 0 112 800 0 FreeSans 448 90 0 0 pcpi_insn[10]
port 2 nsew signal input
flabel metal2 s 672 0 784 800 0 FreeSans 448 90 0 0 pcpi_insn[11]
port 3 nsew signal input
flabel metal2 s 28224 49200 28336 50000 0 FreeSans 448 90 0 0 pcpi_insn[12]
port 4 nsew signal input
flabel metal2 s 28896 49200 29008 50000 0 FreeSans 448 90 0 0 pcpi_insn[13]
port 5 nsew signal input
flabel metal2 s 29568 49200 29680 50000 0 FreeSans 448 90 0 0 pcpi_insn[14]
port 6 nsew signal input
flabel metal2 s 1344 0 1456 800 0 FreeSans 448 90 0 0 pcpi_insn[15]
port 7 nsew signal input
flabel metal2 s 2016 0 2128 800 0 FreeSans 448 90 0 0 pcpi_insn[16]
port 8 nsew signal input
flabel metal2 s 2688 0 2800 800 0 FreeSans 448 90 0 0 pcpi_insn[17]
port 9 nsew signal input
flabel metal2 s 3360 0 3472 800 0 FreeSans 448 90 0 0 pcpi_insn[18]
port 10 nsew signal input
flabel metal2 s 4032 0 4144 800 0 FreeSans 448 90 0 0 pcpi_insn[19]
port 11 nsew signal input
flabel metal3 s 59200 32256 60000 32368 0 FreeSans 448 0 0 0 pcpi_insn[1]
port 12 nsew signal input
flabel metal2 s 4704 0 4816 800 0 FreeSans 448 90 0 0 pcpi_insn[20]
port 13 nsew signal input
flabel metal2 s 5376 0 5488 800 0 FreeSans 448 90 0 0 pcpi_insn[21]
port 14 nsew signal input
flabel metal2 s 6048 0 6160 800 0 FreeSans 448 90 0 0 pcpi_insn[22]
port 15 nsew signal input
flabel metal2 s 6720 0 6832 800 0 FreeSans 448 90 0 0 pcpi_insn[23]
port 16 nsew signal input
flabel metal2 s 7392 0 7504 800 0 FreeSans 448 90 0 0 pcpi_insn[24]
port 17 nsew signal input
flabel metal3 s 59200 35616 60000 35728 0 FreeSans 448 0 0 0 pcpi_insn[25]
port 18 nsew signal input
flabel metal3 s 59200 30912 60000 31024 0 FreeSans 448 0 0 0 pcpi_insn[26]
port 19 nsew signal input
flabel metal3 s 59200 26880 60000 26992 0 FreeSans 448 0 0 0 pcpi_insn[27]
port 20 nsew signal input
flabel metal3 s 59200 30240 60000 30352 0 FreeSans 448 0 0 0 pcpi_insn[28]
port 21 nsew signal input
flabel metal3 s 59200 27552 60000 27664 0 FreeSans 448 0 0 0 pcpi_insn[29]
port 22 nsew signal input
flabel metal3 s 59200 36288 60000 36400 0 FreeSans 448 0 0 0 pcpi_insn[2]
port 23 nsew signal input
flabel metal3 s 59200 32928 60000 33040 0 FreeSans 448 0 0 0 pcpi_insn[30]
port 24 nsew signal input
flabel metal3 s 59200 29568 60000 29680 0 FreeSans 448 0 0 0 pcpi_insn[31]
port 25 nsew signal input
flabel metal3 s 59200 33600 60000 33712 0 FreeSans 448 0 0 0 pcpi_insn[3]
port 26 nsew signal input
flabel metal3 s 59200 34944 60000 35056 0 FreeSans 448 0 0 0 pcpi_insn[4]
port 27 nsew signal input
flabel metal3 s 59200 34272 60000 34384 0 FreeSans 448 0 0 0 pcpi_insn[5]
port 28 nsew signal input
flabel metal3 s 59200 36960 60000 37072 0 FreeSans 448 0 0 0 pcpi_insn[6]
port 29 nsew signal input
flabel metal2 s 8064 0 8176 800 0 FreeSans 448 90 0 0 pcpi_insn[7]
port 30 nsew signal input
flabel metal2 s 8736 0 8848 800 0 FreeSans 448 90 0 0 pcpi_insn[8]
port 31 nsew signal input
flabel metal2 s 9408 0 9520 800 0 FreeSans 448 90 0 0 pcpi_insn[9]
port 32 nsew signal input
flabel metal3 s 59200 14784 60000 14896 0 FreeSans 448 0 0 0 pcpi_rd[0]
port 33 nsew signal tristate
flabel metal3 s 59200 16128 60000 16240 0 FreeSans 448 0 0 0 pcpi_rd[10]
port 34 nsew signal tristate
flabel metal3 s 59200 20832 60000 20944 0 FreeSans 448 0 0 0 pcpi_rd[11]
port 35 nsew signal tristate
flabel metal3 s 59200 25536 60000 25648 0 FreeSans 448 0 0 0 pcpi_rd[12]
port 36 nsew signal tristate
flabel metal3 s 59200 22176 60000 22288 0 FreeSans 448 0 0 0 pcpi_rd[13]
port 37 nsew signal tristate
flabel metal3 s 59200 21504 60000 21616 0 FreeSans 448 0 0 0 pcpi_rd[14]
port 38 nsew signal tristate
flabel metal2 s 33600 0 33712 800 0 FreeSans 448 90 0 0 pcpi_rd[15]
port 39 nsew signal tristate
flabel metal2 s 28224 0 28336 800 0 FreeSans 448 90 0 0 pcpi_rd[16]
port 40 nsew signal tristate
flabel metal3 s 0 25536 800 25648 0 FreeSans 448 0 0 0 pcpi_rd[17]
port 41 nsew signal tristate
flabel metal3 s 0 26880 800 26992 0 FreeSans 448 0 0 0 pcpi_rd[18]
port 42 nsew signal tristate
flabel metal3 s 0 26208 800 26320 0 FreeSans 448 0 0 0 pcpi_rd[19]
port 43 nsew signal tristate
flabel metal3 s 59200 16800 60000 16912 0 FreeSans 448 0 0 0 pcpi_rd[1]
port 44 nsew signal tristate
flabel metal3 s 0 24864 800 24976 0 FreeSans 448 0 0 0 pcpi_rd[20]
port 45 nsew signal tristate
flabel metal2 s 27552 0 27664 800 0 FreeSans 448 90 0 0 pcpi_rd[21]
port 46 nsew signal tristate
flabel metal2 s 26880 49200 26992 50000 0 FreeSans 448 90 0 0 pcpi_rd[22]
port 47 nsew signal tristate
flabel metal2 s 26208 49200 26320 50000 0 FreeSans 448 90 0 0 pcpi_rd[23]
port 48 nsew signal tristate
flabel metal3 s 0 24192 800 24304 0 FreeSans 448 0 0 0 pcpi_rd[24]
port 49 nsew signal tristate
flabel metal3 s 0 23520 800 23632 0 FreeSans 448 0 0 0 pcpi_rd[25]
port 50 nsew signal tristate
flabel metal3 s 59200 28224 60000 28336 0 FreeSans 448 0 0 0 pcpi_rd[26]
port 51 nsew signal tristate
flabel metal2 s 34272 49200 34384 50000 0 FreeSans 448 90 0 0 pcpi_rd[27]
port 52 nsew signal tristate
flabel metal3 s 59200 28896 60000 29008 0 FreeSans 448 0 0 0 pcpi_rd[28]
port 53 nsew signal tristate
flabel metal3 s 59200 24864 60000 24976 0 FreeSans 448 0 0 0 pcpi_rd[29]
port 54 nsew signal tristate
flabel metal3 s 59200 17472 60000 17584 0 FreeSans 448 0 0 0 pcpi_rd[2]
port 55 nsew signal tristate
flabel metal3 s 59200 24192 60000 24304 0 FreeSans 448 0 0 0 pcpi_rd[30]
port 56 nsew signal tristate
flabel metal3 s 59200 19488 60000 19600 0 FreeSans 448 0 0 0 pcpi_rd[31]
port 57 nsew signal tristate
flabel metal3 s 59200 20160 60000 20272 0 FreeSans 448 0 0 0 pcpi_rd[3]
port 58 nsew signal tristate
flabel metal3 s 59200 18144 60000 18256 0 FreeSans 448 0 0 0 pcpi_rd[4]
port 59 nsew signal tristate
flabel metal2 s 34944 0 35056 800 0 FreeSans 448 90 0 0 pcpi_rd[5]
port 60 nsew signal tristate
flabel metal2 s 28896 0 29008 800 0 FreeSans 448 90 0 0 pcpi_rd[6]
port 61 nsew signal tristate
flabel metal3 s 59200 18816 60000 18928 0 FreeSans 448 0 0 0 pcpi_rd[7]
port 62 nsew signal tristate
flabel metal3 s 59200 22848 60000 22960 0 FreeSans 448 0 0 0 pcpi_rd[8]
port 63 nsew signal tristate
flabel metal3 s 59200 15456 60000 15568 0 FreeSans 448 0 0 0 pcpi_rd[9]
port 64 nsew signal tristate
flabel metal3 s 59200 23520 60000 23632 0 FreeSans 448 0 0 0 pcpi_ready
port 65 nsew signal tristate
flabel metal2 s 34272 0 34384 800 0 FreeSans 448 90 0 0 pcpi_rs1[0]
port 66 nsew signal input
flabel metal3 s 0 9408 800 9520 0 FreeSans 448 0 0 0 pcpi_rs1[10]
port 67 nsew signal input
flabel metal3 s 0 8736 800 8848 0 FreeSans 448 0 0 0 pcpi_rs1[11]
port 68 nsew signal input
flabel metal3 s 0 12768 800 12880 0 FreeSans 448 0 0 0 pcpi_rs1[12]
port 69 nsew signal input
flabel metal3 s 0 13440 800 13552 0 FreeSans 448 0 0 0 pcpi_rs1[13]
port 70 nsew signal input
flabel metal3 s 0 14112 800 14224 0 FreeSans 448 0 0 0 pcpi_rs1[14]
port 71 nsew signal input
flabel metal3 s 0 16128 800 16240 0 FreeSans 448 0 0 0 pcpi_rs1[15]
port 72 nsew signal input
flabel metal2 s 17472 49200 17584 50000 0 FreeSans 448 90 0 0 pcpi_rs1[16]
port 73 nsew signal input
flabel metal2 s 12768 49200 12880 50000 0 FreeSans 448 90 0 0 pcpi_rs1[17]
port 74 nsew signal input
flabel metal2 s 12096 49200 12208 50000 0 FreeSans 448 90 0 0 pcpi_rs1[18]
port 75 nsew signal input
flabel metal3 s 0 43680 800 43792 0 FreeSans 448 0 0 0 pcpi_rs1[19]
port 76 nsew signal input
flabel metal2 s 35616 0 35728 800 0 FreeSans 448 90 0 0 pcpi_rs1[1]
port 77 nsew signal input
flabel metal3 s 0 42336 800 42448 0 FreeSans 448 0 0 0 pcpi_rs1[20]
port 78 nsew signal input
flabel metal3 s 0 41664 800 41776 0 FreeSans 448 0 0 0 pcpi_rs1[21]
port 79 nsew signal input
flabel metal3 s 0 38976 800 39088 0 FreeSans 448 0 0 0 pcpi_rs1[22]
port 80 nsew signal input
flabel metal3 s 0 33600 800 33712 0 FreeSans 448 0 0 0 pcpi_rs1[23]
port 81 nsew signal input
flabel metal2 s 44352 49200 44464 50000 0 FreeSans 448 90 0 0 pcpi_rs1[24]
port 82 nsew signal input
flabel metal2 s 45024 49200 45136 50000 0 FreeSans 448 90 0 0 pcpi_rs1[25]
port 83 nsew signal input
flabel metal2 s 43008 49200 43120 50000 0 FreeSans 448 90 0 0 pcpi_rs1[26]
port 84 nsew signal input
flabel metal2 s 41664 49200 41776 50000 0 FreeSans 448 90 0 0 pcpi_rs1[27]
port 85 nsew signal input
flabel metal2 s 36960 49200 37072 50000 0 FreeSans 448 90 0 0 pcpi_rs1[28]
port 86 nsew signal input
flabel metal2 s 39648 49200 39760 50000 0 FreeSans 448 90 0 0 pcpi_rs1[29]
port 87 nsew signal input
flabel metal2 s 37632 0 37744 800 0 FreeSans 448 90 0 0 pcpi_rs1[2]
port 88 nsew signal input
flabel metal2 s 43680 49200 43792 50000 0 FreeSans 448 90 0 0 pcpi_rs1[30]
port 89 nsew signal input
flabel metal2 s 40320 49200 40432 50000 0 FreeSans 448 90 0 0 pcpi_rs1[31]
port 90 nsew signal input
flabel metal2 s 36960 0 37072 800 0 FreeSans 448 90 0 0 pcpi_rs1[3]
port 91 nsew signal input
flabel metal2 s 30240 0 30352 800 0 FreeSans 448 90 0 0 pcpi_rs1[4]
port 92 nsew signal input
flabel metal2 s 26208 0 26320 800 0 FreeSans 448 90 0 0 pcpi_rs1[5]
port 93 nsew signal input
flabel metal2 s 36288 0 36400 800 0 FreeSans 448 90 0 0 pcpi_rs1[6]
port 94 nsew signal input
flabel metal2 s 32928 0 33040 800 0 FreeSans 448 90 0 0 pcpi_rs1[7]
port 95 nsew signal input
flabel metal3 s 0 11424 800 11536 0 FreeSans 448 0 0 0 pcpi_rs1[8]
port 96 nsew signal input
flabel metal3 s 0 12096 800 12208 0 FreeSans 448 0 0 0 pcpi_rs1[9]
port 97 nsew signal input
flabel metal2 s 30912 0 31024 800 0 FreeSans 448 90 0 0 pcpi_rs2[0]
port 98 nsew signal input
flabel metal3 s 0 17472 800 17584 0 FreeSans 448 0 0 0 pcpi_rs2[10]
port 99 nsew signal input
flabel metal3 s 0 18816 800 18928 0 FreeSans 448 0 0 0 pcpi_rs2[11]
port 100 nsew signal input
flabel metal3 s 0 10752 800 10864 0 FreeSans 448 0 0 0 pcpi_rs2[12]
port 101 nsew signal input
flabel metal3 s 0 10080 800 10192 0 FreeSans 448 0 0 0 pcpi_rs2[13]
port 102 nsew signal input
flabel metal3 s 0 8064 800 8176 0 FreeSans 448 0 0 0 pcpi_rs2[14]
port 103 nsew signal input
flabel metal2 s 14112 0 14224 800 0 FreeSans 448 90 0 0 pcpi_rs2[15]
port 104 nsew signal input
flabel metal3 s 0 39648 800 39760 0 FreeSans 448 0 0 0 pcpi_rs2[16]
port 105 nsew signal input
flabel metal3 s 0 40320 800 40432 0 FreeSans 448 0 0 0 pcpi_rs2[17]
port 106 nsew signal input
flabel metal3 s 0 40992 800 41104 0 FreeSans 448 0 0 0 pcpi_rs2[18]
port 107 nsew signal input
flabel metal3 s 0 35616 800 35728 0 FreeSans 448 0 0 0 pcpi_rs2[19]
port 108 nsew signal input
flabel metal2 s 25536 0 25648 800 0 FreeSans 448 90 0 0 pcpi_rs2[1]
port 109 nsew signal input
flabel metal2 s 10080 49200 10192 50000 0 FreeSans 448 90 0 0 pcpi_rs2[20]
port 110 nsew signal input
flabel metal2 s 9408 49200 9520 50000 0 FreeSans 448 90 0 0 pcpi_rs2[21]
port 111 nsew signal input
flabel metal2 s 16800 49200 16912 50000 0 FreeSans 448 90 0 0 pcpi_rs2[22]
port 112 nsew signal input
flabel metal2 s 18144 49200 18256 50000 0 FreeSans 448 90 0 0 pcpi_rs2[23]
port 113 nsew signal input
flabel metal2 s 38976 49200 39088 50000 0 FreeSans 448 90 0 0 pcpi_rs2[24]
port 114 nsew signal input
flabel metal2 s 38304 49200 38416 50000 0 FreeSans 448 90 0 0 pcpi_rs2[25]
port 115 nsew signal input
flabel metal2 s 37632 49200 37744 50000 0 FreeSans 448 90 0 0 pcpi_rs2[26]
port 116 nsew signal input
flabel metal2 s 30240 49200 30352 50000 0 FreeSans 448 90 0 0 pcpi_rs2[27]
port 117 nsew signal input
flabel metal2 s 40992 49200 41104 50000 0 FreeSans 448 90 0 0 pcpi_rs2[28]
port 118 nsew signal input
flabel metal2 s 42336 49200 42448 50000 0 FreeSans 448 90 0 0 pcpi_rs2[29]
port 119 nsew signal input
flabel metal2 s 26880 0 26992 800 0 FreeSans 448 90 0 0 pcpi_rs2[2]
port 120 nsew signal input
flabel metal2 s 46368 49200 46480 50000 0 FreeSans 448 90 0 0 pcpi_rs2[30]
port 121 nsew signal input
flabel metal2 s 45696 49200 45808 50000 0 FreeSans 448 90 0 0 pcpi_rs2[31]
port 122 nsew signal input
flabel metal2 s 29568 0 29680 800 0 FreeSans 448 90 0 0 pcpi_rs2[3]
port 123 nsew signal input
flabel metal2 s 31584 0 31696 800 0 FreeSans 448 90 0 0 pcpi_rs2[4]
port 124 nsew signal input
flabel metal2 s 32256 0 32368 800 0 FreeSans 448 90 0 0 pcpi_rs2[5]
port 125 nsew signal input
flabel metal2 s 39648 0 39760 800 0 FreeSans 448 90 0 0 pcpi_rs2[6]
port 126 nsew signal input
flabel metal2 s 43008 0 43120 800 0 FreeSans 448 90 0 0 pcpi_rs2[7]
port 127 nsew signal input
flabel metal3 s 0 15456 800 15568 0 FreeSans 448 0 0 0 pcpi_rs2[8]
port 128 nsew signal input
flabel metal3 s 0 14784 800 14896 0 FreeSans 448 0 0 0 pcpi_rs2[9]
port 129 nsew signal input
flabel metal3 s 59200 31584 60000 31696 0 FreeSans 448 0 0 0 pcpi_valid
port 130 nsew signal input
flabel metal2 s 21504 0 21616 800 0 FreeSans 448 90 0 0 pcpi_wait
port 131 nsew signal tristate
flabel metal3 s 59200 26208 60000 26320 0 FreeSans 448 0 0 0 pcpi_wr
port 132 nsew signal tristate
flabel metal2 s 10080 0 10192 800 0 FreeSans 448 90 0 0 resetn
port 133 nsew signal input
flabel metal4 s 4448 3076 4768 46316 0 FreeSans 1280 90 0 0 vdd
port 134 nsew power bidirectional
flabel metal4 s 35168 3076 35488 46316 0 FreeSans 1280 90 0 0 vdd
port 134 nsew power bidirectional
flabel metal4 s 19808 3076 20128 46316 0 FreeSans 1280 90 0 0 vss
port 135 nsew ground bidirectional
flabel metal4 s 50528 3076 50848 46316 0 FreeSans 1280 90 0 0 vss
port 135 nsew ground bidirectional
rlabel metal1 29960 46256 29960 46256 0 vdd
rlabel metal1 29960 45472 29960 45472 0 vss
rlabel metal2 40264 19712 40264 19712 0 _0000_
rlabel metal2 43064 17192 43064 17192 0 _0001_
rlabel metal3 48440 17752 48440 17752 0 _0002_
rlabel metal2 47656 20440 47656 20440 0 _0003_
rlabel metal2 45192 18872 45192 18872 0 _0004_
rlabel metal3 33824 17080 33824 17080 0 _0005_
rlabel metal2 29176 17192 29176 17192 0 _0006_
rlabel metal2 36120 19488 36120 19488 0 _0007_
rlabel metal2 45416 23688 45416 23688 0 _0008_
rlabel metal2 42056 23856 42056 23856 0 _0009_
rlabel metal2 47656 23072 47656 23072 0 _0010_
rlabel metal2 45920 20104 45920 20104 0 _0011_
rlabel metal2 42056 25928 42056 25928 0 _0012_
rlabel metal2 37128 22120 37128 22120 0 _0013_
rlabel metal2 33880 21168 33880 21168 0 _0014_
rlabel metal2 31304 19712 31304 19712 0 _0015_
rlabel metal2 29512 21000 29512 21000 0 _0016_
rlabel metal2 11704 26628 11704 26628 0 _0017_
rlabel metal3 11648 25368 11648 25368 0 _0018_
rlabel metal2 14952 25816 14952 25816 0 _0019_
rlabel metal3 23072 26152 23072 26152 0 _0020_
rlabel metal2 26152 21000 26152 21000 0 _0021_
rlabel metal2 25928 25312 25928 25312 0 _0022_
rlabel metal3 25032 28056 25032 28056 0 _0023_
rlabel metal2 18592 24024 18592 24024 0 _0024_
rlabel metal2 23464 24080 23464 24080 0 _0025_
rlabel metal3 35000 27944 35000 27944 0 _0026_
rlabel metal2 32480 27160 32480 27160 0 _0027_
rlabel metal2 39984 27160 39984 27160 0 _0028_
rlabel metal2 34328 25704 34328 25704 0 _0029_
rlabel metal3 35336 24024 35336 24024 0 _0030_
rlabel metal2 39536 20888 39536 20888 0 _0031_
rlabel metal2 3304 30296 3304 30296 0 _0032_
rlabel metal2 3192 35392 3192 35392 0 _0033_
rlabel metal2 4984 34832 4984 34832 0 _0034_
rlabel metal2 4424 29960 4424 29960 0 _0035_
rlabel metal2 7280 34328 7280 34328 0 _0036_
rlabel metal2 2408 30184 2408 30184 0 _0037_
rlabel metal2 12376 31024 12376 31024 0 _0038_
rlabel metal2 3864 31752 3864 31752 0 _0039_
rlabel metal2 2744 31360 2744 31360 0 _0040_
rlabel metal2 2520 30576 2520 30576 0 _0041_
rlabel metal2 10584 39144 10584 39144 0 _0042_
rlabel metal2 16632 34160 16632 34160 0 _0043_
rlabel metal2 6608 30968 6608 30968 0 _0044_
rlabel metal3 6552 32536 6552 32536 0 _0045_
rlabel metal2 6944 31752 6944 31752 0 _0046_
rlabel metal2 6664 32200 6664 32200 0 _0047_
rlabel metal2 7896 32256 7896 32256 0 _0048_
rlabel metal2 7168 31080 7168 31080 0 _0049_
rlabel metal3 4480 30968 4480 30968 0 _0050_
rlabel metal2 4200 29064 4200 29064 0 _0051_
rlabel metal2 20216 28784 20216 28784 0 _0052_
rlabel metal2 22680 41888 22680 41888 0 _0053_
rlabel metal2 19656 41608 19656 41608 0 _0054_
rlabel metal2 15064 44968 15064 44968 0 _0055_
rlabel metal2 21840 45304 21840 45304 0 _0056_
rlabel metal2 21224 45304 21224 45304 0 _0057_
rlabel metal2 19768 44744 19768 44744 0 _0058_
rlabel metal2 19208 42840 19208 42840 0 _0059_
rlabel metal2 13608 42392 13608 42392 0 _0060_
rlabel metal2 13944 43176 13944 43176 0 _0061_
rlabel metal2 7896 43400 7896 43400 0 _0062_
rlabel metal2 8232 43176 8232 43176 0 _0063_
rlabel metal2 12824 43456 12824 43456 0 _0064_
rlabel metal2 11872 44184 11872 44184 0 _0065_
rlabel metal2 11424 43288 11424 43288 0 _0066_
rlabel metal3 12768 44184 12768 44184 0 _0067_
rlabel metal2 15624 43960 15624 43960 0 _0068_
rlabel metal2 19544 43064 19544 43064 0 _0069_
rlabel metal3 21448 41944 21448 41944 0 _0070_
rlabel metal3 21616 41832 21616 41832 0 _0071_
rlabel metal2 21448 28224 21448 28224 0 _0072_
rlabel metal2 21672 28616 21672 28616 0 _0073_
rlabel metal3 21952 27720 21952 27720 0 _0074_
rlabel metal3 26712 27608 26712 27608 0 _0075_
rlabel metal2 16296 31416 16296 31416 0 _0076_
rlabel metal2 16408 30744 16408 30744 0 _0077_
rlabel metal3 19600 28728 19600 28728 0 _0078_
rlabel metal2 30072 22232 30072 22232 0 _0079_
rlabel metal2 25928 20272 25928 20272 0 _0080_
rlabel metal2 30744 20664 30744 20664 0 _0081_
rlabel metal2 13608 26264 13608 26264 0 _0082_
rlabel metal2 28392 27888 28392 27888 0 _0083_
rlabel metal2 19992 26320 19992 26320 0 _0084_
rlabel metal3 4200 30408 4200 30408 0 _0085_
rlabel metal2 3864 29904 3864 29904 0 _0086_
rlabel metal2 4872 29736 4872 29736 0 _0087_
rlabel metal3 6664 29288 6664 29288 0 _0088_
rlabel metal2 7336 29624 7336 29624 0 _0089_
rlabel metal2 9128 30968 9128 30968 0 _0090_
rlabel metal3 7504 31528 7504 31528 0 _0091_
rlabel metal3 11256 34216 11256 34216 0 _0092_
rlabel metal2 8680 31696 8680 31696 0 _0093_
rlabel metal2 8064 30968 8064 30968 0 _0094_
rlabel metal2 8680 30464 8680 30464 0 _0095_
rlabel metal2 6328 30464 6328 30464 0 _0096_
rlabel metal3 7952 30184 7952 30184 0 _0097_
rlabel metal2 8456 29064 8456 29064 0 _0098_
rlabel metal3 11984 27832 11984 27832 0 _0099_
rlabel metal2 17976 38780 17976 38780 0 _0100_
rlabel metal2 19096 39816 19096 39816 0 _0101_
rlabel metal2 22344 39088 22344 39088 0 _0102_
rlabel metal2 23464 40768 23464 40768 0 _0103_
rlabel metal3 22568 40488 22568 40488 0 _0104_
rlabel metal2 13384 42672 13384 42672 0 _0105_
rlabel metal2 12712 41776 12712 41776 0 _0106_
rlabel metal2 16464 42728 16464 42728 0 _0107_
rlabel metal2 16408 41888 16408 41888 0 _0108_
rlabel metal2 14280 39816 14280 39816 0 _0109_
rlabel metal2 16968 41440 16968 41440 0 _0110_
rlabel metal2 18424 40768 18424 40768 0 _0111_
rlabel metal3 13216 41048 13216 41048 0 _0112_
rlabel metal2 9968 41048 9968 41048 0 _0113_
rlabel metal2 10360 41440 10360 41440 0 _0114_
rlabel metal3 12152 41272 12152 41272 0 _0115_
rlabel metal2 13496 42168 13496 42168 0 _0116_
rlabel metal2 14840 41552 14840 41552 0 _0117_
rlabel metal2 17976 40712 17976 40712 0 _0118_
rlabel metal2 22792 40096 22792 40096 0 _0119_
rlabel metal2 21896 39144 21896 39144 0 _0120_
rlabel metal2 23352 38808 23352 38808 0 _0121_
rlabel metal3 22008 38696 22008 38696 0 _0122_
rlabel metal3 16968 27944 16968 27944 0 _0123_
rlabel metal2 21560 26936 21560 26936 0 _0124_
rlabel metal2 18760 27776 18760 27776 0 _0125_
rlabel metal3 18424 27832 18424 27832 0 _0126_
rlabel metal2 18312 26992 18312 26992 0 _0127_
rlabel metal2 16968 30744 16968 30744 0 _0128_
rlabel metal3 16800 31192 16800 31192 0 _0129_
rlabel metal2 17528 28784 17528 28784 0 _0130_
rlabel metal3 17416 28504 17416 28504 0 _0131_
rlabel metal2 18200 28784 18200 28784 0 _0132_
rlabel metal2 17696 28392 17696 28392 0 _0133_
rlabel metal2 18368 25480 18368 25480 0 _0134_
rlabel metal2 18760 26544 18760 26544 0 _0135_
rlabel metal2 12712 25536 12712 25536 0 _0136_
rlabel metal2 8792 29120 8792 29120 0 _0137_
rlabel metal2 7448 28672 7448 28672 0 _0138_
rlabel metal2 10584 28896 10584 28896 0 _0139_
rlabel metal3 17360 32648 17360 32648 0 _0140_
rlabel metal2 10360 30408 10360 30408 0 _0141_
rlabel metal2 9912 30352 9912 30352 0 _0142_
rlabel metal2 10808 29400 10808 29400 0 _0143_
rlabel metal2 12152 28560 12152 28560 0 _0144_
rlabel metal2 23688 40768 23688 40768 0 _0145_
rlabel metal2 22008 39536 22008 39536 0 _0146_
rlabel metal2 22232 38696 22232 38696 0 _0147_
rlabel metal2 17976 39256 17976 39256 0 _0148_
rlabel metal2 14392 41216 14392 41216 0 _0149_
rlabel metal2 14000 40376 14000 40376 0 _0150_
rlabel metal3 16072 40376 16072 40376 0 _0151_
rlabel metal2 18760 37632 18760 37632 0 _0152_
rlabel metal2 13944 39760 13944 39760 0 _0153_
rlabel metal2 12712 40040 12712 40040 0 _0154_
rlabel metal2 12264 39480 12264 39480 0 _0155_
rlabel metal3 11424 38696 11424 38696 0 _0156_
rlabel metal3 12432 38808 12432 38808 0 _0157_
rlabel metal2 14728 39536 14728 39536 0 _0158_
rlabel metal3 17304 38696 17304 38696 0 _0159_
rlabel metal2 20720 38808 20720 38808 0 _0160_
rlabel metal3 16744 28336 16744 28336 0 _0161_
rlabel metal2 14504 28056 14504 28056 0 _0162_
rlabel metal3 21672 28616 21672 28616 0 _0163_
rlabel metal2 22456 27944 22456 27944 0 _0164_
rlabel metal2 15176 27720 15176 27720 0 _0165_
rlabel metal2 14112 27944 14112 27944 0 _0166_
rlabel metal2 14168 27496 14168 27496 0 _0167_
rlabel metal3 16968 25480 16968 25480 0 _0168_
rlabel metal2 14728 31248 14728 31248 0 _0169_
rlabel metal2 13832 30520 13832 30520 0 _0170_
rlabel metal3 15960 30184 15960 30184 0 _0171_
rlabel metal2 17640 29680 17640 29680 0 _0172_
rlabel metal2 16072 29904 16072 29904 0 _0173_
rlabel metal3 16576 29400 16576 29400 0 _0174_
rlabel metal2 17192 25984 17192 25984 0 _0175_
rlabel metal3 16268 25592 16268 25592 0 _0176_
rlabel metal2 15624 25256 15624 25256 0 _0177_
rlabel metal3 12992 28504 12992 28504 0 _0178_
rlabel metal3 13608 28616 13608 28616 0 _0179_
rlabel metal2 18648 29288 18648 29288 0 _0180_
rlabel metal2 10920 28728 10920 28728 0 _0181_
rlabel metal2 19712 30184 19712 30184 0 _0182_
rlabel metal2 19544 37576 19544 37576 0 _0183_
rlabel metal2 21336 36624 21336 36624 0 _0184_
rlabel metal3 21784 36456 21784 36456 0 _0185_
rlabel metal3 18648 36344 18648 36344 0 _0186_
rlabel metal2 16744 33936 16744 33936 0 _0187_
rlabel metal2 13440 37464 13440 37464 0 _0188_
rlabel metal3 16968 37240 16968 37240 0 _0189_
rlabel metal2 16184 37128 16184 37128 0 _0190_
rlabel metal3 17192 37128 17192 37128 0 _0191_
rlabel metal2 17528 36568 17528 36568 0 _0192_
rlabel metal2 18536 36568 18536 36568 0 _0193_
rlabel metal2 14056 35616 14056 35616 0 _0194_
rlabel metal2 14280 36848 14280 36848 0 _0195_
rlabel metal3 10360 34104 10360 34104 0 _0196_
rlabel metal2 9800 35000 9800 35000 0 _0197_
rlabel metal2 14168 36064 14168 36064 0 _0198_
rlabel metal2 17976 35168 17976 35168 0 _0199_
rlabel metal2 21784 36064 21784 36064 0 _0200_
rlabel metal2 22568 36008 22568 36008 0 _0201_
rlabel metal2 22456 36456 22456 36456 0 _0202_
rlabel metal2 21952 31080 21952 31080 0 _0203_
rlabel metal2 19320 29736 19320 29736 0 _0204_
rlabel metal2 18984 29288 18984 29288 0 _0205_
rlabel metal2 18200 27608 18200 27608 0 _0206_
rlabel metal2 11144 32032 11144 32032 0 _0207_
rlabel metal2 11816 31808 11816 31808 0 _0208_
rlabel metal3 12880 31640 12880 31640 0 _0209_
rlabel metal2 12488 30744 12488 30744 0 _0210_
rlabel metal2 13104 30184 13104 30184 0 _0211_
rlabel metal2 13944 31304 13944 31304 0 _0212_
rlabel metal3 21000 30016 21000 30016 0 _0213_
rlabel metal2 14280 30744 14280 30744 0 _0214_
rlabel metal2 17080 28168 17080 28168 0 _0215_
rlabel metal2 17528 26936 17528 26936 0 _0216_
rlabel metal2 15400 25480 15400 25480 0 _0217_
rlabel metal2 21952 30184 21952 30184 0 _0218_
rlabel metal3 20384 35672 20384 35672 0 _0219_
rlabel metal3 21224 34216 21224 34216 0 _0220_
rlabel metal2 22344 33600 22344 33600 0 _0221_
rlabel metal2 19208 34440 19208 34440 0 _0222_
rlabel metal3 14336 35896 14336 35896 0 _0223_
rlabel metal2 14504 35952 14504 35952 0 _0224_
rlabel metal2 15064 35168 15064 35168 0 _0225_
rlabel metal2 17976 34048 17976 34048 0 _0226_
rlabel metal2 16632 33600 16632 33600 0 _0227_
rlabel metal2 12376 34104 12376 34104 0 _0228_
rlabel metal2 13160 34216 13160 34216 0 _0229_
rlabel metal2 15008 33320 15008 33320 0 _0230_
rlabel metal2 15288 33376 15288 33376 0 _0231_
rlabel metal2 22568 32928 22568 32928 0 _0232_
rlabel metal2 23128 31696 23128 31696 0 _0233_
rlabel metal2 22232 30184 22232 30184 0 _0234_
rlabel metal2 24360 30240 24360 30240 0 _0235_
rlabel metal2 22568 30296 22568 30296 0 _0236_
rlabel metal2 22848 30968 22848 30968 0 _0237_
rlabel metal2 36232 30968 36232 30968 0 _0238_
rlabel metal3 23688 30184 23688 30184 0 _0239_
rlabel metal2 24920 35728 24920 35728 0 _0240_
rlabel metal2 23912 36344 23912 36344 0 _0241_
rlabel metal2 24752 30408 24752 30408 0 _0242_
rlabel metal2 24920 30128 24920 30128 0 _0243_
rlabel metal2 23912 26488 23912 26488 0 _0244_
rlabel metal2 26376 25816 26376 25816 0 _0245_
rlabel metal3 25480 24920 25480 24920 0 _0246_
rlabel metal2 23408 24920 23408 24920 0 _0247_
rlabel metal2 24808 24136 24808 24136 0 _0248_
rlabel metal2 23464 26712 23464 26712 0 _0249_
rlabel metal2 17528 33768 17528 33768 0 _0250_
rlabel metal2 18424 34496 18424 34496 0 _0251_
rlabel metal2 21672 34552 21672 34552 0 _0252_
rlabel metal2 20216 32424 20216 32424 0 _0253_
rlabel metal2 19544 31864 19544 31864 0 _0254_
rlabel metal3 18368 33320 18368 33320 0 _0255_
rlabel metal2 17752 32816 17752 32816 0 _0256_
rlabel metal2 13944 33768 13944 33768 0 _0257_
rlabel metal2 17416 33096 17416 33096 0 _0258_
rlabel metal2 19320 31304 19320 31304 0 _0259_
rlabel metal3 23016 30856 23016 30856 0 _0260_
rlabel metal2 26152 30016 26152 30016 0 _0261_
rlabel metal3 25200 30856 25200 30856 0 _0262_
rlabel metal2 26376 30240 26376 30240 0 _0263_
rlabel metal2 27048 33264 27048 33264 0 _0264_
rlabel metal2 27272 20832 27272 20832 0 _0265_
rlabel metal3 27608 21000 27608 21000 0 _0266_
rlabel metal3 28448 20664 28448 20664 0 _0267_
rlabel metal2 19992 31808 19992 31808 0 _0268_
rlabel metal2 20384 31640 20384 31640 0 _0269_
rlabel metal3 22176 31528 22176 31528 0 _0270_
rlabel metal2 23240 32704 23240 32704 0 _0271_
rlabel metal3 23576 32424 23576 32424 0 _0272_
rlabel metal2 26040 31584 26040 31584 0 _0273_
rlabel metal2 26264 31864 26264 31864 0 _0274_
rlabel metal2 26152 32256 26152 32256 0 _0275_
rlabel metal2 26656 32536 26656 32536 0 _0276_
rlabel metal2 26712 33544 26712 33544 0 _0277_
rlabel metal2 26040 25900 26040 25900 0 _0278_
rlabel metal2 25760 22456 25760 22456 0 _0279_
rlabel metal2 27776 26880 27776 26880 0 _0280_
rlabel metal2 26488 25816 26488 25816 0 _0281_
rlabel metal2 25368 31696 25368 31696 0 _0282_
rlabel metal3 24808 34104 24808 34104 0 _0283_
rlabel metal2 25480 33432 25480 33432 0 _0284_
rlabel metal2 25144 32536 25144 32536 0 _0285_
rlabel metal2 25480 29792 25480 29792 0 _0286_
rlabel metal2 24920 27832 24920 27832 0 _0287_
rlabel metal2 25704 28336 25704 28336 0 _0288_
rlabel metal3 19600 24808 19600 24808 0 _0289_
rlabel metal2 45080 40432 45080 40432 0 _0290_
rlabel metal2 45976 35448 45976 35448 0 _0291_
rlabel metal3 46816 38920 46816 38920 0 _0292_
rlabel metal2 46760 36848 46760 36848 0 _0293_
rlabel metal2 43456 42056 43456 42056 0 _0294_
rlabel metal3 42392 45080 42392 45080 0 _0295_
rlabel metal2 43064 40600 43064 40600 0 _0296_
rlabel metal2 40712 44688 40712 44688 0 _0297_
rlabel metal2 43624 41440 43624 41440 0 _0298_
rlabel metal2 49000 43008 49000 43008 0 _0299_
rlabel metal2 42280 41608 42280 41608 0 _0300_
rlabel metal2 43848 40600 43848 40600 0 _0301_
rlabel metal2 43736 39088 43736 39088 0 _0302_
rlabel metal2 42896 41272 42896 41272 0 _0303_
rlabel metal3 46200 41384 46200 41384 0 _0304_
rlabel metal2 41944 44128 41944 44128 0 _0305_
rlabel metal2 44464 44408 44464 44408 0 _0306_
rlabel metal2 45416 43176 45416 43176 0 _0307_
rlabel metal2 45976 41664 45976 41664 0 _0308_
rlabel metal2 45248 41720 45248 41720 0 _0309_
rlabel metal2 45752 41944 45752 41944 0 _0310_
rlabel metal2 47096 42448 47096 42448 0 _0311_
rlabel metal2 45864 43932 45864 43932 0 _0312_
rlabel metal3 47544 43176 47544 43176 0 _0313_
rlabel metal2 46312 45360 46312 45360 0 _0314_
rlabel metal2 49112 45472 49112 45472 0 _0315_
rlabel metal3 41776 43960 41776 43960 0 _0316_
rlabel metal2 47656 45024 47656 45024 0 _0317_
rlabel metal2 47656 43400 47656 43400 0 _0318_
rlabel metal2 48104 43932 48104 43932 0 _0319_
rlabel metal2 46816 39592 46816 39592 0 _0320_
rlabel metal3 48328 37912 48328 37912 0 _0321_
rlabel metal2 29400 38976 29400 38976 0 _0322_
rlabel metal2 48328 37576 48328 37576 0 _0323_
rlabel metal2 48888 44352 48888 44352 0 _0324_
rlabel metal2 47208 43064 47208 43064 0 _0325_
rlabel metal2 49784 42112 49784 42112 0 _0326_
rlabel metal3 50064 44072 50064 44072 0 _0327_
rlabel metal3 51856 44968 51856 44968 0 _0328_
rlabel metal2 50120 45192 50120 45192 0 _0329_
rlabel metal2 50008 45360 50008 45360 0 _0330_
rlabel metal2 49896 45416 49896 45416 0 _0331_
rlabel metal2 49672 44744 49672 44744 0 _0332_
rlabel metal2 49560 37520 49560 37520 0 _0333_
rlabel metal3 48272 38696 48272 38696 0 _0334_
rlabel metal2 37688 40432 37688 40432 0 _0335_
rlabel metal2 41552 39368 41552 39368 0 _0336_
rlabel metal3 37520 42728 37520 42728 0 _0337_
rlabel metal3 47600 39592 47600 39592 0 _0338_
rlabel metal3 45864 39368 45864 39368 0 _0339_
rlabel metal2 38920 44408 38920 44408 0 _0340_
rlabel metal2 41160 40656 41160 40656 0 _0341_
rlabel metal2 39144 44240 39144 44240 0 _0342_
rlabel metal2 39312 44184 39312 44184 0 _0343_
rlabel metal2 39704 38584 39704 38584 0 _0344_
rlabel metal2 40376 39424 40376 39424 0 _0345_
rlabel metal2 37912 40824 37912 40824 0 _0346_
rlabel metal3 38080 41048 38080 41048 0 _0347_
rlabel metal2 37688 41608 37688 41608 0 _0348_
rlabel metal2 37408 41944 37408 41944 0 _0349_
rlabel metal2 38584 41664 38584 41664 0 _0350_
rlabel metal2 37632 42504 37632 42504 0 _0351_
rlabel metal2 36344 44800 36344 44800 0 _0352_
rlabel metal2 37520 42728 37520 42728 0 _0353_
rlabel metal2 39928 40208 39928 40208 0 _0354_
rlabel metal2 37240 38920 37240 38920 0 _0355_
rlabel metal3 37184 38696 37184 38696 0 _0356_
rlabel metal3 29344 38920 29344 38920 0 _0357_
rlabel metal2 50624 35896 50624 35896 0 _0358_
rlabel metal2 28840 40376 28840 40376 0 _0359_
rlabel metal2 40264 37968 40264 37968 0 _0360_
rlabel metal2 40376 37968 40376 37968 0 _0361_
rlabel metal2 38864 38808 38864 38808 0 _0362_
rlabel metal2 39480 38024 39480 38024 0 _0363_
rlabel metal2 35112 38724 35112 38724 0 _0364_
rlabel metal2 35224 39088 35224 39088 0 _0365_
rlabel metal2 34776 43008 34776 43008 0 _0366_
rlabel metal2 34552 37912 34552 37912 0 _0367_
rlabel metal2 29736 41440 29736 41440 0 _0368_
rlabel metal2 32424 36736 32424 36736 0 _0369_
rlabel metal2 33992 37968 33992 37968 0 _0370_
rlabel metal2 30744 42448 30744 42448 0 _0371_
rlabel metal2 31976 42616 31976 42616 0 _0372_
rlabel metal3 33936 43400 33936 43400 0 _0373_
rlabel metal2 31080 41552 31080 41552 0 _0374_
rlabel metal2 46760 39312 46760 39312 0 _0375_
rlabel metal2 39032 42840 39032 42840 0 _0376_
rlabel metal2 37128 43176 37128 43176 0 _0377_
rlabel metal2 29848 41216 29848 41216 0 _0378_
rlabel metal2 33432 42224 33432 42224 0 _0379_
rlabel metal2 33208 42280 33208 42280 0 _0380_
rlabel metal2 34104 44128 34104 44128 0 _0381_
rlabel metal2 33656 43932 33656 43932 0 _0382_
rlabel metal2 34440 37688 34440 37688 0 _0383_
rlabel metal2 37184 33208 37184 33208 0 _0384_
rlabel metal2 44128 33208 44128 33208 0 _0385_
rlabel metal2 52808 34272 52808 34272 0 _0386_
rlabel metal3 36848 33432 36848 33432 0 _0387_
rlabel metal3 29848 35728 29848 35728 0 _0388_
rlabel metal2 36904 36008 36904 36008 0 _0389_
rlabel metal2 37912 35952 37912 35952 0 _0390_
rlabel metal2 44184 36064 44184 36064 0 _0391_
rlabel metal2 40152 35952 40152 35952 0 _0392_
rlabel metal2 41496 36960 41496 36960 0 _0393_
rlabel metal2 42168 38920 42168 38920 0 _0394_
rlabel metal2 41832 37520 41832 37520 0 _0395_
rlabel metal2 42392 37408 42392 37408 0 _0396_
rlabel metal2 41272 35840 41272 35840 0 _0397_
rlabel metal2 39592 35728 39592 35728 0 _0398_
rlabel metal2 38752 34328 38752 34328 0 _0399_
rlabel metal2 37464 35112 37464 35112 0 _0400_
rlabel metal2 38136 35728 38136 35728 0 _0401_
rlabel metal2 38024 35280 38024 35280 0 _0402_
rlabel metal2 37352 34440 37352 34440 0 _0403_
rlabel metal2 38584 33600 38584 33600 0 _0404_
rlabel metal2 39032 32760 39032 32760 0 _0405_
rlabel metal2 38584 32032 38584 32032 0 _0406_
rlabel metal2 37240 31416 37240 31416 0 _0407_
rlabel metal2 35224 31808 35224 31808 0 _0408_
rlabel metal2 33096 36736 33096 36736 0 _0409_
rlabel metal2 33768 36288 33768 36288 0 _0410_
rlabel metal3 42504 36904 42504 36904 0 _0411_
rlabel metal2 34552 34944 34552 34944 0 _0412_
rlabel metal2 46592 40376 46592 40376 0 _0413_
rlabel metal3 35224 40376 35224 40376 0 _0414_
rlabel metal2 33880 41048 33880 41048 0 _0415_
rlabel metal2 33712 34216 33712 34216 0 _0416_
rlabel metal2 30072 40768 30072 40768 0 _0417_
rlabel metal3 30968 40376 30968 40376 0 _0418_
rlabel metal2 43400 39312 43400 39312 0 _0419_
rlabel metal2 43792 39704 43792 39704 0 _0420_
rlabel metal2 31192 40880 31192 40880 0 _0421_
rlabel metal2 31304 39816 31304 39816 0 _0422_
rlabel metal2 29064 39984 29064 39984 0 _0423_
rlabel metal2 29512 39648 29512 39648 0 _0424_
rlabel metal2 36344 40656 36344 40656 0 _0425_
rlabel metal2 35896 40040 35896 40040 0 _0426_
rlabel metal2 31080 40040 31080 40040 0 _0427_
rlabel metal2 31864 39144 31864 39144 0 _0428_
rlabel metal3 41244 37800 41244 37800 0 _0429_
rlabel metal2 31472 38920 31472 38920 0 _0430_
rlabel metal2 31752 39984 31752 39984 0 _0431_
rlabel metal2 32872 40096 32872 40096 0 _0432_
rlabel metal2 32088 39172 32088 39172 0 _0433_
rlabel metal2 34328 34608 34328 34608 0 _0434_
rlabel metal2 35336 35000 35336 35000 0 _0435_
rlabel metal2 34888 32704 34888 32704 0 _0436_
rlabel metal3 32312 31864 32312 31864 0 _0437_
rlabel metal3 28896 37352 28896 37352 0 _0438_
rlabel metal3 28336 34216 28336 34216 0 _0439_
rlabel metal2 28056 33600 28056 33600 0 _0440_
rlabel metal2 20104 25424 20104 25424 0 _0441_
rlabel metal2 18984 24976 18984 24976 0 _0442_
rlabel metal2 24472 24024 24472 24024 0 _0443_
rlabel metal2 39032 33880 39032 33880 0 _0444_
rlabel metal2 37576 33096 37576 33096 0 _0445_
rlabel metal2 38696 33768 38696 33768 0 _0446_
rlabel metal3 42224 32536 42224 32536 0 _0447_
rlabel metal2 45864 34552 45864 34552 0 _0448_
rlabel metal3 44072 34216 44072 34216 0 _0449_
rlabel metal2 42952 35784 42952 35784 0 _0450_
rlabel metal2 43176 35448 43176 35448 0 _0451_
rlabel metal2 45416 35672 45416 35672 0 _0452_
rlabel metal2 43344 34888 43344 34888 0 _0453_
rlabel metal2 43624 35280 43624 35280 0 _0454_
rlabel metal2 43400 34328 43400 34328 0 _0455_
rlabel metal2 41272 34888 41272 34888 0 _0456_
rlabel metal2 39984 34216 39984 34216 0 _0457_
rlabel metal2 41048 33544 41048 33544 0 _0458_
rlabel metal2 41608 32984 41608 32984 0 _0459_
rlabel metal2 42504 31864 42504 31864 0 _0460_
rlabel metal2 50680 38248 50680 38248 0 _0461_
rlabel metal2 50456 37464 50456 37464 0 _0462_
rlabel metal2 54432 36344 54432 36344 0 _0463_
rlabel metal2 54488 40488 54488 40488 0 _0464_
rlabel metal2 49448 41216 49448 41216 0 _0465_
rlabel metal2 50064 42616 50064 42616 0 _0466_
rlabel metal2 50176 41160 50176 41160 0 _0467_
rlabel metal2 50344 41664 50344 41664 0 _0468_
rlabel metal2 54712 41888 54712 41888 0 _0469_
rlabel metal2 53480 42280 53480 42280 0 _0470_
rlabel metal2 53144 43512 53144 43512 0 _0471_
rlabel metal2 52920 42392 52920 42392 0 _0472_
rlabel metal2 50680 44240 50680 44240 0 _0473_
rlabel metal3 47544 43064 47544 43064 0 _0474_
rlabel metal2 52528 41720 52528 41720 0 _0475_
rlabel metal2 55160 41104 55160 41104 0 _0476_
rlabel metal2 55160 37744 55160 37744 0 _0477_
rlabel metal2 54600 37184 54600 37184 0 _0478_
rlabel metal2 42840 31080 42840 31080 0 _0479_
rlabel metal2 43120 30968 43120 30968 0 _0480_
rlabel metal3 41888 30072 41888 30072 0 _0481_
rlabel metal2 37912 29736 37912 29736 0 _0482_
rlabel metal2 37016 31472 37016 31472 0 _0483_
rlabel metal2 37688 30464 37688 30464 0 _0484_
rlabel metal2 37352 29568 37352 29568 0 _0485_
rlabel metal2 27720 26432 27720 26432 0 _0486_
rlabel metal2 29848 37632 29848 37632 0 _0487_
rlabel metal2 29064 38780 29064 38780 0 _0488_
rlabel metal2 28224 33544 28224 33544 0 _0489_
rlabel metal2 28504 34104 28504 34104 0 _0490_
rlabel metal2 28000 29960 28000 29960 0 _0491_
rlabel metal2 22680 25088 22680 25088 0 _0492_
rlabel metal3 41776 34104 41776 34104 0 _0493_
rlabel metal2 41944 34104 41944 34104 0 _0494_
rlabel metal2 42728 32872 42728 32872 0 _0495_
rlabel metal3 44296 32536 44296 32536 0 _0496_
rlabel metal3 49280 33208 49280 33208 0 _0497_
rlabel metal2 45304 33768 45304 33768 0 _0498_
rlabel metal3 44128 34104 44128 34104 0 _0499_
rlabel metal2 45864 32984 45864 32984 0 _0500_
rlabel metal2 44632 31752 44632 31752 0 _0501_
rlabel metal2 55384 39928 55384 39928 0 _0502_
rlabel metal2 55944 38640 55944 38640 0 _0503_
rlabel metal2 54488 37072 54488 37072 0 _0504_
rlabel metal2 56504 37072 56504 37072 0 _0505_
rlabel metal2 53816 38584 53816 38584 0 _0506_
rlabel metal2 51632 41384 51632 41384 0 _0507_
rlabel metal2 53200 41944 53200 41944 0 _0508_
rlabel metal2 54040 40656 54040 40656 0 _0509_
rlabel metal2 51688 40712 51688 40712 0 _0510_
rlabel metal2 51408 41272 51408 41272 0 _0511_
rlabel metal2 43960 26852 43960 26852 0 _0512_
rlabel metal2 52024 40656 52024 40656 0 _0513_
rlabel metal2 49560 40600 49560 40600 0 _0514_
rlabel metal3 47152 40264 47152 40264 0 _0515_
rlabel metal2 51800 40768 51800 40768 0 _0516_
rlabel metal2 54264 39928 54264 39928 0 _0517_
rlabel metal2 57120 37240 57120 37240 0 _0518_
rlabel metal3 51016 31472 51016 31472 0 _0519_
rlabel metal2 39816 31920 39816 31920 0 _0520_
rlabel metal2 41384 31416 41384 31416 0 _0521_
rlabel metal2 41720 29680 41720 29680 0 _0522_
rlabel metal3 44016 28056 44016 28056 0 _0523_
rlabel metal3 37408 29400 37408 29400 0 _0524_
rlabel metal3 31248 34104 31248 34104 0 _0525_
rlabel metal2 29344 36456 29344 36456 0 _0526_
rlabel metal2 28280 36232 28280 36232 0 _0527_
rlabel metal2 30352 34104 30352 34104 0 _0528_
rlabel metal2 31080 34272 31080 34272 0 _0529_
rlabel metal2 33320 30576 33320 30576 0 _0530_
rlabel metal2 33544 29064 33544 29064 0 _0531_
rlabel metal2 32088 25144 32088 25144 0 _0532_
rlabel metal2 32760 25424 32760 25424 0 _0533_
rlabel metal3 44352 27944 44352 27944 0 _0534_
rlabel metal3 33152 28392 33152 28392 0 _0535_
rlabel metal2 38360 28224 38360 28224 0 _0536_
rlabel metal3 44408 30296 44408 30296 0 _0537_
rlabel metal2 44072 30744 44072 30744 0 _0538_
rlabel metal2 54936 38864 54936 38864 0 _0539_
rlabel metal2 55272 36344 55272 36344 0 _0540_
rlabel metal3 56112 33880 56112 33880 0 _0541_
rlabel metal2 51240 35616 51240 35616 0 _0542_
rlabel metal3 52304 34776 52304 34776 0 _0543_
rlabel metal2 44184 26320 44184 26320 0 _0544_
rlabel metal2 51464 37240 51464 37240 0 _0545_
rlabel metal2 52248 39872 52248 39872 0 _0546_
rlabel metal2 53256 38304 53256 38304 0 _0547_
rlabel metal2 53480 36680 53480 36680 0 _0548_
rlabel metal2 52248 36512 52248 36512 0 _0549_
rlabel metal2 51240 38192 51240 38192 0 _0550_
rlabel metal2 52472 37128 52472 37128 0 _0551_
rlabel via2 45080 36456 45080 36456 0 _0552_
rlabel metal2 43736 37184 43736 37184 0 _0553_
rlabel metal2 51912 36624 51912 36624 0 _0554_
rlabel metal2 44408 26600 44408 26600 0 _0555_
rlabel metal2 53760 35672 53760 35672 0 _0556_
rlabel metal2 55216 33880 55216 33880 0 _0557_
rlabel metal2 54712 31752 54712 31752 0 _0558_
rlabel metal3 53816 31640 53816 31640 0 _0559_
rlabel metal2 46312 31584 46312 31584 0 _0560_
rlabel metal3 45976 32760 45976 32760 0 _0561_
rlabel metal3 46144 31752 46144 31752 0 _0562_
rlabel metal2 45640 30856 45640 30856 0 _0563_
rlabel metal2 46424 30576 46424 30576 0 _0564_
rlabel metal2 44296 30072 44296 30072 0 _0565_
rlabel metal2 46424 26040 46424 26040 0 _0566_
rlabel metal2 43848 29736 43848 29736 0 _0567_
rlabel metal3 40936 30240 40936 30240 0 _0568_
rlabel metal3 31752 30072 31752 30072 0 _0569_
rlabel metal2 29848 38304 29848 38304 0 _0570_
rlabel metal2 29624 37800 29624 37800 0 _0571_
rlabel metal3 30856 34888 30856 34888 0 _0572_
rlabel metal2 30072 35616 30072 35616 0 _0573_
rlabel metal2 31416 35672 31416 35672 0 _0574_
rlabel metal2 31304 35168 31304 35168 0 _0575_
rlabel metal3 32144 34776 32144 34776 0 _0576_
rlabel metal2 44296 25200 44296 25200 0 _0577_
rlabel metal2 32424 31304 32424 31304 0 _0578_
rlabel metal2 33320 28504 33320 28504 0 _0579_
rlabel metal2 33040 24920 33040 24920 0 _0580_
rlabel metal2 33824 27944 33824 27944 0 _0581_
rlabel metal3 40264 27944 40264 27944 0 _0582_
rlabel metal2 40040 25872 40040 25872 0 _0583_
rlabel metal2 44856 30968 44856 30968 0 _0584_
rlabel metal2 45360 29624 45360 29624 0 _0585_
rlabel metal2 53368 34496 53368 34496 0 _0586_
rlabel metal3 20720 24696 20720 24696 0 _0587_
rlabel metal2 53704 31584 53704 31584 0 _0588_
rlabel metal2 54824 31248 54824 31248 0 _0589_
rlabel metal2 51912 32816 51912 32816 0 _0590_
rlabel metal2 52024 35952 52024 35952 0 _0591_
rlabel metal2 52696 35896 52696 35896 0 _0592_
rlabel metal2 51800 34832 51800 34832 0 _0593_
rlabel metal2 49000 34272 49000 34272 0 _0594_
rlabel metal2 47768 34552 47768 34552 0 _0595_
rlabel metal3 46760 35672 46760 35672 0 _0596_
rlabel metal2 47376 35672 47376 35672 0 _0597_
rlabel metal2 48440 35560 48440 35560 0 _0598_
rlabel metal3 52472 33320 52472 33320 0 _0599_
rlabel metal2 53928 31248 53928 31248 0 _0600_
rlabel metal2 53592 30408 53592 30408 0 _0601_
rlabel metal3 39144 28392 39144 28392 0 _0602_
rlabel metal2 38696 29344 38696 29344 0 _0603_
rlabel metal2 38472 28224 38472 28224 0 _0604_
rlabel metal2 32312 32424 32312 32424 0 _0605_
rlabel metal2 32648 32816 32648 32816 0 _0606_
rlabel metal2 38920 29008 38920 29008 0 _0607_
rlabel metal2 36232 28840 36232 28840 0 _0608_
rlabel metal2 39536 26264 39536 26264 0 _0609_
rlabel metal2 39816 26516 39816 26516 0 _0610_
rlabel metal2 50848 32536 50848 32536 0 _0611_
rlabel metal2 51352 30800 51352 30800 0 _0612_
rlabel metal2 52920 31024 52920 31024 0 _0613_
rlabel metal2 49448 32032 49448 32032 0 _0614_
rlabel metal2 49224 34888 49224 34888 0 _0615_
rlabel metal2 47208 33600 47208 33600 0 _0616_
rlabel metal2 47992 31976 47992 31976 0 _0617_
rlabel metal2 30408 29792 30408 29792 0 _0618_
rlabel metal3 48832 34104 48832 34104 0 _0619_
rlabel metal3 50232 34104 50232 34104 0 _0620_
rlabel metal2 50792 31836 50792 31836 0 _0621_
rlabel metal2 51576 31304 51576 31304 0 _0622_
rlabel metal3 51436 31080 51436 31080 0 _0623_
rlabel metal2 50344 30968 50344 30968 0 _0624_
rlabel metal2 39200 29400 39200 29400 0 _0625_
rlabel metal3 36624 30184 36624 30184 0 _0626_
rlabel metal2 39144 29848 39144 29848 0 _0627_
rlabel metal2 36120 30408 36120 30408 0 _0628_
rlabel metal3 30632 28616 30632 28616 0 _0629_
rlabel metal2 34104 31864 34104 31864 0 _0630_
rlabel metal2 34944 26488 34944 26488 0 _0631_
rlabel metal2 33880 25144 33880 25144 0 _0632_
rlabel metal2 37072 25704 37072 25704 0 _0633_
rlabel metal2 48776 32256 48776 32256 0 _0634_
rlabel metal2 49448 31248 49448 31248 0 _0635_
rlabel metal3 49504 33320 49504 33320 0 _0636_
rlabel metal3 48888 31080 48888 31080 0 _0637_
rlabel metal2 47656 30352 47656 30352 0 _0638_
rlabel metal2 29064 30576 29064 30576 0 _0639_
rlabel metal3 48328 30296 48328 30296 0 _0640_
rlabel metal2 39368 29904 39368 29904 0 _0641_
rlabel metal2 35000 30072 35000 30072 0 _0642_
rlabel metal2 35336 29568 35336 29568 0 _0643_
rlabel metal2 33152 39368 33152 39368 0 _0644_
rlabel metal2 33824 34776 33824 34776 0 _0645_
rlabel metal2 35784 25396 35784 25396 0 _0646_
rlabel metal2 35336 23912 35336 23912 0 _0647_
rlabel metal2 36232 24192 36232 24192 0 _0648_
rlabel metal2 29848 29904 29848 29904 0 _0649_
rlabel metal2 39256 30352 39256 30352 0 _0650_
rlabel metal2 34720 33320 34720 33320 0 _0651_
rlabel metal3 35448 34888 35448 34888 0 _0652_
rlabel metal2 35784 33992 35784 33992 0 _0653_
rlabel metal3 35000 33320 35000 33320 0 _0654_
rlabel metal2 39928 30184 39928 30184 0 _0655_
rlabel metal2 39984 24584 39984 24584 0 _0656_
rlabel metal3 33880 19880 33880 19880 0 _0657_
rlabel metal2 37632 21000 37632 21000 0 _0658_
rlabel metal2 40488 22232 40488 22232 0 _0659_
rlabel metal2 35784 18032 35784 18032 0 _0660_
rlabel metal3 39032 17416 39032 17416 0 _0661_
rlabel metal2 38696 11816 38696 11816 0 _0662_
rlabel metal2 39032 13496 39032 13496 0 _0663_
rlabel metal2 41160 7392 41160 7392 0 _0664_
rlabel metal2 39256 14112 39256 14112 0 _0665_
rlabel metal2 38920 14392 38920 14392 0 _0666_
rlabel metal2 39144 16744 39144 16744 0 _0667_
rlabel metal2 29624 12208 29624 12208 0 _0668_
rlabel metal2 26656 5992 26656 5992 0 _0669_
rlabel metal2 29288 9744 29288 9744 0 _0670_
rlabel metal2 49672 8848 49672 8848 0 _0671_
rlabel metal3 27104 11256 27104 11256 0 _0672_
rlabel metal2 26824 6720 26824 6720 0 _0673_
rlabel metal2 27496 8624 27496 8624 0 _0674_
rlabel metal2 30352 8456 30352 8456 0 _0675_
rlabel metal2 31416 7728 31416 7728 0 _0676_
rlabel metal2 31864 7392 31864 7392 0 _0677_
rlabel metal2 32200 7056 32200 7056 0 _0678_
rlabel metal2 32536 7448 32536 7448 0 _0679_
rlabel metal2 31416 9072 31416 9072 0 _0680_
rlabel metal2 25704 10976 25704 10976 0 _0681_
rlabel metal2 24696 8120 24696 8120 0 _0682_
rlabel metal2 24472 7056 24472 7056 0 _0683_
rlabel metal2 24696 6720 24696 6720 0 _0684_
rlabel metal2 24360 7504 24360 7504 0 _0685_
rlabel metal2 25816 9128 25816 9128 0 _0686_
rlabel metal2 28280 7392 28280 7392 0 _0687_
rlabel metal2 45528 6384 45528 6384 0 _0688_
rlabel metal3 28560 8008 28560 8008 0 _0689_
rlabel metal2 38808 11032 38808 11032 0 _0690_
rlabel metal2 29288 7560 29288 7560 0 _0691_
rlabel metal2 25928 8680 25928 8680 0 _0692_
rlabel metal2 25256 7896 25256 7896 0 _0693_
rlabel metal2 26040 8904 26040 8904 0 _0694_
rlabel metal2 26600 11032 26600 11032 0 _0695_
rlabel metal2 26824 11620 26824 11620 0 _0696_
rlabel metal2 41608 12376 41608 12376 0 _0697_
rlabel metal3 36344 6440 36344 6440 0 _0698_
rlabel metal2 42280 6384 42280 6384 0 _0699_
rlabel metal2 45304 10472 45304 10472 0 _0700_
rlabel metal2 27664 6104 27664 6104 0 _0701_
rlabel metal2 27048 6384 27048 6384 0 _0702_
rlabel metal2 30576 12152 30576 12152 0 _0703_
rlabel metal2 28392 12600 28392 12600 0 _0704_
rlabel metal2 27160 12040 27160 12040 0 _0705_
rlabel metal2 26768 11928 26768 11928 0 _0706_
rlabel metal2 25928 13832 25928 13832 0 _0707_
rlabel metal2 26936 12488 26936 12488 0 _0708_
rlabel metal2 27944 13440 27944 13440 0 _0709_
rlabel metal2 47544 13048 47544 13048 0 _0710_
rlabel metal2 27384 10976 27384 10976 0 _0711_
rlabel metal2 26488 10192 26488 10192 0 _0712_
rlabel metal2 27496 11872 27496 11872 0 _0713_
rlabel metal3 33880 12264 33880 12264 0 _0714_
rlabel metal3 38640 7728 38640 7728 0 _0715_
rlabel metal2 33376 11368 33376 11368 0 _0716_
rlabel metal2 41048 10640 41048 10640 0 _0717_
rlabel metal2 40600 10976 40600 10976 0 _0718_
rlabel metal2 32312 9856 32312 9856 0 _0719_
rlabel metal2 34216 11032 34216 11032 0 _0720_
rlabel metal2 33096 12712 33096 12712 0 _0721_
rlabel metal2 40264 9408 40264 9408 0 _0722_
rlabel metal2 36400 10584 36400 10584 0 _0723_
rlabel metal3 35672 9128 35672 9128 0 _0724_
rlabel metal3 35672 9688 35672 9688 0 _0725_
rlabel metal2 38976 8120 38976 8120 0 _0726_
rlabel metal2 35336 9576 35336 9576 0 _0727_
rlabel metal2 33992 7952 33992 7952 0 _0728_
rlabel metal2 35896 10416 35896 10416 0 _0729_
rlabel metal2 35112 11032 35112 11032 0 _0730_
rlabel metal2 34776 13160 34776 13160 0 _0731_
rlabel metal2 35560 14504 35560 14504 0 _0732_
rlabel metal2 46424 9576 46424 9576 0 _0733_
rlabel metal2 44520 10920 44520 10920 0 _0734_
rlabel metal2 44296 10080 44296 10080 0 _0735_
rlabel metal2 34664 5488 34664 5488 0 _0736_
rlabel metal2 35896 5600 35896 5600 0 _0737_
rlabel metal2 38248 5488 38248 5488 0 _0738_
rlabel metal3 40600 5096 40600 5096 0 _0739_
rlabel metal2 33992 5152 33992 5152 0 _0740_
rlabel metal2 36568 9184 36568 9184 0 _0741_
rlabel metal2 38472 5432 38472 5432 0 _0742_
rlabel metal2 38248 8624 38248 8624 0 _0743_
rlabel metal2 36792 6440 36792 6440 0 _0744_
rlabel metal2 33320 6384 33320 6384 0 _0745_
rlabel metal3 36624 6776 36624 6776 0 _0746_
rlabel metal2 37912 7448 37912 7448 0 _0747_
rlabel metal3 37352 6664 37352 6664 0 _0748_
rlabel metal2 39144 7056 39144 7056 0 _0749_
rlabel metal2 41048 6552 41048 6552 0 _0750_
rlabel metal2 46088 5880 46088 5880 0 _0751_
rlabel metal2 40264 10192 40264 10192 0 _0752_
rlabel metal2 40432 6440 40432 6440 0 _0753_
rlabel metal3 42560 4872 42560 4872 0 _0754_
rlabel metal2 38696 5376 38696 5376 0 _0755_
rlabel metal2 38920 5488 38920 5488 0 _0756_
rlabel metal2 40152 5600 40152 5600 0 _0757_
rlabel metal2 39816 5768 39816 5768 0 _0758_
rlabel metal2 41272 5992 41272 5992 0 _0759_
rlabel metal2 43960 9352 43960 9352 0 _0760_
rlabel metal2 44072 9968 44072 9968 0 _0761_
rlabel metal2 42616 8260 42616 8260 0 _0762_
rlabel metal2 40936 6160 40936 6160 0 _0763_
rlabel metal2 40040 5992 40040 5992 0 _0764_
rlabel metal2 44184 6664 44184 6664 0 _0765_
rlabel metal2 44296 5320 44296 5320 0 _0766_
rlabel metal2 37240 4088 37240 4088 0 _0767_
rlabel metal3 36120 4312 36120 4312 0 _0768_
rlabel metal2 44632 3920 44632 3920 0 _0769_
rlabel metal3 44464 4200 44464 4200 0 _0770_
rlabel metal2 39312 4312 39312 4312 0 _0771_
rlabel metal2 39088 4200 39088 4200 0 _0772_
rlabel metal3 41216 4312 41216 4312 0 _0773_
rlabel metal2 43624 7784 43624 7784 0 _0774_
rlabel metal2 43960 8204 43960 8204 0 _0775_
rlabel metal2 43176 13104 43176 13104 0 _0776_
rlabel metal2 42616 10416 42616 10416 0 _0777_
rlabel metal3 28672 14392 28672 14392 0 _0778_
rlabel metal2 30184 14952 30184 14952 0 _0779_
rlabel metal2 31192 12656 31192 12656 0 _0780_
rlabel metal3 32256 14504 32256 14504 0 _0781_
rlabel metal2 39984 9800 39984 9800 0 _0782_
rlabel metal2 39368 9800 39368 9800 0 _0783_
rlabel metal2 38360 9856 38360 9856 0 _0784_
rlabel metal2 33544 13832 33544 13832 0 _0785_
rlabel metal3 47992 11256 47992 11256 0 _0786_
rlabel metal2 37912 11088 37912 11088 0 _0787_
rlabel metal2 30632 10360 30632 10360 0 _0788_
rlabel metal2 31192 10304 31192 10304 0 _0789_
rlabel metal2 32088 10192 32088 10192 0 _0790_
rlabel metal2 32536 11032 32536 11032 0 _0791_
rlabel metal2 38416 11480 38416 11480 0 _0792_
rlabel metal2 41160 16464 41160 16464 0 _0793_
rlabel metal2 34216 14392 34216 14392 0 _0794_
rlabel metal2 34608 15512 34608 15512 0 _0795_
rlabel metal3 32368 15288 32368 15288 0 _0796_
rlabel metal3 29680 14504 29680 14504 0 _0797_
rlabel metal2 38136 7728 38136 7728 0 _0798_
rlabel metal2 32312 14056 32312 14056 0 _0799_
rlabel metal2 31640 16464 31640 16464 0 _0800_
rlabel metal2 32144 14728 32144 14728 0 _0801_
rlabel metal2 30520 15344 30520 15344 0 _0802_
rlabel metal2 29512 15008 29512 15008 0 _0803_
rlabel metal2 37016 15344 37016 15344 0 _0804_
rlabel metal2 39424 17640 39424 17640 0 _0805_
rlabel metal2 29624 29344 29624 29344 0 _0806_
rlabel metal2 37688 28784 37688 28784 0 _0807_
rlabel metal2 37240 18032 37240 18032 0 _0808_
rlabel metal2 39984 17640 39984 17640 0 _0809_
rlabel metal2 39256 18144 39256 18144 0 _0810_
rlabel metal3 41440 25368 41440 25368 0 _0811_
rlabel metal2 44856 21336 44856 21336 0 _0812_
rlabel metal2 40936 22400 40936 22400 0 _0813_
rlabel metal3 41720 18424 41720 18424 0 _0814_
rlabel metal2 39928 12712 39928 12712 0 _0815_
rlabel metal2 39816 12880 39816 12880 0 _0816_
rlabel metal2 40824 16520 40824 16520 0 _0817_
rlabel metal2 40488 16072 40488 16072 0 _0818_
rlabel metal3 36064 11592 36064 11592 0 _0819_
rlabel metal2 35448 11480 35448 11480 0 _0820_
rlabel metal2 36008 11872 36008 11872 0 _0821_
rlabel metal2 44632 13384 44632 13384 0 _0822_
rlabel metal2 41720 11256 41720 11256 0 _0823_
rlabel metal2 44072 12376 44072 12376 0 _0824_
rlabel metal2 40936 11480 40936 11480 0 _0825_
rlabel metal2 41608 10472 41608 10472 0 _0826_
rlabel metal2 40936 10472 40936 10472 0 _0827_
rlabel metal2 41384 10584 41384 10584 0 _0828_
rlabel metal2 42056 11760 42056 11760 0 _0829_
rlabel metal2 42616 11984 42616 11984 0 _0830_
rlabel metal2 36680 11480 36680 11480 0 _0831_
rlabel metal2 43736 12488 43736 12488 0 _0832_
rlabel metal2 44296 12488 44296 12488 0 _0833_
rlabel metal2 45360 14952 45360 14952 0 _0834_
rlabel metal2 44632 7980 44632 7980 0 _0835_
rlabel metal3 44016 8904 44016 8904 0 _0836_
rlabel metal2 46984 9184 46984 9184 0 _0837_
rlabel metal3 46928 9128 46928 9128 0 _0838_
rlabel metal2 45192 4032 45192 4032 0 _0839_
rlabel metal2 46984 5040 46984 5040 0 _0840_
rlabel metal3 44240 5096 44240 5096 0 _0841_
rlabel metal2 44968 5488 44968 5488 0 _0842_
rlabel metal2 44408 5600 44408 5600 0 _0843_
rlabel metal2 47432 6496 47432 6496 0 _0844_
rlabel metal3 46984 5096 46984 5096 0 _0845_
rlabel metal2 45752 3640 45752 3640 0 _0846_
rlabel metal2 45976 3920 45976 3920 0 _0847_
rlabel metal2 46312 6272 46312 6272 0 _0848_
rlabel metal2 46536 4536 46536 4536 0 _0849_
rlabel metal2 47488 5096 47488 5096 0 _0850_
rlabel metal2 47936 6664 47936 6664 0 _0851_
rlabel metal2 47432 8204 47432 8204 0 _0852_
rlabel metal2 45304 15568 45304 15568 0 _0853_
rlabel metal3 36960 14504 36960 14504 0 _0854_
rlabel metal3 36120 14280 36120 14280 0 _0855_
rlabel metal3 45024 14504 45024 14504 0 _0856_
rlabel metal2 41160 15848 41160 15848 0 _0857_
rlabel metal2 41664 15960 41664 15960 0 _0858_
rlabel metal2 41440 16184 41440 16184 0 _0859_
rlabel metal2 48888 18424 48888 18424 0 _0860_
rlabel metal2 44408 17528 44408 17528 0 _0861_
rlabel metal2 38808 13104 38808 13104 0 _0862_
rlabel metal2 38248 12656 38248 12656 0 _0863_
rlabel metal2 39816 13440 39816 13440 0 _0864_
rlabel metal2 40264 14448 40264 14448 0 _0865_
rlabel metal2 47936 12376 47936 12376 0 _0866_
rlabel metal2 47656 11928 47656 11928 0 _0867_
rlabel metal3 46760 12376 46760 12376 0 _0868_
rlabel metal3 46704 12936 46704 12936 0 _0869_
rlabel metal2 47264 12824 47264 12824 0 _0870_
rlabel metal2 46984 13776 46984 13776 0 _0871_
rlabel metal2 44800 12152 44800 12152 0 _0872_
rlabel metal2 43624 12824 43624 12824 0 _0873_
rlabel metal3 45920 13608 45920 13608 0 _0874_
rlabel metal2 47320 13832 47320 13832 0 _0875_
rlabel metal2 47712 7560 47712 7560 0 _0876_
rlabel metal2 48048 10584 48048 10584 0 _0877_
rlabel metal2 47544 10192 47544 10192 0 _0878_
rlabel metal2 49224 10864 49224 10864 0 _0879_
rlabel metal2 47544 9296 47544 9296 0 _0880_
rlabel metal3 47768 5208 47768 5208 0 _0881_
rlabel metal2 48216 3808 48216 3808 0 _0882_
rlabel metal2 48216 5992 48216 5992 0 _0883_
rlabel metal2 48328 7420 48328 7420 0 _0884_
rlabel metal2 50232 8176 50232 8176 0 _0885_
rlabel metal2 50792 7672 50792 7672 0 _0886_
rlabel metal2 49224 5880 49224 5880 0 _0887_
rlabel metal2 49336 5824 49336 5824 0 _0888_
rlabel metal2 48776 7728 48776 7728 0 _0889_
rlabel metal2 49000 7000 49000 7000 0 _0890_
rlabel metal2 50344 5600 50344 5600 0 _0891_
rlabel metal2 49616 7000 49616 7000 0 _0892_
rlabel metal2 49728 10472 49728 10472 0 _0893_
rlabel metal2 47768 14728 47768 14728 0 _0894_
rlabel metal2 46200 14840 46200 14840 0 _0895_
rlabel metal2 45192 15176 45192 15176 0 _0896_
rlabel metal3 47264 14616 47264 14616 0 _0897_
rlabel metal2 40376 17416 40376 17416 0 _0898_
rlabel metal2 49112 17192 49112 17192 0 _0899_
rlabel metal2 50008 17752 50008 17752 0 _0900_
rlabel metal2 48664 13440 48664 13440 0 _0901_
rlabel metal3 48440 13720 48440 13720 0 _0902_
rlabel metal3 49448 13832 49448 13832 0 _0903_
rlabel metal2 49896 11760 49896 11760 0 _0904_
rlabel metal2 50456 10640 50456 10640 0 _0905_
rlabel metal2 50232 11648 50232 11648 0 _0906_
rlabel metal3 48552 11928 48552 11928 0 _0907_
rlabel metal2 49728 12040 49728 12040 0 _0908_
rlabel metal2 55944 8904 55944 8904 0 _0909_
rlabel metal2 52808 6160 52808 6160 0 _0910_
rlabel metal3 51352 6664 51352 6664 0 _0911_
rlabel metal2 50232 7056 50232 7056 0 _0912_
rlabel metal2 51128 6888 51128 6888 0 _0913_
rlabel metal2 50848 7336 50848 7336 0 _0914_
rlabel metal2 57288 7616 57288 7616 0 _0915_
rlabel metal2 53480 7952 53480 7952 0 _0916_
rlabel metal2 49336 7896 49336 7896 0 _0917_
rlabel metal2 53592 6720 53592 6720 0 _0918_
rlabel metal2 40376 8316 40376 8316 0 _0919_
rlabel metal2 39536 8232 39536 8232 0 _0920_
rlabel metal3 43680 7056 43680 7056 0 _0921_
rlabel metal2 56672 8232 56672 8232 0 _0922_
rlabel metal2 50680 11984 50680 11984 0 _0923_
rlabel metal3 50204 13720 50204 13720 0 _0924_
rlabel metal2 48552 14784 48552 14784 0 _0925_
rlabel metal2 47600 14504 47600 14504 0 _0926_
rlabel metal2 49224 14840 49224 14840 0 _0927_
rlabel metal2 42728 19096 42728 19096 0 _0928_
rlabel metal2 39592 11872 39592 11872 0 _0929_
rlabel metal2 39872 11368 39872 11368 0 _0930_
rlabel metal2 40040 13496 40040 13496 0 _0931_
rlabel metal2 41160 14504 41160 14504 0 _0932_
rlabel metal2 41384 13944 41384 13944 0 _0933_
rlabel metal2 41944 15288 41944 15288 0 _0934_
rlabel metal3 39900 15400 39900 15400 0 _0935_
rlabel metal2 42504 15344 42504 15344 0 _0936_
rlabel metal2 42168 15792 42168 15792 0 _0937_
rlabel metal3 43176 16184 43176 16184 0 _0938_
rlabel metal3 49000 19992 49000 19992 0 _0939_
rlabel metal2 40152 16072 40152 16072 0 _0940_
rlabel metal2 50456 14168 50456 14168 0 _0941_
rlabel metal2 51296 13944 51296 13944 0 _0942_
rlabel metal2 53144 15680 53144 15680 0 _0943_
rlabel metal2 56336 9016 56336 9016 0 _0944_
rlabel metal2 55440 12712 55440 12712 0 _0945_
rlabel metal2 50120 12544 50120 12544 0 _0946_
rlabel metal2 55608 13104 55608 13104 0 _0947_
rlabel metal3 54040 11256 54040 11256 0 _0948_
rlabel metal2 54264 8120 54264 8120 0 _0949_
rlabel metal2 53872 8232 53872 8232 0 _0950_
rlabel metal2 54600 7784 54600 7784 0 _0951_
rlabel metal2 55608 10472 55608 10472 0 _0952_
rlabel metal2 56056 10136 56056 10136 0 _0953_
rlabel metal3 53368 9800 53368 9800 0 _0954_
rlabel metal2 40936 9744 40936 9744 0 _0955_
rlabel metal2 53704 9744 53704 9744 0 _0956_
rlabel metal2 57512 10640 57512 10640 0 _0957_
rlabel metal2 57288 13272 57288 13272 0 _0958_
rlabel metal2 52920 15624 52920 15624 0 _0959_
rlabel metal2 52808 16464 52808 16464 0 _0960_
rlabel metal3 43736 16744 43736 16744 0 _0961_
rlabel metal3 45864 18424 45864 18424 0 _0962_
rlabel metal2 34384 16184 34384 16184 0 _0963_
rlabel metal2 55832 12712 55832 12712 0 _0964_
rlabel metal2 56728 13048 56728 13048 0 _0965_
rlabel metal2 54488 13104 54488 13104 0 _0966_
rlabel metal2 52248 13104 52248 13104 0 _0967_
rlabel metal2 53368 10864 53368 10864 0 _0968_
rlabel metal2 53424 11368 53424 11368 0 _0969_
rlabel metal2 54936 10080 54936 10080 0 _0970_
rlabel metal2 55104 11256 55104 11256 0 _0971_
rlabel metal2 55944 10696 55944 10696 0 _0972_
rlabel metal2 54600 10864 54600 10864 0 _0973_
rlabel metal2 55720 11424 55720 11424 0 _0974_
rlabel metal2 53536 12936 53536 12936 0 _0975_
rlabel metal2 54264 14056 54264 14056 0 _0976_
rlabel metal2 52024 14560 52024 14560 0 _0977_
rlabel metal2 53368 14392 53368 14392 0 _0978_
rlabel metal2 52136 19040 52136 19040 0 _0979_
rlabel metal2 51744 15960 51744 15960 0 _0980_
rlabel metal2 38696 19628 38696 19628 0 _0981_
rlabel metal2 35280 15960 35280 15960 0 _0982_
rlabel metal2 35168 16184 35168 16184 0 _0983_
rlabel metal2 43176 20720 43176 20720 0 _0984_
rlabel metal3 33712 16856 33712 16856 0 _0985_
rlabel metal2 32536 16464 32536 16464 0 _0986_
rlabel metal2 32144 16072 32144 16072 0 _0987_
rlabel metal2 51856 17416 51856 17416 0 _0988_
rlabel metal2 52024 16576 52024 16576 0 _0989_
rlabel metal3 51744 16856 51744 16856 0 _0990_
rlabel metal3 33712 15176 33712 15176 0 _0991_
rlabel metal3 32256 16184 32256 16184 0 _0992_
rlabel metal2 30184 17528 30184 17528 0 _0993_
rlabel metal2 52248 18312 52248 18312 0 _0994_
rlabel metal2 51240 18088 51240 18088 0 _0995_
rlabel metal2 51688 18088 51688 18088 0 _0996_
rlabel metal2 39032 18256 39032 18256 0 _0997_
rlabel metal2 29176 15736 29176 15736 0 _0998_
rlabel metal2 29848 16128 29848 16128 0 _0999_
rlabel metal2 29288 16464 29288 16464 0 _1000_
rlabel metal2 37968 18648 37968 18648 0 _1001_
rlabel metal3 36792 19096 36792 19096 0 _1002_
rlabel metal3 41496 22344 41496 22344 0 _1003_
rlabel metal2 46088 22904 46088 22904 0 _1004_
rlabel metal2 29400 26180 29400 26180 0 _1005_
rlabel metal2 30072 23800 30072 23800 0 _1006_
rlabel metal2 26264 20272 26264 20272 0 _1007_
rlabel metal2 26824 21784 26824 21784 0 _1008_
rlabel metal2 6440 11984 6440 11984 0 _1009_
rlabel metal2 14280 12152 14280 12152 0 _1010_
rlabel metal2 13944 11200 13944 11200 0 _1011_
rlabel metal2 5880 12208 5880 12208 0 _1012_
rlabel metal2 6552 12376 6552 12376 0 _1013_
rlabel metal2 3640 12376 3640 12376 0 _1014_
rlabel metal2 7560 12544 7560 12544 0 _1015_
rlabel metal3 6720 11368 6720 11368 0 _1016_
rlabel metal2 6888 13496 6888 13496 0 _1017_
rlabel metal2 7448 12712 7448 12712 0 _1018_
rlabel metal2 7784 12712 7784 12712 0 _1019_
rlabel metal2 8344 13272 8344 13272 0 _1020_
rlabel metal2 8848 12376 8848 12376 0 _1021_
rlabel metal3 10080 12824 10080 12824 0 _1022_
rlabel metal3 8008 11984 8008 11984 0 _1023_
rlabel metal2 10360 12600 10360 12600 0 _1024_
rlabel metal2 11480 10248 11480 10248 0 _1025_
rlabel metal2 11368 13328 11368 13328 0 _1026_
rlabel metal2 11704 12432 11704 12432 0 _1027_
rlabel metal2 4536 7896 4536 7896 0 _1028_
rlabel metal2 3864 9856 3864 9856 0 _1029_
rlabel metal2 7336 8316 7336 8316 0 _1030_
rlabel metal2 8064 7448 8064 7448 0 _1031_
rlabel metal2 7000 9856 7000 9856 0 _1032_
rlabel metal2 9800 10136 9800 10136 0 _1033_
rlabel metal2 9912 10528 9912 10528 0 _1034_
rlabel metal2 10136 13048 10136 13048 0 _1035_
rlabel metal2 11088 11144 11088 11144 0 _1036_
rlabel metal2 12488 10864 12488 10864 0 _1037_
rlabel metal3 11256 10024 11256 10024 0 _1038_
rlabel metal2 11816 10416 11816 10416 0 _1039_
rlabel metal2 13776 10360 13776 10360 0 _1040_
rlabel metal2 10024 23744 10024 23744 0 _1041_
rlabel metal2 8344 18760 8344 18760 0 _1042_
rlabel metal2 18536 18760 18536 18760 0 _1043_
rlabel metal2 4984 14448 4984 14448 0 _1044_
rlabel metal2 6552 14392 6552 14392 0 _1045_
rlabel metal2 4312 21448 4312 21448 0 _1046_
rlabel metal2 2184 15568 2184 15568 0 _1047_
rlabel metal2 2632 14896 2632 14896 0 _1048_
rlabel metal2 3080 17752 3080 17752 0 _1049_
rlabel metal2 3528 14560 3528 14560 0 _1050_
rlabel metal2 2968 15344 2968 15344 0 _1051_
rlabel metal2 2856 17472 2856 17472 0 _1052_
rlabel metal2 7392 15512 7392 15512 0 _1053_
rlabel metal3 5880 13944 5880 13944 0 _1054_
rlabel metal2 4872 16296 4872 16296 0 _1055_
rlabel metal2 3304 9576 3304 9576 0 _1056_
rlabel metal2 5656 17528 5656 17528 0 _1057_
rlabel metal2 10472 16240 10472 16240 0 _1058_
rlabel metal2 5544 16184 5544 16184 0 _1059_
rlabel metal2 3080 18984 3080 18984 0 _1060_
rlabel metal2 2856 19152 2856 19152 0 _1061_
rlabel metal2 3248 20888 3248 20888 0 _1062_
rlabel metal2 2352 17640 2352 17640 0 _1063_
rlabel metal2 2968 16800 2968 16800 0 _1064_
rlabel metal3 8288 16072 8288 16072 0 _1065_
rlabel metal2 3416 16800 3416 16800 0 _1066_
rlabel metal2 3192 21672 3192 21672 0 _1067_
rlabel metal3 2576 22344 2576 22344 0 _1068_
rlabel metal2 3080 23184 3080 23184 0 _1069_
rlabel metal2 3416 22792 3416 22792 0 _1070_
rlabel metal2 3976 20496 3976 20496 0 _1071_
rlabel metal2 3640 20048 3640 20048 0 _1072_
rlabel metal2 4256 20776 4256 20776 0 _1073_
rlabel metal2 15960 18088 15960 18088 0 _1074_
rlabel metal2 4536 17360 4536 17360 0 _1075_
rlabel metal2 6216 17696 6216 17696 0 _1076_
rlabel metal2 5880 17416 5880 17416 0 _1077_
rlabel metal2 7784 19376 7784 19376 0 _1078_
rlabel metal2 7448 19824 7448 19824 0 _1079_
rlabel metal2 6384 20776 6384 20776 0 _1080_
rlabel metal3 5152 19992 5152 19992 0 _1081_
rlabel metal2 5040 20104 5040 20104 0 _1082_
rlabel metal3 5376 22456 5376 22456 0 _1083_
rlabel metal2 10136 23968 10136 23968 0 _1084_
rlabel metal2 10864 23800 10864 23800 0 _1085_
rlabel metal3 11480 23688 11480 23688 0 _1086_
rlabel metal2 15848 20608 15848 20608 0 _1087_
rlabel metal2 15456 20104 15456 20104 0 _1088_
rlabel metal2 12712 14252 12712 14252 0 _1089_
rlabel metal2 14504 20160 14504 20160 0 _1090_
rlabel metal2 17528 20048 17528 20048 0 _1091_
rlabel metal2 14672 20216 14672 20216 0 _1092_
rlabel metal3 16184 21112 16184 21112 0 _1093_
rlabel metal2 15960 22064 15960 22064 0 _1094_
rlabel metal2 16296 17248 16296 17248 0 _1095_
rlabel metal2 15400 16632 15400 16632 0 _1096_
rlabel metal2 16296 18144 16296 18144 0 _1097_
rlabel metal2 10136 17920 10136 17920 0 _1098_
rlabel metal2 13608 17696 13608 17696 0 _1099_
rlabel metal2 4984 18032 4984 18032 0 _1100_
rlabel metal2 17640 19432 17640 19432 0 _1101_
rlabel metal2 11256 14728 11256 14728 0 _1102_
rlabel metal2 15064 17920 15064 17920 0 _1103_
rlabel metal2 15288 18088 15288 18088 0 _1104_
rlabel metal2 15624 18704 15624 18704 0 _1105_
rlabel metal2 14112 20888 14112 20888 0 _1106_
rlabel metal2 15400 21560 15400 21560 0 _1107_
rlabel metal2 14616 22288 14616 22288 0 _1108_
rlabel metal3 14168 22344 14168 22344 0 _1109_
rlabel metal2 10696 12992 10696 12992 0 _1110_
rlabel metal2 11032 13496 11032 13496 0 _1111_
rlabel metal2 11032 22120 11032 22120 0 _1112_
rlabel metal2 12152 22680 12152 22680 0 _1113_
rlabel metal2 11480 22344 11480 22344 0 _1114_
rlabel metal2 12040 23912 12040 23912 0 _1115_
rlabel metal2 10920 24248 10920 24248 0 _1116_
rlabel metal2 15512 23240 15512 23240 0 _1117_
rlabel via2 6664 23688 6664 23688 0 _1118_
rlabel metal2 3976 22064 3976 22064 0 _1119_
rlabel metal2 4984 23184 4984 23184 0 _1120_
rlabel metal2 7896 23072 7896 23072 0 _1121_
rlabel metal3 18424 15400 18424 15400 0 _1122_
rlabel metal2 8904 22288 8904 22288 0 _1123_
rlabel metal2 3640 17248 3640 17248 0 _1124_
rlabel metal2 7224 21112 7224 21112 0 _1125_
rlabel metal2 5992 23072 5992 23072 0 _1126_
rlabel metal2 12824 14448 12824 14448 0 _1127_
rlabel metal2 18872 16744 18872 16744 0 _1128_
rlabel metal2 8904 20832 8904 20832 0 _1129_
rlabel metal3 9072 16968 9072 16968 0 _1130_
rlabel metal2 11816 15960 11816 15960 0 _1131_
rlabel metal2 10024 16968 10024 16968 0 _1132_
rlabel metal2 9576 16576 9576 16576 0 _1133_
rlabel metal2 8792 18872 8792 18872 0 _1134_
rlabel metal2 7280 22344 7280 22344 0 _1135_
rlabel metal2 8344 23520 8344 23520 0 _1136_
rlabel metal3 11424 23800 11424 23800 0 _1137_
rlabel metal2 14056 10920 14056 10920 0 _1138_
rlabel metal3 13384 10360 13384 10360 0 _1139_
rlabel metal2 11144 10136 11144 10136 0 _1140_
rlabel metal3 13216 8232 13216 8232 0 _1141_
rlabel metal2 8344 8176 8344 8176 0 _1142_
rlabel metal2 6216 10024 6216 10024 0 _1143_
rlabel metal2 6328 10696 6328 10696 0 _1144_
rlabel metal2 7560 7616 7560 7616 0 _1145_
rlabel metal2 8008 8624 8008 8624 0 _1146_
rlabel metal3 5376 8232 5376 8232 0 _1147_
rlabel metal2 5712 7448 5712 7448 0 _1148_
rlabel metal2 7112 8176 7112 8176 0 _1149_
rlabel metal3 11928 8344 11928 8344 0 _1150_
rlabel metal2 14392 10696 14392 10696 0 _1151_
rlabel metal2 14504 12432 14504 12432 0 _1152_
rlabel metal2 15512 24696 15512 24696 0 _1153_
rlabel metal2 15288 23576 15288 23576 0 _1154_
rlabel metal2 20440 24248 20440 24248 0 _1155_
rlabel metal2 24808 23464 24808 23464 0 _1156_
rlabel metal2 16968 20328 16968 20328 0 _1157_
rlabel metal2 25704 20944 25704 20944 0 _1158_
rlabel metal2 28280 31640 28280 31640 0 _1159_
rlabel metal2 25480 24304 25480 24304 0 _1160_
rlabel metal2 29176 24192 29176 24192 0 _1161_
rlabel metal2 29736 24416 29736 24416 0 _1162_
rlabel metal3 29120 27048 29120 27048 0 _1163_
rlabel metal3 29848 24808 29848 24808 0 _1164_
rlabel metal2 41496 22176 41496 22176 0 _1165_
rlabel metal2 39312 22344 39312 22344 0 _1166_
rlabel metal3 43568 23912 43568 23912 0 _1167_
rlabel metal2 39480 23184 39480 23184 0 _1168_
rlabel metal2 26376 24360 26376 24360 0 _1169_
rlabel metal2 10136 21056 10136 21056 0 _1170_
rlabel metal2 8456 22456 8456 22456 0 _1171_
rlabel metal2 9016 22848 9016 22848 0 _1172_
rlabel metal2 12376 21616 12376 21616 0 _1173_
rlabel metal2 11144 19768 11144 19768 0 _1174_
rlabel metal2 11368 17360 11368 17360 0 _1175_
rlabel metal2 17752 16912 17752 16912 0 _1176_
rlabel metal2 11592 17528 11592 17528 0 _1177_
rlabel metal2 10752 18424 10752 18424 0 _1178_
rlabel metal2 10808 17976 10808 17976 0 _1179_
rlabel metal2 11144 18536 11144 18536 0 _1180_
rlabel metal3 11984 19208 11984 19208 0 _1181_
rlabel metal2 9912 22008 9912 22008 0 _1182_
rlabel metal2 12040 19936 12040 19936 0 _1183_
rlabel metal2 12488 21112 12488 21112 0 _1184_
rlabel metal2 21672 22008 21672 22008 0 _1185_
rlabel metal2 14504 8848 14504 8848 0 _1186_
rlabel metal2 15064 10136 15064 10136 0 _1187_
rlabel metal2 21000 9408 21000 9408 0 _1188_
rlabel metal2 18760 9408 18760 9408 0 _1189_
rlabel metal2 13944 7336 13944 7336 0 _1190_
rlabel metal2 13608 7168 13608 7168 0 _1191_
rlabel metal3 10024 7672 10024 7672 0 _1192_
rlabel metal3 11816 7448 11816 7448 0 _1193_
rlabel metal2 11928 7728 11928 7728 0 _1194_
rlabel metal2 18872 7728 18872 7728 0 _1195_
rlabel metal2 14952 8568 14952 8568 0 _1196_
rlabel metal3 7196 7224 7196 7224 0 _1197_
rlabel metal2 15064 6720 15064 6720 0 _1198_
rlabel metal2 3752 11536 3752 11536 0 _1199_
rlabel metal2 3864 11760 3864 11760 0 _1200_
rlabel metal2 14840 7728 14840 7728 0 _1201_
rlabel metal2 19880 9184 19880 9184 0 _1202_
rlabel metal2 20944 9800 20944 9800 0 _1203_
rlabel metal2 21336 21336 21336 21336 0 _1204_
rlabel metal3 15456 23912 15456 23912 0 _1205_
rlabel metal3 19600 23128 19600 23128 0 _1206_
rlabel metal2 26152 23408 26152 23408 0 _1207_
rlabel metal2 18368 22344 18368 22344 0 _1208_
rlabel metal2 17416 22176 17416 22176 0 _1209_
rlabel metal2 19096 23184 19096 23184 0 _1210_
rlabel metal2 27832 24416 27832 24416 0 _1211_
rlabel metal2 27720 24528 27720 24528 0 _1212_
rlabel metal2 39256 23240 39256 23240 0 _1213_
rlabel metal2 39032 22848 39032 22848 0 _1214_
rlabel metal3 40936 23016 40936 23016 0 _1215_
rlabel metal2 42616 23520 42616 23520 0 _1216_
rlabel metal2 32648 23632 32648 23632 0 _1217_
rlabel metal2 11592 21056 11592 21056 0 _1218_
rlabel metal2 10472 21784 10472 21784 0 _1219_
rlabel metal2 21448 20776 21448 20776 0 _1220_
rlabel metal2 22120 17976 22120 17976 0 _1221_
rlabel metal2 20440 19376 20440 19376 0 _1222_
rlabel metal2 20552 19656 20552 19656 0 _1223_
rlabel metal2 21560 20272 21560 20272 0 _1224_
rlabel metal2 23128 21168 23128 21168 0 _1225_
rlabel metal2 19712 8120 19712 8120 0 _1226_
rlabel metal2 22120 8792 22120 8792 0 _1227_
rlabel metal2 22008 9240 22008 9240 0 _1228_
rlabel metal2 22344 9912 22344 9912 0 _1229_
rlabel metal2 21784 12992 21784 12992 0 _1230_
rlabel metal2 21112 11704 21112 11704 0 _1231_
rlabel metal2 15736 8344 15736 8344 0 _1232_
rlabel metal3 15512 7336 15512 7336 0 _1233_
rlabel metal2 16520 8344 16520 8344 0 _1234_
rlabel metal2 20328 10976 20328 10976 0 _1235_
rlabel metal2 18368 17640 18368 17640 0 _1236_
rlabel metal2 18312 12376 18312 12376 0 _1237_
rlabel metal3 10052 11480 10052 11480 0 _1238_
rlabel metal3 17136 10472 17136 10472 0 _1239_
rlabel metal2 12936 13608 12936 13608 0 _1240_
rlabel metal2 12656 13720 12656 13720 0 _1241_
rlabel metal2 13608 12600 13608 12600 0 _1242_
rlabel metal2 21448 11760 21448 11760 0 _1243_
rlabel metal2 22792 10808 22792 10808 0 _1244_
rlabel metal2 23352 20748 23352 20748 0 _1245_
rlabel metal2 22232 21840 22232 21840 0 _1246_
rlabel metal2 22120 21672 22120 21672 0 _1247_
rlabel metal2 22680 22792 22680 22792 0 _1248_
rlabel metal2 25032 23296 25032 23296 0 _1249_
rlabel metal2 17192 21000 17192 21000 0 _1250_
rlabel metal2 17640 21000 17640 21000 0 _1251_
rlabel metal2 19208 21280 19208 21280 0 _1252_
rlabel metal2 18760 25200 18760 25200 0 _1253_
rlabel metal2 38136 23016 38136 23016 0 _1254_
rlabel metal3 43736 23464 43736 23464 0 _1255_
rlabel metal2 47096 24024 47096 24024 0 _1256_
rlabel metal2 20104 18648 20104 18648 0 _1257_
rlabel metal2 19880 18592 19880 18592 0 _1258_
rlabel metal2 22792 18760 22792 18760 0 _1259_
rlabel metal3 22176 16072 22176 16072 0 _1260_
rlabel metal2 22288 12264 22288 12264 0 _1261_
rlabel metal2 23128 13888 23128 13888 0 _1262_
rlabel metal2 23240 11956 23240 11956 0 _1263_
rlabel metal2 23688 13216 23688 13216 0 _1264_
rlabel metal2 19712 12376 19712 12376 0 _1265_
rlabel metal2 15064 14112 15064 14112 0 _1266_
rlabel metal2 14616 13664 14616 13664 0 _1267_
rlabel metal2 17192 11480 17192 11480 0 _1268_
rlabel metal2 17640 11256 17640 11256 0 _1269_
rlabel metal2 18536 11872 18536 11872 0 _1270_
rlabel metal2 18760 12320 18760 12320 0 _1271_
rlabel metal2 16184 14056 16184 14056 0 _1272_
rlabel metal2 14504 13944 14504 13944 0 _1273_
rlabel metal2 15680 15848 15680 15848 0 _1274_
rlabel metal2 13720 15680 13720 15680 0 _1275_
rlabel metal2 13104 15288 13104 15288 0 _1276_
rlabel metal2 17416 13720 17416 13720 0 _1277_
rlabel metal3 18760 14616 18760 14616 0 _1278_
rlabel metal3 22008 12936 22008 12936 0 _1279_
rlabel metal2 23576 18032 23576 18032 0 _1280_
rlabel metal3 23912 20104 23912 20104 0 _1281_
rlabel metal2 24136 20216 24136 20216 0 _1282_
rlabel metal3 25592 19096 25592 19096 0 _1283_
rlabel metal2 26488 22064 26488 22064 0 _1284_
rlabel metal2 18872 18872 18872 18872 0 _1285_
rlabel metal2 16968 18928 16968 18928 0 _1286_
rlabel metal2 17528 19488 17528 19488 0 _1287_
rlabel metal2 18200 18928 18200 18928 0 _1288_
rlabel metal2 18760 19152 18760 19152 0 _1289_
rlabel metal2 19320 20552 19320 20552 0 _1290_
rlabel metal2 19152 25704 19152 25704 0 _1291_
rlabel metal2 18760 29176 18760 29176 0 _1292_
rlabel metal3 28728 22176 28728 22176 0 _1293_
rlabel metal2 43064 21000 43064 21000 0 _1294_
rlabel metal2 44184 21616 44184 21616 0 _1295_
rlabel metal2 39480 25424 39480 25424 0 _1296_
rlabel metal2 16688 25256 16688 25256 0 _1297_
rlabel metal2 42056 25424 42056 25424 0 _1298_
rlabel metal2 38696 30352 38696 30352 0 _1299_
rlabel metal3 16688 26376 16688 26376 0 _1300_
rlabel metal2 23688 19320 23688 19320 0 _1301_
rlabel metal2 22792 19712 22792 19712 0 _1302_
rlabel metal2 23240 19600 23240 19600 0 _1303_
rlabel metal2 20160 14392 20160 14392 0 _1304_
rlabel metal3 22736 14280 22736 14280 0 _1305_
rlabel metal3 24360 13720 24360 13720 0 _1306_
rlabel metal2 25256 14504 25256 14504 0 _1307_
rlabel metal3 22120 14392 22120 14392 0 _1308_
rlabel metal2 16856 16408 16856 16408 0 _1309_
rlabel metal2 15176 14224 15176 14224 0 _1310_
rlabel metal3 17864 13720 17864 13720 0 _1311_
rlabel metal3 21504 15512 21504 15512 0 _1312_
rlabel metal2 18536 17192 18536 17192 0 _1313_
rlabel metal2 17752 15624 17752 15624 0 _1314_
rlabel metal2 16072 16520 16072 16520 0 _1315_
rlabel metal2 20664 15456 20664 15456 0 _1316_
rlabel metal3 21784 15288 21784 15288 0 _1317_
rlabel metal2 25704 14560 25704 14560 0 _1318_
rlabel metal2 26376 15148 26376 15148 0 _1319_
rlabel metal2 40376 25984 40376 25984 0 _1320_
rlabel metal2 23072 24920 23072 24920 0 _1321_
rlabel metal3 28952 26376 28952 26376 0 _1322_
rlabel metal3 18872 28056 18872 28056 0 _1323_
rlabel metal2 29736 25928 29736 25928 0 _1324_
rlabel metal2 41608 25144 41608 25144 0 _1325_
rlabel metal2 41944 25536 41944 25536 0 _1326_
rlabel metal3 29008 20776 29008 20776 0 _1327_
rlabel metal2 32424 24584 32424 24584 0 _1328_
rlabel metal2 28280 19376 28280 19376 0 _1329_
rlabel metal2 23296 15288 23296 15288 0 _1330_
rlabel metal2 25928 15680 25928 15680 0 _1331_
rlabel metal2 25648 16632 25648 16632 0 _1332_
rlabel metal2 26376 16352 26376 16352 0 _1333_
rlabel metal2 24024 15904 24024 15904 0 _1334_
rlabel metal3 22904 17640 22904 17640 0 _1335_
rlabel metal2 24024 16912 24024 16912 0 _1336_
rlabel metal2 17640 16632 17640 16632 0 _1337_
rlabel metal3 17640 16632 17640 16632 0 _1338_
rlabel metal2 18424 15792 18424 15792 0 _1339_
rlabel metal2 18200 16408 18200 16408 0 _1340_
rlabel metal2 23800 16520 23800 16520 0 _1341_
rlabel metal2 26208 15512 26208 15512 0 _1342_
rlabel metal2 27048 18704 27048 18704 0 _1343_
rlabel metal2 32088 23800 32088 23800 0 _1344_
rlabel metal2 15288 22232 15288 22232 0 _1345_
rlabel metal2 16520 22344 16520 22344 0 _1346_
rlabel metal3 18648 22792 18648 22792 0 _1347_
rlabel metal2 33544 32032 33544 32032 0 _1348_
rlabel metal2 31640 25088 31640 25088 0 _1349_
rlabel metal2 37576 23128 37576 23128 0 _1350_
rlabel metal2 38360 21168 38360 21168 0 _1351_
rlabel metal2 38248 22176 38248 22176 0 _1352_
rlabel metal2 38360 22512 38360 22512 0 _1353_
rlabel metal2 29064 19600 29064 19600 0 _1354_
rlabel metal2 24528 16968 24528 16968 0 _1355_
rlabel metal2 26600 17304 26600 17304 0 _1356_
rlabel metal2 26208 15288 26208 15288 0 _1357_
rlabel metal2 26824 17360 26824 17360 0 _1358_
rlabel metal2 26488 17472 26488 17472 0 _1359_
rlabel metal2 28840 19376 28840 19376 0 _1360_
rlabel metal3 31472 23800 31472 23800 0 _1361_
rlabel metal2 23912 22064 23912 22064 0 _1362_
rlabel metal2 33488 21000 33488 21000 0 _1363_
rlabel metal2 35952 20888 35952 20888 0 _1364_
rlabel metal3 34384 20776 34384 20776 0 _1365_
rlabel metal2 34104 21560 34104 21560 0 _1366_
rlabel metal2 26600 18200 26600 18200 0 _1367_
rlabel metal2 29624 19208 29624 19208 0 _1368_
rlabel metal3 31920 20552 31920 20552 0 _1369_
rlabel metal2 24696 24640 24696 24640 0 _1370_
rlabel metal2 25368 23856 25368 23856 0 _1371_
rlabel metal2 34328 20216 34328 20216 0 _1372_
rlabel metal2 32648 19992 32648 19992 0 _1373_
rlabel metal2 19320 41104 19320 41104 0 _1374_
rlabel metal2 18872 40824 18872 40824 0 _1375_
rlabel metal3 21336 41160 21336 41160 0 _1376_
rlabel metal2 11144 45136 11144 45136 0 _1377_
rlabel metal2 13832 45584 13832 45584 0 _1378_
rlabel metal2 16856 45248 16856 45248 0 _1379_
rlabel metal2 14280 45248 14280 45248 0 _1380_
rlabel metal2 22232 45080 22232 45080 0 _1381_
rlabel metal3 13104 44072 13104 44072 0 _1382_
rlabel metal2 11928 42280 11928 42280 0 _1383_
rlabel metal2 10472 42168 10472 42168 0 _1384_
rlabel metal2 11256 39200 11256 39200 0 _1385_
rlabel metal3 10920 42728 10920 42728 0 _1386_
rlabel metal2 11144 42784 11144 42784 0 _1387_
rlabel metal2 11704 42224 11704 42224 0 _1388_
rlabel metal2 21000 43064 21000 43064 0 _1389_
rlabel metal2 22792 43736 22792 43736 0 _1390_
rlabel metal3 24920 38920 24920 38920 0 _1391_
rlabel metal2 23296 44296 23296 44296 0 _1392_
rlabel metal2 22120 44240 22120 44240 0 _1393_
rlabel metal2 22232 43792 22232 43792 0 _1394_
rlabel metal3 17192 45192 17192 45192 0 _1395_
rlabel metal2 18200 45192 18200 45192 0 _1396_
rlabel metal2 8008 44296 8008 44296 0 _1397_
rlabel metal3 11368 44408 11368 44408 0 _1398_
rlabel metal2 12488 44632 12488 44632 0 _1399_
rlabel metal3 17304 45080 17304 45080 0 _1400_
rlabel metal3 21168 44296 21168 44296 0 _1401_
rlabel metal2 23128 42616 23128 42616 0 _1402_
rlabel metal2 24024 39844 24024 39844 0 _1403_
rlabel metal3 5096 38808 5096 38808 0 _1404_
rlabel metal2 6384 38920 6384 38920 0 _1405_
rlabel metal2 6440 41216 6440 41216 0 _1406_
rlabel metal2 6608 38920 6608 38920 0 _1407_
rlabel metal2 6440 38248 6440 38248 0 _1408_
rlabel metal2 5880 39256 5880 39256 0 _1409_
rlabel metal2 7672 41888 7672 41888 0 _1410_
rlabel metal2 5768 38752 5768 38752 0 _1411_
rlabel metal2 6104 38472 6104 38472 0 _1412_
rlabel metal3 7112 39704 7112 39704 0 _1413_
rlabel metal2 8512 38024 8512 38024 0 _1414_
rlabel metal2 9576 31472 9576 31472 0 _1415_
rlabel metal3 11144 40376 11144 40376 0 _1416_
rlabel metal2 12264 40432 12264 40432 0 _1417_
rlabel metal2 8848 37352 8848 37352 0 _1418_
rlabel metal2 8792 36512 8792 36512 0 _1419_
rlabel metal2 8232 40264 8232 40264 0 _1420_
rlabel metal2 7112 36008 7112 36008 0 _1421_
rlabel metal2 5208 40096 5208 40096 0 _1422_
rlabel metal2 4424 39704 4424 39704 0 _1423_
rlabel metal2 5376 39592 5376 39592 0 _1424_
rlabel metal2 4760 39368 4760 39368 0 _1425_
rlabel metal3 4648 41160 4648 41160 0 _1426_
rlabel metal2 2632 40768 2632 40768 0 _1427_
rlabel metal2 3192 41160 3192 41160 0 _1428_
rlabel metal2 4648 38976 4648 38976 0 _1429_
rlabel metal2 7448 35728 7448 35728 0 _1430_
rlabel metal3 8456 35784 8456 35784 0 _1431_
rlabel metal2 11704 30912 11704 30912 0 _1432_
rlabel metal2 8792 39144 8792 39144 0 _1433_
rlabel metal2 8232 34328 8232 34328 0 _1434_
rlabel metal2 4200 35112 4200 35112 0 _1435_
rlabel metal2 16520 37520 16520 37520 0 _1436_
rlabel metal3 5544 35784 5544 35784 0 _1437_
rlabel metal2 7112 40096 7112 40096 0 _1438_
rlabel metal2 2744 39088 2744 39088 0 _1439_
rlabel metal2 2968 37576 2968 37576 0 _1440_
rlabel metal2 2184 39144 2184 39144 0 _1441_
rlabel metal2 2744 37016 2744 37016 0 _1442_
rlabel metal2 2856 36512 2856 36512 0 _1443_
rlabel metal2 2632 35952 2632 35952 0 _1444_
rlabel metal2 2408 34888 2408 34888 0 _1445_
rlabel metal2 2744 33208 2744 33208 0 _1446_
rlabel metal2 7000 33992 7000 33992 0 _1447_
rlabel metal2 3752 33376 3752 33376 0 _1448_
rlabel metal2 3304 34552 3304 34552 0 _1449_
rlabel metal2 4424 35000 4424 35000 0 _1450_
rlabel metal2 22400 34888 22400 34888 0 _1451_
rlabel metal2 22792 34944 22792 34944 0 _1452_
rlabel metal2 23688 43064 23688 43064 0 _1453_
rlabel metal2 24136 43288 24136 43288 0 _1454_
rlabel metal2 24472 35392 24472 35392 0 _1455_
rlabel metal2 26096 34888 26096 34888 0 _1456_
rlabel metal3 24584 38024 24584 38024 0 _1457_
rlabel metal2 11648 40376 11648 40376 0 _1458_
rlabel metal2 10248 40432 10248 40432 0 _1459_
rlabel metal2 16856 39256 16856 39256 0 _1460_
rlabel metal2 23912 37912 23912 37912 0 _1461_
rlabel metal2 25592 38360 25592 38360 0 _1462_
rlabel metal2 25928 37632 25928 37632 0 _1463_
rlabel metal3 8400 36344 8400 36344 0 _1464_
rlabel metal2 10360 36960 10360 36960 0 _1465_
rlabel metal2 10248 37072 10248 37072 0 _1466_
rlabel metal2 10640 38024 10640 38024 0 _1467_
rlabel metal2 10136 38360 10136 38360 0 _1468_
rlabel metal2 11592 37576 11592 37576 0 _1469_
rlabel metal2 23576 37352 23576 37352 0 _1470_
rlabel metal3 21840 37240 21840 37240 0 _1471_
rlabel metal2 24584 36848 24584 36848 0 _1472_
rlabel metal2 24472 37576 24472 37576 0 _1473_
rlabel metal2 26040 36344 26040 36344 0 _1474_
rlabel metal3 25088 35672 25088 35672 0 _1475_
rlabel metal2 25536 34328 25536 34328 0 _1476_
rlabel metal2 23464 35168 23464 35168 0 _1477_
rlabel metal3 23128 28504 23128 28504 0 _1478_
rlabel metal2 3528 36736 3528 36736 0 _1479_
rlabel metal2 3864 36792 3864 36792 0 _1480_
rlabel metal2 4088 35000 4088 35000 0 _1481_
rlabel metal2 44968 24472 44968 24472 0 active
rlabel metal2 15288 27160 15288 27160 0 clk
rlabel metal1 26712 25256 26712 25256 0 clknet_0_clk
rlabel metal2 25368 21616 25368 21616 0 clknet_2_0__leaf_clk
rlabel metal2 17864 25088 17864 25088 0 clknet_2_1__leaf_clk
rlabel metal2 38808 19712 38808 19712 0 clknet_2_2__leaf_clk
rlabel metal2 38696 23520 38696 23520 0 clknet_2_3__leaf_clk
rlabel metal2 54936 32424 54936 32424 0 net1
rlabel metal2 57848 27608 57848 27608 0 net10
rlabel metal2 21336 24192 21336 24192 0 net100
rlabel metal2 38136 28336 38136 28336 0 net101
rlabel metal2 36904 45360 36904 45360 0 net102
rlabel metal2 54040 30072 54040 30072 0 net103
rlabel metal2 55160 24808 55160 24808 0 net104
rlabel metal2 49672 16352 49672 16352 0 net105
rlabel metal2 53480 24528 53480 24528 0 net106
rlabel metal2 53704 20440 53704 20440 0 net107
rlabel metal2 49672 19488 49672 19488 0 net108
rlabel metal2 47768 18872 47768 18872 0 net109
rlabel metal3 51016 37520 51016 37520 0 net11
rlabel metal2 39704 6384 39704 6384 0 net110
rlabel metal2 31304 16800 31304 16800 0 net111
rlabel metal3 50568 17808 50568 17808 0 net112
rlabel metal2 53480 23072 53480 23072 0 net113
rlabel metal3 45584 19880 45584 19880 0 net114
rlabel metal2 52136 24304 52136 24304 0 net115
rlabel metal2 55608 26768 55608 26768 0 net116
rlabel metal2 21560 2030 21560 2030 0 net117
rlabel metal2 57736 32536 57736 32536 0 net12
rlabel metal2 52136 29008 52136 29008 0 net13
rlabel metal3 56896 34216 56896 34216 0 net14
rlabel metal3 57232 35784 57232 35784 0 net15
rlabel metal2 52584 31696 52584 31696 0 net16
rlabel metal2 45528 26236 45528 26236 0 net17
rlabel metal2 38920 3528 38920 3528 0 net18
rlabel metal3 3192 9128 3192 9128 0 net19
rlabel metal2 27832 42140 27832 42140 0 net2
rlabel metal2 4536 8260 4536 8260 0 net20
rlabel metal2 3528 11088 3528 11088 0 net21
rlabel metal2 3976 13608 3976 13608 0 net22
rlabel metal2 7336 14224 7336 14224 0 net23
rlabel metal2 7896 15960 7896 15960 0 net24
rlabel metal2 13608 44968 13608 44968 0 net25
rlabel metal3 12936 45752 12936 45752 0 net26
rlabel metal2 11592 45808 11592 45808 0 net27
rlabel metal2 7112 43904 7112 43904 0 net28
rlabel metal2 35000 5208 35000 5208 0 net29
rlabel metal2 29176 43876 29176 43876 0 net3
rlabel metal3 5152 42504 5152 42504 0 net30
rlabel metal2 4424 42224 4424 42224 0 net31
rlabel metal2 7000 39256 7000 39256 0 net32
rlabel metal2 6216 34272 6216 34272 0 net33
rlabel metal3 47712 45080 47712 45080 0 net34
rlabel metal3 45864 43512 45864 43512 0 net35
rlabel metal3 44184 43652 44184 43652 0 net36
rlabel metal2 47432 45976 47432 45976 0 net37
rlabel metal2 40264 45136 40264 45136 0 net38
rlabel metal2 40656 41160 40656 41160 0 net39
rlabel metal2 30352 45192 30352 45192 0 net4
rlabel metal2 38920 6776 38920 6776 0 net40
rlabel metal2 48216 45640 48216 45640 0 net41
rlabel metal2 40040 43876 40040 43876 0 net42
rlabel metal3 39592 5152 39592 5152 0 net43
rlabel metal3 29400 5040 29400 5040 0 net44
rlabel metal2 26488 5936 26488 5936 0 net45
rlabel metal2 40712 4088 40712 4088 0 net46
rlabel metal2 33096 7672 33096 7672 0 net47
rlabel metal2 3976 10864 3976 10864 0 net48
rlabel metal3 3808 12264 3808 12264 0 net49
rlabel metal2 43624 30688 43624 30688 0 net5
rlabel metal2 31192 6776 31192 6776 0 net50
rlabel metal2 2072 17808 2072 17808 0 net51
rlabel metal3 5040 19096 5040 19096 0 net52
rlabel metal2 2856 11088 2856 11088 0 net53
rlabel metal2 2296 10528 2296 10528 0 net54
rlabel metal2 2072 7728 2072 7728 0 net55
rlabel metal2 14728 4648 14728 4648 0 net56
rlabel metal2 3752 39200 3752 39200 0 net57
rlabel metal2 4424 41944 4424 41944 0 net58
rlabel metal3 4984 41048 4984 41048 0 net59
rlabel metal3 57064 36232 57064 36232 0 net6
rlabel metal2 2072 36120 2072 36120 0 net60
rlabel metal2 25704 6104 25704 6104 0 net61
rlabel metal2 8344 43876 8344 43876 0 net62
rlabel metal2 9912 44352 9912 44352 0 net63
rlabel metal2 17472 44296 17472 44296 0 net64
rlabel metal2 19096 40600 19096 40600 0 net65
rlabel metal2 39816 44660 39816 44660 0 net66
rlabel metal2 38864 45640 38864 45640 0 net67
rlabel metal2 37576 44296 37576 44296 0 net68
rlabel metal3 30744 42616 30744 42616 0 net69
rlabel metal3 57848 31360 57848 31360 0 net7
rlabel metal2 46424 45472 46424 45472 0 net70
rlabel metal2 44632 46032 44632 46032 0 net71
rlabel metal2 26488 7336 26488 7336 0 net72
rlabel metal2 48776 43456 48776 43456 0 net73
rlabel metal2 52024 44632 52024 44632 0 net74
rlabel metal2 30632 9352 30632 9352 0 net75
rlabel metal2 32088 5264 32088 5264 0 net76
rlabel metal2 32984 4312 32984 4312 0 net77
rlabel metal2 41048 7728 41048 7728 0 net78
rlabel metal2 44408 3416 44408 3416 0 net79
rlabel metal2 57848 25816 57848 25816 0 net8
rlabel metal2 8120 15848 8120 15848 0 net80
rlabel metal3 2912 14280 2912 14280 0 net81
rlabel metal3 53816 30128 53816 30128 0 net82
rlabel metal2 41832 17920 41832 17920 0 net83
rlabel metal2 53592 19656 53592 19656 0 net84
rlabel metal2 43848 21280 43848 21280 0 net85
rlabel metal2 55608 25704 55608 25704 0 net86
rlabel metal2 55608 20720 55608 20720 0 net87
rlabel metal2 52696 22512 52696 22512 0 net88
rlabel metal2 33432 18928 33432 18928 0 net89
rlabel metal2 52696 28000 52696 28000 0 net9
rlabel metal2 31640 20440 31640 20440 0 net90
rlabel metal2 9576 25816 9576 25816 0 net91
rlabel metal2 8680 26040 8680 26040 0 net92
rlabel metal3 8624 26152 8624 26152 0 net93
rlabel metal2 45192 17192 45192 17192 0 net94
rlabel metal2 20328 25984 20328 25984 0 net95
rlabel metal2 29288 19768 29288 19768 0 net96
rlabel metal2 30408 44688 30408 44688 0 net97
rlabel metal3 27776 45864 27776 45864 0 net98
rlabel metal2 20552 24416 20552 24416 0 net99
rlabel metal2 57512 37800 57512 37800 0 pcpi_insn[0]
rlabel metal2 27608 46424 27608 46424 0 pcpi_insn[12]
rlabel metal2 28840 44408 28840 44408 0 pcpi_insn[13]
rlabel metal2 30072 45752 30072 45752 0 pcpi_insn[14]
rlabel metal2 58184 32424 58184 32424 0 pcpi_insn[1]
rlabel metal2 58240 36344 58240 36344 0 pcpi_insn[25]
rlabel metal2 58240 31528 58240 31528 0 pcpi_insn[26]
rlabel metal2 58184 26600 58184 26600 0 pcpi_insn[27]
rlabel metal2 58184 30632 58184 30632 0 pcpi_insn[28]
rlabel metal2 58184 27720 58184 27720 0 pcpi_insn[29]
rlabel metal2 58184 37184 58184 37184 0 pcpi_insn[2]
rlabel metal2 58184 33096 58184 33096 0 pcpi_insn[30]
rlabel metal2 58184 29568 58184 29568 0 pcpi_insn[31]
rlabel metal2 58184 33880 58184 33880 0 pcpi_insn[3]
rlabel metal2 58184 35336 58184 35336 0 pcpi_insn[4]
rlabel metal2 58184 34552 58184 34552 0 pcpi_insn[5]
rlabel metal2 58072 37520 58072 37520 0 pcpi_insn[6]
rlabel metal2 55384 14952 55384 14952 0 pcpi_rd[0]
rlabel metal2 55384 16408 55384 16408 0 pcpi_rd[10]
rlabel metal2 55384 21112 55384 21112 0 pcpi_rd[11]
rlabel metal3 58618 25592 58618 25592 0 pcpi_rd[12]
rlabel metal2 57960 21616 57960 21616 0 pcpi_rd[13]
rlabel metal2 55048 22008 55048 22008 0 pcpi_rd[14]
rlabel metal3 34272 4088 34272 4088 0 pcpi_rd[15]
rlabel metal2 28280 1414 28280 1414 0 pcpi_rd[16]
rlabel metal3 1358 25592 1358 25592 0 pcpi_rd[17]
rlabel metal3 1358 26936 1358 26936 0 pcpi_rd[18]
rlabel metal3 1358 26264 1358 26264 0 pcpi_rd[19]
rlabel metal2 55048 17304 55048 17304 0 pcpi_rd[1]
rlabel metal3 1358 24920 1358 24920 0 pcpi_rd[20]
rlabel metal2 27608 854 27608 854 0 pcpi_rd[21]
rlabel metal2 26936 48202 26936 48202 0 pcpi_rd[22]
rlabel metal2 26264 47698 26264 47698 0 pcpi_rd[23]
rlabel metal2 1960 24192 1960 24192 0 pcpi_rd[24]
rlabel metal3 1358 23576 1358 23576 0 pcpi_rd[25]
rlabel metal2 57960 28504 57960 28504 0 pcpi_rd[26]
rlabel metal2 34328 47138 34328 47138 0 pcpi_rd[27]
rlabel metal2 57288 29512 57288 29512 0 pcpi_rd[28]
rlabel metal2 57960 24528 57960 24528 0 pcpi_rd[29]
rlabel metal2 57960 16912 57960 16912 0 pcpi_rd[2]
rlabel metal3 55412 24472 55412 24472 0 pcpi_rd[30]
rlabel metal3 55412 19768 55412 19768 0 pcpi_rd[31]
rlabel metal3 58618 20216 58618 20216 0 pcpi_rd[3]
rlabel metal3 57330 18200 57330 18200 0 pcpi_rd[4]
rlabel metal3 35616 3640 35616 3640 0 pcpi_rd[5]
rlabel metal2 28952 854 28952 854 0 pcpi_rd[6]
rlabel metal2 57960 18368 57960 18368 0 pcpi_rd[7]
rlabel metal3 57330 22904 57330 22904 0 pcpi_rd[8]
rlabel metal3 58618 15512 58618 15512 0 pcpi_rd[9]
rlabel metal2 57960 23016 57960 23016 0 pcpi_ready
rlabel metal2 34384 3304 34384 3304 0 pcpi_rs1[0]
rlabel metal2 1848 8036 1848 8036 0 pcpi_rs1[10]
rlabel metal2 2408 8904 2408 8904 0 pcpi_rs1[11]
rlabel metal3 1582 12824 1582 12824 0 pcpi_rs1[12]
rlabel metal2 1736 13216 1736 13216 0 pcpi_rs1[13]
rlabel metal2 2408 14000 2408 14000 0 pcpi_rs1[14]
rlabel metal2 1736 16128 1736 16128 0 pcpi_rs1[15]
rlabel metal2 17640 45864 17640 45864 0 pcpi_rs1[16]
rlabel metal2 12376 46424 12376 46424 0 pcpi_rs1[17]
rlabel metal2 12040 45864 12040 45864 0 pcpi_rs1[18]
rlabel metal2 1736 43960 1736 43960 0 pcpi_rs1[19]
rlabel metal2 41384 8008 41384 8008 0 pcpi_rs1[1]
rlabel metal2 2408 42504 2408 42504 0 pcpi_rs1[20]
rlabel metal2 1848 42224 1848 42224 0 pcpi_rs1[21]
rlabel metal2 1736 38416 1736 38416 0 pcpi_rs1[22]
rlabel metal2 1736 33880 1736 33880 0 pcpi_rs1[23]
rlabel metal2 51464 46368 51464 46368 0 pcpi_rs1[24]
rlabel metal2 45528 46032 45528 46032 0 pcpi_rs1[25]
rlabel metal2 44184 45472 44184 45472 0 pcpi_rs1[26]
rlabel metal2 47768 45192 47768 45192 0 pcpi_rs1[27]
rlabel metal2 37128 45864 37128 45864 0 pcpi_rs1[28]
rlabel metal2 40488 46032 40488 46032 0 pcpi_rs1[29]
rlabel metal2 39256 7112 39256 7112 0 pcpi_rs1[2]
rlabel metal2 48440 45248 48440 45248 0 pcpi_rs1[30]
rlabel metal2 40488 46312 40488 46312 0 pcpi_rs1[31]
rlabel metal3 43960 3528 43960 3528 0 pcpi_rs1[3]
rlabel metal3 29344 3416 29344 3416 0 pcpi_rs1[4]
rlabel metal2 25928 3192 25928 3192 0 pcpi_rs1[5]
rlabel metal2 40936 3752 40936 3752 0 pcpi_rs1[6]
rlabel metal2 33320 3248 33320 3248 0 pcpi_rs1[7]
rlabel metal2 2408 11816 2408 11816 0 pcpi_rs1[8]
rlabel metal2 1736 12544 1736 12544 0 pcpi_rs1[9]
rlabel metal2 31248 3304 31248 3304 0 pcpi_rs2[0]
rlabel metal2 1736 17640 1736 17640 0 pcpi_rs2[10]
rlabel metal2 1736 18984 1736 18984 0 pcpi_rs2[11]
rlabel via2 1736 10808 1736 10808 0 pcpi_rs2[12]
rlabel metal2 1736 9968 1736 9968 0 pcpi_rs2[13]
rlabel metal3 1246 8120 1246 8120 0 pcpi_rs2[14]
rlabel metal2 14168 2086 14168 2086 0 pcpi_rs2[15]
rlabel metal2 1848 39256 1848 39256 0 pcpi_rs2[16]
rlabel metal2 1680 41944 1680 41944 0 pcpi_rs2[17]
rlabel metal2 2408 41496 2408 41496 0 pcpi_rs2[18]
rlabel metal2 1736 36008 1736 36008 0 pcpi_rs2[19]
rlabel metal2 25424 3080 25424 3080 0 pcpi_rs2[1]
rlabel metal3 8316 45752 8316 45752 0 pcpi_rs2[20]
rlabel metal2 8792 46144 8792 46144 0 pcpi_rs2[21]
rlabel metal2 16968 45864 16968 45864 0 pcpi_rs2[22]
rlabel metal2 18648 46368 18648 46368 0 pcpi_rs2[23]
rlabel metal2 40040 45808 40040 45808 0 pcpi_rs2[24]
rlabel metal2 38696 46144 38696 46144 0 pcpi_rs2[25]
rlabel metal2 38136 46424 38136 46424 0 pcpi_rs2[26]
rlabel metal2 31528 46256 31528 46256 0 pcpi_rs2[27]
rlabel metal3 50064 45752 50064 45752 0 pcpi_rs2[28]
rlabel metal2 45024 45864 45024 45864 0 pcpi_rs2[29]
rlabel metal2 27048 3304 27048 3304 0 pcpi_rs2[2]
rlabel metal3 49616 45864 49616 45864 0 pcpi_rs2[30]
rlabel metal2 52136 45528 52136 45528 0 pcpi_rs2[31]
rlabel metal2 29848 5152 29848 5152 0 pcpi_rs2[3]
rlabel metal2 31752 5880 31752 5880 0 pcpi_rs2[4]
rlabel metal2 32704 3304 32704 3304 0 pcpi_rs2[5]
rlabel metal2 43848 4648 43848 4648 0 pcpi_rs2[6]
rlabel metal3 45696 3416 45696 3416 0 pcpi_rs2[7]
rlabel metal3 4032 16072 4032 16072 0 pcpi_rs2[8]
rlabel metal2 1904 13720 1904 13720 0 pcpi_rs2[9]
rlabel metal3 58394 31640 58394 31640 0 pcpi_valid
rlabel metal2 57960 26712 57960 26712 0 pcpi_wr
<< properties >>
string FIXED_BBOX 0 0 60000 50000
<< end >>

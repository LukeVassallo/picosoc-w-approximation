* NGSPICE file created from pcpi_approx_mul.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_4 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_2 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VNW VPW VSS
.ends

.subckt pcpi_approx_mul clk pcpi_insn[0] pcpi_insn[10] pcpi_insn[11] pcpi_insn[12]
+ pcpi_insn[13] pcpi_insn[14] pcpi_insn[15] pcpi_insn[16] pcpi_insn[17] pcpi_insn[18]
+ pcpi_insn[19] pcpi_insn[1] pcpi_insn[20] pcpi_insn[21] pcpi_insn[22] pcpi_insn[23]
+ pcpi_insn[24] pcpi_insn[25] pcpi_insn[26] pcpi_insn[27] pcpi_insn[28] pcpi_insn[29]
+ pcpi_insn[2] pcpi_insn[30] pcpi_insn[31] pcpi_insn[3] pcpi_insn[4] pcpi_insn[5]
+ pcpi_insn[6] pcpi_insn[7] pcpi_insn[8] pcpi_insn[9] pcpi_rd[0] pcpi_rd[10] pcpi_rd[11]
+ pcpi_rd[12] pcpi_rd[13] pcpi_rd[14] pcpi_rd[15] pcpi_rd[16] pcpi_rd[17] pcpi_rd[18]
+ pcpi_rd[19] pcpi_rd[1] pcpi_rd[20] pcpi_rd[21] pcpi_rd[22] pcpi_rd[23] pcpi_rd[24]
+ pcpi_rd[25] pcpi_rd[26] pcpi_rd[27] pcpi_rd[28] pcpi_rd[29] pcpi_rd[2] pcpi_rd[30]
+ pcpi_rd[31] pcpi_rd[3] pcpi_rd[4] pcpi_rd[5] pcpi_rd[6] pcpi_rd[7] pcpi_rd[8] pcpi_rd[9]
+ pcpi_ready pcpi_rs1[0] pcpi_rs1[10] pcpi_rs1[11] pcpi_rs1[12] pcpi_rs1[13] pcpi_rs1[14]
+ pcpi_rs1[15] pcpi_rs1[16] pcpi_rs1[17] pcpi_rs1[18] pcpi_rs1[19] pcpi_rs1[1] pcpi_rs1[20]
+ pcpi_rs1[21] pcpi_rs1[22] pcpi_rs1[23] pcpi_rs1[24] pcpi_rs1[25] pcpi_rs1[26] pcpi_rs1[27]
+ pcpi_rs1[28] pcpi_rs1[29] pcpi_rs1[2] pcpi_rs1[30] pcpi_rs1[31] pcpi_rs1[3] pcpi_rs1[4]
+ pcpi_rs1[5] pcpi_rs1[6] pcpi_rs1[7] pcpi_rs1[8] pcpi_rs1[9] pcpi_rs2[0] pcpi_rs2[10]
+ pcpi_rs2[11] pcpi_rs2[12] pcpi_rs2[13] pcpi_rs2[14] pcpi_rs2[15] pcpi_rs2[16] pcpi_rs2[17]
+ pcpi_rs2[18] pcpi_rs2[19] pcpi_rs2[1] pcpi_rs2[20] pcpi_rs2[21] pcpi_rs2[22] pcpi_rs2[23]
+ pcpi_rs2[24] pcpi_rs2[25] pcpi_rs2[26] pcpi_rs2[27] pcpi_rs2[28] pcpi_rs2[29] pcpi_rs2[2]
+ pcpi_rs2[30] pcpi_rs2[31] pcpi_rs2[3] pcpi_rs2[4] pcpi_rs2[5] pcpi_rs2[6] pcpi_rs2[7]
+ pcpi_rs2[8] pcpi_rs2[9] pcpi_valid pcpi_wait pcpi_wr resetn vdd vss
X_2106_ _1257_ _1258_ _1259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2037_ _1031_ _1145_ _1149_ _1192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_2939_ _0617_ _0621_ _0634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_9_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input73_I pcpi_rs2[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2173__A2 _0960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2655_ net66 _0345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2724_ _0311_ _0413_ _0414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_22_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1606_ _0755_ _0769_ _0770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_6_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2586_ _0274_ _0275_ _0276_ _0277_ _1168_ _0278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_1537_ _0676_ _0673_ _0701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1675__A1 _0700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2440_ net92 _1297_ _0136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2371_ _0061_ _0064_ _0068_ _0069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__2146__A2 _1297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2638_ _0315_ _0324_ _0328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2707_ _0393_ _0395_ _0396_ _0397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_40_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2569_ _0235_ _0260_ _0262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2385__A2 _1297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input36_I pcpi_rs1[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1639__A1 _0777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1871_ _1022_ _1024_ _1026_ _1027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1940_ _1056_ _1096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_16_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2423_ _0102_ _0103_ _0119_ _0120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2285_ _1420_ _1433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2354_ _0035_ _0051_ _0052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_19_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1487__I net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2070_ _1222_ _1223_ _1224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2972_ _0007_ clknet_2_2__leaf_clk net112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_8_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1785_ _0909_ _0944_ _0945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1854_ _1009_ net56 _1010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1923_ _1042_ _1020_ _1079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2406_ _0053_ _0070_ _0103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_12_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2268_ _1388_ _1416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2337_ _1435_ _1450_ _0034_ _0035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2199_ _1328_ _1344_ _1347_ _1349_ _1217_ _1350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XTAP_TAPCELL_ROW_27_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2200__A1 _0979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1570_ _0733_ _0664_ _0734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_49_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2053_ _1157_ _1091_ _1208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2122_ _1127_ _1089_ _1275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2955_ _0416_ _0433_ _0651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_32_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2733__A2 _0371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2886_ _0532_ _1284_ _0533_ _0580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_25_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1837_ _0990_ _0994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1906_ _1060_ _1061_ _1062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_4_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1768_ _0662_ _0786_ _0929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1699_ _0861_ _0001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_35_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput97 net97 pcpi_rd[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput86 net86 pcpi_rd[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_2671_ _0357_ _0358_ _0360_ _0361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2740_ _0422_ _0428_ _0429_ _0430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_41_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1622_ _0688_ _0786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_14_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1484_ net11 _0523_ _0534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_22_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1553_ net72 _0717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_27_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2105_ _1220_ _1224_ _1258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2036_ _1190_ _1191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2938_ _0631_ _0632_ _0633_ _0029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_17_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input66_I pcpi_rs2[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2869_ _0498_ _0499_ _0561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2881__A1 _0291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2723_ _0310_ _0304_ _0308_ _0413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_42_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2654_ _0336_ _0339_ _0343_ _0344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2585_ _1456_ _1474_ _0277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_1_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1605_ _0767_ _0768_ _0754_ _0756_ _0769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_1536_ _0699_ _0700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_10_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2019_ _1043_ _1128_ _1174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_5_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2967__CLK clknet_2_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2370_ _0055_ _0067_ _0068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_24_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_19_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2706_ _0394_ _0360_ _0396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_40_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2637_ _0299_ net73 _0327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2499_ _0036_ _0109_ _0194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2568_ _0235_ _0260_ _0261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1519_ net46 net50 _0683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_12_Right_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2845__A1 net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_21_Right_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_2_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input29_I pcpi_rs1[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output97_I net97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_30_Right_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_45_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_24_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1870_ _1009_ _1025_ _1026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2422_ _0104_ _0111_ _0118_ _0119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2353_ _0037_ _0041_ _0050_ _0051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_10_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2284_ _1415_ _1432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_19_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1999_ _1117_ _1154_ _1155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2818__A1 _0371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2971_ _0006_ clknet_2_0__leaf_clk net111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1922_ _1076_ _1077_ _1057_ _1078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_21_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1784_ _0915_ _0922_ _0944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1853_ net48 _1009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_12_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2405_ _0100_ _1460_ _0101_ _0102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2336_ _1437_ _0032_ _0033_ _0034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_46_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2267_ net60 _1415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2198_ _1348_ _1349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_27_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2200__A2 _0981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1950__A1 _1023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2052_ _1185_ _1204_ _1206_ _1207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_16_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2121_ _1273_ _1266_ _1274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2954_ _0627_ _0641_ _0638_ _1299_ _0650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2885_ _0567_ _0569_ _0578_ _0243_ _0579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_32_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1905_ _1047_ _1048_ _1050_ _1061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_40_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_6_Right_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1767_ _0903_ _0924_ _0927_ _0928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_1836_ _0993_ _0006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1698_ _0859_ net94 _0860_ _0861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2319_ _1405_ _1440_ _1467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input11_I pcpi_insn[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput98 net98 pcpi_rd[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput87 net87 pcpi_rd[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_9_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2670_ net41 _0359_ _0360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1621_ _0739_ _0784_ _0785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1552_ _0697_ _0715_ _0716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input3_I pcpi_insn[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1483_ net5 net1 _0523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2104_ _1222_ _1223_ _1257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2035_ _1030_ _1145_ _1149_ _1190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_9_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2868_ _0540_ _0541_ _0557_ _0560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_32_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2937_ net104 _1352_ _0633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input59_I pcpi_rs2[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2799_ _0322_ _0488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_40_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1819_ _0966_ _0976_ _0978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2890__A2 _1320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2633__A2 _0322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2722_ _0410_ _0411_ _0412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2653_ _0340_ _0342_ _0343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2584_ _1456_ _1474_ _0240_ _0276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_22_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1604_ _0698_ _0736_ _0740_ net29 _0768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_1535_ _0698_ _0699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_10_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2018_ _1121_ _1136_ _1172_ _1173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XPHY_EDGE_ROW_19_Left_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_5_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2636_ _0313_ _0324_ _0325_ _0319_ _0311_ _0326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_4
X_2705_ _0359_ _0394_ _0395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_42_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2498_ _0152_ _0191_ _0192_ _0193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2567_ _0253_ _0254_ _0259_ _0260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_1518_ net72 _0669_ _0682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_4_Left_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_18_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2836__A2 _0375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_24_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2421_ _0112_ _0115_ _0117_ _0118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_2283_ _1421_ _1430_ _1431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2352_ _0044_ _0049_ _0050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_19_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2619_ net73 _0309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_30_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1998_ _1153_ _1154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA_input41_I pcpi_rs1[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2754__A1 net100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1852_ _0807_ _1008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1921_ _1058_ _1044_ _1077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2970_ _0005_ clknet_2_2__leaf_clk net110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1783_ _0941_ _0927_ _0942_ _0943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2404_ _0059_ _0069_ _0101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2266_ _1408_ _1412_ _1413_ _1414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2335_ _1442_ _1443_ _1449_ _0033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_20_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2197_ _1159_ _1348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_35_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1484__A1 net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_7_Left_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2120_ _1240_ _1241_ _1273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2051_ _1117_ _1154_ _1205_ _1206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_16_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2884_ _0572_ _0575_ _0576_ _0578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_32_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2953_ _0646_ _0647_ _0648_ _0030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1769__A2 _0700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1904_ _1055_ _1057_ _1059_ _1060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_17_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1835_ _0992_ net111 _0984_ _0993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1697_ _0812_ _0860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_12_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1766_ _0925_ _0897_ _0926_ _0927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2249_ net28 _1397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2318_ _1415_ _1383_ _1466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_33_Left_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_7_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput99 net99 pcpi_rd[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput88 net88 pcpi_rd[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__1620__B2 _0783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1482_ net16 net15 net17 _0512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_1_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1551_ _0677_ _0715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1620_ _0782_ _0752_ _0664_ _0783_ _0784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2103_ _1256_ _0010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2034_ _1102_ net56 _1189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2798_ _0359_ _0487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2867_ _0558_ _0559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2936_ _0532_ _1344_ _0533_ _0632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1818_ _0966_ _0976_ _0977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_17_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1749_ _0887_ _0881_ _0891_ _0910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_7_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output110_I net110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1841__A1 _0777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2652_ _0341_ net67 _0342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2721_ _0293_ _0320_ _0411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_6_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2583_ _0262_ _0273_ _1299_ _0275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2990__CLK clknet_2_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1534_ net40 _0698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1603_ _0736_ _0737_ net29 net18 _0767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_10_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2017_ _1123_ _1170_ _1171_ _1172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2919_ _0588_ _0559_ _0600_ _0613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_input71_I pcpi_rs2[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1823__A1 _0979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_36_Left_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2000__A1 _1008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_20_Left_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_19_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2635_ _0312_ _0318_ _0325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2704_ net42 _0394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2790__A2 _0478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2497_ _1436_ _0187_ _0189_ _0190_ _0192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_2566_ _0256_ _0258_ _0259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1517_ _0674_ _0675_ _0680_ _0681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_TAPCELL_ROW_2_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_2_2__f_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2420_ _0116_ _0106_ _0117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2282_ _1425_ _1429_ _1430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2351_ _0045_ _0047_ _0048_ _0049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_19_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1997_ _1137_ _1152_ _1153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2618_ _0306_ _0307_ _0308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2549_ _1164_ _0243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input34_I pcpi_rs1[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2754__A2 _0248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1851_ _1006_ _1007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_21_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1920_ _1074_ _1075_ _1076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2403_ _1375_ _0100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_24_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1782_ _0903_ _0924_ _0942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2265_ net59 _1397_ _1413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2334_ _1479_ _1480_ _1481_ _0032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2196_ _1346_ _1347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_47_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_35_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2736__A2 _0374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_51_Left_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2727__A2 _0374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2050_ _1137_ _1152_ _1205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2952_ net106 _1352_ _0648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2883_ _0572_ _0575_ _1348_ _0576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_32_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1903_ _1053_ _1058_ _1054_ _1044_ _1059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_1765_ _0875_ _0894_ _0926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1834_ _0935_ _0986_ _0987_ _0991_ _0809_ _0992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_40_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1696_ _0661_ _0817_ _0818_ _0857_ _0858_ _0859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_2248_ _1382_ net64 _1396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2317_ _1464_ _1420_ _1465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2179_ _1312_ _1317_ _1330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xoutput89 net89 pcpi_rd[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_54_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1550_ _0696_ _0709_ _0713_ _0714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2102_ net84 _1003_ _1255_ _1256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2033_ _1011_ _1040_ _1151_ _1186_ _1187_ _1188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_49_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2935_ _0626_ _0628_ _0630_ _1349_ _1168_ _0631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_2866_ _0540_ _0541_ _0557_ _0558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2797_ _0482_ _0484_ _0485_ _0486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_4_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1748_ _0671_ _0733_ _0909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1817_ _0967_ _0975_ _0976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_13_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1679_ _0840_ _0841_ _0766_ _0842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_43_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2651_ net39 _0341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2720_ _0369_ _0409_ _0382_ _0410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_2582_ _0262_ _0273_ _0274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1602_ _0699_ _0751_ _0766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1533_ _0668_ _0697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2016_ _1125_ _1118_ _1135_ _1171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_45_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2918_ _0590_ _0611_ _0612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_9_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input64_I pcpi_rs2[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2849_ _0509_ _0517_ _0539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2848__B2 _0519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1823__A2 _0981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2634_ _0306_ _0307_ _0314_ _0317_ _0324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_42_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2703_ _0358_ _0356_ _0391_ _0393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2565_ _0227_ _0255_ _0257_ _0250_ _0226_ _0258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_2_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1516_ _0676_ _0677_ _0679_ _0680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_10_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2496_ _1436_ _0187_ _0189_ _0190_ _0191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_2_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2980__CLK clknet_2_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2281_ _1426_ _1427_ _1428_ _1429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_2350_ _0046_ _1447_ _0048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_19_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1996_ _1138_ _1151_ _1152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2617_ net36 net35 _0295_ _0305_ _0307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_2548_ _0240_ _1472_ _0241_ _0242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_30_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input27_I pcpi_rs1[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2935__C _1168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2479_ _0172_ _0174_ _0083_ _0175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_38_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output95_I net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1850_ _1005_ _1006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_4_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1781_ _0903_ _0924_ _0941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2333_ _1445_ _1446_ _1448_ _1481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_2402_ _0088_ _0098_ _0099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_20_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2264_ _1409_ _1411_ _1412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2195_ _1345_ _1107_ _1346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_35_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1979_ _1129_ _1134_ _1135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_15_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2112__A1 _1045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2951_ _0532_ _1361_ _0533_ _0647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_8_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1902_ net81 _1058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_16_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2882_ _0573_ _0574_ _0575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_40_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1764_ _0875_ _0894_ _0925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1833_ _0979_ _0989_ _0990_ _0991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2316_ _1409_ _1464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_40_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1695_ _0808_ _0858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2247_ _1379_ _1380_ _1395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2654__A2 _0339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2178_ _1303_ _1319_ _1329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_31_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_46_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_19_Right_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_28_Right_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_37_Right_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_27_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2101_ _1217_ _0898_ _1254_ _1214_ _1255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2032_ _1139_ _1187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_43_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2865_ _0543_ _0548_ _0556_ _0557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2934_ _0422_ _0605_ _0630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_17_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_46_Right_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_40_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2796_ _0482_ _0484_ _0807_ _0485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_25_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1678_ _0755_ _0769_ _0773_ _0841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_1816_ _0969_ _0974_ _0975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1747_ _0906_ _0907_ _0908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_13_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_51_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2650_ net66 net41 _0340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2581_ _0270_ _0272_ _0273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1601_ _0750_ _0763_ _0764_ _0765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1532_ _0672_ _0681_ _0695_ _0696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA_input1_I pcpi_insn[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2015_ _1125_ _1118_ _1135_ _1170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2917_ _0593_ _0599_ _0611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2848_ _0479_ _0521_ _0501_ _0519_ _0480_ _0538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_5_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2779_ _0374_ _0465_ _0466_ _0467_ _0468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA_input57_I pcpi_rs2[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_5_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2775__A1 _0375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2702_ _0335_ _0391_ _0392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2633_ net74 _0322_ _0323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2495_ _0113_ _0149_ _0157_ _0190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_2564_ _0229_ _0223_ _0228_ _0257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_1515_ net46 _0678_ _0679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_3_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2280_ net31 net58 _1428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_35_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2616_ net34 net35 net71 _0305_ _0306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_51_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1995_ _1139_ _1141_ _1150_ _1151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2547_ _1470_ _1471_ _0241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2478_ _1292_ _0173_ _0174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_38_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2739__A1 _0291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_52_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1780_ _0782_ _0666_ _0792_ _0940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2332_ _1425_ _1429_ _1480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2401_ _0089_ _0095_ _0097_ _0098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_20_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2263_ _1410_ _1411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2194_ _1094_ _1105_ _1345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_47_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_35_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1978_ _1130_ _1132_ _1133_ _1134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2970__CLK clknet_2_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2881_ _0291_ _0385_ _0574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2950_ _0642_ _0643_ _0645_ _1364_ _0646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_32_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1832_ _0867_ _0904_ _0969_ _0974_ _0968_ _0990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_1901_ net51 _1056_ _1057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_52_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1763_ _0908_ _0923_ _0924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1694_ _0834_ _0853_ _0856_ _0857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_2246_ _1390_ _1392_ _1393_ _1394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2315_ _1457_ _1462_ _1463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__2993__CLK clknet_2_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2177_ _0807_ _1328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_43_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2586__C _1168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2100_ _1169_ _1249_ _1253_ _1211_ _1164_ _1254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_43_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2031_ _1141_ _1150_ _1186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2864_ _0549_ _0551_ _0554_ _0556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_2795_ _0407_ _0483_ _0484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2933_ _0238_ _0627_ _0628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1815_ _0952_ _0972_ _0973_ _0974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_17_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1677_ _0839_ _0840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1746_ _0877_ _0878_ _0893_ _0907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_13_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2229_ net63 _1377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_51_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_48_Left_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_54_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2580_ _0271_ _0272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1600_ _0757_ _0758_ _0753_ _0764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_1_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1531_ _0686_ _0694_ _0695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2014_ _0806_ _1169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2778_ _0315_ _0324_ _0331_ _0467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_45_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2847_ _0501_ _0519_ _0537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2916_ _0582_ _0610_ _0028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1729_ _0889_ _0890_ _0891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_0_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_5_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2472__A1 _1300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2701_ net41 _0391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2632_ _0294_ _0322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_42_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2494_ _0188_ _0189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2563_ _0140_ _0187_ _0255_ _0256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1514_ net61 _0678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_2_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_24_Left_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_10_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1994_ _1142_ _1146_ _1149_ _1150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_7_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2615_ net70 _0305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_42_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2546_ _0213_ _0240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2477_ _0128_ _0129_ _0171_ _0173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2381__B1 _0078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_29_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_52_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2400_ _0096_ _0085_ _0097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2262_ net30 _1410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_46_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2331_ _1439_ _1440_ _1441_ _1479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_2193_ _1329_ _1343_ _1344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_35_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1977_ _1131_ _1065_ _1133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2529_ _0154_ _0189_ _0198_ _0223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_30_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input32_I pcpi_rs1[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2896__A1 _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2880_ _0388_ _0488_ _0573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1900_ net20 _1056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1831_ _0988_ _0980_ _0989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_52_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1762_ _0909_ _0915_ _0922_ _0923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_12_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1693_ _0854_ _0804_ _0855_ _0856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2245_ net25 net64 _1393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2314_ _1391_ _1461_ _1462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2887__A1 net102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_27_Left_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2176_ _1214_ _1327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_11_Left_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_28_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_1_Right_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_54_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2030_ _1173_ _1184_ _1185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_2932_ _0603_ _0625_ _0627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_27_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1844__A2 _0997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2863_ _0552_ _0553_ _0554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2794_ _0406_ _0436_ _0483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_4_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_4_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1745_ _0786_ _0904_ _0905_ _0906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1814_ _0953_ _0970_ _0971_ _0973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1676_ _0754_ _0769_ _0773_ _0839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_0_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2228_ _1374_ _1375_ _1376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2159_ _1272_ _1309_ _1310_ _1311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_TAPCELL_ROW_51_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_8_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1530_ _0692_ _0693_ _0694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_38_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2013_ _1163_ _1168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_54_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2915_ active _0583_ _0609_ _0610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2777_ _0315_ _0324_ _0331_ _0466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2846_ _0531_ _0535_ _0536_ _0026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1728_ net46 _0743_ _0890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_5_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1659_ _0714_ _0731_ _0821_ _0822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA_output101_I net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2631_ _0293_ _0320_ _0321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2700_ _0386_ _0388_ _0389_ _0390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_40_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2562_ _0140_ _1458_ _0230_ _0255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_6_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_2_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_10_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2493_ _0113_ _0149_ _0157_ _0188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1513_ net45 _0677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_4_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2215__A2 _0991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input62_I pcpi_rs2[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2829_ _0506_ _0509_ _0517_ _0518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_33_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1993_ _1147_ _1148_ _1149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2614_ _0298_ _0301_ _0303_ _0304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_2545_ _0236_ _0237_ _0238_ _0239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_15_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2476_ _0128_ _0129_ _0171_ _0172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_41_Left_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_38_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2261_ net58 _1409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2330_ _1452_ _1476_ _1477_ _1478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2192_ _1333_ _1342_ _1343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_43_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1976_ _1058_ _1131_ _1132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_53_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2528_ _0036_ _1375_ _0222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input25_I pcpi_rs1[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2459_ _0154_ _0155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_26_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1761_ _0916_ _0918_ _0921_ _0922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_1830_ _0823_ _0904_ _0975_ _0988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2313_ _1374_ _1458_ _1459_ _1460_ _1461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_20_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1692_ _0732_ _0776_ _0855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2244_ _1391_ _1381_ _1392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2175_ _1298_ _1326_ _0012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1959_ _1109_ _1113_ _1114_ _1115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__2878__A2 _0375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_27_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1541__A2 _0688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2931_ _0603_ _0625_ _0626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_0_clk clk clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_2862_ _0394_ _0419_ _0553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2793_ _0479_ _0481_ _0482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1744_ _0884_ _0892_ _0905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1813_ _0970_ _0971_ _0953_ _0972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_13_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1675_ _0700_ net79 _0838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_15_Right_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2227_ net65 _1375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_24_Right_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2089_ _1237_ _1239_ _1242_ _1243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_2158_ _1273_ _1267_ _1277_ _1310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_TAPCELL_ROW_51_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_33_Right_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_42_Right_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_42_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_51_Right_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2012_ _1004_ _1167_ _0008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2914_ _0602_ _0604_ _0607_ _1323_ _0609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2845_ net101 _0280_ _0536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2776_ _0309_ _0465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1727_ _0677_ _0745_ _0889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1658_ _0716_ _0819_ _0820_ _0821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_13_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1589_ _0751_ _0752_ _0753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2630_ _0311_ _0319_ _0320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2492_ _0109_ _0187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2561_ _0043_ _0100_ _0254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1512_ net50 _0676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_49_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2828_ _0510_ _0513_ _0516_ _0517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_45_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2759_ _0391_ _0448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2973__CLK clknet_2_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input55_I pcpi_rs2[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1992_ net21 _1029_ _1148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2613_ _0294_ _0302_ _0300_ _0299_ _0303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2544_ _1299_ _0238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2475_ _0169_ _0170_ _0171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2996__CLK clknet_2_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_21_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2060__A1 _1168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2260_ _1405_ _1407_ _1408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2191_ _1334_ _1336_ _1341_ _1342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_47_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1975_ net24 _1131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2458_ _1423_ net32 _1385_ _1387_ _0154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_2527_ _0220_ _0201_ _0221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2389_ _0040_ _0032_ _0050_ _0086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_TAPCELL_ROW_26_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input18_I pcpi_rs1[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1760_ _0919_ _0920_ _0921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_12_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1691_ _0732_ _0776_ _0854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2312_ _1383_ _1460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2243_ _1379_ _1391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2174_ active _1324_ _1325_ _1326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_31_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1958_ _1111_ _1112_ _1114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1889_ _1044_ _1045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_16_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_45_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2861_ _0391_ _0302_ _0552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2930_ _0623_ _0624_ _0625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2792_ _0480_ _0481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_25_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1674_ _0735_ _0760_ _0775_ _0835_ _0836_ _0837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
X_1812_ _0955_ _0949_ _0954_ _0971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_1743_ _0733_ _0904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2226_ net25 _1374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_21_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2157_ _1273_ _1267_ _1277_ _1309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_2088_ _1240_ _1241_ _1242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_17_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_51_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2011_ active _1162_ _1166_ _1167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_45_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2913_ _1292_ _0605_ _0606_ _0607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2844_ _0532_ _1249_ _0533_ _0535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_5_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2775_ _0375_ _0292_ _0464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1726_ _0887_ _0881_ _0888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_0_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1588_ _0741_ _0752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1657_ _0720_ _0711_ _0730_ _0820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_13_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2209_ _1221_ _1260_ _1336_ _1341_ _1335_ _1359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_48_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_2_0__f_clk clknet_0_clk clknet_2_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_24_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2491_ _1436_ _1375_ _0186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2560_ _0222_ _0251_ _0252_ _0253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1511_ net47 net50 _0675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2827_ _0514_ _0515_ _0516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2758_ _0384_ _0445_ _0446_ _0447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_5_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2689_ _0368_ _0375_ _0378_ _0379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_1_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input48_I pcpi_rs1[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1709_ _0866_ _0869_ _0870_ _0871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_1_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2612_ _0296_ _0302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_42_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1991_ net20 _1028_ _1147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2543_ _0221_ _0232_ _0237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2474_ _0077_ _0038_ _0170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_21_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2190_ _1312_ _1339_ _1340_ _1341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_1974_ _1075_ _1064_ _1127_ _1130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_43_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2457_ _1440_ _0109_ _0153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2526_ _0186_ _0219_ _0220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2388_ _0040_ _0032_ _0050_ _0085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_38_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_26_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_34_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2986__CLK clknet_2_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1690_ _0837_ _0852_ _0853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_12_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2242_ _1379_ _1381_ _1389_ _1390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_2311_ _1387_ _1459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2173_ _1165_ _0960_ _1325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1957_ _1111_ _1112_ _1113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_22_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2509_ _0182_ _0203_ _0204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_31_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1888_ net21 _1044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input30_I pcpi_rs1[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_54_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2860_ _0550_ _0545_ _0551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2791_ _0460_ _0478_ _0480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_4_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1811_ _0955_ _0949_ _0954_ _0970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_7_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1673_ _0762_ _0836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1742_ _0901_ _0902_ _0903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2225_ _1373_ _0015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_5_Right_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_8_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2087_ _1127_ _1018_ _1241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2156_ _1122_ _1230_ _1308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2989_ _0024_ clknet_2_1__leaf_clk net99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input78_I pcpi_rs2[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2484__A2 _0161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2172__A1 _1300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2010_ _1165_ _0805_ _1166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2912_ _0428_ _0429_ _0606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_53_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2774_ _0323_ _0461_ _0462_ _0333_ _0321_ _0463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
X_2843_ _0587_ _0533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1725_ _0848_ _0849_ _0887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_5_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1587_ net78 _0751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1656_ _0720_ _0711_ _0730_ _0819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_13_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2139_ _1159_ _1292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2466__A2 _0122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2208_ _1356_ _1357_ _1358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_4_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2490_ _0146_ _0120_ _0160_ _0185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1510_ net72 _0673_ _0674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_14_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2688_ _0376_ _0377_ _0349_ _0378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_2826_ net41 _0300_ _0515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2757_ _0444_ _0399_ _0403_ _0446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_5_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1708_ _0830_ _0832_ _0829_ _0870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_41_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1639_ _0777_ _0778_ _0803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_18_Left_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_49_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_54_Left_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_36_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2375__A1 _0052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1990_ _1031_ _1145_ _1146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_7_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2611_ _0299_ _0294_ _0296_ _0300_ _0301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_2542_ _0180_ _0218_ _0234_ _0236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2473_ _0076_ _1417_ _0169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1801__B1 _0960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input60_I pcpi_rs2[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2809_ _0452_ _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_14_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_29_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_3_Left_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_37_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1973_ _1128_ _1100_ _1129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2525_ _0193_ _0199_ _0219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_11_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2456_ _0111_ _0118_ _0151_ _0152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2387_ _0083_ _0084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_11_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_34_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2241_ _1383_ _1385_ _1387_ _1388_ _1389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2310_ _1385_ _1458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2172_ _1300_ _1320_ _1322_ _1323_ _1324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_48_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1956_ _1080_ _1081_ _1112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1887_ _1042_ _1043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_7_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2508_ _0201_ _0202_ _0203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2439_ _0082_ _0135_ _0017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input23_I pcpi_rs1[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_6_Left_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2790_ _0460_ _0478_ _0479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_1810_ _0867_ _0885_ _0968_ _0969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1741_ _0871_ _0874_ _0902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_21_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1672_ _0765_ _0774_ _0835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_23_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2224_ _1372_ net89 _1214_ _1373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_0_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2155_ _1305_ _1306_ _1307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2086_ _1054_ _1017_ _1240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2988_ _0023_ clknet_2_1__leaf_clk net98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1939_ _1058_ _1095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_16_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2976__CLK clknet_2_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1508__A2 _0671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_50_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_32_Left_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_11_Right_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_13_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_20_Right_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_54_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2172__A2 _1320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2911_ _0428_ _0429_ _0605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2773_ _0326_ _0332_ _0462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2842_ _1006_ _0532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1724_ _0671_ _0885_ _0886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1586_ _0747_ _0748_ _0749_ _0750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_0_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1655_ _0816_ _0663_ _0815_ _0666_ _0818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_2138_ _1290_ _1291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_2069_ _1181_ _1183_ _1178_ _1223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_14_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2207_ _1331_ _1332_ _1342_ _1357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_44_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_4_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1901__A2 _1056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2825_ _0346_ _0296_ _0514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2687_ _0347_ _0337_ _0377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2756_ _0399_ _0403_ _0444_ _0445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_30_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1707_ _0868_ _0869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1638_ _0796_ _0800_ _0801_ _0802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1569_ net79 _0733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_51_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_19_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_35_Left_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_15_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2610_ _0297_ _0300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2541_ _0180_ _0218_ _0233_ _0234_ _0235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_2472_ _1300_ _0167_ _0168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_2_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1877__A1 _1023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2808_ _0447_ _0459_ _0495_ _0496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_18_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2739_ _0291_ _0419_ _0429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input53_I pcpi_rs2[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1868__A1 _1023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_37_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1940__I _1056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2587__A2 _1362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1972_ _1127_ _1128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_51_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_49_Right_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2455_ _0112_ _0149_ _0150_ _0151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2524_ _0182_ _0203_ _0218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_11_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2386_ _1005_ _0083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_38_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2240_ net27 _1388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2171_ _1006_ _1323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_48_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1886_ net52 _1042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1955_ _1026_ _1110_ _1111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_44_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2507_ _0184_ _0185_ _0200_ _0202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_2438_ _0084_ _1210_ _0127_ _0133_ _0134_ _0135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_11_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2369_ _0065_ _0066_ _1398_ _1399_ _0067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA_input16_I pcpi_insn[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1490__I _0587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1740_ _0868_ _0870_ _0901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1671_ _0822_ _0833_ _0834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_13_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input8_I pcpi_insn[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2478__A1 _1292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2223_ _1364_ _0997_ _1369_ _1371_ _1372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2085_ _1238_ _1232_ _1239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2154_ _1262_ _1263_ _1279_ _1306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_48_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2987_ _0022_ clknet_2_1__leaf_clk net97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1938_ _1088_ _1090_ _1094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1869_ net55 _1025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput80 pcpi_rs2[8] net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_42_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_7_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2841_ _1328_ _0524_ _0530_ _0243_ _0531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2910_ _1008_ _0603_ _0604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2772_ _0326_ _0332_ _0461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_5_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1723_ _0751_ _0885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1654_ _0663_ _0815_ _0666_ _0816_ _0817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_28_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2206_ _1334_ _1355_ _1356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1585_ net78 _0664_ _0749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2137_ _1285_ _1289_ _1290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2068_ _1043_ _1221_ _1222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_10_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2853__A1 _0339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2824_ _0511_ _0507_ _0513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_5_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2966__CLK clknet_2_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2686_ net66 _0341_ _0376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2755_ _0387_ _0444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_26_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1706_ _0710_ _0867_ _0868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1637_ _0797_ _0799_ _0801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1499_ _0662_ _0663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1568_ _0714_ _0731_ _0732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_49_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2540_ _0182_ _0203_ _0234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2471_ _0144_ _0161_ _0166_ _0167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_2_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2738_ _0423_ _0424_ _0427_ _0428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_2807_ _0493_ _0494_ _0449_ _0495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_33_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2172__C _1323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2669_ _0347_ _0359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input46_I pcpi_rs1[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1971_ net23 _1127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_51_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2454_ _0116_ _0106_ _0115_ _0150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_2523_ _0177_ _0217_ _0019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2385_ net91 _1297_ _0082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput1 pcpi_insn[0] net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_36_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_0_clk_I clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2170_ _1160_ _1321_ _1322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1954_ _1022_ _1024_ _1110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_51_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1885_ _1011_ _1040_ _1041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2368_ _1388_ _1382_ _1384_ _1386_ _0066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_2506_ _0184_ _0185_ _0200_ _0201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2437_ _0587_ _0134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2299_ net32 _1409_ _1447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_53_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1670_ _0824_ _0830_ _0832_ _0833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2222_ _1160_ _1370_ _1212_ _1371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_21_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2084_ _1199_ _1200_ _1238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2153_ _1265_ _1304_ _1305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_33_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2986_ _0021_ clknet_2_0__leaf_clk net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1937_ _1023_ _1087_ _1092_ _1093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
Xinput70 pcpi_rs2[28] net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1868_ _1023_ _1019_ _1024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput81 pcpi_rs2[9] net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1799_ _0947_ _0958_ _0959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2469__A2 _0122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_42_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_50_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_7_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2840_ _0525_ _0528_ _0529_ _0530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2771_ _0447_ _0459_ _0460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1722_ _0844_ _0851_ _0883_ _0884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1584_ _0739_ _0742_ _0748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_9_Right_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1653_ _0690_ _0816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_13_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2205_ _1336_ _1341_ _1355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_48_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2136_ _1286_ _1287_ _1288_ _1289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_8_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2067_ _1176_ _1221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_2969_ _0004_ clknet_2_2__leaf_clk net109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input76_I pcpi_rs2[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2823_ _0473_ _0474_ _0511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2754_ net100 _0248_ _0443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1705_ _0827_ _0867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2685_ _0374_ _0375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1567_ _0716_ _0721_ _0730_ _0731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_1636_ _0797_ _0799_ _0800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1498_ net50 _0662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2119_ _1122_ _1236_ _1272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_15_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2470_ _0162_ _0164_ _0165_ _0166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XPHY_EDGE_ROW_50_Left_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2668_ _0341_ _0358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2737_ _0425_ _0426_ _0427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_41_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2806_ _0456_ _0457_ _0455_ _0494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_14_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input39_I pcpi_rs1[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2599_ net99 _0248_ _0289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1619_ _0745_ _0783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_49_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1556__A2 _0715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1774__I _0660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1970_ _1125_ _1068_ _1126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2522_ _0084_ _1291_ _0206_ _0216_ _0134_ _0217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_2453_ _0116_ _0105_ _0115_ _0149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2384_ _1327_ _0079_ _0080_ _0081_ _0016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
Xinput2 pcpi_insn[12] net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_36_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1483__A1 net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2979__CLK clknet_2_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_31_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1953_ _1093_ _1108_ _1109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_7_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1884_ _1027_ _1039_ _1040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2505_ _0186_ _0193_ _0199_ _0200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__2717__A1 _0334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2367_ net25 _1382_ _1377_ _1378_ _0065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_2298_ _1404_ net33 _1446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_2436_ _0130_ _0132_ _1323_ _0133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_19_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_53_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2221_ _1086_ _1115_ _1370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2152_ _1271_ _1278_ _1304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_17_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2083_ _1045_ _1236_ _1237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_16_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2985_ _0020_ clknet_2_1__leaf_clk net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1936_ _1088_ _1089_ _1090_ _1091_ _1092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1867_ _1015_ _1023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput71 pcpi_rs2[29] net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput60 pcpi_rs2[19] net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput82 pcpi_valid net82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_31_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1798_ _0948_ _0952_ _0957_ _0958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_12_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2419_ _0062_ _0063_ _0116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA_input21_I pcpi_rs1[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2770_ _0449_ _0455_ _0458_ _0459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__1840__A1 _0979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1721_ _0845_ _0881_ _0882_ _0883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA_clkbuf_2_1__f_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1583_ _0739_ _0742_ _0746_ _0747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_0_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1652_ _0752_ _0815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_21_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2204_ _1303_ _1319_ _1343_ _1354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_2135_ _1095_ _1102_ _1288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2066_ _1174_ _1218_ _1219_ _1184_ _1173_ _1220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_8_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input69_I pcpi_rs2[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2899_ _0549_ _0591_ _0592_ _0556_ _0548_ _0593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
X_2968_ _0003_ clknet_2_2__leaf_clk net108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1919_ _1049_ _1075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_40_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2684_ _0299_ _0374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2822_ _0338_ _0309_ _0510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2753_ _0289_ _0442_ _0024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1704_ _0710_ _0866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_39_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1635_ _0798_ _0749_ _0799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1566_ _0723_ _0729_ _0730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1497_ _0660_ _0661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_49_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2049_ _1188_ _1203_ _1204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_2118_ _1235_ _1269_ _1270_ _1271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_44_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2914__C _1323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2599__A2 _0248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_15_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2805_ _0456_ _0457_ _0455_ _0493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_54_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2667_ _0345_ _0357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2736_ _0335_ _0374_ _0426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1618_ _0743_ _0782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_14_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2598_ _0286_ _0287_ _0288_ _0023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_5_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1549_ _0710_ _0671_ _0711_ _0712_ _0713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_49_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2202__A1 net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_39_Left_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1492__A2 net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_23_Left_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2521_ _1323_ _0215_ _0216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2452_ _1433_ net65 _0148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2383_ net90 _0813_ _0081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_18_Right_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xinput3 pcpi_insn[13] net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1483__A2 net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_27_Right_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_52_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2719_ _0363_ _0367_ _0409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XPHY_EDGE_ROW_36_Right_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input51_I pcpi_rs2[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_45_Right_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_54_Right_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_52_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1952_ _1094_ _1105_ _1107_ _1108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_7_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1883_ _1037_ _1038_ _1039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_51_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2504_ _0194_ _0195_ _0198_ _0199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_2435_ _1292_ _0131_ _0132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2366_ _0062_ _0063_ _0064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_47_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2297_ _1423_ _1438_ _1445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_45_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2151_ _1281_ _1301_ _1282_ _1302_ _1303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_2220_ _1354_ _1360_ _1368_ _1008_ _1369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2082_ _1025_ _1236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2984_ _0019_ clknet_2_1__leaf_clk net93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2969__CLK clknet_2_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_26_Left_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1935_ _1035_ _1091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput50 pcpi_rs2[0] net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput61 pcpi_rs2[1] net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput72 pcpi_rs2[2] net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1797_ _0953_ _0954_ _0956_ _0957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_1866_ _1015_ _1019_ _1021_ _1022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_2418_ _0113_ _0114_ _0115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XPHY_EDGE_ROW_10_Left_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input14_I pcpi_insn[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2349_ _1464_ _0046_ _0047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_EDGE_ROW_0_Right_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_38_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1651_ _0814_ _0000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1720_ _0846_ _0840_ _0850_ _0882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_1582_ _0698_ _0743_ _0741_ _0745_ _0746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_0_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2856__A1 _0339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input6_I pcpi_insn[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2203_ _1327_ _1350_ _1351_ _1353_ _0013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2065_ _1182_ _1170_ _1180_ _1219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2134_ _1091_ _1101_ _1287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2967_ _0002_ clknet_2_2__leaf_clk net105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_44_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2898_ _0551_ _0554_ _0592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1849_ _0608_ _0618_ _1005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_4_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1918_ _1053_ _1074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_54_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2821_ _0470_ _0507_ _0508_ _0476_ _0469_ _0509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XTAP_TAPCELL_ROW_18_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2683_ _0351_ _0353_ _0373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2799__I _0322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2752_ _0084_ _1155_ _0441_ _0134_ _0442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_26_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1634_ _0747_ _0748_ _0798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1703_ _0862_ _0863_ _0864_ _0865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_1496_ _0629_ _0649_ _0660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1565_ _0725_ _0727_ _0728_ _0729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_1_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2048_ _1189_ _1195_ _1202_ _1203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2117_ _1237_ _1267_ _1268_ _1270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_36_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input81_I pcpi_rs2[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_23_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2804_ _0443_ _0492_ _0025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2735_ _0357_ _0338_ _0425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2666_ _0345_ net42 _0356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_2597_ net98 _0280_ _0288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1617_ _0703_ _0780_ _0781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1548_ _0681_ _0686_ _0694_ _0712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_37_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2451_ _0146_ _0120_ _0147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2520_ _0209_ _0212_ _0214_ _0215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_23_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput4 pcpi_insn[14] net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_39_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2382_ _1157_ _1158_ _1007_ _0080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_46_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_34_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_2_1__f_clk clknet_0_clk clknet_2_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_19_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2718_ _0406_ _0407_ _0408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_34_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_34_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2649_ _0338_ _0339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_40_Left_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input44_I pcpi_rs1[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_48_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_31_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1951_ _1087_ _1106_ _1107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_22_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1882_ _1036_ _1033_ _1034_ _1038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_51_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2365_ net30 net62 _0063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_47_Left_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2503_ _0196_ _0197_ _0198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2434_ _0128_ _0129_ _0078_ _0131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2296_ _1442_ _1443_ _1444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2150_ _1259_ _1280_ _1302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2081_ _1195_ _1202_ _1234_ _1235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_48_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2983_ _0018_ clknet_2_1__leaf_clk net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1934_ _1018_ _1090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput73 pcpi_rs2[30] net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput62 pcpi_rs2[20] net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_31_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput40 pcpi_rs1[2] net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1796_ _0955_ _0949_ _0956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1865_ _1012_ _1017_ _1018_ _1020_ _1021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xinput51 pcpi_rs2[10] net51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2417_ _1410_ _1384_ _1386_ _1406_ _0114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2348_ net33 _0046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_35_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2279_ net57 net32 _1427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1834__B1 _0991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1650_ _0810_ net83 _0813_ _0814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1581_ _0744_ _0745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_5_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2202_ net87 _1352_ _1353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_21_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2064_ _1181_ _1183_ _1218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2133_ _1074_ _1096_ _1286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2897_ _0550_ _0545_ _0554_ _0591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1917_ _1062_ _1071_ _1072_ _1073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_8_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2966_ _0001_ clknet_2_2__leaf_clk net94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1848_ net113 _1003_ _1004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1779_ _0939_ _0003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2847__A2 _0519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2820_ _0472_ _0475_ _0508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_38_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2751_ _1300_ _0437_ _0440_ _0083_ _0441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_30_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2682_ net69 _0371_ _0372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1564_ _0726_ _0679_ _0728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1633_ _0705_ _0706_ _0704_ _0797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_1702_ _0816_ _0815_ _0864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1495_ net4 _0639_ net3 _0649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_49_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2047_ _1196_ _1198_ _1201_ _1202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XTAP_TAPCELL_ROW_1_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2116_ _1267_ _1268_ _1237_ _1269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA_input74_I pcpi_rs2[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2949_ _0240_ _0433_ _0644_ _0645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_32_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_23_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2734_ _0368_ _0322_ _0424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2803_ _0245_ _1207_ _0486_ _0491_ _0246_ _0492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_26_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2665_ _0346_ net68 _0355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2596_ _0245_ _1370_ _0246_ _0287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1547_ _0686_ _0694_ _0681_ _0711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1616_ _0668_ _0699_ _0780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1486__A1 net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2910__A1 _1008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2450_ _0104_ _0145_ _0146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2381_ _1328_ _0075_ _0078_ _1349_ _1217_ _0079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_23_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput5 pcpi_insn[1] net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_34_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2717_ _0334_ _0405_ _0407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1943__A2 _1045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input37_I pcpi_rs1[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2648_ _0337_ _0338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2579_ _0140_ _0100_ _0256_ _0258_ _0255_ _0271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_10_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1950_ _1023_ _1092_ _1106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2502_ _0046_ _1459_ _0197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_31_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1881_ _1033_ _1034_ _1036_ _1037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2364_ net28 net63 _0062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_51_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2433_ _0077_ _0128_ _0129_ _0076_ _0130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_11_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2295_ _1425_ _1429_ _1443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_34_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2992__CLK clknet_2_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2080_ _1196_ _1232_ _1233_ _1234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_17_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2982_ _0017_ clknet_2_1__leaf_clk net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1933_ _1017_ _1089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput74 pcpi_rs2[31] net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput41 pcpi_rs1[30] net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput63 pcpi_rs2[21] net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput30 pcpi_rs1[20] net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput52 pcpi_rs2[11] net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1864_ _1016_ _1020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1795_ _0827_ _0782_ _0919_ _0955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_12_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2416_ _1406_ _1410_ _1384_ _1386_ _0113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_2278_ net59 net30 _1426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2347_ _1407_ _1446_ _0042_ _0045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_50_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1580_ net77 _0744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_13_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2201_ _1296_ _1352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_28_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2132_ _1088_ _1043_ _1285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2063_ _1163_ _1217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2896_ _0386_ _0542_ _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1847_ _0812_ _1003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2965_ _0000_ clknet_2_2__leaf_clk net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1916_ _1060_ _1061_ _1072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_8_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1778_ _0938_ net108 _0860_ _0939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_4_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2681_ _0316_ _0371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2750_ _0438_ _0439_ _1211_ _0440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_38_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1701_ _0718_ _0665_ _0863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1494_ net2 _0639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1563_ _0726_ _0690_ _0727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1632_ _0781_ _0785_ _0795_ _0796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_1_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2115_ _1238_ _1232_ _1242_ _1268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_2046_ _1199_ _1200_ _1201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA_input67_I pcpi_rs2[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2948_ _0431_ _0432_ _0644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2879_ _0570_ _0571_ _0572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_44_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2664_ _0351_ _0353_ _0354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2733_ _0359_ _0371_ _0423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2802_ _0240_ _0489_ _0490_ _0083_ _0491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2595_ _0282_ _0275_ _0285_ _0243_ _0286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_5_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1546_ _0697_ _0710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1615_ _0777_ _0778_ _0779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_49_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_37_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2435__A1 _1292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2029_ _1174_ _1181_ _1183_ _1184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_9_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2380_ _0076_ _0077_ _0078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xinput6 pcpi_insn[25] net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_36_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2647_ net38 _0337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_42_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2716_ _0334_ _0405_ _0406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2578_ _0253_ _0268_ _0269_ _0270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1529_ _0682_ _0683_ _0684_ _0693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_10_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_14_Right_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_output98_I net98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_23_Right_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_32_Right_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_31_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1880_ _1035_ _1025_ _1036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2501_ _0042_ _1458_ _0196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2363_ _1388_ _0060_ _0061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2294_ _1439_ _1440_ _1441_ _1442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_EDGE_ROW_41_Right_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2432_ _1460_ _0129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_50_Right_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_42_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_30_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput31 pcpi_rs1[21] net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2981_ _0016_ clknet_2_0__leaf_clk net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput20 pcpi_rs1[11] net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1863_ _1012_ _1016_ _1017_ _1018_ _1019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_1932_ _1009_ _1088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput64 pcpi_rs2[22] net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput42 pcpi_rs1[31] net42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2415_ _1420_ _0060_ _0112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput75 pcpi_rs2[3] net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1794_ _0827_ _0783_ _0954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput53 pcpi_rs2[12] net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2277_ _1422_ _1413_ _1424_ _1425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2346_ _1438_ _0043_ _0044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2062_ _1216_ _0009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2200_ _0979_ _0981_ _1007_ _1351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2131_ _1259_ _1280_ _1283_ _1284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_29_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2964_ _1003_ _0656_ _0658_ _0659_ _0031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XPHY_EDGE_ROW_14_Left_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_44_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2895_ _0588_ _0558_ _0589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1846_ _1002_ _0007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1915_ net52 _1056_ _1071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1777_ _0858_ _0928_ _0937_ _0938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_40_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_4_Right_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2329_ _1403_ _1451_ _1477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input12_I pcpi_insn[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2471__A2 _0161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_18_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2680_ _0363_ _0367_ _0369_ _0370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_30_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2223__A2 _0997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1700_ _0663_ _0700_ _0862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1631_ _0793_ _0794_ _0795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_39_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1493_ _0608_ _0618_ _0629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1562_ net47 _0726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input4_I pcpi_insn[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2045_ _1049_ _1014_ _1200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2114_ _1266_ _1267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2947_ _0627_ _0641_ _0238_ _0643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_17_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2878_ _0487_ _0375_ _0571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1829_ _0796_ _0800_ _0987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_40_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2437__I _0587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2801_ _0439_ _0487_ _0488_ _0438_ _0490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_39_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2663_ _0352_ _0340_ _0342_ _0353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_2732_ _0378_ _0417_ _0421_ _0422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_41_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2594_ _1476_ _0283_ _0284_ _0285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1614_ _0696_ _0709_ _0778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_5_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1545_ _0704_ _0707_ _0708_ _0709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_37_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2028_ _1182_ _1170_ _1183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_49_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_17_Left_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_32_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2426__A2 _0122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1937__A1 _1023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput7 pcpi_insn[26] net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_52_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2646_ _0335_ _0336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2715_ _0384_ _0387_ _0404_ _0405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2577_ _0254_ _0259_ _0269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1528_ _0687_ _0689_ _0691_ _0692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_37_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_33_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_2_Left_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2500_ _0154_ _0188_ _0195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2431_ _1464_ _0128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_3_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2362_ net64 _0060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_47_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2293_ _1427_ _1428_ _1441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_2_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_44_Left_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2629_ _0312_ _0313_ _0318_ _0319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA_input42_I pcpi_rs1[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2877__A2 _0371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1704__I _0710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1540__A2 _0700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2980_ _0015_ clknet_2_0__leaf_clk net89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput32 pcpi_rs1[22] net32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput10 pcpi_insn[29] net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1931_ _1078_ _1079_ _1087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
Xinput43 pcpi_rs1[3] net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput54 pcpi_rs2[13] net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1793_ _0823_ _0885_ _0953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xinput21 pcpi_rs1[12] net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1862_ _1014_ _1018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput65 pcpi_rs2[23] net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2414_ _0059_ _0108_ _0110_ _0111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
Xinput76 pcpi_rs2[4] net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2276_ _1404_ _1423_ _1409_ _1411_ _1424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_2345_ _0042_ _0043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_50_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_5_Left_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2710__A1 _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2061_ net114 _1003_ _1215_ _1216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2130_ _1281_ _1282_ _1283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_44_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2963_ net107 _0813_ _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1914_ _1068_ _1069_ _1070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_52_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2894_ _0543_ _0586_ _0588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1845_ _1001_ net112 _0984_ _1002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_12_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1776_ _0931_ _0934_ _0936_ _0937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2328_ _1456_ _1474_ _1475_ _1476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_33_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_4_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2259_ _1406_ _1407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_7_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_31_Left_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_26_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1630_ _0781_ _0785_ _0794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_39_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1492_ net4 net2 _0618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1561_ _0724_ _0677_ _0722_ _0725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_1_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2044_ net21 _1013_ _1199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2113_ _1238_ _1232_ _1242_ _1266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2877_ _0357_ _0371_ _0570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2946_ _0627_ _0641_ _0642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_44_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1759_ _0726_ _0743_ _0920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1828_ _0796_ _0800_ _0986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_50_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2913__A1 _1292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2972__CLK clknet_2_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1622__I _0688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2731_ _0298_ _0420_ _0421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_41_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2800_ _0438_ _0439_ _0487_ _0488_ _0489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_26_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2662_ net68 net38 _0352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2593_ _1476_ _0283_ _1211_ _0284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1613_ _0734_ _0760_ _0777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1544_ _0705_ _0706_ _0708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_5_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_37_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2027_ _1129_ _1134_ _1182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_9_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2929_ _0612_ _0613_ _0622_ _0624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_32_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input72_I pcpi_rs2[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2995__CLK clknet_2_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput8 pcpi_insn[27] net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_36_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2714_ _0399_ _0403_ _0404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_34_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2645_ net68 _0335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2576_ _0254_ _0259_ _0268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1527_ _0690_ _0676_ _0673_ _0670_ _0691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_9_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2592__A2 _1451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2041__A1 _1056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2361_ _1394_ _1401_ _0058_ _0059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2430_ _0123_ _0125_ _0126_ _0127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2292_ _1411_ _1440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_47_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2628_ _0315_ _0317_ _0318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input35_I pcpi_rs1[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2559_ _0220_ _0201_ _0232_ _0252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_33_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1930_ _1085_ _1086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
Xinput66 pcpi_rs2[24] net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput11 pcpi_insn[2] net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput33 pcpi_rs1[23] net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput55 pcpi_rs2[14] net55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput77 pcpi_rs2[5] net77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput44 pcpi_rs1[4] net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1792_ _0915_ _0922_ _0951_ _0952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
Xinput22 pcpi_rs1[13] net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1861_ _1013_ _1017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2413_ _1416_ _0109_ _0106_ _0107_ _0110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_2344_ net32 _0042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_20_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2275_ net31 _1423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_50_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_53_Left_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2060_ _1168_ _0857_ _1213_ _1214_ _1215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2893_ _0548_ _0556_ _0586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_29_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2962_ _1364_ _0657_ _0658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1913_ _1067_ _1052_ _1062_ _1069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_1844_ _0858_ _0997_ _1000_ _1001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_12_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1775_ _0931_ _0934_ _0935_ _0936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2258_ net31 _1406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2327_ _1454_ _1455_ _1475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_4_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2189_ _1313_ _1337_ _1338_ _1340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_7_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1560_ _0662_ _0724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1491_ net3 _0608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2112_ _1045_ _1230_ _1265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2043_ _1197_ _1190_ _1198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_17_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2945_ _0638_ _0640_ _0641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2876_ _1300_ _0568_ _0569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_32_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1827_ _0985_ _0005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1689_ _0838_ _0844_ _0851_ _0852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_1758_ _0722_ _0783_ _0919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output104_I net104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2661_ _0348_ _0349_ _0350_ _0351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2730_ _0290_ _0302_ _0419_ _0322_ _0420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_39_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2592_ _1403_ _1451_ _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_22_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1612_ _0761_ _0775_ _0776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1543_ _0705_ _0706_ _0707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_37_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2026_ _1180_ _1181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_9_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input65_I pcpi_rs2[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2859_ _0514_ _0515_ _0550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2928_ _0612_ _0613_ _0622_ _0623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_32_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2831__A1 _0334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput9 pcpi_insn[28] net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_52_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2644_ _0321_ _0333_ _0334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_42_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2713_ _0400_ _0401_ _0402_ _0403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_27_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2575_ _1327_ _0265_ _0266_ _0267_ _0021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_22_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1526_ _0678_ _0690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_10_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2009_ _1164_ _1165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_9_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2360_ _0056_ _0057_ _1396_ _0058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_51_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2291_ _1438_ _1439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_11_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_47_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_10_Right_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_30_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2627_ net36 _0295_ _0297_ _0316_ _0317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_30_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput110 net110 pcpi_rd[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_15_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input28_I pcpi_rs1[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2489_ _1433_ _0100_ _0183_ _0184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2558_ _0226_ _0250_ _0251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1509_ net45 _0673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_2_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_53_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1860_ net19 _1016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput34 pcpi_rs1[24] net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput67 pcpi_rs2[25] net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput12 pcpi_insn[30] net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput56 pcpi_rs2[15] net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput45 pcpi_rs1[5] net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput78 pcpi_rs2[6] net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1791_ _0916_ _0949_ _0950_ _0951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_12_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput23 pcpi_rs1[14] net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2412_ _0060_ _0109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2274_ _1404_ _1406_ net58 _1410_ _1422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_42_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2343_ _0040_ _0032_ _0041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_50_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1989_ _1143_ _1144_ _1030_ _1032_ _1145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_15_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1755__A1 _0715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2180__A1 _1122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2483__A2 _0161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2892_ _0537_ _0538_ _0563_ _0584_ _0585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1912_ _1052_ _1062_ _1067_ _1068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2961_ _1354_ _1360_ _1368_ _0657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1843_ _0802_ _0998_ _0999_ _1000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_17_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1774_ _0660_ _0935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2326_ _1463_ _1472_ _1473_ _1474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2257_ _1404_ _1405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_47_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2188_ _1337_ _1338_ _1313_ _1339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_19_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_14_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1490_ _0587_ active vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2042_ _1147_ _1148_ _1197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2111_ _1262_ _1263_ _1264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XPHY_EDGE_ROW_8_Right_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_17_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2944_ _0635_ _0623_ _0637_ _0640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_2875_ _0537_ _0538_ _0565_ _0568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_4_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1826_ _0983_ net110 _0984_ _0985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_17_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_39_Right_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2383__A1 net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1757_ _0917_ _0910_ _0918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1688_ _0845_ _0847_ _0850_ _0851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_2309_ _1414_ _1418_ _1457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA_input10_I pcpi_insn[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_48_Right_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2374__A1 _0052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2660_ _0345_ _0346_ _0347_ _0337_ _0350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_41_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1611_ _0762_ _0765_ _0774_ _0775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2591_ _0270_ _0272_ _0282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1542_ _0692_ _0693_ _0706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA_input2_I pcpi_insn[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2025_ _1178_ _1179_ _1180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2927_ _0614_ _0617_ _0621_ _0622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_2789_ _0463_ _0477_ _0478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2858_ _0358_ _0465_ _0549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1809_ _0867_ _0783_ _0956_ _0968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA_input58_I pcpi_rs2[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_54_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2643_ _0323_ _0326_ _0332_ _0333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_42_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2712_ _0392_ _0397_ _0402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2574_ net96 _0813_ _0267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2889__A2 _0248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1525_ net72 _0688_ _0689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2008_ _1163_ _1164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_33_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1552__A2 _0715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2290_ net59 _1438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_2_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_30_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2626_ net37 _0316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_42_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2557_ _0227_ _0228_ _0230_ _0250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
Xoutput100 net100 pcpi_rd[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput111 net111 pcpi_rd[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_2488_ _0152_ _0159_ _0183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_37_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1508_ _0668_ _0671_ _0672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_53_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1525__A2 _0688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput13 pcpi_insn[31] net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_33_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1790_ _0917_ _0911_ _0921_ _0950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
Xinput35 pcpi_rs1[25] net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput68 pcpi_rs2[26] net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2411_ _1416_ _0060_ _0106_ _0107_ _0108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xinput57 pcpi_rs2[16] net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_20_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput46 pcpi_rs1[6] net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput79 pcpi_rs2[7] net79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput24 pcpi_rs1[15] net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2273_ net60 _1420_ _1421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2342_ _0036_ _0038_ _0039_ _0040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_47_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1988_ net49 _1016_ _1013_ _1014_ _1144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_2609_ net36 _0299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_2_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input40_I pcpi_rs1[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_2_2__f_clk clknet_0_clk clknet_2_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_41_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2843__I _0587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2975__CLK clknet_2_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2960_ _1168_ _0650_ _0655_ _0656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_29_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1682__A1 _0688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2891_ _0562_ _0559_ _0560_ _0584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1773_ _0932_ _0933_ _0934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1842_ _0802_ _0998_ _0935_ _0999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1911_ _1063_ _1064_ _1066_ _1067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_12_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2325_ _1391_ _1457_ _1461_ _1473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2256_ net57 _1404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2187_ _1315_ _1309_ _1314_ _1338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_47_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_9_Left_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_38_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1967__A2 _1122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2041_ _1056_ _1025_ _1196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2110_ _1227_ _1228_ _1244_ _1263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2943_ _0635_ _0623_ _0637_ _0638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_29_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2874_ _0537_ _0538_ _0565_ _0567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1825_ _0812_ _0984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_4_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1756_ _0889_ _0890_ _0917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2308_ _1454_ _1455_ _1456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_31_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1687_ _0848_ _0849_ _0850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_0_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2239_ _1386_ _1387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_45_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2590_ _0278_ _0279_ _0281_ _0022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1610_ _0766_ _0770_ _0773_ _0774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_1541_ _0668_ _0688_ _0705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2024_ _1101_ _1130_ _1132_ _1179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_45_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2857_ _0509_ _0517_ _0547_ _0548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2926_ _0593_ _0599_ _0620_ _0621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_9_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2788_ _0464_ _0469_ _0476_ _0477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_20_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1739_ _0900_ _0002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1808_ _0823_ _0904_ _0967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_36_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2711_ _0365_ _0366_ _0364_ _0401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2642_ _0327_ _0328_ _0331_ _0332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_2573_ _1007_ _1347_ _0266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1524_ net43 _0688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_10_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2007_ _0629_ _1163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_26_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input70_I pcpi_rs2[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2909_ _0585_ _0601_ _0603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_33_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2329__A2 _1451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_38_Left_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_24_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_22_Left_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2625_ _0314_ _0315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_42_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2487_ _0141_ _0142_ _0181_ _0182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
Xoutput101 net101 pcpi_rd[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_2556_ _0244_ _0247_ _0249_ _0020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_23_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1507_ _0670_ _0671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xoutput112 net112 pcpi_rd[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__1845__I1 net112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput36 pcpi_rs1[26] net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput25 pcpi_rs1[16] net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput14 pcpi_insn[3] net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput69 pcpi_rs2[27] net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2410_ _0055_ _0067_ _0064_ _0107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
Xinput58 pcpi_rs2[17] net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2341_ _1446_ _1448_ _0039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xinput47 pcpi_rs1[7] net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2272_ _1397_ _1420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_23_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1987_ net49 net48 _1028_ _1029_ _1143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_15_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2608_ _0290_ _0294_ _0296_ _0297_ _0298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_2539_ _0221_ _0232_ _0233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA_input33_I pcpi_rs1[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_6_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2890_ _1165_ _1320_ _0583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1910_ _1053_ _1054_ _1065_ _1066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_4_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1772_ _0710_ _0665_ _0933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1841_ _0777_ _0778_ _0998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2324_ _1470_ _1471_ _1472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2255_ _1376_ _1402_ _1403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XPHY_EDGE_ROW_25_Left_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2186_ _1315_ _1309_ _1314_ _1337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_18_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2040_ _1141_ _1193_ _1194_ _1195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_44_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2942_ _0497_ _0542_ _0616_ _0636_ _0637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_2873_ _0563_ _0564_ _0565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_29_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1686_ net45 _0740_ _0849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1755_ _0715_ _0885_ _0916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1824_ _0935_ _0795_ _0963_ _0982_ _0809_ _0983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_2238_ net62 _1386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2307_ _1419_ _1431_ _1455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_48_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2169_ _1094_ _1105_ _1321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_24_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2965__CLK clknet_2_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1540_ _0697_ _0700_ _0703_ _0704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_10_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2023_ _1175_ _1177_ _1178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2856_ _0339_ _0465_ _0545_ _0546_ _0547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_2925_ _0448_ _0594_ _0615_ _0619_ _0620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_1807_ _0948_ _0964_ _0965_ _0966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_15_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2787_ _0470_ _0472_ _0475_ _0476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_40_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1669_ _0831_ _0819_ _0832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1738_ _0899_ net105 _0860_ _0900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_28_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output102_I net102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2710_ _0386_ _0388_ _0389_ _0400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_27_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2641_ _0329_ _0330_ _0331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2572_ _0261_ _0263_ _0264_ _1160_ _1212_ _0265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_22_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1523_ _0676_ _0673_ _0670_ _0678_ _0687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_10_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_33_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2006_ _1007_ _1156_ _1161_ _1162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_18_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input63_I pcpi_rs2[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2839_ _0525_ _0528_ _1348_ _0529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_33_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2908_ _0585_ _0601_ _0602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_5_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2624_ net37 net36 net71 _0305_ _0314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_42_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput102 net102 pcpi_rd[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_2486_ _0139_ _0143_ _0181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2555_ net95 _0248_ _0249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput113 net113 pcpi_rd[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_1506_ _0669_ _0670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_18_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput37 pcpi_rs1[27] net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput26 pcpi_rs1[17] net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput59 pcpi_rs2[18] net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput15 pcpi_insn[4] net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput48 pcpi_rs1[8] net48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2271_ _1414_ _1418_ _1419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2340_ _1438_ _0038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_32_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1986_ _1020_ net55 _1142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_7_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2607_ net70 _0297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_15_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input26_I pcpi_rs1[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2538_ _0222_ _0226_ _0231_ _0232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2469_ _0099_ _0122_ _0165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_46_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2156__A1 _1122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1840_ _0979_ _0995_ _0996_ _0997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_12_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1771_ _0718_ _0815_ _0932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2254_ _1394_ _1401_ _1402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2323_ _1374_ _1459_ _1471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2185_ _1221_ _1236_ _1335_ _1336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_43_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1969_ _1100_ _1075_ _1124_ _1125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__2689__A2 _0375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2941_ _0497_ _0594_ _0616_ _0621_ _0636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2872_ _0562_ _0559_ _0560_ _0564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_25_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1823_ _0979_ _0981_ _0982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_20_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1685_ _0669_ _0745_ _0848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1754_ _0884_ _0913_ _0914_ _0915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2306_ _1393_ _1453_ _1454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2237_ _1384_ _1385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_29_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2099_ _1250_ _1251_ _1252_ _1253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_2168_ _1303_ _1319_ _1320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_0_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_17_Right_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_26_Right_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_39_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2834__A2 _0519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_35_Right_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_44_Right_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_53_Right_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2589__A1 net97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2022_ _1100_ _1176_ _1177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2786_ _0473_ _0474_ _0475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_2855_ _0511_ _0507_ _0516_ _0546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_2924_ _0597_ _0591_ _0596_ _0619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_31_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1806_ _0945_ _0946_ _0958_ _0965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_17_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1599_ _0753_ _0757_ _0758_ _0763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1668_ _0723_ _0729_ _0831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1737_ _0661_ _0865_ _0898_ _0809_ _0899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__2685__I _0374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2640_ net38 _0305_ _0330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1794__A2 _0783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2571_ _1463_ _1472_ _0264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_22_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1522_ _0682_ _0685_ _0686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2005_ _1157_ _1158_ _1160_ _1161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2907_ _0589_ _0600_ _0601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_33_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1482__A1 net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2838_ _0526_ _0527_ _0528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_41_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2769_ _0456_ _0457_ _0458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_5_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input56_I pcpi_rs2[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1494__I net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2978__CLK clknet_2_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1700__A2 _0700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2623_ net35 net73 _0313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__2716__A1 _0334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput103 net103 pcpi_rd[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_30_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2554_ _1296_ _0248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_12_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput114 net114 pcpi_rd[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_2485_ _0178_ _0166_ _0179_ _0180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_2_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1505_ net44 _0669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_10_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_2_0__f_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1758__A2 _0783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_44_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput38 pcpi_rs1[28] net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput27 pcpi_rs1[18] net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_52_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput16 pcpi_insn[5] net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput49 pcpi_rs1[9] net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2270_ _1415_ _1417_ _1418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_9_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2937__A1 net104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1985_ _1027_ _1140_ _1037_ _1141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_15_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2606_ _0295_ _0296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2537_ _0227_ _0228_ _0230_ _0231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_47_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2399_ _0044_ _0049_ _0096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2468_ _1478_ _0073_ _0163_ _0164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_3_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_41_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input19_I pcpi_rs1[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output87_I net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1770_ _0929_ _0930_ _0931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_8_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2253_ _1395_ _1396_ _1400_ _1401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2322_ _1465_ _1466_ _1469_ _1470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_2184_ _1221_ _1089_ _1316_ _1335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_34_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2083__A1 _1045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1899_ _1053_ _1054_ _1044_ net81 _1055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1968_ _1064_ _1066_ _1124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_43_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_3_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2940_ _0614_ _0634_ _0635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2871_ _0559_ _0560_ _0562_ _0563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_20_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1753_ _0886_ _0911_ _0912_ _0914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_13_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1822_ _0943_ _0959_ _0980_ _0978_ _0981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_17_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1684_ _0846_ _0839_ _0847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2305_ _1390_ _1392_ _1453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2236_ net63 _1384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_0_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2167_ _1307_ _1318_ _1319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_48_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2098_ _1158_ _1101_ _1252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_39_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_14_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1497__I _0660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2021_ _1131_ _1176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_49_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2923_ _0497_ _0594_ _0616_ _0617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_53_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2785_ _0341_ _0297_ _0474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2854_ _0511_ _0507_ _0516_ _0545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1805_ _0952_ _0957_ _0964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1736_ _0875_ _0894_ _0897_ _0898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__2513__A2 _1417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1598_ net79 _0752_ _0762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1667_ _0825_ _0826_ _0829_ _0830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_28_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2219_ _1358_ _1367_ _1368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_51_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_46_Left_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_36_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2570_ _0238_ _0262_ _0263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1521_ _0683_ _0684_ _0685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2004_ _1159_ _1160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_45_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2906_ _0590_ _0593_ _0599_ _0600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_TAPCELL_ROW_33_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1482__A2 net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2734__A2 _0322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2699_ _0356_ _0361_ _0389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2768_ _0400_ _0401_ _0402_ _0457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2837_ _0439_ _0388_ _0527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1719_ _0846_ _0840_ _0850_ _0881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_13_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input49_I pcpi_rs1[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_47_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2622_ _0306_ _0307_ _0312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2553_ _0245_ _1321_ _0246_ _0247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput104 net104 pcpi_rd[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput115 net115 pcpi_ready vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_23_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1504_ net75 _0668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2484_ _0144_ _0161_ _0179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_52_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput39 pcpi_rs1[29] net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput28 pcpi_rs1[19] net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput17 pcpi_insn[6] net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_32_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1984_ _1036_ _1033_ _1034_ _1140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_15_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2605_ net71 _0295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2536_ _0229_ _0223_ _0230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2467_ _0052_ _0071_ _0163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2398_ _0090_ _0091_ _0094_ _0095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_41_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2968__CLK clknet_2_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2321_ _1467_ _1468_ _1469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2252_ _1398_ _1399_ _1400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2183_ _1128_ _1260_ _1334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1967_ _1042_ _1122_ _1123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1898_ net22 _1054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input31_I pcpi_rs1[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2519_ _0209_ _0212_ _0213_ _0214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_54_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2870_ _0496_ _0500_ _0561_ _0562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_44_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_29_Left_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_25_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1752_ _0911_ _0912_ _0886_ _0913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1683_ _0771_ _0772_ _0846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1821_ _0977_ _0980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2304_ _1403_ _1451_ _1452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_13_Left_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2235_ _1382_ _1383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_45_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2097_ _1091_ _1095_ _1251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_0_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2166_ _1308_ _1312_ _1317_ _1318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2999_ net115 net116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_3_Right_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input79_I pcpi_rs2[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_39_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2020_ _1130_ _1132_ _1175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2853_ _0339_ _0542_ _0543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2922_ _0615_ _0616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_17_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2784_ net38 _0295_ _0473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1549__A1 _0710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1666_ _0826_ _0828_ _0829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1735_ _0895_ _0856_ _0896_ _0897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1804_ _0793_ _0794_ _0963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1597_ _0735_ _0760_ _0761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_36_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2149_ _1259_ _1280_ _1301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2218_ _1359_ _1367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_8_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1788__A1 _0715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2440__A2 _1297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1520_ net61 net45 _0684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2003_ _0649_ _1159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1482__A3 net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2836_ _0438_ _0375_ _0526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2905_ _0595_ _0596_ _0598_ _0599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_9_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2698_ _0335_ _0388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_41_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2767_ _0392_ _0397_ _0456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1649_ _0812_ _0813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1718_ _0786_ net79 _0880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_16_Left_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_output100_I net100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2621_ _0304_ _0308_ _0310_ _0311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_50_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2483_ _0144_ _0161_ _0178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput116 net116 pcpi_wr vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_2552_ _0587_ _0246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_10_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1503_ _0663_ _0666_ _0667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput105 net105 pcpi_rd[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_37_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2819_ _0471_ _0466_ _0475_ _0507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_33_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input61_I pcpi_rs2[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_1_Left_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_52_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput18 pcpi_rs1[0] net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_32_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput29 pcpi_rs1[1] net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_9_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2604_ net35 _0294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_7_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1983_ _1035_ net56 _1139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2535_ _0092_ _1459_ _0196_ _0229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2466_ _0099_ _0122_ _0162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_43_Left_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2397_ _0091_ _0093_ _0094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_41_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2251_ net27 _1377_ _1378_ _1397_ _1399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_2320_ _1439_ _1416_ _1468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2182_ _1331_ _1332_ _1333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_18_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1966_ _1075_ _1122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_43_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1897_ net80 _1053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2449_ _0111_ _0118_ _0145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2518_ net4 _0639_ _0608_ _0213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA_input24_I pcpi_rs1[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1820_ _0943_ _0959_ _0977_ _0978_ _0979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_2
XTAP_TAPCELL_ROW_17_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1751_ _0887_ _0881_ _0891_ _0912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_1682_ _0688_ _0751_ _0845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2234_ net26 _1382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2303_ _1435_ _1450_ _1451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_0_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2096_ _1157_ _1102_ _1250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_0_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2165_ _1313_ _1314_ _1316_ _1317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_48_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2213__B1 _1362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1949_ _1097_ _1104_ _1105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_31_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_30_Left_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_22_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_13_Right_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_53_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2783_ _0471_ _0466_ _0472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2852_ _0292_ _0542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2921_ _0597_ _0591_ _0596_ _0615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_31_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_22_Right_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1803_ _0962_ _0004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_9_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1596_ _0750_ _0753_ _0759_ _0760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_1665_ _0717_ _0827_ _0828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1549__A2 _0671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1734_ _0834_ _0853_ _0896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_31_Right_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2217_ _1327_ _1363_ _1365_ _1366_ _0014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_48_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_36_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2148_ _1299_ _1300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__1485__A1 net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2079_ _1197_ _1191_ _1201_ _1233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_48_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_40_Right_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_8_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2002_ _1088_ _1158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_18_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2904_ _0597_ _0591_ _0598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2766_ _0450_ _0451_ _0454_ _0455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2835_ _0487_ _0488_ _0525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2697_ _0385_ _0386_ _0387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1648_ _0811_ _0812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_6_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1579_ _0740_ _0743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1717_ _0877_ _0878_ _0879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_47_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2620_ _0290_ _0309_ _0310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_27_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2482_ net93 _1297_ _0177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput106 net106 pcpi_rd[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_2551_ _1006_ _0245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_2_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1502_ _0665_ _0666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_18_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2818_ _0371_ _0292_ _0506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2749_ _0291_ _0439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1915__A2 _1056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input54_I pcpi_rs2[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput19 pcpi_rs1[10] net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2991__CLK clknet_2_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1982_ _1011_ _1040_ _1138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2603_ _0291_ _0292_ _0293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2534_ _0092_ _1458_ _0228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2465_ _0147_ _0160_ _0161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2396_ _1439_ _0092_ _0093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_38_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1833__A1 _0979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2250_ _1397_ net27 net63 net62 _1398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__2304__A2 _1451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2181_ _1305_ _1306_ _1318_ _1332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_47_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1965_ _1119_ _1083_ _1120_ _1121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_7_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2791__A2 _0478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2517_ _0210_ _0211_ _0212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_11_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1896_ _1047_ _1051_ _1052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2379_ _1374_ _0077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2448_ _0139_ _0143_ _0144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_54_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input17_I pcpi_insn[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1750_ _0910_ _0911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_17_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_52_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1681_ _0765_ _0842_ _0843_ _0844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2233_ _1380_ _1381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2302_ _1437_ _1444_ _1449_ _1450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA_input9_I pcpi_insn[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2164_ _1315_ _1309_ _1316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_48_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2095_ _1225_ _1245_ _1248_ _1249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_TAPCELL_ROW_0_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2997_ active clknet_2_3__leaf_clk net115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1879_ _1012_ _1035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1948_ _1098_ _1099_ _1103_ _1104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_3_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_22_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2920_ _0448_ _0542_ _0614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_2_3__f_clk clknet_0_clk clknet_2_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_2782_ _0329_ _0330_ _0471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_45_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2851_ _0503_ _0504_ _0518_ _0541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_40_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1802_ _0961_ net109 _0860_ _0962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1733_ _0834_ _0853_ _0895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1595_ _0757_ _0758_ _0759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1664_ _0726_ _0827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2147_ _0618_ _1299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2216_ net88 _1352_ _1366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_2_3__f_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2078_ _1197_ _1191_ _1201_ _1232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_27_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2001_ _1074_ _1157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2903_ _0452_ _0419_ _0552_ _0597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_9_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2696_ _0358_ _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2765_ _0451_ _0453_ _0454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2834_ _0501_ _0519_ _0522_ _0524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_26_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1716_ _0837_ _0852_ _0878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1647_ _0544_ _0555_ _0577_ _0811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_6_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1578_ _0698_ _0736_ _0740_ _0741_ _0742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_13_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2407__A1 _1417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2550_ _0235_ _0239_ _0242_ _0243_ _0244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_30_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput107 net107 pcpi_rd[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_2_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2481_ _0136_ _0176_ _0018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1501_ _0664_ _0665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_46_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2817_ _0503_ _0504_ _0505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2679_ _0368_ _0339_ _0369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2748_ _0357_ _0438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_41_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_14_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2876__A1 _1300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input47_I pcpi_rs1[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_52_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1981_ _1121_ _1136_ _1137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_23_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2602_ net74 _0292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2533_ _0043_ _0187_ _0227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2464_ _0148_ _0152_ _0159_ _0160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2395_ _0046_ _0092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_46_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2180_ _1122_ _1260_ _1330_ _1331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_34_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1964_ _1046_ _1118_ _1069_ _1120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_7_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1895_ _1048_ _1050_ _1051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2516_ _0077_ _1432_ _0211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2447_ _0141_ _0142_ _0143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_3_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_54_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2378_ _1405_ _0076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2981__CLK clknet_2_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2301_ _1445_ _1446_ _1448_ _1449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_20_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1680_ _0766_ _0840_ _0841_ _0843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2232_ net27 net26 _1377_ _1378_ _1380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_45_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_0_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2163_ _1176_ _1090_ _1275_ _1315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_48_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2094_ _1246_ _1206_ _1247_ _1248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_31_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2996_ _0031_ clknet_2_3__leaf_clk net107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1947_ _1101_ _1102_ _1103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1878_ _1015_ _1019_ _1031_ _1032_ _1034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_2
XFILLER_0_16_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1724__A1 _0671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2140__A1 _1008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2140__B2 _1292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2850_ _0506_ _0539_ _0540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_15_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2781_ _0316_ _0309_ _0470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1663_ _0725_ _0727_ _0826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1732_ _0879_ _0893_ _0894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_13_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1801_ _0661_ _0793_ _0940_ _0960_ _0858_ _0961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_1594_ _0738_ _0742_ _0755_ _0756_ _0758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_0_0_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_7_Right_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1706__A1 _0710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2682__A2 _0371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2146_ net86 _1297_ _1298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2215_ _1364_ _0991_ _1365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2077_ _1096_ _1230_ _1231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2979_ _0014_ clknet_2_0__leaf_clk net88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_8_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input77_I pcpi_rs2[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_27_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2000_ _1008_ _1155_ _1156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2902_ _0452_ _0302_ _0596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2833_ _0479_ _0521_ _0480_ _0522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_53_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2764_ _0336_ _0452_ _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2695_ _0368_ _0385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_41_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1715_ _0838_ _0876_ _0877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1646_ _0661_ _0667_ _0805_ _0809_ _0810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1577_ net29 _0741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2129_ _1246_ _1206_ _1225_ _1245_ _1247_ _1282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_44_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_30_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2480_ _0084_ _1253_ _0168_ _0175_ _0134_ _0176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_23_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput108 net108 pcpi_rd[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_1500_ net18 _0664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_12_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput90 net90 pcpi_rd[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_37_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2816_ _0463_ _0477_ _0504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_33_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_52_Left_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2678_ net69 _0368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2747_ _0408_ _0436_ _0437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_1_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1629_ _0782_ _0665_ _0792_ _0793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_TAPCELL_ROW_52_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1980_ _1123_ _1126_ _1135_ _1136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_23_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2601_ _0290_ _0291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2463_ _0153_ _0157_ _0158_ _0159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2532_ _0193_ _0199_ _0225_ _0226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__2555__A1 net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2394_ _0045_ _0047_ _0091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1963_ _1118_ _1069_ _1046_ _1119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_3_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1894_ net81 _1049_ _1050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2515_ _0038_ _1460_ _0210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2446_ _0095_ _0097_ _0094_ _0142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_54_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2700__A1 _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2377_ _1478_ _0074_ _0075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_34_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_25_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2231_ net25 net26 _1377_ _1378_ _1379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_40_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2300_ _1405_ _1407_ _1447_ _1448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_0_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2093_ _1185_ _1204_ _1247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_0_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2162_ _1176_ _1089_ _1314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2995_ _0030_ clknet_2_3__leaf_clk net106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1877_ _1023_ _1019_ _1031_ _1032_ _1033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_1946_ _1020_ _1102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2429_ _0123_ _0125_ _1169_ _0126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1488__A1 net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input22_I pcpi_rs1[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output90_I net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_8_Left_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1800_ _0943_ _0959_ _0960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2780_ _0326_ _0332_ _0468_ _0469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_40_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1731_ _0880_ _0884_ _0892_ _0893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_1662_ _0718_ _0825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2214_ _1164_ _1364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1593_ _0739_ _0742_ _0755_ _0756_ _0757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__2971__CLK clknet_2_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2145_ _1296_ _1297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2076_ net56 _1230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2434__A3 _0078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1929_ _1041_ _1084_ _1085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2978_ _0013_ clknet_2_2__leaf_clk net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_8_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_34_Left_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_54_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_27_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2994__CLK clknet_2_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2763_ _0394_ _0452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_42_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2901_ _0448_ _0594_ _0595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2832_ _0406_ _0436_ _0520_ _0521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_33_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2694_ _0370_ _0382_ _0383_ _0384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1576_ net76 _0740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1714_ _0844_ _0851_ _0876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_13_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1645_ _0808_ _0809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_6_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2059_ _0811_ _1214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2128_ _1225_ _1245_ _1281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1615__A1 _0777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput109 net109 pcpi_rd[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_37_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput91 net91 pcpi_rd[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_46_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2815_ _0464_ _0502_ _0503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2746_ _0412_ _0434_ _0435_ _0436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_18_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2677_ _0364_ _0365_ _0366_ _0367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_41_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1559_ _0722_ _0717_ _0723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1628_ _0787_ _0791_ _0792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_52_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_43_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_37_Left_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2600_ net34 _0290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_21_Left_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2462_ _0113_ _0149_ _0158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2531_ _0194_ _0223_ _0224_ _0225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2393_ _0038_ _0090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2555__A2 _0248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2729_ _0300_ _0419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_10_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input52_I pcpi_rs2[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_29_Right_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_52_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_38_Right_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_47_Right_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1962_ _1068_ _1118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_50_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1893_ net22 _1049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2514_ _0207_ _0208_ _0209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2445_ _1432_ _0140_ _0141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2376_ _0072_ _0073_ _0074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_3_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_54_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_25_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2230_ net62 _1378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_45_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2092_ _1185_ _1204_ _1246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_0_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2161_ _1128_ _1236_ _1313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_43_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2994_ _0029_ clknet_2_3__leaf_clk net104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1945_ _1100_ _1101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1876_ _1016_ _1028_ _1029_ net20 _1032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_2359_ _1379_ _1381_ _0055_ _1399_ _0057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_0_43_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2428_ _0072_ _0124_ _0125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input15_I pcpi_insn[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1730_ _0886_ _0888_ _0891_ _0892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_1592_ net40 _0744_ _0737_ net43 _0756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_0_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1661_ _0697_ _0823_ _0824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input7_I pcpi_insn[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2144_ _0811_ _1296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2213_ _1328_ _1361_ _1362_ _1349_ _1217_ _1363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_48_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1642__A2 net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2075_ _1227_ _1228_ _1229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1890__A2 _1045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2977_ _0012_ clknet_2_3__leaf_clk net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1928_ _1046_ _1070_ _1083_ _1084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_1859_ _1012_ _1009_ _1013_ _1014_ _1015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_35_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2900_ _0465_ _0594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_45_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2762_ _0393_ _0395_ _0451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2831_ _0334_ _0405_ _0520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_33_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1713_ _0871_ _0874_ _0875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2693_ _0369_ _0363_ _0367_ _0383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1644_ _0608_ _0807_ _0808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1575_ _0738_ _0739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_49_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2127_ _1264_ _1279_ _1280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_36_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2058_ _1169_ _1207_ _1210_ _1211_ _1212_ _1213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_8_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input82_I pcpi_valid vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput92 net92 pcpi_rd[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_53_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2270__A2 _1417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2676_ _0351_ _0353_ _0366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2814_ _0469_ _0476_ _0502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2745_ _0410_ _0411_ _0435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_26_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1489_ _0544_ _0555_ _0577_ _0587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_1558_ net46 _0722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1627_ _0788_ _0789_ _0790_ _0791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_49_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1772__A1 _0710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2530_ _0154_ _0189_ _0198_ _0224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_48_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2461_ _0155_ _0156_ _0157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2392_ _1432_ _0043_ _0089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2659_ net68 _0316_ _0349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2728_ _0378_ _0417_ _0418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA_input45_I pcpi_rs1[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2482__A2 _1297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1809__A2 _0783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2552__I _0587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2220__C _1008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2473__A2 _1417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1961_ _1086_ _1115_ _1116_ _1117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_1892_ net80 net23 _1048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2513_ _1464_ _1417_ _0208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2444_ _0092_ _0140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2375_ _0052_ _0071_ _0073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_3_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_54_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_49_Left_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_46_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2160_ _1271_ _1278_ _1311_ _1312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_48_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2091_ _1229_ _1244_ _1245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_TAPCELL_ROW_16_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2993_ _0028_ clknet_2_3__leaf_clk net103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1875_ _1030_ _1031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1944_ net51 _1100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2427_ _1478_ _0073_ _0124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_10_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2358_ _1391_ _1381_ _0055_ _1399_ _0056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2289_ net60 _1436_ _1437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_36_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1488__A3 net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1591_ _0754_ _0755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1660_ _0722_ _0823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2143_ _1295_ _0011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2212_ _1109_ _1113_ _1362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_36_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2074_ _1188_ _1203_ _1228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1927_ _1073_ _1082_ _1083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2976_ _0011_ clknet_2_2__leaf_clk net85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1858_ net53 _1014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1789_ _0917_ _0911_ _0921_ _0949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA_output114_I net114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2830_ _0505_ _0518_ _0519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_53_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2692_ _0366_ _0372_ _0373_ _0381_ _0382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_41_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2761_ _0336_ _0450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_38_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1643_ _0806_ _0807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_5_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1712_ _0824_ _0872_ _0873_ _0833_ _0822_ _0874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_6_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1574_ _0736_ _0737_ net29 net18 _0738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XTAP_TAPCELL_ROW_49_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2057_ _1163_ _1212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2126_ _1265_ _1271_ _1278_ _1279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2959_ _0651_ _0653_ _0654_ _0655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_32_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input75_I pcpi_rs2[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_35_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput93 net93 pcpi_rd[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_46_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2813_ _0496_ _0500_ _0501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_2675_ _0336_ _0338_ _0343_ _0365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_41_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2744_ _0416_ _0433_ _0434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1626_ _0717_ _0699_ _0790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2730__B2 _0322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1488_ net7 _0566_ net9 net8 _0577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_1557_ _0720_ _0711_ _0721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2109_ _1096_ _1260_ _1261_ _1262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_9_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2460_ _1423_ _1385_ _1387_ _0042_ _0156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2960__A1 _1168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2391_ _0035_ _0051_ _0087_ _0088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__2779__A1 _0374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2727_ net69 _0374_ _0417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2658_ _0345_ _0346_ _0347_ _0337_ _0348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2589_ net97 _0280_ _0281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1609_ _0771_ _0772_ _0773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_input38_I pcpi_rs1[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1960_ _1041_ _1084_ _1116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_7_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1891_ net51 net21 _1047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_52_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2512_ _0076_ _1433_ _0207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2443_ _0089_ _0137_ _0138_ _0098_ _0088_ _0139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XANTENNA__2974__CLK clknet_2_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2374_ _0052_ _0071_ _0072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_54_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_19_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2997__CLK clknet_2_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2090_ _1231_ _1235_ _1243_ _1244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_45_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2992_ _0027_ clknet_2_0__leaf_clk net102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_8_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1874_ net20 net19 _1028_ _1029_ _1030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_12_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1943_ _1074_ _1045_ _1099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2426_ _0099_ _0122_ _0123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_3_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2357_ _1398_ _0055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2288_ _1411_ _1436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_39_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2061__A1 net114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1590_ net43 net40 _0744_ _0737_ _0754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_0_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2142_ _1294_ net85 _0984_ _1295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2211_ _1354_ _1360_ _1361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2073_ _1189_ _1226_ _1227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2975_ _0010_ clknet_2_2__leaf_clk net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1926_ _1080_ _1081_ _1082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1857_ net54 _1013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1788_ _0715_ _0733_ _0948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2409_ _0105_ _0106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input20_I pcpi_rs1[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2691_ _0379_ _0380_ _0381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2760_ _0385_ _0448_ _0449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1642_ net4 net2 _0806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_26_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1711_ _0830_ _0832_ _0873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1573_ net76 _0737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_49_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2056_ _1159_ _1211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2125_ _1272_ _1274_ _1277_ _1278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_2958_ _0651_ _0653_ _1348_ _0654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_8_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1909_ net81 net23 _1065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input68_I pcpi_rs2[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2889_ net103 _0248_ _0582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput83 net83 pcpi_rd[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput94 net94 pcpi_rd[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_46_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2743_ _0431_ _0432_ _0433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2812_ _0498_ _0499_ _0500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_26_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2674_ _0355_ _0356_ _0361_ _0364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_41_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1625_ _0662_ _0670_ _0789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1556_ _0718_ _0715_ _0719_ _0720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_1487_ net6 _0566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_49_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2039_ _1142_ _1191_ _1192_ _1194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_2108_ _1235_ _1243_ _1261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_32_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_43_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2390_ _0037_ _0085_ _0086_ _0087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__1826__I1 net110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2726_ _0414_ _0415_ _0416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_13_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2657_ net67 _0347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2588_ _1296_ _0280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1608_ net44 net76 _0772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1539_ _0701_ _0702_ _0689_ _0703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_14_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2467__A1 _0052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_34_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_16_Right_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_50_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_25_Right_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1890_ _1043_ _1045_ _1046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2373_ _0053_ _0070_ _0071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2511_ _0180_ _0204_ _0205_ _0206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2442_ _0095_ _0097_ _0138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_11_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_34_Right_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_46_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_43_Right_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2709_ _0390_ _0363_ _0398_ _0399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_40_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_52_Right_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input50_I pcpi_rs2[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2603__A1 _0291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2991_ _0026_ clknet_2_3__leaf_clk net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1942_ _1035_ _1042_ _1098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_16_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1873_ net53 _1029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_10_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2356_ net65 _1383_ _0054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2425_ _0120_ _0121_ _0122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_2287_ _1419_ _1431_ _1434_ _1435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_42_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2749__I _0291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2210_ _1358_ _1359_ _1360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_28_Left_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2141_ _1165_ _0928_ _1293_ _1294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2072_ _1195_ _1202_ _1226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_44_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2974_ _0009_ clknet_2_3__leaf_clk net114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1925_ _1060_ _1061_ _1071_ _1081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_8_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_12_Left_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1856_ net49 _1012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1787_ _0945_ _0946_ _0947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2408_ _1398_ _0067_ _0064_ _0105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_41_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2339_ _1415_ _0036_ _0037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_2_Right_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_47_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input13_I pcpi_insn[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2690_ _0351_ _0353_ _0372_ _0380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_41_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1572_ net77 _0736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1710_ _0830_ _0832_ _0872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1641_ _0732_ _0776_ _0804_ _0805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA_input5_I pcpi_insn[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2124_ _1275_ _1276_ _1277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_49_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2055_ _1208_ _1209_ _1210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_44_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2957_ _0412_ _0652_ _0653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_32_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2888_ _0579_ _0580_ _0581_ _0027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_29_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1908_ net80 net24 _1064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_17_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1839_ _0988_ _0980_ _0994_ _0996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_37_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput95 net95 pcpi_rd[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput84 net84 pcpi_rd[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_46_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2742_ _0414_ _0415_ _0432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2811_ _0455_ _0458_ _0454_ _0499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2673_ _0344_ _0354_ _0362_ _0363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_41_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xpcpi_approx_mul_117 pcpi_wait vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_1_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1555_ _0675_ _0680_ _0719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1624_ net75 _0741_ _0788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1486_ net12 net10 net13 _0555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_2107_ _1230_ _1260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_49_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2038_ _1191_ _1192_ _1142_ _1193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XPHY_EDGE_ROW_15_Left_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input80_I pcpi_rs2[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1748__A1 _0671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_11_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2725_ _0379_ _0380_ _0415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2656_ net39 _0346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_42_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2587_ _0245_ _1362_ _0246_ _0279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1538_ _0678_ _0669_ _0702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1607_ net43 _0744_ _0771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_0_Left_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_13_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2510_ _0180_ _0204_ _1169_ _0205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_11_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2372_ _0054_ _0059_ _0069_ _0070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__2697__A2 _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2441_ _0095_ _0097_ _0137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2436__B _1323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2639_ net37 net71 _0329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_42_Left_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2708_ _0392_ _0397_ _0398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_6_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_2_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input43_I pcpi_rs1[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2679__A2 _0339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_45_Left_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_43_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2990_ _0025_ clknet_2_0__leaf_clk net100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_8_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1872_ net54 _1028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_16_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1941_ _1095_ _1096_ _1097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2119__A1 _1122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2355_ _1376_ _1402_ _0053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2424_ _0102_ _0103_ _0119_ _0121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_43_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2286_ _1432_ _1433_ _1430_ _1434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_47_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2597__A1 net98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2521__A1 _1323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2140_ _1008_ _1284_ _1291_ _1292_ _1212_ _1293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_2071_ _1220_ _1224_ _1225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_29_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2973_ _0008_ clknet_2_3__leaf_clk net113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1924_ _1078_ _1079_ _1080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1855_ _1010_ _1011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_24_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1786_ _0906_ _0907_ _0923_ _0946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2407_ _1417_ net65 _0104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2269_ _1416_ _1417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2338_ _1407_ _0036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_27_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2751__A1 _1300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1571_ _0734_ _0735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1640_ _0779_ _0802_ _0803_ _0804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_49_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2123_ _1131_ _1090_ _1276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2054_ _1095_ _1158_ _1209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2956_ _0410_ _0411_ _0652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_32_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2887_ net102 _0280_ _0581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1838_ _0988_ _0980_ _0994_ _0995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1907_ net51 _1049_ _1063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1769_ _0816_ _0700_ _0930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output112_I net112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput85 net85 pcpi_rd[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput96 net96 pcpi_rd[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_46_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2741_ _0418_ _0421_ _0430_ _0431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2672_ _0355_ _0356_ _0361_ _0362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2810_ _0385_ _0497_ _0498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1485_ net14 net82 _0512_ _0534_ _0544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__2977__CLK clknet_2_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1623_ _0690_ _0786_ _0787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1554_ _0717_ _0718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
.ends

